magic
tech sky130A
magscale 1 2
timestamp 1638662845
<< locali >>
rect 10517 8959 10551 9061
rect 12633 3927 12667 4029
rect 3525 3383 3559 3621
rect 10701 3451 10735 3689
rect 12081 1955 12115 2057
<< viali >>
rect 7297 10761 7331 10795
rect 10425 10761 10459 10795
rect 12081 10761 12115 10795
rect 14013 10761 14047 10795
rect 18153 10761 18187 10795
rect 7849 10693 7883 10727
rect 9045 10693 9079 10727
rect 17877 10693 17911 10727
rect 1501 10625 1535 10659
rect 3893 10625 3927 10659
rect 7481 10625 7515 10659
rect 7665 10625 7699 10659
rect 8861 10625 8895 10659
rect 9689 10625 9723 10659
rect 10609 10625 10643 10659
rect 11253 10625 11287 10659
rect 12449 10625 12483 10659
rect 13737 10625 13771 10659
rect 14197 10625 14231 10659
rect 15117 10625 15151 10659
rect 15669 10625 15703 10659
rect 16957 10625 16991 10659
rect 18061 10625 18095 10659
rect 18245 10625 18279 10659
rect 18521 10625 18555 10659
rect 3801 10557 3835 10591
rect 9137 10557 9171 10591
rect 11069 10557 11103 10591
rect 11161 10557 11195 10591
rect 12541 10557 12575 10591
rect 12725 10557 12759 10591
rect 8309 10489 8343 10523
rect 13277 10489 13311 10523
rect 18337 10489 18371 10523
rect 1501 10421 1535 10455
rect 3249 10421 3283 10455
rect 4261 10421 4295 10455
rect 8585 10421 8619 10455
rect 10333 10421 10367 10455
rect 11621 10421 11655 10455
rect 13553 10421 13587 10455
rect 14473 10421 14507 10455
rect 15025 10421 15059 10455
rect 16313 10421 16347 10455
rect 16957 10421 16991 10455
rect 3525 10217 3559 10251
rect 12817 10217 12851 10251
rect 15163 10217 15197 10251
rect 17831 10217 17865 10251
rect 8769 10149 8803 10183
rect 10701 10149 10735 10183
rect 12173 10149 12207 10183
rect 1317 10081 1351 10115
rect 1685 10081 1719 10115
rect 4721 10081 4755 10115
rect 5825 10081 5859 10115
rect 8953 10081 8987 10115
rect 13369 10081 13403 10115
rect 13737 10081 13771 10115
rect 16037 10081 16071 10115
rect 3341 10013 3375 10047
rect 3525 10013 3559 10047
rect 3709 10013 3743 10047
rect 4261 10013 4295 10047
rect 4445 10013 4479 10047
rect 4629 10013 4663 10047
rect 4813 10013 4847 10047
rect 4905 10013 4939 10047
rect 5089 10013 5123 10047
rect 5365 10013 5399 10047
rect 5549 10013 5583 10047
rect 6101 10013 6135 10047
rect 6469 10013 6503 10047
rect 8677 10013 8711 10047
rect 12909 10013 12943 10047
rect 16405 10013 16439 10047
rect 18245 10013 18279 10047
rect 18521 10013 18555 10047
rect 3111 9945 3145 9979
rect 4997 9945 5031 9979
rect 9229 9945 9263 9979
rect 10885 9945 10919 9979
rect 4445 9877 4479 9911
rect 5641 9877 5675 9911
rect 7895 9877 7929 9911
rect 8493 9877 8527 9911
rect 15761 9877 15795 9911
rect 15945 9877 15979 9911
rect 18337 9877 18371 9911
rect 2053 9673 2087 9707
rect 5457 9673 5491 9707
rect 5825 9673 5859 9707
rect 9321 9673 9355 9707
rect 12449 9673 12483 9707
rect 2605 9605 2639 9639
rect 2789 9605 2823 9639
rect 2973 9605 3007 9639
rect 3157 9605 3191 9639
rect 5365 9605 5399 9639
rect 5733 9605 5767 9639
rect 5917 9605 5951 9639
rect 6193 9605 6227 9639
rect 7297 9605 7331 9639
rect 8208 9605 8242 9639
rect 10057 9605 10091 9639
rect 14013 9605 14047 9639
rect 17509 9605 17543 9639
rect 2145 9537 2179 9571
rect 2329 9537 2363 9571
rect 2513 9537 2547 9571
rect 2881 9537 2915 9571
rect 3249 9537 3283 9571
rect 3433 9537 3467 9571
rect 4169 9537 4203 9571
rect 5181 9537 5215 9571
rect 5457 9537 5491 9571
rect 5641 9537 5675 9571
rect 6285 9537 6319 9571
rect 7757 9537 7791 9571
rect 10149 9537 10183 9571
rect 14841 9537 14875 9571
rect 15209 9537 15243 9571
rect 16635 9537 16669 9571
rect 16865 9537 16899 9571
rect 305 9469 339 9503
rect 581 9469 615 9503
rect 2237 9469 2271 9503
rect 4261 9469 4295 9503
rect 7941 9469 7975 9503
rect 10425 9469 10459 9503
rect 11897 9469 11931 9503
rect 14289 9469 14323 9503
rect 2513 9401 2547 9435
rect 3341 9401 3375 9435
rect 3617 9401 3651 9435
rect 3065 9333 3099 9367
rect 4445 9333 4479 9367
rect 6009 9333 6043 9367
rect 9781 9333 9815 9367
rect 12541 9333 12575 9367
rect 14657 9333 14691 9367
rect 1409 9129 1443 9163
rect 3065 9129 3099 9163
rect 10701 9129 10735 9163
rect 13277 9129 13311 9163
rect 10057 9061 10091 9095
rect 10517 9061 10551 9095
rect 1961 8993 1995 9027
rect 4629 8993 4663 9027
rect 5549 8993 5583 9027
rect 10885 8993 10919 9027
rect 13737 8993 13771 9027
rect 15485 8993 15519 9027
rect 15761 8993 15795 9027
rect 1501 8925 1535 8959
rect 2973 8925 3007 8959
rect 3157 8925 3191 8959
rect 4445 8925 4479 8959
rect 5365 8925 5399 8959
rect 6837 8925 6871 8959
rect 7104 8925 7138 8959
rect 8677 8925 8711 8959
rect 10149 8925 10183 8959
rect 10425 8925 10459 8959
rect 10517 8925 10551 8959
rect 11253 8925 11287 8959
rect 13461 8925 13495 8959
rect 16129 8925 16163 8959
rect 5457 8857 5491 8891
rect 8944 8857 8978 8891
rect 10241 8857 10275 8891
rect 4077 8789 4111 8823
rect 4537 8789 4571 8823
rect 4997 8789 5031 8823
rect 8217 8789 8251 8823
rect 10149 8789 10183 8823
rect 12679 8789 12713 8823
rect 17877 8789 17911 8823
rect 2145 8585 2179 8619
rect 4169 8585 4203 8619
rect 4905 8585 4939 8619
rect 5273 8585 5307 8619
rect 8953 8585 8987 8619
rect 9505 8585 9539 8619
rect 11069 8585 11103 8619
rect 11529 8585 11563 8619
rect 11621 8585 11655 8619
rect 14657 8585 14691 8619
rect 14887 8585 14921 8619
rect 18337 8585 18371 8619
rect 2513 8517 2547 8551
rect 3433 8517 3467 8551
rect 4261 8517 4295 8551
rect 6000 8517 6034 8551
rect 10977 8517 11011 8551
rect 13001 8517 13035 8551
rect 2145 8449 2179 8483
rect 2329 8449 2363 8483
rect 2697 8449 2731 8483
rect 2789 8449 2823 8483
rect 3341 8449 3375 8483
rect 7389 8449 7423 8483
rect 7573 8449 7607 8483
rect 7757 8449 7791 8483
rect 8493 8449 8527 8483
rect 9045 8449 9079 8483
rect 10793 8449 10827 8483
rect 11069 8449 11103 8483
rect 12265 8449 12299 8483
rect 12725 8449 12759 8483
rect 13369 8449 13403 8483
rect 14013 8449 14047 8483
rect 14197 8449 14231 8483
rect 16313 8449 16347 8483
rect 18521 8449 18555 8483
rect 305 8381 339 8415
rect 581 8381 615 8415
rect 2513 8381 2547 8415
rect 3617 8381 3651 8415
rect 4445 8381 4479 8415
rect 5365 8381 5399 8415
rect 5457 8381 5491 8415
rect 5733 8381 5767 8415
rect 7481 8381 7515 8415
rect 8033 8381 8067 8415
rect 11805 8381 11839 8415
rect 12541 8381 12575 8415
rect 13277 8381 13311 8415
rect 16681 8381 16715 8415
rect 18245 8381 18279 8415
rect 2053 8313 2087 8347
rect 3801 8313 3835 8347
rect 7113 8313 7147 8347
rect 11161 8313 11195 8347
rect 2973 8245 3007 8279
rect 7849 8245 7883 8279
rect 7941 8245 7975 8279
rect 8585 8245 8619 8279
rect 9321 8245 9355 8279
rect 12173 8245 12207 8279
rect 14013 8245 14047 8279
rect 2237 8041 2271 8075
rect 12449 8041 12483 8075
rect 13737 8041 13771 8075
rect 15117 8041 15151 8075
rect 15669 8041 15703 8075
rect 1869 7973 1903 8007
rect 5457 7973 5491 8007
rect 7665 7973 7699 8007
rect 7941 7973 7975 8007
rect 11897 7973 11931 8007
rect 2513 7905 2547 7939
rect 3249 7905 3283 7939
rect 5273 7905 5307 7939
rect 7297 7905 7331 7939
rect 7849 7905 7883 7939
rect 8493 7905 8527 7939
rect 11437 7905 11471 7939
rect 14289 7905 14323 7939
rect 15853 7905 15887 7939
rect 1961 7837 1995 7871
rect 2145 7837 2179 7871
rect 2329 7837 2363 7871
rect 2973 7837 3007 7871
rect 5549 7837 5583 7871
rect 6469 7837 6503 7871
rect 7481 7837 7515 7871
rect 8125 7837 8159 7871
rect 11529 7837 11563 7871
rect 12081 7837 12115 7871
rect 12173 7837 12207 7871
rect 12265 7837 12299 7871
rect 13001 7837 13035 7871
rect 14105 7837 14139 7871
rect 14565 7837 14599 7871
rect 14841 7837 14875 7871
rect 15025 7837 15059 7871
rect 5273 7769 5307 7803
rect 6193 7769 6227 7803
rect 6377 7769 6411 7803
rect 6653 7769 6687 7803
rect 8769 7769 8803 7803
rect 10517 7769 10551 7803
rect 13093 7769 13127 7803
rect 14197 7769 14231 7803
rect 16129 7769 16163 7803
rect 17877 7769 17911 7803
rect 2605 7701 2639 7735
rect 3065 7701 3099 7735
rect 8309 7701 8343 7735
rect 14657 7701 14691 7735
rect 15025 7701 15059 7735
rect 2237 7497 2271 7531
rect 4721 7497 4755 7531
rect 8953 7497 8987 7531
rect 10701 7497 10735 7531
rect 11345 7497 11379 7531
rect 11713 7497 11747 7531
rect 13737 7497 13771 7531
rect 13921 7497 13955 7531
rect 2605 7429 2639 7463
rect 2789 7429 2823 7463
rect 10609 7429 10643 7463
rect 14289 7429 14323 7463
rect 14519 7429 14553 7463
rect 2145 7361 2179 7395
rect 2329 7361 2363 7395
rect 3433 7361 3467 7395
rect 4077 7361 4111 7395
rect 4261 7361 4295 7395
rect 4353 7361 4387 7395
rect 4445 7361 4479 7395
rect 5089 7361 5123 7395
rect 5365 7361 5399 7395
rect 5457 7361 5491 7395
rect 5825 7361 5859 7395
rect 7757 7361 7791 7395
rect 7849 7361 7883 7395
rect 8861 7361 8895 7395
rect 10241 7361 10275 7395
rect 10425 7361 10459 7395
rect 10885 7361 10919 7395
rect 11161 7361 11195 7395
rect 11437 7361 11471 7395
rect 11621 7361 11655 7395
rect 11897 7361 11931 7395
rect 13461 7361 13495 7395
rect 13645 7361 13679 7395
rect 13735 7383 13769 7417
rect 13829 7361 13863 7395
rect 14105 7361 14139 7395
rect 305 7293 339 7327
rect 581 7293 615 7327
rect 2973 7293 3007 7327
rect 5733 7293 5767 7327
rect 6193 7293 6227 7327
rect 8033 7293 8067 7327
rect 9045 7293 9079 7327
rect 10333 7293 10367 7327
rect 15945 7293 15979 7327
rect 16313 7293 16347 7327
rect 2053 7225 2087 7259
rect 10149 7225 10183 7259
rect 5549 7157 5583 7191
rect 7389 7157 7423 7191
rect 8309 7157 8343 7191
rect 8493 7157 8527 7191
rect 10977 7157 11011 7191
rect 2145 6953 2179 6987
rect 6929 6953 6963 6987
rect 15945 6953 15979 6987
rect 16129 6953 16163 6987
rect 17619 6953 17653 6987
rect 18337 6953 18371 6987
rect 3985 6885 4019 6919
rect 3433 6817 3467 6851
rect 4629 6817 4663 6851
rect 6561 6817 6595 6851
rect 7573 6817 7607 6851
rect 8217 6817 8251 6851
rect 8493 6817 8527 6851
rect 11437 6817 11471 6851
rect 11713 6817 11747 6851
rect 13829 6817 13863 6851
rect 14657 6817 14691 6851
rect 15393 6817 15427 6851
rect 2697 6749 2731 6783
rect 2881 6749 2915 6783
rect 3065 6749 3099 6783
rect 3157 6749 3191 6783
rect 3341 6749 3375 6783
rect 4261 6749 4295 6783
rect 4813 6749 4847 6783
rect 5089 6749 5123 6783
rect 5641 6749 5675 6783
rect 5733 6749 5767 6783
rect 6653 6749 6687 6783
rect 8125 6749 8159 6783
rect 10241 6749 10275 6783
rect 10609 6749 10643 6783
rect 11805 6749 11839 6783
rect 12725 6749 12759 6783
rect 14381 6749 14415 6783
rect 15117 6749 15151 6783
rect 17877 6749 17911 6783
rect 18245 6749 18279 6783
rect 18521 6749 18555 6783
rect 2789 6681 2823 6715
rect 5917 6681 5951 6715
rect 7297 6681 7331 6715
rect 10333 6681 10367 6715
rect 10517 6681 10551 6715
rect 11345 6681 11379 6715
rect 13645 6681 13679 6715
rect 2513 6613 2547 6647
rect 5825 6613 5859 6647
rect 6193 6613 6227 6647
rect 6837 6613 6871 6647
rect 7389 6613 7423 6647
rect 7757 6613 7791 6647
rect 10425 6613 10459 6647
rect 10885 6613 10919 6647
rect 11253 6613 11287 6647
rect 12541 6613 12575 6647
rect 13277 6613 13311 6647
rect 13737 6613 13771 6647
rect 14749 6613 14783 6647
rect 15209 6613 15243 6647
rect 2145 6409 2179 6443
rect 2881 6409 2915 6443
rect 3709 6409 3743 6443
rect 5273 6409 5307 6443
rect 5917 6409 5951 6443
rect 6653 6409 6687 6443
rect 6745 6409 6779 6443
rect 10333 6409 10367 6443
rect 11897 6409 11931 6443
rect 14565 6409 14599 6443
rect 15393 6409 15427 6443
rect 16865 6409 16899 6443
rect 17233 6409 17267 6443
rect 17693 6409 17727 6443
rect 18061 6409 18095 6443
rect 5825 6341 5859 6375
rect 9505 6341 9539 6375
rect 11437 6341 11471 6375
rect 12357 6341 12391 6375
rect 14013 6341 14047 6375
rect 2605 6273 2639 6307
rect 2789 6273 2823 6307
rect 3249 6273 3283 6307
rect 3433 6273 3467 6307
rect 3617 6273 3651 6307
rect 4169 6273 4203 6307
rect 5733 6273 5767 6307
rect 6009 6273 6043 6307
rect 9689 6273 9723 6307
rect 9873 6273 9907 6307
rect 12081 6273 12115 6307
rect 14289 6273 14323 6307
rect 14565 6273 14599 6307
rect 14749 6273 14783 6307
rect 15301 6273 15335 6307
rect 15761 6273 15795 6307
rect 16681 6273 16715 6307
rect 305 6205 339 6239
rect 581 6205 615 6239
rect 2053 6205 2087 6239
rect 3065 6205 3099 6239
rect 3157 6205 3191 6239
rect 5365 6205 5399 6239
rect 5457 6205 5491 6239
rect 6561 6205 6595 6239
rect 10149 6205 10183 6239
rect 10241 6205 10275 6239
rect 10977 6205 11011 6239
rect 11069 6205 11103 6239
rect 13829 6205 13863 6239
rect 15669 6205 15703 6239
rect 17325 6205 17359 6239
rect 17509 6205 17543 6239
rect 18153 6205 18187 6239
rect 18337 6205 18371 6239
rect 2789 6137 2823 6171
rect 4905 6137 4939 6171
rect 7113 6137 7147 6171
rect 9873 6137 9907 6171
rect 10701 6137 10735 6171
rect 14197 6137 14231 6171
rect 3893 6069 3927 6103
rect 4077 6069 4111 6103
rect 8217 6069 8251 6103
rect 10793 6069 10827 6103
rect 14105 6069 14139 6103
rect 16497 6069 16531 6103
rect 2421 5865 2455 5899
rect 3525 5865 3559 5899
rect 3893 5865 3927 5899
rect 4340 5865 4374 5899
rect 5825 5865 5859 5899
rect 7895 5865 7929 5899
rect 8217 5865 8251 5899
rect 8953 5865 8987 5899
rect 11437 5865 11471 5899
rect 15853 5865 15887 5899
rect 17831 5865 17865 5899
rect 18245 5865 18279 5899
rect 3433 5797 3467 5831
rect 3709 5729 3743 5763
rect 4077 5729 4111 5763
rect 6101 5729 6135 5763
rect 6469 5729 6503 5763
rect 10425 5729 10459 5763
rect 10701 5729 10735 5763
rect 11161 5729 11195 5763
rect 14289 5729 14323 5763
rect 14749 5729 14783 5763
rect 16405 5729 16439 5763
rect 949 5661 983 5695
rect 2605 5661 2639 5695
rect 2881 5661 2915 5695
rect 3065 5661 3099 5695
rect 3985 5661 4019 5695
rect 8217 5661 8251 5695
rect 11069 5661 11103 5695
rect 14381 5661 14415 5695
rect 16037 5661 16071 5695
rect 18061 5661 18095 5695
rect 581 5593 615 5627
rect 2789 5525 2823 5559
rect 3709 5525 3743 5559
rect 8769 5525 8803 5559
rect 2513 5321 2547 5355
rect 2881 5321 2915 5355
rect 9781 5321 9815 5355
rect 10425 5321 10459 5355
rect 12081 5321 12115 5355
rect 6653 5253 6687 5287
rect 10333 5253 10367 5287
rect 10701 5253 10735 5287
rect 11897 5253 11931 5287
rect 13553 5253 13587 5287
rect 14841 5253 14875 5287
rect 489 5185 523 5219
rect 2283 5185 2317 5219
rect 2789 5185 2823 5219
rect 6469 5185 6503 5219
rect 7573 5185 7607 5219
rect 10609 5185 10643 5219
rect 10793 5185 10827 5219
rect 14933 5185 14967 5219
rect 18245 5185 18279 5219
rect 18521 5185 18555 5219
rect 857 5117 891 5151
rect 7849 5117 7883 5151
rect 13829 5117 13863 5151
rect 15209 5117 15243 5151
rect 18337 5049 18371 5083
rect 3617 4981 3651 5015
rect 3893 4981 3927 5015
rect 5917 4981 5951 5015
rect 7389 4981 7423 5015
rect 9321 4981 9355 5015
rect 16681 4981 16715 5015
rect 13277 4777 13311 4811
rect 3433 4709 3467 4743
rect 10885 4709 10919 4743
rect 15669 4709 15703 4743
rect 2973 4641 3007 4675
rect 3709 4641 3743 4675
rect 7113 4641 7147 4675
rect 8953 4641 8987 4675
rect 9413 4641 9447 4675
rect 11345 4641 11379 4675
rect 11437 4641 11471 4675
rect 14749 4641 14783 4675
rect 15025 4641 15059 4675
rect 16129 4641 16163 4675
rect 17877 4641 17911 4675
rect 3065 4573 3099 4607
rect 4077 4573 4111 4607
rect 6285 4573 6319 4607
rect 6377 4573 6411 4607
rect 7021 4573 7055 4607
rect 9045 4573 9079 4607
rect 11713 4573 11747 4607
rect 15117 4573 15151 4607
rect 15853 4573 15887 4607
rect 5503 4505 5537 4539
rect 11253 4505 11287 4539
rect 11958 4505 11992 4539
rect 15228 4505 15262 4539
rect 15393 4505 15427 4539
rect 6101 4437 6135 4471
rect 6745 4437 6779 4471
rect 7389 4437 7423 4471
rect 13093 4437 13127 4471
rect 15117 4437 15151 4471
rect 2329 4233 2363 4267
rect 2973 4233 3007 4267
rect 7665 4233 7699 4267
rect 8585 4233 8619 4267
rect 9137 4233 9171 4267
rect 9689 4233 9723 4267
rect 10057 4233 10091 4267
rect 11253 4233 11287 4267
rect 12725 4233 12759 4267
rect 13553 4233 13587 4267
rect 14289 4233 14323 4267
rect 3433 4165 3467 4199
rect 2605 4097 2639 4131
rect 2697 4097 2731 4131
rect 2789 4097 2823 4131
rect 3985 4097 4019 4131
rect 4905 4097 4939 4131
rect 6699 4097 6733 4131
rect 8493 4097 8527 4131
rect 8677 4097 8711 4131
rect 10149 4097 10183 4131
rect 11161 4097 11195 4131
rect 11345 4097 11379 4131
rect 12909 4097 12943 4131
rect 13185 4097 13219 4131
rect 13369 4097 13403 4131
rect 13829 4097 13863 4131
rect 18245 4097 18279 4131
rect 18521 4097 18555 4131
rect 305 4029 339 4063
rect 673 4029 707 4063
rect 2145 4029 2179 4063
rect 3525 4029 3559 4063
rect 3617 4029 3651 4063
rect 5273 4029 5307 4063
rect 7757 4029 7791 4063
rect 7941 4029 7975 4063
rect 9229 4029 9263 4063
rect 9413 4029 9447 4063
rect 10241 4029 10275 4063
rect 12633 4029 12667 4063
rect 13093 4029 13127 4063
rect 14657 4029 14691 4063
rect 14841 4029 14875 4063
rect 15209 4029 15243 4063
rect 3893 3961 3927 3995
rect 14473 3961 14507 3995
rect 18337 3961 18371 3995
rect 3065 3893 3099 3927
rect 4629 3893 4663 3927
rect 7297 3893 7331 3927
rect 8769 3893 8803 3927
rect 12633 3893 12667 3927
rect 13185 3893 13219 3927
rect 14105 3893 14139 3927
rect 16635 3893 16669 3927
rect 857 3689 891 3723
rect 6285 3689 6319 3723
rect 8493 3689 8527 3723
rect 10701 3689 10735 3723
rect 13645 3689 13679 3723
rect 15209 3689 15243 3723
rect 15393 3689 15427 3723
rect 3525 3621 3559 3655
rect 5917 3621 5951 3655
rect 2237 3553 2271 3587
rect 1041 3485 1075 3519
rect 1961 3485 1995 3519
rect 3065 3485 3099 3519
rect 3249 3485 3283 3519
rect 2053 3417 2087 3451
rect 6745 3553 6779 3587
rect 6929 3553 6963 3587
rect 8769 3553 8803 3587
rect 5917 3485 5951 3519
rect 6653 3485 6687 3519
rect 8677 3485 8711 3519
rect 9229 3485 9263 3519
rect 9597 3485 9631 3519
rect 9781 3485 9815 3519
rect 10241 3485 10275 3519
rect 10517 3485 10551 3519
rect 11253 3621 11287 3655
rect 12449 3621 12483 3655
rect 13001 3621 13035 3655
rect 12265 3553 12299 3587
rect 13093 3553 13127 3587
rect 16129 3553 16163 3587
rect 17509 3553 17543 3587
rect 12541 3485 12575 3519
rect 12817 3485 12851 3519
rect 13461 3485 13495 3519
rect 13737 3485 13771 3519
rect 13829 3485 13863 3519
rect 15761 3485 15795 3519
rect 18245 3485 18279 3519
rect 5641 3417 5675 3451
rect 5825 3417 5859 3451
rect 9321 3417 9355 3451
rect 9505 3417 9539 3451
rect 10333 3417 10367 3451
rect 10701 3417 10735 3451
rect 10885 3417 10919 3451
rect 11529 3417 11563 3451
rect 13277 3417 13311 3451
rect 14096 3417 14130 3451
rect 18061 3417 18095 3451
rect 1593 3349 1627 3383
rect 2421 3349 2455 3383
rect 3157 3349 3191 3383
rect 3433 3349 3467 3383
rect 3525 3349 3559 3383
rect 7297 3349 7331 3383
rect 9137 3349 9171 3383
rect 9229 3349 9263 3383
rect 9689 3349 9723 3383
rect 10241 3349 10275 3383
rect 11345 3349 11379 3383
rect 12265 3349 12299 3383
rect 12633 3349 12667 3383
rect 2237 3145 2271 3179
rect 3157 3145 3191 3179
rect 3709 3145 3743 3179
rect 5549 3145 5583 3179
rect 5641 3145 5675 3179
rect 6745 3145 6779 3179
rect 7297 3145 7331 3179
rect 7757 3145 7791 3179
rect 8585 3145 8619 3179
rect 10425 3145 10459 3179
rect 12081 3145 12115 3179
rect 15853 3145 15887 3179
rect 15945 3145 15979 3179
rect 5273 3077 5307 3111
rect 5457 3077 5491 3111
rect 6837 3077 6871 3111
rect 12541 3077 12575 3111
rect 14718 3077 14752 3111
rect 16497 3077 16531 3111
rect 305 3009 339 3043
rect 2789 3009 2823 3043
rect 3617 3009 3651 3043
rect 5549 3009 5583 3043
rect 7665 3009 7699 3043
rect 8125 3009 8159 3043
rect 8309 3009 8343 3043
rect 8861 3009 8895 3043
rect 9045 3009 9079 3043
rect 10057 3009 10091 3043
rect 10241 3009 10275 3043
rect 10609 3009 10643 3043
rect 10701 3009 10735 3043
rect 10793 3009 10827 3043
rect 11161 3009 11195 3043
rect 11437 3009 11471 3043
rect 11897 3009 11931 3043
rect 12265 3009 12299 3043
rect 14473 3009 14507 3043
rect 16405 3009 16439 3043
rect 581 2941 615 2975
rect 2697 2941 2731 2975
rect 3801 2941 3835 2975
rect 6009 2941 6043 2975
rect 6101 2941 6135 2975
rect 7021 2941 7055 2975
rect 7941 2941 7975 2975
rect 8953 2941 8987 2975
rect 11713 2941 11747 2975
rect 14289 2941 14323 2975
rect 3249 2873 3283 2907
rect 6377 2873 6411 2907
rect 2053 2805 2087 2839
rect 6285 2805 6319 2839
rect 16129 2805 16163 2839
rect 765 2601 799 2635
rect 2789 2601 2823 2635
rect 3157 2601 3191 2635
rect 3341 2601 3375 2635
rect 4169 2601 4203 2635
rect 7113 2601 7147 2635
rect 11069 2601 11103 2635
rect 2605 2533 2639 2567
rect 8769 2533 8803 2567
rect 11345 2533 11379 2567
rect 11529 2533 11563 2567
rect 15669 2533 15703 2567
rect 2053 2465 2087 2499
rect 2237 2465 2271 2499
rect 2421 2465 2455 2499
rect 5917 2465 5951 2499
rect 8861 2465 8895 2499
rect 15209 2465 15243 2499
rect 15853 2465 15887 2499
rect 17877 2465 17911 2499
rect 949 2397 983 2431
rect 2697 2397 2731 2431
rect 2789 2397 2823 2431
rect 2973 2397 3007 2431
rect 6377 2397 6411 2431
rect 9229 2397 9263 2431
rect 10885 2397 10919 2431
rect 11069 2397 11103 2431
rect 11437 2397 11471 2431
rect 15025 2397 15059 2431
rect 15393 2397 15427 2431
rect 18245 2397 18279 2431
rect 18521 2397 18555 2431
rect 1961 2329 1995 2363
rect 3985 2329 4019 2363
rect 5641 2329 5675 2363
rect 7205 2329 7239 2363
rect 8585 2329 8619 2363
rect 10655 2329 10689 2363
rect 16129 2329 16163 2363
rect 1593 2261 1627 2295
rect 2697 2261 2731 2295
rect 6193 2261 6227 2295
rect 8309 2261 8343 2295
rect 14565 2261 14599 2295
rect 14933 2261 14967 2295
rect 18337 2261 18371 2295
rect 2053 2057 2087 2091
rect 9137 2057 9171 2091
rect 11437 2057 11471 2091
rect 12081 2057 12115 2091
rect 12265 2057 12299 2091
rect 12633 2057 12667 2091
rect 13093 2057 13127 2091
rect 13553 2057 13587 2091
rect 16681 2057 16715 2091
rect 17325 2057 17359 2091
rect 18153 2057 18187 2091
rect 6101 1989 6135 2023
rect 9781 1989 9815 2023
rect 10057 1989 10091 2023
rect 15209 1989 15243 2023
rect 2881 1921 2915 1955
rect 3525 1921 3559 1955
rect 3709 1921 3743 1955
rect 4721 1921 4755 1955
rect 5273 1921 5307 1955
rect 5365 1921 5399 1955
rect 5457 1921 5491 1955
rect 6561 1921 6595 1955
rect 6745 1921 6779 1955
rect 6837 1921 6871 1955
rect 7297 1921 7331 1955
rect 7481 1921 7515 1955
rect 7573 1921 7607 1955
rect 8953 1921 8987 1955
rect 9229 1921 9263 1955
rect 9865 1911 9899 1945
rect 9965 1921 9999 1955
rect 10149 1921 10183 1955
rect 11069 1921 11103 1955
rect 11713 1921 11747 1955
rect 11897 1921 11931 1955
rect 12081 1921 12115 1955
rect 12725 1921 12759 1955
rect 13461 1921 13495 1955
rect 13921 1921 13955 1955
rect 14105 1921 14139 1955
rect 14289 1921 14323 1955
rect 14841 1921 14875 1955
rect 17233 1921 17267 1955
rect 18245 1921 18279 1955
rect 305 1853 339 1887
rect 581 1853 615 1887
rect 2513 1853 2547 1887
rect 2789 1853 2823 1887
rect 3985 1853 4019 1887
rect 10977 1853 11011 1887
rect 12817 1853 12851 1887
rect 13737 1853 13771 1887
rect 14197 1853 14231 1887
rect 14565 1853 14599 1887
rect 14933 1853 14967 1887
rect 17417 1853 17451 1887
rect 4353 1785 4387 1819
rect 8401 1785 8435 1819
rect 14657 1785 14691 1819
rect 16865 1785 16899 1819
rect 2237 1717 2271 1751
rect 3249 1717 3283 1751
rect 4445 1717 4479 1751
rect 4629 1717 4663 1751
rect 5641 1717 5675 1751
rect 8677 1717 8711 1751
rect 11805 1717 11839 1751
rect 14749 1717 14783 1751
rect 10609 1513 10643 1547
rect 14565 1513 14599 1547
rect 14749 1513 14783 1547
rect 3525 1445 3559 1479
rect 7205 1445 7239 1479
rect 7941 1445 7975 1479
rect 2053 1377 2087 1411
rect 3709 1377 3743 1411
rect 3893 1377 3927 1411
rect 3985 1377 4019 1411
rect 5181 1377 5215 1411
rect 8493 1377 8527 1411
rect 15301 1377 15335 1411
rect 1777 1309 1811 1343
rect 4905 1309 4939 1343
rect 5457 1309 5491 1343
rect 5641 1309 5675 1343
rect 5917 1309 5951 1343
rect 7021 1309 7055 1343
rect 7205 1309 7239 1343
rect 7481 1309 7515 1343
rect 8861 1309 8895 1343
rect 10287 1309 10321 1343
rect 12633 1309 12667 1343
rect 13369 1309 13403 1343
rect 13553 1309 13587 1343
rect 14473 1309 14507 1343
rect 15117 1309 15151 1343
rect 15209 1309 15243 1343
rect 15761 1309 15795 1343
rect 15945 1309 15979 1343
rect 16037 1309 16071 1343
rect 16405 1309 16439 1343
rect 4537 1241 4571 1275
rect 6837 1241 6871 1275
rect 12357 1241 12391 1275
rect 17877 1241 17911 1275
rect 4353 1173 4387 1207
rect 5365 1173 5399 1207
rect 5825 1173 5859 1207
rect 8217 1173 8251 1207
rect 10885 1173 10919 1207
rect 13369 1173 13403 1207
rect 15853 1173 15887 1207
rect 4307 969 4341 1003
rect 4997 969 5031 1003
rect 7113 969 7147 1003
rect 7389 969 7423 1003
rect 9413 969 9447 1003
rect 11805 969 11839 1003
rect 12265 969 12299 1003
rect 14565 969 14599 1003
rect 16681 969 16715 1003
rect 17049 969 17083 1003
rect 17509 969 17543 1003
rect 18337 969 18371 1003
rect 9137 901 9171 935
rect 11529 901 11563 935
rect 15025 901 15059 935
rect 2513 833 2547 867
rect 4629 833 4663 867
rect 4721 833 4755 867
rect 4905 833 4939 867
rect 5089 833 5123 867
rect 5365 833 5399 867
rect 7297 833 7331 867
rect 7481 833 7515 867
rect 7573 833 7607 867
rect 7757 833 7791 867
rect 8217 833 8251 867
rect 8493 833 8527 867
rect 8769 833 8803 867
rect 9045 833 9079 867
rect 9321 833 9355 867
rect 9965 833 9999 867
rect 10149 833 10183 867
rect 10425 833 10459 867
rect 11713 833 11747 867
rect 11805 833 11839 867
rect 12081 833 12115 867
rect 12265 833 12299 867
rect 12541 833 12575 867
rect 13001 833 13035 867
rect 13185 833 13219 867
rect 13737 833 13771 867
rect 17417 833 17451 867
rect 18245 833 18279 867
rect 18521 833 18555 867
rect 2881 765 2915 799
rect 4445 765 4479 799
rect 5641 765 5675 799
rect 12633 765 12667 799
rect 14289 765 14323 799
rect 14749 765 14783 799
rect 17601 765 17635 799
rect 4537 697 4571 731
rect 7757 697 7791 731
rect 8033 697 8067 731
rect 8585 697 8619 731
rect 9689 697 9723 731
rect 10333 697 10367 731
rect 12909 697 12943 731
rect 2329 629 2363 663
rect 5273 629 5307 663
rect 9229 629 9263 663
rect 9965 629 9999 663
rect 16497 629 16531 663
rect 5549 425 5583 459
rect 6193 425 6227 459
rect 9137 425 9171 459
rect 13461 425 13495 459
rect 13553 425 13587 459
rect 15669 425 15703 459
rect 16221 425 16255 459
rect 17325 425 17359 459
rect 5457 357 5491 391
rect 12265 357 12299 391
rect 15945 357 15979 391
rect 16957 289 16991 323
rect 5365 221 5399 255
rect 5917 221 5951 255
rect 6101 221 6135 255
rect 6285 221 6319 255
rect 9137 221 9171 255
rect 9229 221 9263 255
rect 12081 221 12115 255
rect 12357 221 12391 255
rect 13277 221 13311 255
rect 13461 221 13495 255
rect 13553 221 13587 255
rect 13737 221 13771 255
rect 15853 221 15887 255
rect 16037 221 16071 255
rect 16221 221 16255 255
rect 17049 221 17083 255
rect 9413 153 9447 187
rect 12173 153 12207 187
rect 5825 85 5859 119
<< metal1 >>
rect 0 10906 18860 10928
rect 0 10854 4660 10906
rect 4712 10854 4724 10906
rect 4776 10854 4788 10906
rect 4840 10854 4852 10906
rect 4904 10854 4916 10906
rect 4968 10854 7760 10906
rect 7812 10854 7824 10906
rect 7876 10854 7888 10906
rect 7940 10854 7952 10906
rect 8004 10854 8016 10906
rect 8068 10854 10860 10906
rect 10912 10854 10924 10906
rect 10976 10854 10988 10906
rect 11040 10854 11052 10906
rect 11104 10854 11116 10906
rect 11168 10854 13960 10906
rect 14012 10854 14024 10906
rect 14076 10854 14088 10906
rect 14140 10854 14152 10906
rect 14204 10854 14216 10906
rect 14268 10854 17060 10906
rect 17112 10854 17124 10906
rect 17176 10854 17188 10906
rect 17240 10854 17252 10906
rect 17304 10854 17316 10906
rect 17368 10854 18860 10906
rect 0 10832 18860 10854
rect 7098 10752 7104 10804
rect 7156 10792 7162 10804
rect 7285 10795 7343 10801
rect 7285 10792 7297 10795
rect 7156 10764 7297 10792
rect 7156 10752 7162 10764
rect 7285 10761 7297 10764
rect 7331 10761 7343 10795
rect 7285 10755 7343 10761
rect 7484 10764 9904 10792
rect 290 10616 296 10668
rect 348 10656 354 10668
rect 1489 10659 1547 10665
rect 1489 10656 1501 10659
rect 348 10628 1501 10656
rect 348 10616 354 10628
rect 1489 10625 1501 10628
rect 1535 10625 1547 10659
rect 1489 10619 1547 10625
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10656 3939 10659
rect 4154 10656 4160 10668
rect 3927 10628 4160 10656
rect 3927 10625 3939 10628
rect 3881 10619 3939 10625
rect 4154 10616 4160 10628
rect 4212 10616 4218 10668
rect 7484 10665 7512 10764
rect 7837 10727 7895 10733
rect 7837 10693 7849 10727
rect 7883 10724 7895 10727
rect 9033 10727 9091 10733
rect 9033 10724 9045 10727
rect 7883 10696 9045 10724
rect 7883 10693 7895 10696
rect 7837 10687 7895 10693
rect 9033 10693 9045 10696
rect 9079 10693 9091 10727
rect 9876 10724 9904 10764
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10413 10795 10471 10801
rect 10413 10792 10425 10795
rect 10008 10764 10425 10792
rect 10008 10752 10014 10764
rect 10413 10761 10425 10764
rect 10459 10761 10471 10795
rect 12069 10795 12127 10801
rect 12069 10792 12081 10795
rect 10413 10755 10471 10761
rect 10520 10764 12081 10792
rect 10520 10724 10548 10764
rect 12069 10761 12081 10764
rect 12115 10792 12127 10795
rect 12115 10764 12434 10792
rect 12115 10761 12127 10764
rect 12069 10755 12127 10761
rect 11330 10724 11336 10736
rect 9876 10696 10548 10724
rect 10612 10696 11336 10724
rect 9033 10687 9091 10693
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10625 7527 10659
rect 7650 10656 7656 10668
rect 7611 10628 7656 10656
rect 7469 10619 7527 10625
rect 7650 10616 7656 10628
rect 7708 10616 7714 10668
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10656 8907 10659
rect 8938 10656 8944 10668
rect 8895 10628 8944 10656
rect 8895 10625 8907 10628
rect 8849 10619 8907 10625
rect 8938 10616 8944 10628
rect 8996 10656 9002 10668
rect 10612 10665 10640 10696
rect 11330 10684 11336 10696
rect 11388 10684 11394 10736
rect 12406 10724 12434 10764
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 14001 10795 14059 10801
rect 14001 10792 14013 10795
rect 12860 10764 14013 10792
rect 12860 10752 12866 10764
rect 14001 10761 14013 10764
rect 14047 10761 14059 10795
rect 18141 10795 18199 10801
rect 18141 10792 18153 10795
rect 14001 10755 14059 10761
rect 14200 10764 18153 10792
rect 12406 10696 13768 10724
rect 9677 10659 9735 10665
rect 9677 10656 9689 10659
rect 8996 10628 9689 10656
rect 8996 10616 9002 10628
rect 9677 10625 9689 10628
rect 9723 10625 9735 10659
rect 9677 10619 9735 10625
rect 10597 10659 10655 10665
rect 10597 10625 10609 10659
rect 10643 10625 10655 10659
rect 11238 10656 11244 10668
rect 11199 10628 11244 10656
rect 10597 10619 10655 10625
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 13740 10665 13768 10696
rect 14200 10665 14228 10764
rect 18141 10761 18153 10764
rect 18187 10761 18199 10795
rect 18141 10755 18199 10761
rect 17865 10727 17923 10733
rect 17865 10693 17877 10727
rect 17911 10724 17923 10727
rect 17911 10696 18552 10724
rect 17911 10693 17923 10696
rect 17865 10687 17923 10693
rect 12437 10659 12495 10665
rect 12437 10656 12449 10659
rect 11624 10628 12449 10656
rect 3510 10548 3516 10600
rect 3568 10588 3574 10600
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 3568 10560 3801 10588
rect 3568 10548 3574 10560
rect 3789 10557 3801 10560
rect 3835 10557 3847 10591
rect 8754 10588 8760 10600
rect 3789 10551 3847 10557
rect 8312 10560 8760 10588
rect 2682 10480 2688 10532
rect 2740 10520 2746 10532
rect 7006 10520 7012 10532
rect 2740 10480 2774 10520
rect 1302 10412 1308 10464
rect 1360 10452 1366 10464
rect 1489 10455 1547 10461
rect 1489 10452 1501 10455
rect 1360 10424 1501 10452
rect 1360 10412 1366 10424
rect 1489 10421 1501 10424
rect 1535 10421 1547 10455
rect 2746 10452 2774 10480
rect 3252 10492 7012 10520
rect 3252 10461 3280 10492
rect 7006 10480 7012 10492
rect 7064 10520 7070 10532
rect 8312 10529 8340 10560
rect 8754 10548 8760 10560
rect 8812 10588 8818 10600
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 8812 10560 9137 10588
rect 8812 10548 8818 10560
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 11054 10588 11060 10600
rect 11015 10560 11060 10588
rect 9125 10551 9183 10557
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 11149 10591 11207 10597
rect 11149 10557 11161 10591
rect 11195 10557 11207 10591
rect 11149 10551 11207 10557
rect 8297 10523 8355 10529
rect 8297 10520 8309 10523
rect 7064 10492 8309 10520
rect 7064 10480 7070 10492
rect 8297 10489 8309 10492
rect 8343 10489 8355 10523
rect 8297 10483 8355 10489
rect 10686 10480 10692 10532
rect 10744 10520 10750 10532
rect 11164 10520 11192 10551
rect 10744 10492 11192 10520
rect 10744 10480 10750 10492
rect 3237 10455 3295 10461
rect 3237 10452 3249 10455
rect 2746 10424 3249 10452
rect 1489 10415 1547 10421
rect 3237 10421 3249 10424
rect 3283 10421 3295 10455
rect 3237 10415 3295 10421
rect 4249 10455 4307 10461
rect 4249 10421 4261 10455
rect 4295 10452 4307 10455
rect 4430 10452 4436 10464
rect 4295 10424 4436 10452
rect 4295 10421 4307 10424
rect 4249 10415 4307 10421
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 8573 10455 8631 10461
rect 8573 10421 8585 10455
rect 8619 10452 8631 10455
rect 8662 10452 8668 10464
rect 8619 10424 8668 10452
rect 8619 10421 8631 10424
rect 8573 10415 8631 10421
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 10321 10455 10379 10461
rect 10321 10452 10333 10455
rect 9272 10424 10333 10452
rect 9272 10412 9278 10424
rect 10321 10421 10333 10424
rect 10367 10421 10379 10455
rect 10321 10415 10379 10421
rect 11514 10412 11520 10464
rect 11572 10452 11578 10464
rect 11624 10461 11652 10628
rect 12437 10625 12449 10628
rect 12483 10625 12495 10659
rect 12437 10619 12495 10625
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10625 13783 10659
rect 13725 10619 13783 10625
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10625 14243 10659
rect 14185 10619 14243 10625
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 12529 10591 12587 10597
rect 12529 10557 12541 10591
rect 12575 10557 12587 10591
rect 12529 10551 12587 10557
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10588 12771 10591
rect 12802 10588 12808 10600
rect 12759 10560 12808 10588
rect 12759 10557 12771 10560
rect 12713 10551 12771 10557
rect 12544 10520 12572 10551
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 13740 10588 13768 10619
rect 15120 10588 15148 10619
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 15657 10659 15715 10665
rect 15657 10656 15669 10659
rect 15252 10628 15669 10656
rect 15252 10616 15258 10628
rect 15657 10625 15669 10628
rect 15703 10625 15715 10659
rect 15657 10619 15715 10625
rect 16945 10659 17003 10665
rect 16945 10625 16957 10659
rect 16991 10625 17003 10659
rect 18046 10656 18052 10668
rect 18007 10628 18052 10656
rect 16945 10619 17003 10625
rect 16960 10588 16988 10619
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 18524 10665 18552 10696
rect 18233 10659 18291 10665
rect 18233 10625 18245 10659
rect 18279 10656 18291 10659
rect 18509 10659 18567 10665
rect 18279 10628 18368 10656
rect 18279 10625 18291 10628
rect 18233 10619 18291 10625
rect 13740 10560 16988 10588
rect 13170 10520 13176 10532
rect 12544 10492 13176 10520
rect 13170 10480 13176 10492
rect 13228 10480 13234 10532
rect 13265 10523 13323 10529
rect 13265 10489 13277 10523
rect 13311 10520 13323 10523
rect 14366 10520 14372 10532
rect 13311 10492 14372 10520
rect 13311 10489 13323 10492
rect 13265 10483 13323 10489
rect 14366 10480 14372 10492
rect 14424 10480 14430 10532
rect 18340 10529 18368 10628
rect 18509 10625 18521 10659
rect 18555 10656 18567 10659
rect 18782 10656 18788 10668
rect 18555 10628 18788 10656
rect 18555 10625 18567 10628
rect 18509 10619 18567 10625
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 18325 10523 18383 10529
rect 18325 10489 18337 10523
rect 18371 10489 18383 10523
rect 18325 10483 18383 10489
rect 11609 10455 11667 10461
rect 11609 10452 11621 10455
rect 11572 10424 11621 10452
rect 11572 10412 11578 10424
rect 11609 10421 11621 10424
rect 11655 10421 11667 10455
rect 11609 10415 11667 10421
rect 13354 10412 13360 10464
rect 13412 10452 13418 10464
rect 13541 10455 13599 10461
rect 13541 10452 13553 10455
rect 13412 10424 13553 10452
rect 13412 10412 13418 10424
rect 13541 10421 13553 10424
rect 13587 10421 13599 10455
rect 14458 10452 14464 10464
rect 14419 10424 14464 10452
rect 13541 10415 13599 10421
rect 14458 10412 14464 10424
rect 14516 10412 14522 10464
rect 14826 10412 14832 10464
rect 14884 10452 14890 10464
rect 15013 10455 15071 10461
rect 15013 10452 15025 10455
rect 14884 10424 15025 10452
rect 14884 10412 14890 10424
rect 15013 10421 15025 10424
rect 15059 10421 15071 10455
rect 15013 10415 15071 10421
rect 15286 10412 15292 10464
rect 15344 10452 15350 10464
rect 16301 10455 16359 10461
rect 16301 10452 16313 10455
rect 15344 10424 16313 10452
rect 15344 10412 15350 10424
rect 16301 10421 16313 10424
rect 16347 10421 16359 10455
rect 16942 10452 16948 10464
rect 16903 10424 16948 10452
rect 16301 10415 16359 10421
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 0 10362 18860 10384
rect 0 10310 3110 10362
rect 3162 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 6210 10362
rect 6262 10310 6274 10362
rect 6326 10310 6338 10362
rect 6390 10310 6402 10362
rect 6454 10310 6466 10362
rect 6518 10310 9310 10362
rect 9362 10310 9374 10362
rect 9426 10310 9438 10362
rect 9490 10310 9502 10362
rect 9554 10310 9566 10362
rect 9618 10310 12410 10362
rect 12462 10310 12474 10362
rect 12526 10310 12538 10362
rect 12590 10310 12602 10362
rect 12654 10310 12666 10362
rect 12718 10310 15510 10362
rect 15562 10310 15574 10362
rect 15626 10310 15638 10362
rect 15690 10310 15702 10362
rect 15754 10310 15766 10362
rect 15818 10310 18860 10362
rect 0 10288 18860 10310
rect 3510 10248 3516 10260
rect 3471 10220 3516 10248
rect 3510 10208 3516 10220
rect 3568 10208 3574 10260
rect 7650 10208 7656 10260
rect 7708 10248 7714 10260
rect 7708 10220 10824 10248
rect 7708 10208 7714 10220
rect 4338 10180 4344 10192
rect 3712 10152 4344 10180
rect 1302 10112 1308 10124
rect 1263 10084 1308 10112
rect 1302 10072 1308 10084
rect 1360 10072 1366 10124
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 2590 10112 2596 10124
rect 1719 10084 2596 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 2590 10072 2596 10084
rect 2648 10072 2654 10124
rect 3712 10112 3740 10152
rect 4338 10140 4344 10152
rect 4396 10180 4402 10192
rect 4890 10180 4896 10192
rect 4396 10152 4896 10180
rect 4396 10140 4402 10152
rect 4890 10140 4896 10152
rect 4948 10140 4954 10192
rect 8754 10180 8760 10192
rect 8715 10152 8760 10180
rect 8754 10140 8760 10152
rect 8812 10140 8818 10192
rect 10686 10180 10692 10192
rect 10647 10152 10692 10180
rect 10686 10140 10692 10152
rect 10744 10140 10750 10192
rect 10796 10180 10824 10220
rect 11238 10208 11244 10260
rect 11296 10248 11302 10260
rect 12805 10251 12863 10257
rect 12805 10248 12817 10251
rect 11296 10220 12817 10248
rect 11296 10208 11302 10220
rect 12805 10217 12817 10220
rect 12851 10217 12863 10251
rect 12805 10211 12863 10217
rect 13170 10208 13176 10260
rect 13228 10248 13234 10260
rect 14918 10248 14924 10260
rect 13228 10220 14924 10248
rect 13228 10208 13234 10220
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 15194 10257 15200 10260
rect 15151 10251 15200 10257
rect 15151 10217 15163 10251
rect 15197 10217 15200 10251
rect 15151 10211 15200 10217
rect 15194 10208 15200 10211
rect 15252 10208 15258 10260
rect 17819 10251 17877 10257
rect 17819 10217 17831 10251
rect 17865 10248 17877 10251
rect 18046 10248 18052 10260
rect 17865 10220 18052 10248
rect 17865 10217 17877 10220
rect 17819 10211 17877 10217
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 12161 10183 12219 10189
rect 12161 10180 12173 10183
rect 10796 10152 12173 10180
rect 12161 10149 12173 10152
rect 12207 10180 12219 10183
rect 12207 10152 12434 10180
rect 12207 10149 12219 10152
rect 12161 10143 12219 10149
rect 2976 10084 3740 10112
rect 2682 9936 2688 9988
rect 2740 9936 2746 9988
rect 2222 9868 2228 9920
rect 2280 9908 2286 9920
rect 2976 9908 3004 10084
rect 3712 10053 3740 10084
rect 4154 10072 4160 10124
rect 4212 10112 4218 10124
rect 4709 10115 4767 10121
rect 4212 10084 4476 10112
rect 4212 10072 4218 10084
rect 4448 10053 4476 10084
rect 4709 10081 4721 10115
rect 4755 10112 4767 10115
rect 4755 10084 5120 10112
rect 4755 10081 4767 10084
rect 4709 10075 4767 10081
rect 3329 10047 3387 10053
rect 3329 10013 3341 10047
rect 3375 10013 3387 10047
rect 3329 10007 3387 10013
rect 3513 10047 3571 10053
rect 3513 10013 3525 10047
rect 3559 10044 3571 10047
rect 3697 10047 3755 10053
rect 3697 10044 3709 10047
rect 3559 10016 3709 10044
rect 3559 10013 3571 10016
rect 3513 10007 3571 10013
rect 3697 10013 3709 10016
rect 3743 10013 3755 10047
rect 3697 10007 3755 10013
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10044 4491 10047
rect 4617 10047 4675 10053
rect 4617 10044 4629 10047
rect 4479 10016 4629 10044
rect 4479 10013 4491 10016
rect 4433 10007 4491 10013
rect 4617 10013 4629 10016
rect 4663 10013 4675 10047
rect 4617 10007 4675 10013
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 3099 9979 3157 9985
rect 3099 9945 3111 9979
rect 3145 9976 3157 9979
rect 3344 9976 3372 10007
rect 4062 9976 4068 9988
rect 3145 9948 4068 9976
rect 3145 9945 3157 9948
rect 3099 9939 3157 9945
rect 4062 9936 4068 9948
rect 4120 9976 4126 9988
rect 4264 9976 4292 10007
rect 4816 9976 4844 10007
rect 4890 10004 4896 10056
rect 4948 10044 4954 10056
rect 5092 10053 5120 10084
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 5813 10115 5871 10121
rect 5813 10112 5825 10115
rect 5500 10084 5825 10112
rect 5500 10072 5506 10084
rect 5813 10081 5825 10084
rect 5859 10112 5871 10115
rect 6362 10112 6368 10124
rect 5859 10084 6368 10112
rect 5859 10081 5871 10084
rect 5813 10075 5871 10081
rect 6362 10072 6368 10084
rect 6420 10072 6426 10124
rect 5077 10047 5135 10053
rect 4948 10016 4993 10044
rect 4948 10004 4954 10016
rect 5077 10013 5089 10047
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 5353 10047 5411 10053
rect 5353 10013 5365 10047
rect 5399 10013 5411 10047
rect 5534 10044 5540 10056
rect 5495 10016 5540 10044
rect 5353 10007 5411 10013
rect 4120 9948 4844 9976
rect 4985 9979 5043 9985
rect 4120 9936 4126 9948
rect 4985 9945 4997 9979
rect 5031 9976 5043 9979
rect 5368 9976 5396 10007
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 6089 10047 6147 10053
rect 6089 10013 6101 10047
rect 6135 10044 6147 10047
rect 6178 10044 6184 10056
rect 6135 10016 6184 10044
rect 6135 10013 6147 10016
rect 6089 10007 6147 10013
rect 6178 10004 6184 10016
rect 6236 10004 6242 10056
rect 6454 10044 6460 10056
rect 6415 10016 6460 10044
rect 6454 10004 6460 10016
rect 6512 10004 6518 10056
rect 8662 10044 8668 10056
rect 8623 10016 8668 10044
rect 8662 10004 8668 10016
rect 8720 10004 8726 10056
rect 5031 9948 5396 9976
rect 5031 9945 5043 9948
rect 4985 9939 5043 9945
rect 7006 9936 7012 9988
rect 7064 9936 7070 9988
rect 2280 9880 3004 9908
rect 4433 9911 4491 9917
rect 2280 9868 2286 9880
rect 4433 9877 4445 9911
rect 4479 9908 4491 9911
rect 4522 9908 4528 9920
rect 4479 9880 4528 9908
rect 4479 9877 4491 9880
rect 4433 9871 4491 9877
rect 4522 9868 4528 9880
rect 4580 9868 4586 9920
rect 5629 9911 5687 9917
rect 5629 9877 5641 9911
rect 5675 9908 5687 9911
rect 5718 9908 5724 9920
rect 5675 9880 5724 9908
rect 5675 9877 5687 9880
rect 5629 9871 5687 9877
rect 5718 9868 5724 9880
rect 5776 9868 5782 9920
rect 7650 9868 7656 9920
rect 7708 9908 7714 9920
rect 7883 9911 7941 9917
rect 7883 9908 7895 9911
rect 7708 9880 7895 9908
rect 7708 9868 7714 9880
rect 7883 9877 7895 9880
rect 7929 9877 7941 9911
rect 8478 9908 8484 9920
rect 8439 9880 8484 9908
rect 7883 9871 7941 9877
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 8772 9908 8800 10140
rect 8941 10115 8999 10121
rect 8941 10081 8953 10115
rect 8987 10112 8999 10115
rect 9950 10112 9956 10124
rect 8987 10084 9956 10112
rect 8987 10081 8999 10084
rect 8941 10075 8999 10081
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 12406 10044 12434 10152
rect 13354 10112 13360 10124
rect 13315 10084 13360 10112
rect 13354 10072 13360 10084
rect 13412 10072 13418 10124
rect 13725 10115 13783 10121
rect 13725 10081 13737 10115
rect 13771 10112 13783 10115
rect 14458 10112 14464 10124
rect 13771 10084 14464 10112
rect 13771 10081 13783 10084
rect 13725 10075 13783 10081
rect 14458 10072 14464 10084
rect 14516 10072 14522 10124
rect 16025 10115 16083 10121
rect 16025 10081 16037 10115
rect 16071 10112 16083 10115
rect 16942 10112 16948 10124
rect 16071 10084 16948 10112
rect 16071 10081 16083 10084
rect 16025 10075 16083 10081
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 12897 10047 12955 10053
rect 12897 10044 12909 10047
rect 12406 10016 12909 10044
rect 12897 10013 12909 10016
rect 12943 10013 12955 10047
rect 12897 10007 12955 10013
rect 16393 10047 16451 10053
rect 16393 10013 16405 10047
rect 16439 10044 16451 10047
rect 16482 10044 16488 10056
rect 16439 10016 16488 10044
rect 16439 10013 16451 10016
rect 16393 10007 16451 10013
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 18233 10047 18291 10053
rect 18233 10013 18245 10047
rect 18279 10044 18291 10047
rect 18509 10047 18567 10053
rect 18509 10044 18521 10047
rect 18279 10016 18521 10044
rect 18279 10013 18291 10016
rect 18233 10007 18291 10013
rect 18509 10013 18521 10016
rect 18555 10044 18567 10047
rect 18598 10044 18604 10056
rect 18555 10016 18604 10044
rect 18555 10013 18567 10016
rect 18509 10007 18567 10013
rect 18598 10004 18604 10016
rect 18656 10004 18662 10056
rect 9214 9976 9220 9988
rect 9175 9948 9220 9976
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 9674 9936 9680 9988
rect 9732 9936 9738 9988
rect 10873 9979 10931 9985
rect 10873 9976 10885 9979
rect 10520 9948 10885 9976
rect 9692 9908 9720 9936
rect 8772 9880 9720 9908
rect 9858 9868 9864 9920
rect 9916 9908 9922 9920
rect 10520 9908 10548 9948
rect 10873 9945 10885 9948
rect 10919 9945 10931 9979
rect 10873 9939 10931 9945
rect 9916 9880 10548 9908
rect 9916 9868 9922 9880
rect 14366 9868 14372 9920
rect 14424 9908 14430 9920
rect 14752 9908 14780 9962
rect 15749 9911 15807 9917
rect 15749 9908 15761 9911
rect 14424 9880 15761 9908
rect 14424 9868 14430 9880
rect 15749 9877 15761 9880
rect 15795 9908 15807 9911
rect 15933 9911 15991 9917
rect 15933 9908 15945 9911
rect 15795 9880 15945 9908
rect 15795 9877 15807 9880
rect 15749 9871 15807 9877
rect 15933 9877 15945 9880
rect 15979 9908 15991 9911
rect 16776 9908 16804 9962
rect 18322 9908 18328 9920
rect 15979 9880 16804 9908
rect 18283 9880 18328 9908
rect 15979 9877 15991 9880
rect 15933 9871 15991 9877
rect 18322 9868 18328 9880
rect 18380 9868 18386 9920
rect 0 9818 18860 9840
rect 0 9766 4660 9818
rect 4712 9766 4724 9818
rect 4776 9766 4788 9818
rect 4840 9766 4852 9818
rect 4904 9766 4916 9818
rect 4968 9766 7760 9818
rect 7812 9766 7824 9818
rect 7876 9766 7888 9818
rect 7940 9766 7952 9818
rect 8004 9766 8016 9818
rect 8068 9766 10860 9818
rect 10912 9766 10924 9818
rect 10976 9766 10988 9818
rect 11040 9766 11052 9818
rect 11104 9766 11116 9818
rect 11168 9766 13960 9818
rect 14012 9766 14024 9818
rect 14076 9766 14088 9818
rect 14140 9766 14152 9818
rect 14204 9766 14216 9818
rect 14268 9766 17060 9818
rect 17112 9766 17124 9818
rect 17176 9766 17188 9818
rect 17240 9766 17252 9818
rect 17304 9766 17316 9818
rect 17368 9766 18860 9818
rect 0 9744 18860 9766
rect 2041 9707 2099 9713
rect 2041 9673 2053 9707
rect 2087 9704 2099 9707
rect 4154 9704 4160 9716
rect 2087 9676 4160 9704
rect 2087 9673 2099 9676
rect 2041 9667 2099 9673
rect 1946 9636 1952 9648
rect 1794 9608 1952 9636
rect 1946 9596 1952 9608
rect 2004 9596 2010 9648
rect 2593 9639 2651 9645
rect 2593 9605 2605 9639
rect 2639 9636 2651 9639
rect 2682 9636 2688 9648
rect 2639 9608 2688 9636
rect 2639 9605 2651 9608
rect 2593 9599 2651 9605
rect 2682 9596 2688 9608
rect 2740 9596 2746 9648
rect 2792 9645 2820 9676
rect 4154 9664 4160 9676
rect 4212 9664 4218 9716
rect 5445 9707 5503 9713
rect 5445 9673 5457 9707
rect 5491 9704 5503 9707
rect 5813 9707 5871 9713
rect 5491 9676 5580 9704
rect 5491 9673 5503 9676
rect 5445 9667 5503 9673
rect 2777 9639 2835 9645
rect 2777 9605 2789 9639
rect 2823 9605 2835 9639
rect 2777 9599 2835 9605
rect 2961 9639 3019 9645
rect 2961 9605 2973 9639
rect 3007 9636 3019 9639
rect 3050 9636 3056 9648
rect 3007 9608 3056 9636
rect 3007 9605 3019 9608
rect 2961 9599 3019 9605
rect 3050 9596 3056 9608
rect 3108 9596 3114 9648
rect 3145 9639 3203 9645
rect 3145 9605 3157 9639
rect 3191 9636 3203 9639
rect 4062 9636 4068 9648
rect 3191 9608 4068 9636
rect 3191 9605 3203 9608
rect 3145 9599 3203 9605
rect 4062 9596 4068 9608
rect 4120 9636 4126 9648
rect 5350 9636 5356 9648
rect 4120 9608 4200 9636
rect 5311 9608 5356 9636
rect 4120 9596 4126 9608
rect 2130 9568 2136 9580
rect 2091 9540 2136 9568
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9537 2375 9571
rect 2498 9568 2504 9580
rect 2459 9540 2504 9568
rect 2317 9531 2375 9537
rect 290 9500 296 9512
rect 251 9472 296 9500
rect 290 9460 296 9472
rect 348 9460 354 9512
rect 569 9503 627 9509
rect 569 9469 581 9503
rect 615 9500 627 9503
rect 2225 9503 2283 9509
rect 2225 9500 2237 9503
rect 615 9472 2237 9500
rect 615 9469 627 9472
rect 569 9463 627 9469
rect 2225 9469 2237 9472
rect 2271 9469 2283 9503
rect 2332 9500 2360 9531
rect 2498 9528 2504 9540
rect 2556 9568 2562 9580
rect 4172 9577 4200 9608
rect 5350 9596 5356 9608
rect 5408 9596 5414 9648
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 2556 9540 2881 9568
rect 2556 9528 2562 9540
rect 2869 9537 2881 9540
rect 2915 9537 2927 9571
rect 2869 9531 2927 9537
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9537 3295 9571
rect 3237 9531 3295 9537
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9537 4215 9571
rect 4157 9531 4215 9537
rect 2332 9472 2544 9500
rect 2225 9463 2283 9469
rect 2516 9441 2544 9472
rect 3050 9460 3056 9512
rect 3108 9500 3114 9512
rect 3252 9500 3280 9531
rect 3108 9472 3280 9500
rect 3108 9460 3114 9472
rect 2501 9435 2559 9441
rect 2501 9401 2513 9435
rect 2547 9401 2559 9435
rect 3329 9435 3387 9441
rect 3329 9432 3341 9435
rect 2501 9395 2559 9401
rect 2976 9404 3341 9432
rect 2682 9324 2688 9376
rect 2740 9364 2746 9376
rect 2976 9364 3004 9404
rect 3329 9401 3341 9404
rect 3375 9401 3387 9435
rect 3329 9395 3387 9401
rect 2740 9336 3004 9364
rect 3053 9367 3111 9373
rect 2740 9324 2746 9336
rect 3053 9333 3065 9367
rect 3099 9364 3111 9367
rect 3436 9364 3464 9531
rect 4522 9528 4528 9580
rect 4580 9568 4586 9580
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 4580 9540 5181 9568
rect 4580 9528 4586 9540
rect 5169 9537 5181 9540
rect 5215 9537 5227 9571
rect 5442 9568 5448 9580
rect 5403 9540 5448 9568
rect 5169 9531 5227 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 5552 9568 5580 9676
rect 5813 9673 5825 9707
rect 5859 9704 5871 9707
rect 6454 9704 6460 9716
rect 5859 9676 6460 9704
rect 5859 9673 5871 9676
rect 5813 9667 5871 9673
rect 6454 9664 6460 9676
rect 6512 9664 6518 9716
rect 8938 9664 8944 9716
rect 8996 9704 9002 9716
rect 9309 9707 9367 9713
rect 9309 9704 9321 9707
rect 8996 9676 9321 9704
rect 8996 9664 9002 9676
rect 9309 9673 9321 9676
rect 9355 9673 9367 9707
rect 9309 9667 9367 9673
rect 12437 9707 12495 9713
rect 12437 9673 12449 9707
rect 12483 9704 12495 9707
rect 14366 9704 14372 9716
rect 12483 9676 14372 9704
rect 12483 9673 12495 9676
rect 12437 9667 12495 9673
rect 5718 9636 5724 9648
rect 5679 9608 5724 9636
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 5905 9639 5963 9645
rect 5905 9605 5917 9639
rect 5951 9636 5963 9639
rect 6178 9636 6184 9648
rect 5951 9608 6031 9636
rect 6139 9608 6184 9636
rect 5951 9605 5963 9608
rect 5905 9599 5963 9605
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5552 9540 5641 9568
rect 5629 9537 5641 9540
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 6003 9512 6031 9608
rect 6178 9596 6184 9608
rect 6236 9596 6242 9648
rect 6362 9596 6368 9648
rect 6420 9636 6426 9648
rect 7285 9639 7343 9645
rect 7285 9636 7297 9639
rect 6420 9608 7297 9636
rect 6420 9596 6426 9608
rect 7285 9605 7297 9608
rect 7331 9605 7343 9639
rect 7285 9599 7343 9605
rect 8196 9639 8254 9645
rect 8196 9605 8208 9639
rect 8242 9636 8254 9639
rect 8478 9636 8484 9648
rect 8242 9608 8484 9636
rect 8242 9605 8254 9608
rect 8196 9599 8254 9605
rect 8478 9596 8484 9608
rect 8536 9596 8542 9648
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 10042 9636 10048 9648
rect 9732 9608 10048 9636
rect 9732 9596 9738 9608
rect 10042 9596 10048 9608
rect 10100 9636 10106 9648
rect 10686 9636 10692 9648
rect 10100 9608 10692 9636
rect 10100 9596 10106 9608
rect 10686 9596 10692 9608
rect 10744 9636 10750 9648
rect 10744 9608 10902 9636
rect 10744 9596 10750 9608
rect 6086 9528 6092 9580
rect 6144 9568 6150 9580
rect 6273 9571 6331 9577
rect 6273 9568 6285 9571
rect 6144 9540 6285 9568
rect 6144 9528 6150 9540
rect 6273 9537 6285 9540
rect 6319 9537 6331 9571
rect 6273 9531 6331 9537
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 7745 9571 7803 9577
rect 7745 9568 7757 9571
rect 7708 9540 7757 9568
rect 7708 9528 7714 9540
rect 7745 9537 7757 9540
rect 7791 9568 7803 9571
rect 7791 9540 8984 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9500 4307 9503
rect 4338 9500 4344 9512
rect 4295 9472 4344 9500
rect 4295 9469 4307 9472
rect 4249 9463 4307 9469
rect 4338 9460 4344 9472
rect 4396 9460 4402 9512
rect 5994 9460 6000 9512
rect 6052 9500 6058 9512
rect 6052 9472 6145 9500
rect 6052 9460 6058 9472
rect 3602 9392 3608 9444
rect 3660 9432 3666 9444
rect 3660 9404 5396 9432
rect 3660 9392 3666 9404
rect 3099 9336 3464 9364
rect 4433 9367 4491 9373
rect 3099 9333 3111 9336
rect 3053 9327 3111 9333
rect 4433 9333 4445 9367
rect 4479 9364 4491 9367
rect 5258 9364 5264 9376
rect 4479 9336 5264 9364
rect 4479 9333 4491 9336
rect 4433 9327 4491 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5368 9364 5396 9404
rect 5997 9367 6055 9373
rect 5997 9364 6009 9367
rect 5368 9336 6009 9364
rect 5997 9333 6009 9336
rect 6043 9333 6055 9367
rect 6104 9364 6132 9472
rect 7558 9460 7564 9512
rect 7616 9500 7622 9512
rect 7929 9503 7987 9509
rect 7929 9500 7941 9503
rect 7616 9472 7941 9500
rect 7616 9460 7622 9472
rect 7929 9469 7941 9472
rect 7975 9469 7987 9503
rect 8956 9500 8984 9540
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10137 9571 10195 9577
rect 10137 9568 10149 9571
rect 10008 9540 10149 9568
rect 10008 9528 10014 9540
rect 10137 9537 10149 9540
rect 10183 9537 10195 9571
rect 10137 9531 10195 9537
rect 11790 9528 11796 9580
rect 11848 9568 11854 9580
rect 12452 9568 12480 9667
rect 13556 9622 13584 9676
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 14458 9664 14464 9716
rect 14516 9704 14522 9716
rect 14516 9676 15608 9704
rect 14516 9664 14522 9676
rect 14001 9639 14059 9645
rect 14001 9605 14013 9639
rect 14047 9636 14059 9639
rect 14047 9608 14688 9636
rect 15580 9622 15608 9676
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 16632 9676 17540 9704
rect 16632 9664 16638 9676
rect 17512 9645 17540 9676
rect 17497 9639 17555 9645
rect 14047 9605 14059 9608
rect 14001 9599 14059 9605
rect 11848 9540 12480 9568
rect 11848 9528 11854 9540
rect 10413 9503 10471 9509
rect 8956 9472 10088 9500
rect 7929 9463 7987 9469
rect 9674 9432 9680 9444
rect 8864 9404 9680 9432
rect 8864 9364 8892 9404
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 9766 9364 9772 9376
rect 6104 9336 8892 9364
rect 9727 9336 9772 9364
rect 5997 9327 6055 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 10060 9364 10088 9472
rect 10413 9469 10425 9503
rect 10459 9500 10471 9503
rect 11146 9500 11152 9512
rect 10459 9472 11152 9500
rect 10459 9469 10471 9472
rect 10413 9463 10471 9469
rect 11146 9460 11152 9472
rect 11204 9500 11210 9512
rect 11606 9500 11612 9512
rect 11204 9472 11612 9500
rect 11204 9460 11210 9472
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9500 11943 9503
rect 12802 9500 12808 9512
rect 11931 9472 12808 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 14277 9503 14335 9509
rect 14277 9469 14289 9503
rect 14323 9469 14335 9503
rect 14660 9500 14688 9608
rect 17497 9605 17509 9639
rect 17543 9605 17555 9639
rect 17497 9599 17555 9605
rect 14826 9568 14832 9580
rect 14787 9540 14832 9568
rect 14826 9528 14832 9540
rect 14884 9528 14890 9580
rect 15197 9571 15255 9577
rect 15197 9537 15209 9571
rect 15243 9568 15255 9571
rect 15286 9568 15292 9580
rect 15243 9540 15292 9568
rect 15243 9537 15255 9540
rect 15197 9531 15255 9537
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 16623 9571 16681 9577
rect 16623 9537 16635 9571
rect 16669 9568 16681 9571
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16669 9540 16865 9568
rect 16669 9537 16681 9540
rect 16623 9531 16681 9537
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 18322 9500 18328 9512
rect 14660 9472 18328 9500
rect 14277 9463 14335 9469
rect 14292 9432 14320 9463
rect 18322 9460 18328 9472
rect 18380 9460 18386 9512
rect 14292 9404 14780 9432
rect 11422 9364 11428 9376
rect 10060 9336 11428 9364
rect 11422 9324 11428 9336
rect 11480 9324 11486 9376
rect 12529 9367 12587 9373
rect 12529 9333 12541 9367
rect 12575 9364 12587 9367
rect 13354 9364 13360 9376
rect 12575 9336 13360 9364
rect 12575 9333 12587 9336
rect 12529 9327 12587 9333
rect 13354 9324 13360 9336
rect 13412 9324 13418 9376
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 14292 9364 14320 9404
rect 13504 9336 14320 9364
rect 13504 9324 13510 9336
rect 14458 9324 14464 9376
rect 14516 9364 14522 9376
rect 14645 9367 14703 9373
rect 14645 9364 14657 9367
rect 14516 9336 14657 9364
rect 14516 9324 14522 9336
rect 14645 9333 14657 9336
rect 14691 9333 14703 9367
rect 14752 9364 14780 9404
rect 16666 9364 16672 9376
rect 14752 9336 16672 9364
rect 14645 9327 14703 9333
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 0 9274 18860 9296
rect 0 9222 3110 9274
rect 3162 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 6210 9274
rect 6262 9222 6274 9274
rect 6326 9222 6338 9274
rect 6390 9222 6402 9274
rect 6454 9222 6466 9274
rect 6518 9222 9310 9274
rect 9362 9222 9374 9274
rect 9426 9222 9438 9274
rect 9490 9222 9502 9274
rect 9554 9222 9566 9274
rect 9618 9222 12410 9274
rect 12462 9222 12474 9274
rect 12526 9222 12538 9274
rect 12590 9222 12602 9274
rect 12654 9222 12666 9274
rect 12718 9222 15510 9274
rect 15562 9222 15574 9274
rect 15626 9222 15638 9274
rect 15690 9222 15702 9274
rect 15754 9222 15766 9274
rect 15818 9222 18860 9274
rect 0 9200 18860 9222
rect 1394 9160 1400 9172
rect 1355 9132 1400 9160
rect 1394 9120 1400 9132
rect 1452 9120 1458 9172
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 3053 9163 3111 9169
rect 3053 9160 3065 9163
rect 3016 9132 3065 9160
rect 3016 9120 3022 9132
rect 3053 9129 3065 9132
rect 3099 9129 3111 9163
rect 10686 9160 10692 9172
rect 10647 9132 10692 9160
rect 3053 9123 3111 9129
rect 10686 9120 10692 9132
rect 10744 9160 10750 9172
rect 11790 9160 11796 9172
rect 10744 9132 11796 9160
rect 10744 9120 10750 9132
rect 11790 9120 11796 9132
rect 11848 9160 11854 9172
rect 13265 9163 13323 9169
rect 13265 9160 13277 9163
rect 11848 9132 13277 9160
rect 11848 9120 11854 9132
rect 13265 9129 13277 9132
rect 13311 9160 13323 9163
rect 14182 9160 14188 9172
rect 13311 9132 14188 9160
rect 13311 9129 13323 9132
rect 13265 9123 13323 9129
rect 14182 9120 14188 9132
rect 14240 9160 14246 9172
rect 14458 9160 14464 9172
rect 14240 9132 14464 9160
rect 14240 9120 14246 9132
rect 14458 9120 14464 9132
rect 14516 9120 14522 9172
rect 10045 9095 10103 9101
rect 10045 9061 10057 9095
rect 10091 9092 10103 9095
rect 10505 9095 10563 9101
rect 10505 9092 10517 9095
rect 10091 9064 10517 9092
rect 10091 9061 10103 9064
rect 10045 9055 10103 9061
rect 10505 9061 10517 9064
rect 10551 9061 10563 9095
rect 10505 9055 10563 9061
rect 1946 9024 1952 9036
rect 1907 8996 1952 9024
rect 1946 8984 1952 8996
rect 2004 8984 2010 9036
rect 4522 8984 4528 9036
rect 4580 9024 4586 9036
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 4580 8996 4629 9024
rect 4580 8984 4586 8996
rect 4617 8993 4629 8996
rect 4663 9024 4675 9027
rect 5537 9027 5595 9033
rect 5537 9024 5549 9027
rect 4663 8996 5549 9024
rect 4663 8993 4675 8996
rect 4617 8987 4675 8993
rect 5537 8993 5549 8996
rect 5583 8993 5595 9027
rect 10686 9024 10692 9036
rect 5537 8987 5595 8993
rect 10060 8996 10692 9024
rect 1394 8916 1400 8968
rect 1452 8956 1458 8968
rect 1489 8959 1547 8965
rect 1489 8956 1501 8959
rect 1452 8928 1501 8956
rect 1452 8916 1458 8928
rect 1489 8925 1501 8928
rect 1535 8925 1547 8959
rect 1489 8919 1547 8925
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 2961 8959 3019 8965
rect 2961 8956 2973 8959
rect 2740 8928 2973 8956
rect 2740 8916 2746 8928
rect 2961 8925 2973 8928
rect 3007 8925 3019 8959
rect 2961 8919 3019 8925
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 4430 8956 4436 8968
rect 4391 8928 4436 8956
rect 3145 8919 3203 8925
rect 3160 8888 3188 8919
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 4982 8916 4988 8968
rect 5040 8916 5046 8968
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 5316 8928 5365 8956
rect 5316 8916 5322 8928
rect 5353 8925 5365 8928
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 6086 8916 6092 8968
rect 6144 8956 6150 8968
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 6144 8928 6837 8956
rect 6144 8916 6150 8928
rect 6825 8925 6837 8928
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 7092 8959 7150 8965
rect 7092 8925 7104 8959
rect 7138 8956 7150 8959
rect 8386 8956 8392 8968
rect 7138 8928 8392 8956
rect 7138 8925 7150 8928
rect 7092 8919 7150 8925
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 8665 8959 8723 8965
rect 8665 8956 8677 8959
rect 8536 8928 8677 8956
rect 8536 8916 8542 8928
rect 8665 8925 8677 8928
rect 8711 8956 8723 8959
rect 10060 8956 10088 8996
rect 10686 8984 10692 8996
rect 10744 9024 10750 9036
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 10744 8996 10885 9024
rect 10744 8984 10750 8996
rect 10873 8993 10885 8996
rect 10919 8993 10931 9027
rect 10873 8987 10931 8993
rect 10980 8996 12020 9024
rect 8711 8928 10088 8956
rect 8711 8925 8723 8928
rect 8665 8919 8723 8925
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 10413 8959 10471 8965
rect 10192 8928 10237 8956
rect 10192 8916 10198 8928
rect 10413 8925 10425 8959
rect 10459 8956 10471 8959
rect 10505 8959 10563 8965
rect 10505 8956 10517 8959
rect 10459 8928 10517 8956
rect 10459 8925 10471 8928
rect 10413 8919 10471 8925
rect 10505 8925 10517 8928
rect 10551 8925 10563 8959
rect 10505 8919 10563 8925
rect 10778 8916 10784 8968
rect 10836 8956 10842 8968
rect 10980 8956 11008 8996
rect 11238 8956 11244 8968
rect 10836 8928 11008 8956
rect 11199 8928 11244 8956
rect 10836 8916 10842 8928
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 11992 8956 12020 8996
rect 13354 8984 13360 9036
rect 13412 9024 13418 9036
rect 13725 9027 13783 9033
rect 13725 9024 13737 9027
rect 13412 8996 13737 9024
rect 13412 8984 13418 8996
rect 13725 8993 13737 8996
rect 13771 8993 13783 9027
rect 13725 8987 13783 8993
rect 14458 8984 14464 9036
rect 14516 9024 14522 9036
rect 15473 9027 15531 9033
rect 15473 9024 15485 9027
rect 14516 8996 15485 9024
rect 14516 8984 14522 8996
rect 15473 8993 15485 8996
rect 15519 8993 15531 9027
rect 15473 8987 15531 8993
rect 15749 9027 15807 9033
rect 15749 8993 15761 9027
rect 15795 9024 15807 9027
rect 16666 9024 16672 9036
rect 15795 8996 16672 9024
rect 15795 8993 15807 8996
rect 15749 8987 15807 8993
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 13446 8956 13452 8968
rect 11992 8928 12434 8956
rect 13407 8928 13452 8956
rect 4338 8888 4344 8900
rect 3160 8860 4344 8888
rect 4338 8848 4344 8860
rect 4396 8848 4402 8900
rect 5000 8888 5028 8916
rect 5445 8891 5503 8897
rect 5445 8888 5457 8891
rect 5000 8860 5457 8888
rect 5445 8857 5457 8860
rect 5491 8857 5503 8891
rect 5445 8851 5503 8857
rect 8294 8848 8300 8900
rect 8352 8888 8358 8900
rect 8932 8891 8990 8897
rect 8352 8860 8708 8888
rect 8352 8848 8358 8860
rect 1946 8780 1952 8832
rect 2004 8820 2010 8832
rect 2498 8820 2504 8832
rect 2004 8792 2504 8820
rect 2004 8780 2010 8792
rect 2498 8780 2504 8792
rect 2556 8820 2562 8832
rect 3602 8820 3608 8832
rect 2556 8792 3608 8820
rect 2556 8780 2562 8792
rect 3602 8780 3608 8792
rect 3660 8780 3666 8832
rect 4065 8823 4123 8829
rect 4065 8789 4077 8823
rect 4111 8820 4123 8823
rect 4154 8820 4160 8832
rect 4111 8792 4160 8820
rect 4111 8789 4123 8792
rect 4065 8783 4123 8789
rect 4154 8780 4160 8792
rect 4212 8780 4218 8832
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4488 8792 4537 8820
rect 4488 8780 4494 8792
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 4525 8783 4583 8789
rect 4985 8823 5043 8829
rect 4985 8789 4997 8823
rect 5031 8820 5043 8823
rect 5258 8820 5264 8832
rect 5031 8792 5264 8820
rect 5031 8789 5043 8792
rect 4985 8783 5043 8789
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 8205 8823 8263 8829
rect 8205 8789 8217 8823
rect 8251 8820 8263 8823
rect 8570 8820 8576 8832
rect 8251 8792 8576 8820
rect 8251 8789 8263 8792
rect 8205 8783 8263 8789
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 8680 8820 8708 8860
rect 8932 8857 8944 8891
rect 8978 8888 8990 8891
rect 9122 8888 9128 8900
rect 8978 8860 9128 8888
rect 8978 8857 8990 8860
rect 8932 8851 8990 8857
rect 9122 8848 9128 8860
rect 9180 8848 9186 8900
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 10229 8891 10287 8897
rect 10229 8888 10241 8891
rect 9548 8860 10241 8888
rect 9548 8848 9554 8860
rect 10229 8857 10241 8860
rect 10275 8857 10287 8891
rect 10229 8851 10287 8857
rect 11790 8848 11796 8900
rect 11848 8848 11854 8900
rect 12406 8888 12434 8928
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 16117 8959 16175 8965
rect 16117 8956 16129 8959
rect 15896 8928 16129 8956
rect 15896 8916 15902 8928
rect 16117 8925 16129 8928
rect 16163 8925 16175 8959
rect 16117 8919 16175 8925
rect 12406 8860 14136 8888
rect 10137 8823 10195 8829
rect 10137 8820 10149 8823
rect 8680 8792 10149 8820
rect 10137 8789 10149 8792
rect 10183 8789 10195 8823
rect 10137 8783 10195 8789
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 12667 8823 12725 8829
rect 12667 8820 12679 8823
rect 12032 8792 12679 8820
rect 12032 8780 12038 8792
rect 12667 8789 12679 8792
rect 12713 8789 12725 8823
rect 14108 8820 14136 8860
rect 14182 8848 14188 8900
rect 14240 8848 14246 8900
rect 16482 8848 16488 8900
rect 16540 8848 16546 8900
rect 14366 8820 14372 8832
rect 14108 8792 14372 8820
rect 12667 8783 12725 8789
rect 14366 8780 14372 8792
rect 14424 8820 14430 8832
rect 17865 8823 17923 8829
rect 17865 8820 17877 8823
rect 14424 8792 17877 8820
rect 14424 8780 14430 8792
rect 17865 8789 17877 8792
rect 17911 8820 17923 8823
rect 18046 8820 18052 8832
rect 17911 8792 18052 8820
rect 17911 8789 17923 8792
rect 17865 8783 17923 8789
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 0 8730 18860 8752
rect 0 8678 4660 8730
rect 4712 8678 4724 8730
rect 4776 8678 4788 8730
rect 4840 8678 4852 8730
rect 4904 8678 4916 8730
rect 4968 8678 7760 8730
rect 7812 8678 7824 8730
rect 7876 8678 7888 8730
rect 7940 8678 7952 8730
rect 8004 8678 8016 8730
rect 8068 8678 10860 8730
rect 10912 8678 10924 8730
rect 10976 8678 10988 8730
rect 11040 8678 11052 8730
rect 11104 8678 11116 8730
rect 11168 8678 13960 8730
rect 14012 8678 14024 8730
rect 14076 8678 14088 8730
rect 14140 8678 14152 8730
rect 14204 8678 14216 8730
rect 14268 8678 17060 8730
rect 17112 8678 17124 8730
rect 17176 8678 17188 8730
rect 17240 8678 17252 8730
rect 17304 8678 17316 8730
rect 17368 8678 18860 8730
rect 0 8656 18860 8678
rect 2130 8616 2136 8628
rect 2091 8588 2136 8616
rect 2130 8576 2136 8588
rect 2188 8576 2194 8628
rect 4154 8616 4160 8628
rect 4115 8588 4160 8616
rect 4154 8576 4160 8588
rect 4212 8576 4218 8628
rect 4338 8576 4344 8628
rect 4396 8616 4402 8628
rect 4893 8619 4951 8625
rect 4893 8616 4905 8619
rect 4396 8588 4905 8616
rect 4396 8576 4402 8588
rect 4893 8585 4905 8588
rect 4939 8585 4951 8619
rect 5258 8616 5264 8628
rect 5219 8588 5264 8616
rect 4893 8579 4951 8585
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 8941 8619 8999 8625
rect 8941 8585 8953 8619
rect 8987 8585 8999 8619
rect 9490 8616 9496 8628
rect 9451 8588 9496 8616
rect 8941 8579 8999 8585
rect 1946 8548 1952 8560
rect 1794 8520 1952 8548
rect 1946 8508 1952 8520
rect 2004 8508 2010 8560
rect 2501 8551 2559 8557
rect 2501 8548 2513 8551
rect 2240 8520 2513 8548
rect 2130 8480 2136 8492
rect 2091 8452 2136 8480
rect 2130 8440 2136 8452
rect 2188 8440 2194 8492
rect 290 8412 296 8424
rect 251 8384 296 8412
rect 290 8372 296 8384
rect 348 8372 354 8424
rect 569 8415 627 8421
rect 569 8381 581 8415
rect 615 8412 627 8415
rect 2240 8412 2268 8520
rect 2501 8517 2513 8520
rect 2547 8517 2559 8551
rect 2501 8511 2559 8517
rect 3421 8551 3479 8557
rect 3421 8517 3433 8551
rect 3467 8548 3479 8551
rect 4062 8548 4068 8560
rect 3467 8520 4068 8548
rect 3467 8517 3479 8520
rect 3421 8511 3479 8517
rect 4062 8508 4068 8520
rect 4120 8508 4126 8560
rect 4249 8551 4307 8557
rect 4249 8517 4261 8551
rect 4295 8548 4307 8551
rect 4430 8548 4436 8560
rect 4295 8520 4436 8548
rect 4295 8517 4307 8520
rect 4249 8511 4307 8517
rect 4430 8508 4436 8520
rect 4488 8548 4494 8560
rect 5350 8548 5356 8560
rect 4488 8520 5356 8548
rect 4488 8508 4494 8520
rect 5350 8508 5356 8520
rect 5408 8548 5414 8560
rect 5988 8551 6046 8557
rect 5988 8548 6000 8551
rect 5408 8520 6000 8548
rect 5408 8508 5414 8520
rect 5988 8517 6000 8520
rect 6034 8548 6046 8551
rect 7466 8548 7472 8560
rect 6034 8520 7472 8548
rect 6034 8517 6046 8520
rect 5988 8511 6046 8517
rect 7466 8508 7472 8520
rect 7524 8548 7530 8560
rect 8956 8548 8984 8579
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 11057 8619 11115 8625
rect 9732 8588 10640 8616
rect 9732 8576 9738 8588
rect 10612 8560 10640 8588
rect 11057 8585 11069 8619
rect 11103 8616 11115 8619
rect 11238 8616 11244 8628
rect 11103 8588 11244 8616
rect 11103 8585 11115 8588
rect 11057 8579 11115 8585
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 11514 8616 11520 8628
rect 11475 8588 11520 8616
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11609 8619 11667 8625
rect 11609 8585 11621 8619
rect 11655 8616 11667 8619
rect 11655 8588 13032 8616
rect 11655 8585 11667 8588
rect 11609 8579 11667 8585
rect 10134 8548 10140 8560
rect 7524 8520 7604 8548
rect 8956 8520 10140 8548
rect 7524 8508 7530 8520
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2682 8480 2688 8492
rect 2643 8452 2688 8480
rect 2317 8443 2375 8449
rect 615 8384 2268 8412
rect 615 8381 627 8384
rect 569 8375 627 8381
rect 2041 8347 2099 8353
rect 2041 8313 2053 8347
rect 2087 8344 2099 8347
rect 2222 8344 2228 8356
rect 2087 8316 2228 8344
rect 2087 8313 2099 8316
rect 2041 8307 2099 8313
rect 2222 8304 2228 8316
rect 2280 8304 2286 8356
rect 2332 8344 2360 8443
rect 2682 8440 2688 8452
rect 2740 8440 2746 8492
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 3329 8483 3387 8489
rect 3329 8480 3341 8483
rect 2832 8452 3341 8480
rect 2832 8440 2838 8452
rect 3329 8449 3341 8452
rect 3375 8449 3387 8483
rect 4522 8480 4528 8492
rect 3329 8443 3387 8449
rect 3620 8452 4528 8480
rect 2406 8372 2412 8424
rect 2464 8412 2470 8424
rect 3620 8421 3648 8452
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 7282 8480 7288 8492
rect 7116 8452 7288 8480
rect 2501 8415 2559 8421
rect 2501 8412 2513 8415
rect 2464 8384 2513 8412
rect 2464 8372 2470 8384
rect 2501 8381 2513 8384
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 3605 8415 3663 8421
rect 3605 8381 3617 8415
rect 3651 8381 3663 8415
rect 3605 8375 3663 8381
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 3789 8347 3847 8353
rect 3789 8344 3801 8347
rect 2332 8316 3801 8344
rect 3789 8313 3801 8316
rect 3835 8313 3847 8347
rect 4448 8344 4476 8375
rect 4982 8372 4988 8424
rect 5040 8412 5046 8424
rect 5353 8415 5411 8421
rect 5353 8412 5365 8415
rect 5040 8384 5365 8412
rect 5040 8372 5046 8384
rect 5353 8381 5365 8384
rect 5399 8381 5411 8415
rect 5353 8375 5411 8381
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8381 5503 8415
rect 5445 8375 5503 8381
rect 5721 8415 5779 8421
rect 5721 8381 5733 8415
rect 5767 8381 5779 8415
rect 5721 8375 5779 8381
rect 5166 8344 5172 8356
rect 4448 8316 5172 8344
rect 3789 8307 3847 8313
rect 5166 8304 5172 8316
rect 5224 8344 5230 8356
rect 5460 8344 5488 8375
rect 5224 8316 5488 8344
rect 5224 8304 5230 8316
rect 2958 8276 2964 8288
rect 2919 8248 2964 8276
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 5736 8276 5764 8375
rect 7116 8353 7144 8452
rect 7282 8440 7288 8452
rect 7340 8480 7346 8492
rect 7576 8489 7604 8520
rect 10134 8508 10140 8520
rect 10192 8508 10198 8560
rect 10594 8508 10600 8560
rect 10652 8548 10658 8560
rect 10965 8551 11023 8557
rect 10965 8548 10977 8551
rect 10652 8520 10977 8548
rect 10652 8508 10658 8520
rect 10965 8517 10977 8520
rect 11011 8517 11023 8551
rect 12894 8548 12900 8560
rect 10965 8511 11023 8517
rect 11072 8520 12900 8548
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 7340 8452 7389 8480
rect 7340 8440 7346 8452
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8449 7619 8483
rect 7561 8443 7619 8449
rect 7745 8483 7803 8489
rect 7745 8449 7757 8483
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8412 7527 8415
rect 7760 8412 7788 8443
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 8481 8483 8539 8489
rect 8481 8480 8493 8483
rect 8444 8452 8493 8480
rect 8444 8440 8450 8452
rect 8481 8449 8493 8452
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 7515 8384 7788 8412
rect 8021 8415 8079 8421
rect 7515 8381 7527 8384
rect 7469 8375 7527 8381
rect 8021 8381 8033 8415
rect 8067 8381 8079 8415
rect 8496 8412 8524 8443
rect 8570 8440 8576 8492
rect 8628 8480 8634 8492
rect 11072 8489 11100 8520
rect 12894 8508 12900 8520
rect 12952 8508 12958 8560
rect 13004 8557 13032 8588
rect 14550 8576 14556 8628
rect 14608 8616 14614 8628
rect 14645 8619 14703 8625
rect 14645 8616 14657 8619
rect 14608 8588 14657 8616
rect 14608 8576 14614 8588
rect 14645 8585 14657 8588
rect 14691 8585 14703 8619
rect 14645 8579 14703 8585
rect 14875 8619 14933 8625
rect 14875 8585 14887 8619
rect 14921 8616 14933 8619
rect 15838 8616 15844 8628
rect 14921 8588 15844 8616
rect 14921 8585 14933 8588
rect 14875 8579 14933 8585
rect 12989 8551 13047 8557
rect 12989 8517 13001 8551
rect 13035 8548 13047 8551
rect 13446 8548 13452 8560
rect 13035 8520 13452 8548
rect 13035 8517 13047 8520
rect 12989 8511 13047 8517
rect 13446 8508 13452 8520
rect 13504 8508 13510 8560
rect 14660 8548 14688 8579
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 18325 8619 18383 8625
rect 18325 8585 18337 8619
rect 18371 8585 18383 8619
rect 18325 8579 18383 8585
rect 15102 8548 15108 8560
rect 14660 8520 15108 8548
rect 15102 8508 15108 8520
rect 15160 8548 15166 8560
rect 15160 8520 15318 8548
rect 15160 8508 15166 8520
rect 9033 8483 9091 8489
rect 9033 8480 9045 8483
rect 8628 8452 9045 8480
rect 8628 8440 8634 8452
rect 9033 8449 9045 8452
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 8662 8412 8668 8424
rect 8496 8384 8668 8412
rect 8021 8375 8079 8381
rect 7101 8347 7159 8353
rect 7101 8313 7113 8347
rect 7147 8313 7159 8347
rect 8036 8344 8064 8375
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 10796 8412 10824 8443
rect 11974 8440 11980 8492
rect 12032 8480 12038 8492
rect 12253 8483 12311 8489
rect 12253 8480 12265 8483
rect 12032 8452 12265 8480
rect 12032 8440 12038 8452
rect 12253 8449 12265 8452
rect 12299 8449 12311 8483
rect 12253 8443 12311 8449
rect 12713 8483 12771 8489
rect 12713 8449 12725 8483
rect 12759 8480 12771 8483
rect 12802 8480 12808 8492
rect 12759 8452 12808 8480
rect 12759 8449 12771 8452
rect 12713 8443 12771 8449
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 13354 8480 13360 8492
rect 13315 8452 13360 8480
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 14185 8483 14243 8489
rect 14185 8449 14197 8483
rect 14231 8480 14243 8483
rect 14366 8480 14372 8492
rect 14231 8452 14372 8480
rect 14231 8449 14243 8452
rect 14185 8443 14243 8449
rect 11698 8412 11704 8424
rect 10796 8384 11704 8412
rect 11698 8372 11704 8384
rect 11756 8372 11762 8424
rect 11793 8415 11851 8421
rect 11793 8381 11805 8415
rect 11839 8381 11851 8415
rect 11793 8375 11851 8381
rect 11149 8347 11207 8353
rect 8036 8316 11100 8344
rect 7101 8307 7159 8313
rect 6086 8276 6092 8288
rect 5736 8248 6092 8276
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 7837 8279 7895 8285
rect 7837 8276 7849 8279
rect 7708 8248 7849 8276
rect 7708 8236 7714 8248
rect 7837 8245 7849 8248
rect 7883 8245 7895 8279
rect 7837 8239 7895 8245
rect 7926 8236 7932 8288
rect 7984 8276 7990 8288
rect 8570 8276 8576 8288
rect 7984 8248 8029 8276
rect 8531 8248 8576 8276
rect 7984 8236 7990 8248
rect 8570 8236 8576 8248
rect 8628 8236 8634 8288
rect 8662 8236 8668 8288
rect 8720 8276 8726 8288
rect 9309 8279 9367 8285
rect 9309 8276 9321 8279
rect 8720 8248 9321 8276
rect 8720 8236 8726 8248
rect 9309 8245 9321 8248
rect 9355 8276 9367 8279
rect 10778 8276 10784 8288
rect 9355 8248 10784 8276
rect 9355 8245 9367 8248
rect 9309 8239 9367 8245
rect 10778 8236 10784 8248
rect 10836 8236 10842 8288
rect 11072 8276 11100 8316
rect 11149 8313 11161 8347
rect 11195 8344 11207 8347
rect 11330 8344 11336 8356
rect 11195 8316 11336 8344
rect 11195 8313 11207 8316
rect 11149 8307 11207 8313
rect 11330 8304 11336 8316
rect 11388 8304 11394 8356
rect 11808 8344 11836 8375
rect 12158 8372 12164 8424
rect 12216 8412 12222 8424
rect 12529 8415 12587 8421
rect 12529 8412 12541 8415
rect 12216 8384 12541 8412
rect 12216 8372 12222 8384
rect 12529 8381 12541 8384
rect 12575 8381 12587 8415
rect 13262 8412 13268 8424
rect 13223 8384 13268 8412
rect 12529 8375 12587 8381
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 14016 8412 14044 8443
rect 14366 8440 14372 8452
rect 14424 8440 14430 8492
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8480 16359 8483
rect 18340 8480 18368 8579
rect 16347 8452 18368 8480
rect 18509 8483 18567 8489
rect 16347 8449 16359 8452
rect 16301 8443 16359 8449
rect 18509 8449 18521 8483
rect 18555 8480 18567 8483
rect 18598 8480 18604 8492
rect 18555 8452 18604 8480
rect 18555 8449 18567 8452
rect 18509 8443 18567 8449
rect 14458 8412 14464 8424
rect 14016 8384 14464 8412
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 16666 8412 16672 8424
rect 16579 8384 16672 8412
rect 16666 8372 16672 8384
rect 16724 8412 16730 8424
rect 17862 8412 17868 8424
rect 16724 8384 17868 8412
rect 16724 8372 16730 8384
rect 17862 8372 17868 8384
rect 17920 8372 17926 8424
rect 18233 8415 18291 8421
rect 18233 8381 18245 8415
rect 18279 8412 18291 8415
rect 18524 8412 18552 8443
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 18279 8384 18552 8412
rect 18279 8381 18291 8384
rect 18233 8375 18291 8381
rect 12710 8344 12716 8356
rect 11808 8316 12716 8344
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 11238 8276 11244 8288
rect 11072 8248 11244 8276
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 12161 8279 12219 8285
rect 12161 8245 12173 8279
rect 12207 8276 12219 8279
rect 12250 8276 12256 8288
rect 12207 8248 12256 8276
rect 12207 8245 12219 8248
rect 12161 8239 12219 8245
rect 12250 8236 12256 8248
rect 12308 8236 12314 8288
rect 14001 8279 14059 8285
rect 14001 8245 14013 8279
rect 14047 8276 14059 8279
rect 14274 8276 14280 8288
rect 14047 8248 14280 8276
rect 14047 8245 14059 8248
rect 14001 8239 14059 8245
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 0 8186 18860 8208
rect 0 8134 3110 8186
rect 3162 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 6210 8186
rect 6262 8134 6274 8186
rect 6326 8134 6338 8186
rect 6390 8134 6402 8186
rect 6454 8134 6466 8186
rect 6518 8134 9310 8186
rect 9362 8134 9374 8186
rect 9426 8134 9438 8186
rect 9490 8134 9502 8186
rect 9554 8134 9566 8186
rect 9618 8134 12410 8186
rect 12462 8134 12474 8186
rect 12526 8134 12538 8186
rect 12590 8134 12602 8186
rect 12654 8134 12666 8186
rect 12718 8134 15510 8186
rect 15562 8134 15574 8186
rect 15626 8134 15638 8186
rect 15690 8134 15702 8186
rect 15754 8134 15766 8186
rect 15818 8134 18860 8186
rect 0 8112 18860 8134
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2188 8044 2237 8072
rect 2188 8032 2194 8044
rect 2225 8041 2237 8044
rect 2271 8072 2283 8075
rect 2682 8072 2688 8084
rect 2271 8044 2688 8072
rect 2271 8041 2283 8044
rect 2225 8035 2283 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 9766 8072 9772 8084
rect 4304 8044 9772 8072
rect 4304 8032 4310 8044
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 12437 8075 12495 8081
rect 12437 8041 12449 8075
rect 12483 8072 12495 8075
rect 12894 8072 12900 8084
rect 12483 8044 12900 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 13725 8075 13783 8081
rect 13725 8072 13737 8075
rect 13412 8044 13737 8072
rect 13412 8032 13418 8044
rect 13725 8041 13737 8044
rect 13771 8041 13783 8075
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 13725 8035 13783 8041
rect 15102 8032 15108 8044
rect 15160 8072 15166 8084
rect 15657 8075 15715 8081
rect 15657 8072 15669 8075
rect 15160 8044 15669 8072
rect 15160 8032 15166 8044
rect 15657 8041 15669 8044
rect 15703 8072 15715 8075
rect 16482 8072 16488 8084
rect 15703 8044 16488 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 1857 8007 1915 8013
rect 1857 7973 1869 8007
rect 1903 8004 1915 8007
rect 2774 8004 2780 8016
rect 1903 7976 2780 8004
rect 1903 7973 1915 7976
rect 1857 7967 1915 7973
rect 2774 7964 2780 7976
rect 2832 7964 2838 8016
rect 5074 7964 5080 8016
rect 5132 8004 5138 8016
rect 5350 8004 5356 8016
rect 5132 7976 5356 8004
rect 5132 7964 5138 7976
rect 5350 7964 5356 7976
rect 5408 8004 5414 8016
rect 5445 8007 5503 8013
rect 5445 8004 5457 8007
rect 5408 7976 5457 8004
rect 5408 7964 5414 7976
rect 5445 7973 5457 7976
rect 5491 7973 5503 8007
rect 7650 8004 7656 8016
rect 7611 7976 7656 8004
rect 5445 7967 5503 7973
rect 7650 7964 7656 7976
rect 7708 7964 7714 8016
rect 7926 8004 7932 8016
rect 7887 7976 7932 8004
rect 7926 7964 7932 7976
rect 7984 7964 7990 8016
rect 11330 8004 11336 8016
rect 9784 7976 11336 8004
rect 2222 7936 2228 7948
rect 1964 7908 2228 7936
rect 1964 7877 1992 7908
rect 2222 7896 2228 7908
rect 2280 7896 2286 7948
rect 2498 7936 2504 7948
rect 2459 7908 2504 7936
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 3237 7939 3295 7945
rect 3237 7905 3249 7939
rect 3283 7936 3295 7939
rect 3510 7936 3516 7948
rect 3283 7908 3516 7936
rect 3283 7905 3295 7908
rect 3237 7899 3295 7905
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 5258 7936 5264 7948
rect 5219 7908 5264 7936
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 6638 7936 6644 7948
rect 5552 7908 6644 7936
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7837 2007 7871
rect 2130 7868 2136 7880
rect 2091 7840 2136 7868
rect 1949 7831 2007 7837
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 2314 7868 2320 7880
rect 2275 7840 2320 7868
rect 2314 7828 2320 7840
rect 2372 7828 2378 7880
rect 2958 7868 2964 7880
rect 2919 7840 2964 7868
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 4982 7828 4988 7880
rect 5040 7868 5046 7880
rect 5552 7877 5580 7908
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 7282 7936 7288 7948
rect 7243 7908 7288 7936
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 8294 7936 8300 7948
rect 7883 7908 8300 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 8478 7936 8484 7948
rect 8439 7908 8484 7936
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 9784 7936 9812 7976
rect 11330 7964 11336 7976
rect 11388 8004 11394 8016
rect 11885 8007 11943 8013
rect 11388 7976 11560 8004
rect 11388 7964 11394 7976
rect 11422 7936 11428 7948
rect 9180 7908 9812 7936
rect 11383 7908 11428 7936
rect 9180 7896 9186 7908
rect 11422 7896 11428 7908
rect 11480 7896 11486 7948
rect 11532 7936 11560 7976
rect 11885 7973 11897 8007
rect 11931 8004 11943 8007
rect 12802 8004 12808 8016
rect 11931 7976 12808 8004
rect 11931 7973 11943 7976
rect 11885 7967 11943 7973
rect 12802 7964 12808 7976
rect 12860 7964 12866 8016
rect 13740 7976 14872 8004
rect 13740 7948 13768 7976
rect 11532 7908 12434 7936
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 5040 7840 5549 7868
rect 5040 7828 5046 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 6086 7828 6092 7880
rect 6144 7868 6150 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 6144 7840 6469 7868
rect 6144 7828 6150 7840
rect 6457 7837 6469 7840
rect 6503 7837 6515 7871
rect 7466 7868 7472 7880
rect 7427 7840 7472 7868
rect 6457 7831 6515 7837
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 8110 7868 8116 7880
rect 8071 7840 8116 7868
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7868 11575 7871
rect 11974 7868 11980 7880
rect 11563 7840 11980 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 12069 7871 12127 7877
rect 12069 7837 12081 7871
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12161 7871 12219 7877
rect 12161 7837 12173 7871
rect 12207 7837 12219 7871
rect 12161 7831 12219 7837
rect 5261 7803 5319 7809
rect 5261 7769 5273 7803
rect 5307 7800 5319 7803
rect 5350 7800 5356 7812
rect 5307 7772 5356 7800
rect 5307 7769 5319 7772
rect 5261 7763 5319 7769
rect 5350 7760 5356 7772
rect 5408 7800 5414 7812
rect 6181 7803 6239 7809
rect 6181 7800 6193 7803
rect 5408 7772 6193 7800
rect 5408 7760 5414 7772
rect 6181 7769 6193 7772
rect 6227 7769 6239 7803
rect 6181 7763 6239 7769
rect 6365 7803 6423 7809
rect 6365 7769 6377 7803
rect 6411 7800 6423 7803
rect 6546 7800 6552 7812
rect 6411 7772 6552 7800
rect 6411 7769 6423 7772
rect 6365 7763 6423 7769
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 6641 7803 6699 7809
rect 6641 7769 6653 7803
rect 6687 7800 6699 7803
rect 8386 7800 8392 7812
rect 6687 7772 8392 7800
rect 6687 7769 6699 7772
rect 6641 7763 6699 7769
rect 8386 7760 8392 7772
rect 8444 7760 8450 7812
rect 8757 7803 8815 7809
rect 8757 7769 8769 7803
rect 8803 7769 8815 7803
rect 10042 7800 10048 7812
rect 9982 7772 10048 7800
rect 8757 7763 8815 7769
rect 2498 7692 2504 7744
rect 2556 7732 2562 7744
rect 2593 7735 2651 7741
rect 2593 7732 2605 7735
rect 2556 7704 2605 7732
rect 2556 7692 2562 7704
rect 2593 7701 2605 7704
rect 2639 7701 2651 7735
rect 2593 7695 2651 7701
rect 3053 7735 3111 7741
rect 3053 7701 3065 7735
rect 3099 7732 3111 7735
rect 4154 7732 4160 7744
rect 3099 7704 4160 7732
rect 3099 7701 3111 7704
rect 3053 7695 3111 7701
rect 4154 7692 4160 7704
rect 4212 7692 4218 7744
rect 8297 7735 8355 7741
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 8772 7732 8800 7763
rect 10042 7760 10048 7772
rect 10100 7760 10106 7812
rect 10134 7760 10140 7812
rect 10192 7800 10198 7812
rect 10505 7803 10563 7809
rect 10505 7800 10517 7803
rect 10192 7772 10517 7800
rect 10192 7760 10198 7772
rect 10505 7769 10517 7772
rect 10551 7769 10563 7803
rect 10505 7763 10563 7769
rect 11790 7760 11796 7812
rect 11848 7800 11854 7812
rect 12084 7800 12112 7831
rect 11848 7772 12112 7800
rect 11848 7760 11854 7772
rect 8343 7704 8800 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 11238 7692 11244 7744
rect 11296 7732 11302 7744
rect 12176 7732 12204 7831
rect 12250 7828 12256 7880
rect 12308 7868 12314 7880
rect 12406 7868 12434 7908
rect 13722 7896 13728 7948
rect 13780 7896 13786 7948
rect 14274 7936 14280 7948
rect 14235 7908 14280 7936
rect 14274 7896 14280 7908
rect 14332 7896 14338 7948
rect 12989 7871 13047 7877
rect 12989 7868 13001 7871
rect 12308 7840 12353 7868
rect 12406 7840 13001 7868
rect 12308 7828 12314 7840
rect 12989 7837 13001 7840
rect 13035 7868 13047 7871
rect 13538 7868 13544 7880
rect 13035 7840 13544 7868
rect 13035 7837 13047 7840
rect 12989 7831 13047 7837
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7868 14151 7871
rect 14550 7868 14556 7880
rect 14139 7840 14556 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 14550 7828 14556 7840
rect 14608 7828 14614 7880
rect 14844 7877 14872 7976
rect 15841 7939 15899 7945
rect 15841 7905 15853 7939
rect 15887 7936 15899 7939
rect 16666 7936 16672 7948
rect 15887 7908 16672 7936
rect 15887 7905 15899 7908
rect 15841 7899 15899 7905
rect 16666 7896 16672 7908
rect 16724 7896 16730 7948
rect 14829 7871 14887 7877
rect 14829 7837 14841 7871
rect 14875 7837 14887 7871
rect 14829 7831 14887 7837
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7837 15071 7871
rect 15013 7831 15071 7837
rect 13081 7803 13139 7809
rect 13081 7769 13093 7803
rect 13127 7800 13139 7803
rect 13262 7800 13268 7812
rect 13127 7772 13268 7800
rect 13127 7769 13139 7772
rect 13081 7763 13139 7769
rect 13262 7760 13268 7772
rect 13320 7800 13326 7812
rect 13630 7800 13636 7812
rect 13320 7772 13636 7800
rect 13320 7760 13326 7772
rect 13630 7760 13636 7772
rect 13688 7760 13694 7812
rect 13814 7760 13820 7812
rect 13872 7800 13878 7812
rect 14185 7803 14243 7809
rect 14185 7800 14197 7803
rect 13872 7772 14197 7800
rect 13872 7760 13878 7772
rect 14185 7769 14197 7772
rect 14231 7769 14243 7803
rect 14185 7763 14243 7769
rect 14366 7760 14372 7812
rect 14424 7800 14430 7812
rect 15028 7800 15056 7831
rect 16114 7800 16120 7812
rect 14424 7772 15056 7800
rect 16075 7772 16120 7800
rect 14424 7760 14430 7772
rect 16114 7760 16120 7772
rect 16172 7760 16178 7812
rect 16574 7760 16580 7812
rect 16632 7760 16638 7812
rect 17494 7760 17500 7812
rect 17552 7800 17558 7812
rect 17865 7803 17923 7809
rect 17865 7800 17877 7803
rect 17552 7772 17877 7800
rect 17552 7760 17558 7772
rect 17865 7769 17877 7772
rect 17911 7769 17923 7803
rect 17865 7763 17923 7769
rect 11296 7704 12204 7732
rect 11296 7692 11302 7704
rect 13446 7692 13452 7744
rect 13504 7732 13510 7744
rect 14642 7732 14648 7744
rect 13504 7704 14648 7732
rect 13504 7692 13510 7704
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 15010 7732 15016 7744
rect 14971 7704 15016 7732
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 0 7642 18860 7664
rect 0 7590 4660 7642
rect 4712 7590 4724 7642
rect 4776 7590 4788 7642
rect 4840 7590 4852 7642
rect 4904 7590 4916 7642
rect 4968 7590 7760 7642
rect 7812 7590 7824 7642
rect 7876 7590 7888 7642
rect 7940 7590 7952 7642
rect 8004 7590 8016 7642
rect 8068 7590 10860 7642
rect 10912 7590 10924 7642
rect 10976 7590 10988 7642
rect 11040 7590 11052 7642
rect 11104 7590 11116 7642
rect 11168 7590 13960 7642
rect 14012 7590 14024 7642
rect 14076 7590 14088 7642
rect 14140 7590 14152 7642
rect 14204 7590 14216 7642
rect 14268 7590 17060 7642
rect 17112 7590 17124 7642
rect 17176 7590 17188 7642
rect 17240 7590 17252 7642
rect 17304 7590 17316 7642
rect 17368 7590 18860 7642
rect 0 7568 18860 7590
rect 2130 7488 2136 7540
rect 2188 7488 2194 7540
rect 2225 7531 2283 7537
rect 2225 7497 2237 7531
rect 2271 7528 2283 7531
rect 2406 7528 2412 7540
rect 2271 7500 2412 7528
rect 2271 7497 2283 7500
rect 2225 7491 2283 7497
rect 2406 7488 2412 7500
rect 2464 7488 2470 7540
rect 4709 7531 4767 7537
rect 4709 7497 4721 7531
rect 4755 7528 4767 7531
rect 5442 7528 5448 7540
rect 4755 7500 5448 7528
rect 4755 7497 4767 7500
rect 4709 7491 4767 7497
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 7190 7488 7196 7540
rect 7248 7528 7254 7540
rect 8941 7531 8999 7537
rect 8941 7528 8953 7531
rect 7248 7500 8953 7528
rect 7248 7488 7254 7500
rect 8941 7497 8953 7500
rect 8987 7528 8999 7531
rect 9122 7528 9128 7540
rect 8987 7500 9128 7528
rect 8987 7497 8999 7500
rect 8941 7491 8999 7497
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 10686 7528 10692 7540
rect 10647 7500 10692 7528
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11333 7531 11391 7537
rect 11333 7528 11345 7531
rect 11296 7500 11345 7528
rect 11296 7488 11302 7500
rect 11333 7497 11345 7500
rect 11379 7497 11391 7531
rect 11698 7528 11704 7540
rect 11659 7500 11704 7528
rect 11333 7491 11391 7497
rect 11698 7488 11704 7500
rect 11756 7488 11762 7540
rect 13722 7528 13728 7540
rect 13683 7500 13728 7528
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 13909 7531 13967 7537
rect 13909 7497 13921 7531
rect 13955 7497 13967 7531
rect 13909 7491 13967 7497
rect 1946 7460 1952 7472
rect 1794 7432 1952 7460
rect 1946 7420 1952 7432
rect 2004 7420 2010 7472
rect 2148 7460 2176 7488
rect 2593 7463 2651 7469
rect 2593 7460 2605 7463
rect 2148 7432 2605 7460
rect 2593 7429 2605 7432
rect 2639 7429 2651 7463
rect 2593 7423 2651 7429
rect 2777 7463 2835 7469
rect 2777 7429 2789 7463
rect 2823 7460 2835 7463
rect 2866 7460 2872 7472
rect 2823 7432 2872 7460
rect 2823 7429 2835 7432
rect 2777 7423 2835 7429
rect 2038 7352 2044 7404
rect 2096 7392 2102 7404
rect 2133 7395 2191 7401
rect 2133 7392 2145 7395
rect 2096 7364 2145 7392
rect 2096 7352 2102 7364
rect 2133 7361 2145 7364
rect 2179 7361 2191 7395
rect 2133 7355 2191 7361
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 2498 7392 2504 7404
rect 2363 7364 2504 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 2608 7392 2636 7423
rect 2866 7420 2872 7432
rect 2924 7420 2930 7472
rect 4356 7432 5028 7460
rect 3421 7395 3479 7401
rect 2608 7364 3004 7392
rect 290 7324 296 7336
rect 251 7296 296 7324
rect 290 7284 296 7296
rect 348 7284 354 7336
rect 566 7324 572 7336
rect 527 7296 572 7324
rect 566 7284 572 7296
rect 624 7284 630 7336
rect 2976 7333 3004 7364
rect 3421 7361 3433 7395
rect 3467 7392 3479 7395
rect 3510 7392 3516 7404
rect 3467 7364 3516 7392
rect 3467 7361 3479 7364
rect 3421 7355 3479 7361
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 4062 7392 4068 7404
rect 4023 7364 4068 7392
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4246 7392 4252 7404
rect 4207 7364 4252 7392
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 4356 7401 4384 7432
rect 5000 7404 5028 7432
rect 5258 7420 5264 7472
rect 5316 7460 5322 7472
rect 7208 7460 7236 7488
rect 5316 7432 7236 7460
rect 5316 7420 5322 7432
rect 8386 7420 8392 7472
rect 8444 7460 8450 7472
rect 10597 7463 10655 7469
rect 10597 7460 10609 7463
rect 8444 7432 10609 7460
rect 8444 7420 8450 7432
rect 10597 7429 10609 7432
rect 10643 7429 10655 7463
rect 13924 7460 13952 7491
rect 13998 7460 14004 7472
rect 10597 7423 10655 7429
rect 10796 7432 11652 7460
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 4890 7392 4896 7404
rect 4479 7364 4896 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 4982 7352 4988 7404
rect 5040 7352 5046 7404
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7361 5135 7395
rect 5350 7392 5356 7404
rect 5311 7364 5356 7392
rect 5077 7355 5135 7361
rect 2961 7327 3019 7333
rect 2961 7293 2973 7327
rect 3007 7324 3019 7327
rect 5092 7324 5120 7355
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 5813 7395 5871 7401
rect 5491 7364 5764 7392
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 5626 7324 5632 7336
rect 3007 7296 5632 7324
rect 3007 7293 3019 7296
rect 2961 7287 3019 7293
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 5736 7333 5764 7364
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 6914 7392 6920 7404
rect 5859 7364 6920 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7098 7352 7104 7404
rect 7156 7392 7162 7404
rect 7745 7395 7803 7401
rect 7745 7392 7757 7395
rect 7156 7364 7757 7392
rect 7156 7352 7162 7364
rect 7745 7361 7757 7364
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8662 7392 8668 7404
rect 7883 7364 8668 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7324 5779 7327
rect 5767 7296 5856 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 5828 7268 5856 7296
rect 5902 7284 5908 7336
rect 5960 7324 5966 7336
rect 6181 7327 6239 7333
rect 6181 7324 6193 7327
rect 5960 7296 6193 7324
rect 5960 7284 5966 7296
rect 6181 7293 6193 7296
rect 6227 7293 6239 7327
rect 6181 7287 6239 7293
rect 6638 7284 6644 7336
rect 6696 7324 6702 7336
rect 7852 7324 7880 7355
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 8846 7392 8852 7404
rect 8807 7364 8852 7392
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 9858 7352 9864 7404
rect 9916 7392 9922 7404
rect 10229 7395 10287 7401
rect 10229 7392 10241 7395
rect 9916 7364 10241 7392
rect 9916 7352 9922 7364
rect 10229 7361 10241 7364
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 10413 7395 10471 7401
rect 10413 7361 10425 7395
rect 10459 7392 10471 7395
rect 10502 7392 10508 7404
rect 10459 7364 10508 7392
rect 10459 7361 10471 7364
rect 10413 7355 10471 7361
rect 10502 7352 10508 7364
rect 10560 7352 10566 7404
rect 6696 7296 7880 7324
rect 6696 7284 6702 7296
rect 8018 7284 8024 7336
rect 8076 7324 8082 7336
rect 8076 7296 8294 7324
rect 8076 7284 8082 7296
rect 2041 7259 2099 7265
rect 2041 7225 2053 7259
rect 2087 7256 2099 7259
rect 2087 7228 2774 7256
rect 2087 7225 2099 7228
rect 2041 7219 2099 7225
rect 2746 7188 2774 7228
rect 5810 7216 5816 7268
rect 5868 7216 5874 7268
rect 8266 7256 8294 7296
rect 9030 7284 9036 7336
rect 9088 7324 9094 7336
rect 10321 7327 10379 7333
rect 9088 7296 9133 7324
rect 9088 7284 9094 7296
rect 10321 7293 10333 7327
rect 10367 7324 10379 7327
rect 10796 7324 10824 7432
rect 10870 7352 10876 7404
rect 10928 7392 10934 7404
rect 11149 7395 11207 7401
rect 10928 7364 10973 7392
rect 10928 7352 10934 7364
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11330 7392 11336 7404
rect 11195 7364 11336 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 11624 7401 11652 7432
rect 11425 7395 11483 7401
rect 11425 7361 11437 7395
rect 11471 7361 11483 7395
rect 11425 7355 11483 7361
rect 11609 7395 11667 7401
rect 11609 7361 11621 7395
rect 11655 7392 11667 7395
rect 11790 7392 11796 7404
rect 11655 7364 11796 7392
rect 11655 7361 11667 7364
rect 11609 7355 11667 7361
rect 10367 7296 10824 7324
rect 10367 7293 10379 7296
rect 10321 7287 10379 7293
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 11440 7324 11468 7355
rect 11790 7352 11796 7364
rect 11848 7352 11854 7404
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7392 11943 7395
rect 12250 7392 12256 7404
rect 11931 7364 12256 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 13446 7392 13452 7404
rect 13407 7364 13452 7392
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 13630 7392 13636 7404
rect 13591 7364 13636 7392
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 13722 7386 13728 7438
rect 13780 7386 13786 7438
rect 13924 7432 14004 7460
rect 13998 7420 14004 7432
rect 14056 7420 14062 7472
rect 14277 7463 14335 7469
rect 14277 7429 14289 7463
rect 14323 7460 14335 7463
rect 14366 7460 14372 7472
rect 14323 7432 14372 7460
rect 14323 7429 14335 7432
rect 14277 7423 14335 7429
rect 14366 7420 14372 7432
rect 14424 7420 14430 7472
rect 14550 7469 14556 7472
rect 14507 7463 14556 7469
rect 14507 7429 14519 7463
rect 14553 7429 14556 7463
rect 14507 7423 14556 7429
rect 14550 7420 14556 7423
rect 14608 7420 14614 7472
rect 15102 7420 15108 7472
rect 15160 7420 15166 7472
rect 13817 7395 13875 7401
rect 13723 7383 13735 7386
rect 13769 7383 13781 7386
rect 13723 7377 13781 7383
rect 13817 7361 13829 7395
rect 13863 7390 13875 7395
rect 13906 7390 13912 7404
rect 13863 7362 13912 7390
rect 13863 7361 13875 7362
rect 13817 7355 13875 7361
rect 13906 7352 13912 7362
rect 13964 7352 13970 7404
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7392 14151 7395
rect 14642 7392 14648 7404
rect 14139 7364 14648 7392
rect 14139 7361 14151 7364
rect 14093 7355 14151 7361
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 12158 7324 12164 7336
rect 11112 7296 12164 7324
rect 11112 7284 11118 7296
rect 12158 7284 12164 7296
rect 12216 7284 12222 7336
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 15933 7327 15991 7333
rect 15933 7324 15945 7327
rect 15068 7296 15945 7324
rect 15068 7284 15074 7296
rect 15933 7293 15945 7296
rect 15979 7293 15991 7327
rect 16298 7324 16304 7336
rect 16259 7296 16304 7324
rect 15933 7287 15991 7293
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 10042 7256 10048 7268
rect 8266 7228 10048 7256
rect 10042 7216 10048 7228
rect 10100 7216 10106 7268
rect 10137 7259 10195 7265
rect 10137 7225 10149 7259
rect 10183 7256 10195 7259
rect 10226 7256 10232 7268
rect 10183 7228 10232 7256
rect 10183 7225 10195 7228
rect 10137 7219 10195 7225
rect 10226 7216 10232 7228
rect 10284 7256 10290 7268
rect 10284 7228 14688 7256
rect 10284 7216 10290 7228
rect 2958 7188 2964 7200
rect 2746 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 5534 7188 5540 7200
rect 5495 7160 5540 7188
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 7374 7188 7380 7200
rect 7335 7160 7380 7188
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 8294 7188 8300 7200
rect 8255 7160 8300 7188
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 8478 7188 8484 7200
rect 8439 7160 8484 7188
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 10962 7188 10968 7200
rect 10923 7160 10968 7188
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 13722 7148 13728 7200
rect 13780 7188 13786 7200
rect 13998 7188 14004 7200
rect 13780 7160 14004 7188
rect 13780 7148 13786 7160
rect 13998 7148 14004 7160
rect 14056 7188 14062 7200
rect 14366 7188 14372 7200
rect 14056 7160 14372 7188
rect 14056 7148 14062 7160
rect 14366 7148 14372 7160
rect 14424 7148 14430 7200
rect 14660 7188 14688 7228
rect 18506 7188 18512 7200
rect 14660 7160 18512 7188
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 0 7098 18860 7120
rect 0 7046 3110 7098
rect 3162 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 6210 7098
rect 6262 7046 6274 7098
rect 6326 7046 6338 7098
rect 6390 7046 6402 7098
rect 6454 7046 6466 7098
rect 6518 7046 9310 7098
rect 9362 7046 9374 7098
rect 9426 7046 9438 7098
rect 9490 7046 9502 7098
rect 9554 7046 9566 7098
rect 9618 7046 12410 7098
rect 12462 7046 12474 7098
rect 12526 7046 12538 7098
rect 12590 7046 12602 7098
rect 12654 7046 12666 7098
rect 12718 7046 15510 7098
rect 15562 7046 15574 7098
rect 15626 7046 15638 7098
rect 15690 7046 15702 7098
rect 15754 7046 15766 7098
rect 15818 7046 18860 7098
rect 0 7024 18860 7046
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 2133 6987 2191 6993
rect 2133 6984 2145 6987
rect 2004 6956 2145 6984
rect 2004 6944 2010 6956
rect 2133 6953 2145 6956
rect 2179 6953 2191 6987
rect 6914 6984 6920 6996
rect 6875 6956 6920 6984
rect 2133 6947 2191 6953
rect 6914 6944 6920 6956
rect 6972 6944 6978 6996
rect 7466 6944 7472 6996
rect 7524 6984 7530 6996
rect 10042 6984 10048 6996
rect 7524 6956 10048 6984
rect 7524 6944 7530 6956
rect 10042 6944 10048 6956
rect 10100 6984 10106 6996
rect 10962 6984 10968 6996
rect 10100 6956 10968 6984
rect 10100 6944 10106 6956
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 15102 6944 15108 6996
rect 15160 6984 15166 6996
rect 15838 6984 15844 6996
rect 15160 6956 15844 6984
rect 15160 6944 15166 6956
rect 15838 6944 15844 6956
rect 15896 6984 15902 6996
rect 15933 6987 15991 6993
rect 15933 6984 15945 6987
rect 15896 6956 15945 6984
rect 15896 6944 15902 6956
rect 15933 6953 15945 6956
rect 15979 6953 15991 6987
rect 16114 6984 16120 6996
rect 16075 6956 16120 6984
rect 15933 6947 15991 6953
rect 16114 6944 16120 6956
rect 16172 6944 16178 6996
rect 17607 6987 17665 6993
rect 17607 6953 17619 6987
rect 17653 6984 17665 6987
rect 18325 6987 18383 6993
rect 18325 6984 18337 6987
rect 17653 6956 18337 6984
rect 17653 6953 17665 6956
rect 17607 6947 17665 6953
rect 18325 6953 18337 6956
rect 18371 6953 18383 6987
rect 18325 6947 18383 6953
rect 2314 6876 2320 6928
rect 2372 6916 2378 6928
rect 3973 6919 4031 6925
rect 3973 6916 3985 6919
rect 2372 6888 3985 6916
rect 2372 6876 2378 6888
rect 3973 6885 3985 6888
rect 4019 6885 4031 6919
rect 3973 6879 4031 6885
rect 4246 6876 4252 6928
rect 4304 6916 4310 6928
rect 4304 6888 4660 6916
rect 4304 6876 4310 6888
rect 3421 6851 3479 6857
rect 3421 6848 3433 6851
rect 2700 6820 3433 6848
rect 2700 6789 2728 6820
rect 3421 6817 3433 6820
rect 3467 6848 3479 6851
rect 4062 6848 4068 6860
rect 3467 6820 4068 6848
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 4062 6808 4068 6820
rect 4120 6848 4126 6860
rect 4632 6857 4660 6888
rect 5258 6876 5264 6928
rect 5316 6916 5322 6928
rect 5810 6916 5816 6928
rect 5316 6888 5816 6916
rect 5316 6876 5322 6888
rect 5810 6876 5816 6888
rect 5868 6916 5874 6928
rect 8110 6916 8116 6928
rect 5868 6888 8116 6916
rect 5868 6876 5874 6888
rect 4617 6851 4675 6857
rect 4120 6820 4292 6848
rect 4120 6808 4126 6820
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6749 2743 6783
rect 2866 6780 2872 6792
rect 2827 6752 2872 6780
rect 2685 6743 2743 6749
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 2958 6740 2964 6792
rect 3016 6780 3022 6792
rect 4264 6789 4292 6820
rect 4617 6817 4629 6851
rect 4663 6848 4675 6851
rect 5350 6848 5356 6860
rect 4663 6820 5356 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 3016 6752 3065 6780
rect 3016 6740 3022 6752
rect 3053 6749 3065 6752
rect 3099 6780 3111 6783
rect 3145 6783 3203 6789
rect 3145 6780 3157 6783
rect 3099 6752 3157 6780
rect 3099 6749 3111 6752
rect 3053 6743 3111 6749
rect 3145 6749 3157 6752
rect 3191 6749 3203 6783
rect 3145 6743 3203 6749
rect 3329 6783 3387 6789
rect 3329 6749 3341 6783
rect 3375 6749 3387 6783
rect 3329 6743 3387 6749
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6780 4859 6783
rect 4890 6780 4896 6792
rect 4847 6752 4896 6780
rect 4847 6749 4859 6752
rect 4801 6743 4859 6749
rect 566 6672 572 6724
rect 624 6712 630 6724
rect 624 6684 2544 6712
rect 624 6672 630 6684
rect 2516 6653 2544 6684
rect 2774 6672 2780 6724
rect 2832 6712 2838 6724
rect 3344 6712 3372 6743
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 5074 6780 5080 6792
rect 5035 6752 5080 6780
rect 5074 6740 5080 6752
rect 5132 6740 5138 6792
rect 5626 6780 5632 6792
rect 5587 6752 5632 6780
rect 5626 6740 5632 6752
rect 5684 6740 5690 6792
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 6472 6780 6500 6888
rect 8110 6876 8116 6888
rect 8168 6876 8174 6928
rect 9030 6876 9036 6928
rect 9088 6916 9094 6928
rect 9088 6888 11468 6916
rect 9088 6876 9094 6888
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 7374 6848 7380 6860
rect 6595 6820 7380 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 7561 6851 7619 6857
rect 7561 6848 7573 6851
rect 7524 6820 7573 6848
rect 7524 6808 7530 6820
rect 7561 6817 7573 6820
rect 7607 6848 7619 6851
rect 8018 6848 8024 6860
rect 7607 6820 8024 6848
rect 7607 6817 7619 6820
rect 7561 6811 7619 6817
rect 8018 6808 8024 6820
rect 8076 6808 8082 6860
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6817 8263 6851
rect 8205 6811 8263 6817
rect 6641 6783 6699 6789
rect 6641 6780 6653 6783
rect 5776 6752 5821 6780
rect 6472 6752 6653 6780
rect 5776 6740 5782 6752
rect 6641 6749 6653 6752
rect 6687 6749 6699 6783
rect 7650 6780 7656 6792
rect 6641 6743 6699 6749
rect 7208 6752 7656 6780
rect 2832 6684 2877 6712
rect 3068 6684 3372 6712
rect 5905 6715 5963 6721
rect 2832 6672 2838 6684
rect 2501 6647 2559 6653
rect 2501 6613 2513 6647
rect 2547 6613 2559 6647
rect 2501 6607 2559 6613
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 3068 6644 3096 6684
rect 5905 6681 5917 6715
rect 5951 6712 5963 6715
rect 7208 6712 7236 6752
rect 7650 6740 7656 6752
rect 7708 6780 7714 6792
rect 8113 6783 8171 6789
rect 8113 6780 8125 6783
rect 7708 6752 8125 6780
rect 7708 6740 7714 6752
rect 8113 6749 8125 6752
rect 8159 6749 8171 6783
rect 8220 6780 8248 6811
rect 8386 6808 8392 6860
rect 8444 6848 8450 6860
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 8444 6820 8493 6848
rect 8444 6808 8450 6820
rect 8481 6817 8493 6820
rect 8527 6817 8539 6851
rect 10502 6848 10508 6860
rect 8481 6811 8539 6817
rect 8588 6820 10508 6848
rect 8588 6780 8616 6820
rect 10502 6808 10508 6820
rect 10560 6808 10566 6860
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 10870 6848 10876 6860
rect 10744 6820 10876 6848
rect 10744 6808 10750 6820
rect 10870 6808 10876 6820
rect 10928 6808 10934 6860
rect 11440 6857 11468 6888
rect 13740 6888 13952 6916
rect 11425 6851 11483 6857
rect 11425 6817 11437 6851
rect 11471 6848 11483 6851
rect 11701 6851 11759 6857
rect 11701 6848 11713 6851
rect 11471 6820 11713 6848
rect 11471 6817 11483 6820
rect 11425 6811 11483 6817
rect 11701 6817 11713 6820
rect 11747 6817 11759 6851
rect 13740 6848 13768 6888
rect 11701 6811 11759 6817
rect 12406 6820 13768 6848
rect 13817 6851 13875 6857
rect 10226 6780 10232 6792
rect 8220 6752 8616 6780
rect 10187 6752 10232 6780
rect 8113 6743 8171 6749
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 10410 6740 10416 6792
rect 10468 6780 10474 6792
rect 10597 6783 10655 6789
rect 10597 6780 10609 6783
rect 10468 6752 10609 6780
rect 10468 6740 10474 6752
rect 10597 6749 10609 6752
rect 10643 6780 10655 6783
rect 11054 6780 11060 6792
rect 10643 6752 11060 6780
rect 10643 6749 10655 6752
rect 10597 6743 10655 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11790 6780 11796 6792
rect 11751 6752 11796 6780
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 5951 6684 7236 6712
rect 7285 6715 7343 6721
rect 5951 6681 5963 6684
rect 5905 6675 5963 6681
rect 7285 6681 7297 6715
rect 7331 6712 7343 6715
rect 8478 6712 8484 6724
rect 7331 6684 8484 6712
rect 7331 6681 7343 6684
rect 7285 6675 7343 6681
rect 8478 6672 8484 6684
rect 8536 6672 8542 6724
rect 9674 6672 9680 6724
rect 9732 6712 9738 6724
rect 10321 6715 10379 6721
rect 10321 6712 10333 6715
rect 9732 6684 10333 6712
rect 9732 6672 9738 6684
rect 10321 6681 10333 6684
rect 10367 6681 10379 6715
rect 10321 6675 10379 6681
rect 10505 6715 10563 6721
rect 10505 6681 10517 6715
rect 10551 6712 10563 6715
rect 10778 6712 10784 6724
rect 10551 6684 10784 6712
rect 10551 6681 10563 6684
rect 10505 6675 10563 6681
rect 10778 6672 10784 6684
rect 10836 6672 10842 6724
rect 10962 6672 10968 6724
rect 11020 6712 11026 6724
rect 11333 6715 11391 6721
rect 11333 6712 11345 6715
rect 11020 6684 11345 6712
rect 11020 6672 11026 6684
rect 11333 6681 11345 6684
rect 11379 6712 11391 6715
rect 12406 6712 12434 6820
rect 13817 6817 13829 6851
rect 13863 6817 13875 6851
rect 13924 6848 13952 6888
rect 14458 6848 14464 6860
rect 13924 6820 14464 6848
rect 13817 6811 13875 6817
rect 12713 6783 12771 6789
rect 12713 6749 12725 6783
rect 12759 6780 12771 6783
rect 12759 6752 13308 6780
rect 12759 6749 12771 6752
rect 12713 6743 12771 6749
rect 11379 6684 12434 6712
rect 11379 6681 11391 6684
rect 11333 6675 11391 6681
rect 2648 6616 3096 6644
rect 5813 6647 5871 6653
rect 2648 6604 2654 6616
rect 5813 6613 5825 6647
rect 5859 6644 5871 6647
rect 6181 6647 6239 6653
rect 6181 6644 6193 6647
rect 5859 6616 6193 6644
rect 5859 6613 5871 6616
rect 5813 6607 5871 6613
rect 6181 6613 6193 6616
rect 6227 6613 6239 6647
rect 6822 6644 6828 6656
rect 6783 6616 6828 6644
rect 6181 6607 6239 6613
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7190 6604 7196 6656
rect 7248 6644 7254 6656
rect 7377 6647 7435 6653
rect 7377 6644 7389 6647
rect 7248 6616 7389 6644
rect 7248 6604 7254 6616
rect 7377 6613 7389 6616
rect 7423 6613 7435 6647
rect 7377 6607 7435 6613
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 7745 6647 7803 6653
rect 7745 6644 7757 6647
rect 7524 6616 7757 6644
rect 7524 6604 7530 6616
rect 7745 6613 7757 6616
rect 7791 6613 7803 6647
rect 10410 6644 10416 6656
rect 10371 6616 10416 6644
rect 7745 6607 7803 6613
rect 10410 6604 10416 6616
rect 10468 6604 10474 6656
rect 10594 6604 10600 6656
rect 10652 6644 10658 6656
rect 10873 6647 10931 6653
rect 10873 6644 10885 6647
rect 10652 6616 10885 6644
rect 10652 6604 10658 6616
rect 10873 6613 10885 6616
rect 10919 6613 10931 6647
rect 11238 6644 11244 6656
rect 11199 6616 11244 6644
rect 10873 6607 10931 6613
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 12342 6604 12348 6656
rect 12400 6644 12406 6656
rect 13280 6653 13308 6752
rect 13538 6740 13544 6792
rect 13596 6780 13602 6792
rect 13832 6780 13860 6811
rect 14458 6808 14464 6820
rect 14516 6848 14522 6860
rect 14645 6851 14703 6857
rect 14516 6820 14596 6848
rect 14516 6808 14522 6820
rect 14366 6780 14372 6792
rect 13596 6752 13860 6780
rect 14327 6752 14372 6780
rect 13596 6740 13602 6752
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 14568 6780 14596 6820
rect 14645 6817 14657 6851
rect 14691 6848 14703 6851
rect 15381 6851 15439 6857
rect 15381 6848 15393 6851
rect 14691 6820 15393 6848
rect 14691 6817 14703 6820
rect 14645 6811 14703 6817
rect 15381 6817 15393 6820
rect 15427 6848 15439 6851
rect 18322 6848 18328 6860
rect 15427 6820 18328 6848
rect 15427 6817 15439 6820
rect 15381 6811 15439 6817
rect 18322 6808 18328 6820
rect 18380 6808 18386 6860
rect 15105 6783 15163 6789
rect 15105 6780 15117 6783
rect 14568 6752 15117 6780
rect 15105 6749 15117 6752
rect 15151 6749 15163 6783
rect 15105 6743 15163 6749
rect 17862 6740 17868 6792
rect 17920 6780 17926 6792
rect 18233 6783 18291 6789
rect 17920 6752 17965 6780
rect 17920 6740 17926 6752
rect 18233 6749 18245 6783
rect 18279 6780 18291 6783
rect 18506 6780 18512 6792
rect 18279 6752 18512 6780
rect 18279 6749 18291 6752
rect 18233 6743 18291 6749
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 13633 6715 13691 6721
rect 13633 6681 13645 6715
rect 13679 6712 13691 6715
rect 13679 6684 14780 6712
rect 13679 6681 13691 6684
rect 13633 6675 13691 6681
rect 12529 6647 12587 6653
rect 12529 6644 12541 6647
rect 12400 6616 12541 6644
rect 12400 6604 12406 6616
rect 12529 6613 12541 6616
rect 12575 6613 12587 6647
rect 12529 6607 12587 6613
rect 13265 6647 13323 6653
rect 13265 6613 13277 6647
rect 13311 6613 13323 6647
rect 13722 6644 13728 6656
rect 13683 6616 13728 6644
rect 13265 6607 13323 6613
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 14752 6653 14780 6684
rect 15838 6672 15844 6724
rect 15896 6712 15902 6724
rect 15896 6684 16422 6712
rect 15896 6672 15902 6684
rect 14737 6647 14795 6653
rect 14737 6613 14749 6647
rect 14783 6613 14795 6647
rect 14737 6607 14795 6613
rect 15194 6604 15200 6656
rect 15252 6644 15258 6656
rect 15252 6616 15297 6644
rect 15252 6604 15258 6616
rect 0 6554 18860 6576
rect 0 6502 4660 6554
rect 4712 6502 4724 6554
rect 4776 6502 4788 6554
rect 4840 6502 4852 6554
rect 4904 6502 4916 6554
rect 4968 6502 7760 6554
rect 7812 6502 7824 6554
rect 7876 6502 7888 6554
rect 7940 6502 7952 6554
rect 8004 6502 8016 6554
rect 8068 6502 10860 6554
rect 10912 6502 10924 6554
rect 10976 6502 10988 6554
rect 11040 6502 11052 6554
rect 11104 6502 11116 6554
rect 11168 6502 13960 6554
rect 14012 6502 14024 6554
rect 14076 6502 14088 6554
rect 14140 6502 14152 6554
rect 14204 6502 14216 6554
rect 14268 6502 17060 6554
rect 17112 6502 17124 6554
rect 17176 6502 17188 6554
rect 17240 6502 17252 6554
rect 17304 6502 17316 6554
rect 17368 6502 18860 6554
rect 0 6480 18860 6502
rect 1946 6440 1952 6452
rect 1780 6412 1952 6440
rect 1780 6358 1808 6412
rect 1946 6400 1952 6412
rect 2004 6440 2010 6452
rect 2133 6443 2191 6449
rect 2133 6440 2145 6443
rect 2004 6412 2145 6440
rect 2004 6400 2010 6412
rect 2133 6409 2145 6412
rect 2179 6440 2191 6443
rect 2498 6440 2504 6452
rect 2179 6412 2504 6440
rect 2179 6409 2191 6412
rect 2133 6403 2191 6409
rect 2498 6400 2504 6412
rect 2556 6400 2562 6452
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 2869 6443 2927 6449
rect 2869 6440 2881 6443
rect 2832 6412 2881 6440
rect 2832 6400 2838 6412
rect 2869 6409 2881 6412
rect 2915 6409 2927 6443
rect 2869 6403 2927 6409
rect 2958 6400 2964 6452
rect 3016 6440 3022 6452
rect 3694 6440 3700 6452
rect 3016 6412 3700 6440
rect 3016 6400 3022 6412
rect 3694 6400 3700 6412
rect 3752 6400 3758 6452
rect 5258 6440 5264 6452
rect 5219 6412 5264 6440
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 5718 6400 5724 6452
rect 5776 6400 5782 6452
rect 5902 6440 5908 6452
rect 5863 6412 5908 6440
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 6638 6440 6644 6452
rect 6599 6412 6644 6440
rect 6638 6400 6644 6412
rect 6696 6400 6702 6452
rect 6733 6443 6791 6449
rect 6733 6409 6745 6443
rect 6779 6440 6791 6443
rect 7466 6440 7472 6452
rect 6779 6412 7472 6440
rect 6779 6409 6791 6412
rect 6733 6403 6791 6409
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 10226 6440 10232 6452
rect 7576 6412 10232 6440
rect 3510 6372 3516 6384
rect 3252 6344 3516 6372
rect 2590 6304 2596 6316
rect 2551 6276 2596 6304
rect 2590 6264 2596 6276
rect 2648 6264 2654 6316
rect 3252 6313 3280 6344
rect 3510 6332 3516 6344
rect 3568 6372 3574 6384
rect 5736 6372 5764 6400
rect 5813 6375 5871 6381
rect 5813 6372 5825 6375
rect 3568 6344 4200 6372
rect 5736 6344 5825 6372
rect 3568 6332 3574 6344
rect 2777 6307 2835 6313
rect 2777 6304 2789 6307
rect 2700 6276 2789 6304
rect 290 6236 296 6248
rect 251 6208 296 6236
rect 290 6196 296 6208
rect 348 6196 354 6248
rect 566 6236 572 6248
rect 527 6208 572 6236
rect 566 6196 572 6208
rect 624 6196 630 6248
rect 2041 6239 2099 6245
rect 2041 6205 2053 6239
rect 2087 6236 2099 6239
rect 2700 6236 2728 6276
rect 2777 6273 2789 6276
rect 2823 6273 2835 6307
rect 2777 6267 2835 6273
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6273 3295 6307
rect 3418 6304 3424 6316
rect 3379 6276 3424 6304
rect 3237 6267 3295 6273
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 4172 6313 4200 6344
rect 5813 6341 5825 6344
rect 5859 6341 5871 6375
rect 6546 6372 6552 6384
rect 5813 6335 5871 6341
rect 6472 6344 6552 6372
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6273 3663 6307
rect 3605 6267 3663 6273
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4203 6276 4936 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 2958 6236 2964 6248
rect 2087 6208 2964 6236
rect 2087 6205 2099 6208
rect 2041 6199 2099 6205
rect 2958 6196 2964 6208
rect 3016 6236 3022 6248
rect 3053 6239 3111 6245
rect 3053 6236 3065 6239
rect 3016 6208 3065 6236
rect 3016 6196 3022 6208
rect 3053 6205 3065 6208
rect 3099 6205 3111 6239
rect 3053 6199 3111 6205
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 3436 6236 3464 6264
rect 3191 6208 3464 6236
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 2777 6171 2835 6177
rect 2777 6137 2789 6171
rect 2823 6168 2835 6171
rect 3620 6168 3648 6267
rect 4908 6177 4936 6276
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 5721 6307 5779 6313
rect 5721 6304 5733 6307
rect 5684 6276 5733 6304
rect 5684 6264 5690 6276
rect 5721 6273 5733 6276
rect 5767 6273 5779 6307
rect 5994 6304 6000 6316
rect 5955 6276 6000 6304
rect 5721 6267 5779 6273
rect 5166 6196 5172 6248
rect 5224 6236 5230 6248
rect 5353 6239 5411 6245
rect 5353 6236 5365 6239
rect 5224 6208 5365 6236
rect 5224 6196 5230 6208
rect 5353 6205 5365 6208
rect 5399 6205 5411 6239
rect 5353 6199 5411 6205
rect 2823 6140 3648 6168
rect 4893 6171 4951 6177
rect 2823 6137 2835 6140
rect 2777 6131 2835 6137
rect 4893 6137 4905 6171
rect 4939 6137 4951 6171
rect 5368 6168 5396 6199
rect 5442 6196 5448 6248
rect 5500 6236 5506 6248
rect 5736 6236 5764 6267
rect 5994 6264 6000 6276
rect 6052 6264 6058 6316
rect 6472 6236 6500 6344
rect 6546 6332 6552 6344
rect 6604 6372 6610 6384
rect 7576 6372 7604 6412
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 10321 6443 10379 6449
rect 10321 6409 10333 6443
rect 10367 6440 10379 6443
rect 10594 6440 10600 6452
rect 10367 6412 10600 6440
rect 10367 6409 10379 6412
rect 10321 6403 10379 6409
rect 10594 6400 10600 6412
rect 10652 6400 10658 6452
rect 11882 6440 11888 6452
rect 11843 6412 11888 6440
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 13814 6440 13820 6452
rect 12084 6412 13820 6440
rect 6604 6344 7604 6372
rect 9493 6375 9551 6381
rect 6604 6332 6610 6344
rect 9493 6341 9505 6375
rect 9539 6372 9551 6375
rect 9766 6372 9772 6384
rect 9539 6344 9772 6372
rect 9539 6341 9551 6344
rect 9493 6335 9551 6341
rect 9766 6332 9772 6344
rect 9824 6332 9830 6384
rect 10410 6332 10416 6384
rect 10468 6372 10474 6384
rect 11425 6375 11483 6381
rect 11425 6372 11437 6375
rect 10468 6344 11437 6372
rect 10468 6332 10474 6344
rect 11425 6341 11437 6344
rect 11471 6341 11483 6375
rect 11425 6335 11483 6341
rect 9030 6304 9036 6316
rect 6564 6276 9036 6304
rect 6564 6245 6592 6276
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9674 6304 9680 6316
rect 9635 6276 9680 6304
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 9861 6307 9919 6313
rect 9861 6273 9873 6307
rect 9907 6304 9919 6307
rect 10594 6304 10600 6316
rect 9907 6276 10600 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 5500 6208 5545 6236
rect 5736 6208 6500 6236
rect 6549 6239 6607 6245
rect 5500 6196 5506 6208
rect 6549 6205 6561 6239
rect 6595 6205 6607 6239
rect 7374 6236 7380 6248
rect 6549 6199 6607 6205
rect 6656 6208 7380 6236
rect 6656 6168 6684 6208
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7650 6196 7656 6248
rect 7708 6236 7714 6248
rect 9876 6236 9904 6267
rect 10594 6264 10600 6276
rect 10652 6264 10658 6316
rect 10686 6264 10692 6316
rect 10744 6304 10750 6316
rect 12084 6313 12112 6412
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 14366 6400 14372 6452
rect 14424 6440 14430 6452
rect 14553 6443 14611 6449
rect 14553 6440 14565 6443
rect 14424 6412 14565 6440
rect 14424 6400 14430 6412
rect 14553 6409 14565 6412
rect 14599 6409 14611 6443
rect 14553 6403 14611 6409
rect 15194 6400 15200 6452
rect 15252 6440 15258 6452
rect 15381 6443 15439 6449
rect 15381 6440 15393 6443
rect 15252 6412 15393 6440
rect 15252 6400 15258 6412
rect 15381 6409 15393 6412
rect 15427 6409 15439 6443
rect 15381 6403 15439 6409
rect 16853 6443 16911 6449
rect 16853 6409 16865 6443
rect 16899 6409 16911 6443
rect 16853 6403 16911 6409
rect 17221 6443 17279 6449
rect 17221 6409 17233 6443
rect 17267 6440 17279 6443
rect 17681 6443 17739 6449
rect 17681 6440 17693 6443
rect 17267 6412 17693 6440
rect 17267 6409 17279 6412
rect 17221 6403 17279 6409
rect 17681 6409 17693 6412
rect 17727 6409 17739 6443
rect 18046 6440 18052 6452
rect 18007 6412 18052 6440
rect 17681 6403 17739 6409
rect 12342 6372 12348 6384
rect 12303 6344 12348 6372
rect 12342 6332 12348 6344
rect 12400 6332 12406 6384
rect 13722 6332 13728 6384
rect 13780 6372 13786 6384
rect 14001 6375 14059 6381
rect 14001 6372 14013 6375
rect 13780 6344 14013 6372
rect 13780 6332 13786 6344
rect 14001 6341 14013 6344
rect 14047 6372 14059 6375
rect 14047 6344 15792 6372
rect 14047 6341 14059 6344
rect 14001 6335 14059 6341
rect 12069 6307 12127 6313
rect 12069 6304 12081 6307
rect 10744 6276 12081 6304
rect 10744 6264 10750 6276
rect 12069 6273 12081 6276
rect 12115 6273 12127 6307
rect 12069 6267 12127 6273
rect 10134 6236 10140 6248
rect 7708 6208 9904 6236
rect 10095 6208 10140 6236
rect 7708 6196 7714 6208
rect 10134 6196 10140 6208
rect 10192 6196 10198 6248
rect 10229 6239 10287 6245
rect 10229 6205 10241 6239
rect 10275 6205 10287 6239
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 10229 6199 10287 6205
rect 10336 6208 10977 6236
rect 7098 6168 7104 6180
rect 5368 6140 6684 6168
rect 7059 6140 7104 6168
rect 4893 6131 4951 6137
rect 7098 6128 7104 6140
rect 7156 6128 7162 6180
rect 8110 6128 8116 6180
rect 8168 6168 8174 6180
rect 9858 6168 9864 6180
rect 8168 6140 9260 6168
rect 9819 6140 9864 6168
rect 8168 6128 8174 6140
rect 2866 6060 2872 6112
rect 2924 6100 2930 6112
rect 3881 6103 3939 6109
rect 3881 6100 3893 6103
rect 2924 6072 3893 6100
rect 2924 6060 2930 6072
rect 3881 6069 3893 6072
rect 3927 6100 3939 6103
rect 4065 6103 4123 6109
rect 4065 6100 4077 6103
rect 3927 6072 4077 6100
rect 3927 6069 3939 6072
rect 3881 6063 3939 6069
rect 4065 6069 4077 6072
rect 4111 6069 4123 6103
rect 4065 6063 4123 6069
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6100 8263 6103
rect 9122 6100 9128 6112
rect 8251 6072 9128 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9232 6100 9260 6140
rect 9858 6128 9864 6140
rect 9916 6128 9922 6180
rect 10042 6128 10048 6180
rect 10100 6168 10106 6180
rect 10244 6168 10272 6199
rect 10100 6140 10272 6168
rect 10100 6128 10106 6140
rect 10336 6100 10364 6208
rect 10965 6205 10977 6208
rect 11011 6205 11023 6239
rect 10965 6199 11023 6205
rect 11057 6239 11115 6245
rect 11057 6205 11069 6239
rect 11103 6205 11115 6239
rect 11057 6199 11115 6205
rect 10689 6171 10747 6177
rect 10689 6137 10701 6171
rect 10735 6168 10747 6171
rect 11072 6168 11100 6199
rect 11882 6196 11888 6248
rect 11940 6236 11946 6248
rect 13464 6236 13492 6290
rect 11940 6208 13492 6236
rect 13817 6239 13875 6245
rect 11940 6196 11946 6208
rect 13817 6205 13829 6239
rect 13863 6236 13875 6239
rect 14016 6236 14044 6335
rect 14568 6313 14596 6344
rect 15764 6313 15792 6344
rect 14277 6307 14335 6313
rect 14277 6273 14289 6307
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 14553 6307 14611 6313
rect 14553 6273 14565 6307
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 14737 6307 14795 6313
rect 14737 6273 14749 6307
rect 14783 6273 14795 6307
rect 14737 6267 14795 6273
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6273 15347 6307
rect 15289 6267 15347 6273
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6273 15807 6307
rect 15749 6267 15807 6273
rect 16669 6307 16727 6313
rect 16669 6273 16681 6307
rect 16715 6304 16727 6307
rect 16868 6304 16896 6403
rect 18046 6400 18052 6412
rect 18104 6400 18110 6452
rect 16715 6276 16896 6304
rect 16715 6273 16727 6276
rect 16669 6267 16727 6273
rect 13863 6208 14044 6236
rect 13863 6205 13875 6208
rect 13817 6199 13875 6205
rect 10735 6140 11100 6168
rect 10735 6137 10747 6140
rect 10689 6131 10747 6137
rect 13538 6128 13544 6180
rect 13596 6168 13602 6180
rect 14185 6171 14243 6177
rect 14185 6168 14197 6171
rect 13596 6140 14197 6168
rect 13596 6128 13602 6140
rect 14185 6137 14197 6140
rect 14231 6137 14243 6171
rect 14292 6168 14320 6267
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 14752 6236 14780 6267
rect 14424 6208 14780 6236
rect 15304 6236 15332 6267
rect 15657 6239 15715 6245
rect 15657 6236 15669 6239
rect 15304 6208 15669 6236
rect 14424 6196 14430 6208
rect 15304 6168 15332 6208
rect 15657 6205 15669 6208
rect 15703 6236 15715 6239
rect 17310 6236 17316 6248
rect 15703 6208 17316 6236
rect 15703 6205 15715 6208
rect 15657 6199 15715 6205
rect 17310 6196 17316 6208
rect 17368 6196 17374 6248
rect 17494 6236 17500 6248
rect 17455 6208 17500 6236
rect 17494 6196 17500 6208
rect 17552 6196 17558 6248
rect 18138 6236 18144 6248
rect 18099 6208 18144 6236
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 18322 6236 18328 6248
rect 18283 6208 18328 6236
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 17512 6168 17540 6196
rect 14292 6140 15332 6168
rect 15396 6140 17540 6168
rect 14185 6131 14243 6137
rect 9232 6072 10364 6100
rect 10410 6060 10416 6112
rect 10468 6100 10474 6112
rect 10781 6103 10839 6109
rect 10781 6100 10793 6103
rect 10468 6072 10793 6100
rect 10468 6060 10474 6072
rect 10781 6069 10793 6072
rect 10827 6069 10839 6103
rect 14090 6100 14096 6112
rect 14051 6072 14096 6100
rect 10781 6063 10839 6069
rect 14090 6060 14096 6072
rect 14148 6060 14154 6112
rect 14200 6100 14228 6131
rect 15396 6100 15424 6140
rect 14200 6072 15424 6100
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 16485 6103 16543 6109
rect 16485 6100 16497 6103
rect 16448 6072 16497 6100
rect 16448 6060 16454 6072
rect 16485 6069 16497 6072
rect 16531 6069 16543 6103
rect 16485 6063 16543 6069
rect 0 6010 18860 6032
rect 0 5958 3110 6010
rect 3162 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 6210 6010
rect 6262 5958 6274 6010
rect 6326 5958 6338 6010
rect 6390 5958 6402 6010
rect 6454 5958 6466 6010
rect 6518 5958 9310 6010
rect 9362 5958 9374 6010
rect 9426 5958 9438 6010
rect 9490 5958 9502 6010
rect 9554 5958 9566 6010
rect 9618 5958 12410 6010
rect 12462 5958 12474 6010
rect 12526 5958 12538 6010
rect 12590 5958 12602 6010
rect 12654 5958 12666 6010
rect 12718 5958 15510 6010
rect 15562 5958 15574 6010
rect 15626 5958 15638 6010
rect 15690 5958 15702 6010
rect 15754 5958 15766 6010
rect 15818 5958 18860 6010
rect 0 5936 18860 5958
rect 566 5856 572 5908
rect 624 5896 630 5908
rect 2409 5899 2467 5905
rect 2409 5896 2421 5899
rect 624 5868 2421 5896
rect 624 5856 630 5868
rect 2409 5865 2421 5868
rect 2455 5865 2467 5899
rect 2409 5859 2467 5865
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 3881 5899 3939 5905
rect 3881 5896 3893 5899
rect 3559 5868 3893 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 3881 5865 3893 5868
rect 3927 5865 3939 5899
rect 3881 5859 3939 5865
rect 4328 5899 4386 5905
rect 4328 5865 4340 5899
rect 4374 5896 4386 5899
rect 5534 5896 5540 5908
rect 4374 5868 5540 5896
rect 4374 5865 4386 5868
rect 4328 5859 4386 5865
rect 5534 5856 5540 5868
rect 5592 5856 5598 5908
rect 5813 5899 5871 5905
rect 5813 5865 5825 5899
rect 5859 5896 5871 5899
rect 5994 5896 6000 5908
rect 5859 5868 6000 5896
rect 5859 5865 5871 5868
rect 5813 5859 5871 5865
rect 5994 5856 6000 5868
rect 6052 5896 6058 5908
rect 6052 5868 7236 5896
rect 6052 5856 6058 5868
rect 3418 5828 3424 5840
rect 3379 5800 3424 5828
rect 3418 5788 3424 5800
rect 3476 5788 3482 5840
rect 3620 5800 4108 5828
rect 290 5720 296 5772
rect 348 5760 354 5772
rect 3620 5760 3648 5800
rect 348 5732 3648 5760
rect 348 5720 354 5732
rect 952 5701 980 5732
rect 3694 5720 3700 5772
rect 3752 5760 3758 5772
rect 4080 5769 4108 5800
rect 4065 5763 4123 5769
rect 3752 5732 3797 5760
rect 3752 5720 3758 5732
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 6086 5760 6092 5772
rect 4111 5732 6092 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5760 6515 5763
rect 6822 5760 6828 5772
rect 6503 5732 6828 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 7208 5760 7236 5868
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 7883 5899 7941 5905
rect 7883 5896 7895 5899
rect 7708 5868 7895 5896
rect 7708 5856 7714 5868
rect 7883 5865 7895 5868
rect 7929 5865 7941 5899
rect 7883 5859 7941 5865
rect 8205 5899 8263 5905
rect 8205 5865 8217 5899
rect 8251 5896 8263 5899
rect 8846 5896 8852 5908
rect 8251 5868 8852 5896
rect 8251 5865 8263 5868
rect 8205 5859 8263 5865
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 8941 5899 8999 5905
rect 8941 5865 8953 5899
rect 8987 5896 8999 5899
rect 9674 5896 9680 5908
rect 8987 5868 9680 5896
rect 8987 5865 8999 5868
rect 8941 5859 8999 5865
rect 9674 5856 9680 5868
rect 9732 5896 9738 5908
rect 9732 5868 10824 5896
rect 9732 5856 9738 5868
rect 10042 5760 10048 5772
rect 7208 5732 10048 5760
rect 937 5695 995 5701
rect 937 5661 949 5695
rect 983 5661 995 5695
rect 937 5655 995 5661
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2774 5692 2780 5704
rect 2639 5664 2780 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5692 2927 5695
rect 2958 5692 2964 5704
rect 2915 5664 2964 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 2958 5652 2964 5664
rect 3016 5692 3022 5704
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 3016 5664 3065 5692
rect 3016 5652 3022 5664
rect 3053 5661 3065 5664
rect 3099 5661 3111 5695
rect 3970 5692 3976 5704
rect 3931 5664 3976 5692
rect 3053 5655 3111 5661
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 5442 5652 5448 5704
rect 5500 5652 5506 5704
rect 8220 5701 8248 5732
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 10410 5760 10416 5772
rect 10371 5732 10416 5760
rect 10410 5720 10416 5732
rect 10468 5720 10474 5772
rect 10686 5760 10692 5772
rect 10647 5732 10692 5760
rect 10686 5720 10692 5732
rect 10744 5720 10750 5772
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5661 8263 5695
rect 10796 5692 10824 5868
rect 11238 5856 11244 5908
rect 11296 5896 11302 5908
rect 11425 5899 11483 5905
rect 11425 5896 11437 5899
rect 11296 5868 11437 5896
rect 11296 5856 11302 5868
rect 11425 5865 11437 5868
rect 11471 5865 11483 5899
rect 15838 5896 15844 5908
rect 15799 5868 15844 5896
rect 11425 5859 11483 5865
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 17310 5856 17316 5908
rect 17368 5896 17374 5908
rect 17819 5899 17877 5905
rect 17819 5896 17831 5899
rect 17368 5868 17831 5896
rect 17368 5856 17374 5868
rect 17819 5865 17831 5868
rect 17865 5896 17877 5899
rect 17865 5868 18092 5896
rect 17865 5865 17877 5868
rect 17819 5859 17877 5865
rect 11149 5763 11207 5769
rect 11149 5729 11161 5763
rect 11195 5760 11207 5763
rect 11238 5760 11244 5772
rect 11195 5732 11244 5760
rect 11195 5729 11207 5732
rect 11149 5723 11207 5729
rect 11238 5720 11244 5732
rect 11296 5720 11302 5772
rect 14090 5720 14096 5772
rect 14148 5760 14154 5772
rect 14277 5763 14335 5769
rect 14277 5760 14289 5763
rect 14148 5732 14289 5760
rect 14148 5720 14154 5732
rect 14277 5729 14289 5732
rect 14323 5729 14335 5763
rect 14734 5760 14740 5772
rect 14695 5732 14740 5760
rect 14277 5723 14335 5729
rect 14734 5720 14740 5732
rect 14792 5720 14798 5772
rect 16390 5760 16396 5772
rect 16351 5732 16396 5760
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 11057 5695 11115 5701
rect 11057 5692 11069 5695
rect 10796 5664 11069 5692
rect 8205 5655 8263 5661
rect 11057 5661 11069 5664
rect 11103 5661 11115 5695
rect 14366 5692 14372 5704
rect 14327 5664 14372 5692
rect 11057 5655 11115 5661
rect 14366 5652 14372 5664
rect 14424 5652 14430 5704
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5692 16083 5695
rect 16298 5692 16304 5704
rect 16071 5664 16304 5692
rect 16071 5661 16083 5664
rect 16025 5655 16083 5661
rect 566 5624 572 5636
rect 527 5596 572 5624
rect 566 5584 572 5596
rect 624 5584 630 5636
rect 7006 5584 7012 5636
rect 7064 5584 7070 5636
rect 11882 5624 11888 5636
rect 9982 5596 11888 5624
rect 11882 5584 11888 5596
rect 11940 5584 11946 5636
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 15010 5624 15016 5636
rect 13872 5596 15016 5624
rect 13872 5584 13878 5596
rect 15010 5584 15016 5596
rect 15068 5624 15074 5636
rect 16040 5624 16068 5655
rect 16298 5652 16304 5664
rect 16356 5652 16362 5704
rect 18064 5701 18092 5868
rect 18138 5856 18144 5908
rect 18196 5896 18202 5908
rect 18233 5899 18291 5905
rect 18233 5896 18245 5899
rect 18196 5868 18245 5896
rect 18196 5856 18202 5868
rect 18233 5865 18245 5868
rect 18279 5865 18291 5899
rect 18233 5859 18291 5865
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5661 18107 5695
rect 18049 5655 18107 5661
rect 15068 5596 16068 5624
rect 15068 5584 15074 5596
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5556 2835 5559
rect 2866 5556 2872 5568
rect 2823 5528 2872 5556
rect 2823 5525 2835 5528
rect 2777 5519 2835 5525
rect 2866 5516 2872 5528
rect 2924 5516 2930 5568
rect 3694 5556 3700 5568
rect 3655 5528 3700 5556
rect 3694 5516 3700 5528
rect 3752 5516 3758 5568
rect 8110 5516 8116 5568
rect 8168 5556 8174 5568
rect 8757 5559 8815 5565
rect 8757 5556 8769 5559
rect 8168 5528 8769 5556
rect 8168 5516 8174 5528
rect 8757 5525 8769 5528
rect 8803 5525 8815 5559
rect 8757 5519 8815 5525
rect 9766 5516 9772 5568
rect 9824 5556 9830 5568
rect 15378 5556 15384 5568
rect 9824 5528 15384 5556
rect 9824 5516 9830 5528
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 15838 5516 15844 5568
rect 15896 5556 15902 5568
rect 16776 5556 16804 5610
rect 15896 5528 16804 5556
rect 15896 5516 15902 5528
rect 0 5466 18860 5488
rect 0 5414 4660 5466
rect 4712 5414 4724 5466
rect 4776 5414 4788 5466
rect 4840 5414 4852 5466
rect 4904 5414 4916 5466
rect 4968 5414 7760 5466
rect 7812 5414 7824 5466
rect 7876 5414 7888 5466
rect 7940 5414 7952 5466
rect 8004 5414 8016 5466
rect 8068 5414 10860 5466
rect 10912 5414 10924 5466
rect 10976 5414 10988 5466
rect 11040 5414 11052 5466
rect 11104 5414 11116 5466
rect 11168 5414 13960 5466
rect 14012 5414 14024 5466
rect 14076 5414 14088 5466
rect 14140 5414 14152 5466
rect 14204 5414 14216 5466
rect 14268 5414 17060 5466
rect 17112 5414 17124 5466
rect 17176 5414 17188 5466
rect 17240 5414 17252 5466
rect 17304 5414 17316 5466
rect 17368 5414 18860 5466
rect 0 5392 18860 5414
rect 2498 5352 2504 5364
rect 1872 5324 2504 5352
rect 1872 5270 1900 5324
rect 2498 5312 2504 5324
rect 2556 5312 2562 5364
rect 2869 5355 2927 5361
rect 2869 5321 2881 5355
rect 2915 5352 2927 5355
rect 3970 5352 3976 5364
rect 2915 5324 3976 5352
rect 2915 5321 2927 5324
rect 2869 5315 2927 5321
rect 3970 5312 3976 5324
rect 4028 5312 4034 5364
rect 9766 5352 9772 5364
rect 6656 5324 9168 5352
rect 9727 5324 9772 5352
rect 6656 5293 6684 5324
rect 9140 5296 9168 5324
rect 9766 5312 9772 5324
rect 9824 5312 9830 5364
rect 9950 5312 9956 5364
rect 10008 5352 10014 5364
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 10008 5324 10425 5352
rect 10008 5312 10014 5324
rect 10413 5321 10425 5324
rect 10459 5352 10471 5355
rect 11330 5352 11336 5364
rect 10459 5324 11336 5352
rect 10459 5321 10471 5324
rect 10413 5315 10471 5321
rect 11330 5312 11336 5324
rect 11388 5312 11394 5364
rect 11606 5312 11612 5364
rect 11664 5352 11670 5364
rect 12069 5355 12127 5361
rect 12069 5352 12081 5355
rect 11664 5324 12081 5352
rect 11664 5312 11670 5324
rect 12069 5321 12081 5324
rect 12115 5321 12127 5355
rect 18138 5352 18144 5364
rect 12069 5315 12127 5321
rect 13556 5324 18144 5352
rect 6641 5287 6699 5293
rect 6641 5253 6653 5287
rect 6687 5253 6699 5287
rect 6641 5247 6699 5253
rect 7006 5244 7012 5296
rect 7064 5284 7070 5296
rect 8110 5284 8116 5296
rect 7064 5256 8116 5284
rect 7064 5244 7070 5256
rect 8110 5244 8116 5256
rect 8168 5284 8174 5296
rect 8168 5256 8326 5284
rect 8168 5244 8174 5256
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 10321 5287 10379 5293
rect 10321 5284 10333 5287
rect 9180 5256 10333 5284
rect 9180 5244 9186 5256
rect 10321 5253 10333 5256
rect 10367 5253 10379 5287
rect 10321 5247 10379 5253
rect 10689 5287 10747 5293
rect 10689 5253 10701 5287
rect 10735 5284 10747 5287
rect 11238 5284 11244 5296
rect 10735 5256 11244 5284
rect 10735 5253 10747 5256
rect 10689 5247 10747 5253
rect 11238 5244 11244 5256
rect 11296 5244 11302 5296
rect 11882 5284 11888 5296
rect 11843 5256 11888 5284
rect 11882 5244 11888 5256
rect 11940 5284 11946 5296
rect 13556 5293 13584 5324
rect 18138 5312 18144 5324
rect 18196 5312 18202 5364
rect 13541 5287 13599 5293
rect 11940 5256 12374 5284
rect 11940 5244 11946 5256
rect 13541 5253 13553 5287
rect 13587 5253 13599 5287
rect 13541 5247 13599 5253
rect 14274 5244 14280 5296
rect 14332 5284 14338 5296
rect 14829 5287 14887 5293
rect 14829 5284 14841 5287
rect 14332 5256 14841 5284
rect 14332 5244 14338 5256
rect 14829 5253 14841 5256
rect 14875 5284 14887 5287
rect 15286 5284 15292 5296
rect 14875 5256 15292 5284
rect 14875 5253 14887 5256
rect 14829 5247 14887 5253
rect 15286 5244 15292 5256
rect 15344 5284 15350 5296
rect 15654 5284 15660 5296
rect 15344 5256 15660 5284
rect 15344 5244 15350 5256
rect 15654 5244 15660 5256
rect 15712 5244 15718 5296
rect 15838 5244 15844 5296
rect 15896 5244 15902 5296
rect 477 5219 535 5225
rect 477 5185 489 5219
rect 523 5216 535 5219
rect 566 5216 572 5228
rect 523 5188 572 5216
rect 523 5185 535 5188
rect 477 5179 535 5185
rect 566 5176 572 5188
rect 624 5176 630 5228
rect 2271 5219 2329 5225
rect 2271 5185 2283 5219
rect 2317 5216 2329 5219
rect 2590 5216 2596 5228
rect 2317 5188 2596 5216
rect 2317 5185 2329 5188
rect 2271 5179 2329 5185
rect 2590 5176 2596 5188
rect 2648 5216 2654 5228
rect 2777 5219 2835 5225
rect 2777 5216 2789 5219
rect 2648 5188 2789 5216
rect 2648 5176 2654 5188
rect 2777 5185 2789 5188
rect 2823 5185 2835 5219
rect 2777 5179 2835 5185
rect 5994 5176 6000 5228
rect 6052 5216 6058 5228
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 6052 5188 6469 5216
rect 6052 5176 6058 5188
rect 6457 5185 6469 5188
rect 6503 5216 6515 5219
rect 7558 5216 7564 5228
rect 6503 5188 7564 5216
rect 6503 5185 6515 5188
rect 6457 5179 6515 5185
rect 7558 5176 7564 5188
rect 7616 5176 7622 5228
rect 10594 5216 10600 5228
rect 10555 5188 10600 5216
rect 10594 5176 10600 5188
rect 10652 5176 10658 5228
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 14918 5216 14924 5228
rect 14879 5188 14924 5216
rect 10781 5179 10839 5185
rect 845 5151 903 5157
rect 845 5117 857 5151
rect 891 5148 903 5151
rect 3694 5148 3700 5160
rect 891 5120 3700 5148
rect 891 5117 903 5120
rect 845 5111 903 5117
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5148 7895 5151
rect 8478 5148 8484 5160
rect 7883 5120 8484 5148
rect 7883 5117 7895 5120
rect 7837 5111 7895 5117
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10502 5148 10508 5160
rect 10100 5120 10508 5148
rect 10100 5108 10106 5120
rect 10502 5108 10508 5120
rect 10560 5148 10566 5160
rect 10796 5148 10824 5179
rect 14918 5176 14924 5188
rect 14976 5176 14982 5228
rect 18233 5219 18291 5225
rect 18233 5185 18245 5219
rect 18279 5216 18291 5219
rect 18506 5216 18512 5228
rect 18279 5188 18512 5216
rect 18279 5185 18291 5188
rect 18233 5179 18291 5185
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 13814 5148 13820 5160
rect 10560 5120 10824 5148
rect 13775 5120 13820 5148
rect 10560 5108 10566 5120
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5148 15255 5151
rect 15243 5120 18368 5148
rect 15243 5117 15255 5120
rect 15197 5111 15255 5117
rect 18340 5089 18368 5120
rect 18325 5083 18383 5089
rect 18325 5049 18337 5083
rect 18371 5049 18383 5083
rect 18325 5043 18383 5049
rect 2498 4972 2504 5024
rect 2556 5012 2562 5024
rect 3605 5015 3663 5021
rect 3605 5012 3617 5015
rect 2556 4984 3617 5012
rect 2556 4972 2562 4984
rect 3605 4981 3617 4984
rect 3651 5012 3663 5015
rect 3881 5015 3939 5021
rect 3881 5012 3893 5015
rect 3651 4984 3893 5012
rect 3651 4981 3663 4984
rect 3605 4975 3663 4981
rect 3881 4981 3893 4984
rect 3927 4981 3939 5015
rect 3881 4975 3939 4981
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 5442 5012 5448 5024
rect 4488 4984 5448 5012
rect 4488 4972 4494 4984
rect 5442 4972 5448 4984
rect 5500 5012 5506 5024
rect 5905 5015 5963 5021
rect 5905 5012 5917 5015
rect 5500 4984 5917 5012
rect 5500 4972 5506 4984
rect 5905 4981 5917 4984
rect 5951 5012 5963 5015
rect 7006 5012 7012 5024
rect 5951 4984 7012 5012
rect 5951 4981 5963 4984
rect 5905 4975 5963 4981
rect 7006 4972 7012 4984
rect 7064 5012 7070 5024
rect 7377 5015 7435 5021
rect 7377 5012 7389 5015
rect 7064 4984 7389 5012
rect 7064 4972 7070 4984
rect 7377 4981 7389 4984
rect 7423 4981 7435 5015
rect 7377 4975 7435 4981
rect 9030 4972 9036 5024
rect 9088 5012 9094 5024
rect 9309 5015 9367 5021
rect 9309 5012 9321 5015
rect 9088 4984 9321 5012
rect 9088 4972 9094 4984
rect 9309 4981 9321 4984
rect 9355 4981 9367 5015
rect 16666 5012 16672 5024
rect 16627 4984 16672 5012
rect 9309 4975 9367 4981
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 0 4922 18860 4944
rect 0 4870 3110 4922
rect 3162 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 6210 4922
rect 6262 4870 6274 4922
rect 6326 4870 6338 4922
rect 6390 4870 6402 4922
rect 6454 4870 6466 4922
rect 6518 4870 9310 4922
rect 9362 4870 9374 4922
rect 9426 4870 9438 4922
rect 9490 4870 9502 4922
rect 9554 4870 9566 4922
rect 9618 4870 12410 4922
rect 12462 4870 12474 4922
rect 12526 4870 12538 4922
rect 12590 4870 12602 4922
rect 12654 4870 12666 4922
rect 12718 4870 15510 4922
rect 15562 4870 15574 4922
rect 15626 4870 15638 4922
rect 15690 4870 15702 4922
rect 15754 4870 15766 4922
rect 15818 4870 18860 4922
rect 0 4848 18860 4870
rect 13265 4811 13323 4817
rect 13265 4777 13277 4811
rect 13311 4808 13323 4811
rect 14366 4808 14372 4820
rect 13311 4780 14372 4808
rect 13311 4777 13323 4780
rect 13265 4771 13323 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 14550 4768 14556 4820
rect 14608 4808 14614 4820
rect 14608 4780 17908 4808
rect 14608 4768 14614 4780
rect 3421 4743 3479 4749
rect 3421 4709 3433 4743
rect 3467 4709 3479 4743
rect 3421 4703 3479 4709
rect 10873 4743 10931 4749
rect 10873 4709 10885 4743
rect 10919 4740 10931 4743
rect 11238 4740 11244 4752
rect 10919 4712 11244 4740
rect 10919 4709 10931 4712
rect 10873 4703 10931 4709
rect 2958 4672 2964 4684
rect 2919 4644 2964 4672
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4573 3111 4607
rect 3436 4604 3464 4703
rect 11238 4700 11244 4712
rect 11296 4700 11302 4752
rect 15286 4700 15292 4752
rect 15344 4740 15350 4752
rect 15657 4743 15715 4749
rect 15657 4740 15669 4743
rect 15344 4712 15669 4740
rect 15344 4700 15350 4712
rect 15657 4709 15669 4712
rect 15703 4709 15715 4743
rect 15657 4703 15715 4709
rect 3697 4675 3755 4681
rect 3697 4641 3709 4675
rect 3743 4672 3755 4675
rect 5994 4672 6000 4684
rect 3743 4644 6000 4672
rect 3743 4641 3755 4644
rect 3697 4635 3755 4641
rect 5994 4632 6000 4644
rect 6052 4632 6058 4684
rect 7101 4675 7159 4681
rect 7101 4641 7113 4675
rect 7147 4672 7159 4675
rect 8294 4672 8300 4684
rect 7147 4644 8300 4672
rect 7147 4641 7159 4644
rect 7101 4635 7159 4641
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8938 4672 8944 4684
rect 8899 4644 8944 4672
rect 8938 4632 8944 4644
rect 8996 4632 9002 4684
rect 9401 4675 9459 4681
rect 9401 4641 9413 4675
rect 9447 4672 9459 4675
rect 10042 4672 10048 4684
rect 9447 4644 10048 4672
rect 9447 4641 9459 4644
rect 9401 4635 9459 4641
rect 10042 4632 10048 4644
rect 10100 4632 10106 4684
rect 11330 4672 11336 4684
rect 11291 4644 11336 4672
rect 11330 4632 11336 4644
rect 11388 4632 11394 4684
rect 11422 4632 11428 4684
rect 11480 4672 11486 4684
rect 14734 4672 14740 4684
rect 11480 4644 11525 4672
rect 14695 4644 14740 4672
rect 11480 4632 11486 4644
rect 14734 4632 14740 4644
rect 14792 4632 14798 4684
rect 15010 4672 15016 4684
rect 14971 4644 15016 4672
rect 15010 4632 15016 4644
rect 15068 4632 15074 4684
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 3436 4576 4077 4604
rect 3053 4567 3111 4573
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 3068 4468 3096 4567
rect 6178 4564 6184 4616
rect 6236 4604 6242 4616
rect 6273 4607 6331 4613
rect 6273 4604 6285 4607
rect 6236 4576 6285 4604
rect 6236 4564 6242 4576
rect 6273 4573 6285 4576
rect 6319 4573 6331 4607
rect 6273 4567 6331 4573
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4604 6423 4607
rect 6546 4604 6552 4616
rect 6411 4576 6552 4604
rect 6411 4573 6423 4576
rect 6365 4567 6423 4573
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 7006 4604 7012 4616
rect 6967 4576 7012 4604
rect 7006 4564 7012 4576
rect 7064 4564 7070 4616
rect 9030 4604 9036 4616
rect 8991 4576 9036 4604
rect 9030 4564 9036 4576
rect 9088 4564 9094 4616
rect 11348 4604 11376 4632
rect 11701 4607 11759 4613
rect 11701 4604 11713 4607
rect 11348 4576 11713 4604
rect 11701 4573 11713 4576
rect 11747 4604 11759 4607
rect 12250 4604 12256 4616
rect 11747 4576 12256 4604
rect 11747 4573 11759 4576
rect 11701 4567 11759 4573
rect 12250 4564 12256 4576
rect 12308 4564 12314 4616
rect 15105 4607 15163 4613
rect 15105 4573 15117 4607
rect 15151 4573 15163 4607
rect 15105 4567 15163 4573
rect 4430 4496 4436 4548
rect 4488 4496 4494 4548
rect 5491 4539 5549 4545
rect 5491 4536 5503 4539
rect 5184 4508 5503 4536
rect 5184 4468 5212 4508
rect 5491 4505 5503 4508
rect 5537 4536 5549 4539
rect 11241 4539 11299 4545
rect 11241 4536 11253 4539
rect 5537 4508 11253 4536
rect 5537 4505 5549 4508
rect 5491 4499 5549 4505
rect 11241 4505 11253 4508
rect 11287 4505 11299 4539
rect 11241 4499 11299 4505
rect 11330 4496 11336 4548
rect 11388 4536 11394 4548
rect 11946 4539 12004 4545
rect 11946 4536 11958 4539
rect 11388 4508 11958 4536
rect 11388 4496 11394 4508
rect 11946 4505 11958 4508
rect 11992 4505 12004 4539
rect 11946 4499 12004 4505
rect 14274 4496 14280 4548
rect 14332 4496 14338 4548
rect 14642 4496 14648 4548
rect 14700 4536 14706 4548
rect 15120 4536 15148 4567
rect 15216 4539 15274 4545
rect 15216 4536 15228 4539
rect 14700 4508 15148 4536
rect 14700 4496 14706 4508
rect 15212 4505 15228 4536
rect 15262 4505 15274 4539
rect 15378 4536 15384 4548
rect 15339 4508 15384 4536
rect 15212 4499 15274 4505
rect 6086 4468 6092 4480
rect 3068 4440 5212 4468
rect 6047 4440 6092 4468
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 6730 4468 6736 4480
rect 6691 4440 6736 4468
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 7377 4471 7435 4477
rect 7377 4437 7389 4471
rect 7423 4468 7435 4471
rect 7650 4468 7656 4480
rect 7423 4440 7656 4468
rect 7423 4437 7435 4440
rect 7377 4431 7435 4437
rect 7650 4428 7656 4440
rect 7708 4428 7714 4480
rect 13081 4471 13139 4477
rect 13081 4437 13093 4471
rect 13127 4468 13139 4471
rect 13170 4468 13176 4480
rect 13127 4440 13176 4468
rect 13127 4437 13139 4440
rect 13081 4431 13139 4437
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 13722 4428 13728 4480
rect 13780 4468 13786 4480
rect 14292 4468 14320 4496
rect 13780 4440 14320 4468
rect 13780 4428 13786 4440
rect 14458 4428 14464 4480
rect 14516 4468 14522 4480
rect 15105 4471 15163 4477
rect 15105 4468 15117 4471
rect 14516 4440 15117 4468
rect 14516 4428 14522 4440
rect 15105 4437 15117 4440
rect 15151 4437 15163 4471
rect 15212 4468 15240 4499
rect 15378 4496 15384 4508
rect 15436 4496 15442 4548
rect 15672 4536 15700 4703
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4672 16175 4675
rect 16666 4672 16672 4684
rect 16163 4644 16672 4672
rect 16163 4641 16175 4644
rect 16117 4635 16175 4641
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 17880 4681 17908 4780
rect 17865 4675 17923 4681
rect 17865 4641 17877 4675
rect 17911 4641 17923 4675
rect 17865 4635 17923 4641
rect 15838 4604 15844 4616
rect 15799 4576 15844 4604
rect 15838 4564 15844 4576
rect 15896 4564 15902 4616
rect 15746 4536 15752 4548
rect 15659 4508 15752 4536
rect 15746 4496 15752 4508
rect 15804 4536 15810 4548
rect 16574 4536 16580 4548
rect 15804 4508 16580 4536
rect 15804 4496 15810 4508
rect 16574 4496 16580 4508
rect 16632 4496 16638 4548
rect 15930 4468 15936 4480
rect 15212 4440 15936 4468
rect 15105 4431 15163 4437
rect 15930 4428 15936 4440
rect 15988 4428 15994 4480
rect 0 4378 18860 4400
rect 0 4326 4660 4378
rect 4712 4326 4724 4378
rect 4776 4326 4788 4378
rect 4840 4326 4852 4378
rect 4904 4326 4916 4378
rect 4968 4326 7760 4378
rect 7812 4326 7824 4378
rect 7876 4326 7888 4378
rect 7940 4326 7952 4378
rect 8004 4326 8016 4378
rect 8068 4326 10860 4378
rect 10912 4326 10924 4378
rect 10976 4326 10988 4378
rect 11040 4326 11052 4378
rect 11104 4326 11116 4378
rect 11168 4326 13960 4378
rect 14012 4326 14024 4378
rect 14076 4326 14088 4378
rect 14140 4326 14152 4378
rect 14204 4326 14216 4378
rect 14268 4326 17060 4378
rect 17112 4326 17124 4378
rect 17176 4326 17188 4378
rect 17240 4326 17252 4378
rect 17304 4326 17316 4378
rect 17368 4326 18860 4378
rect 0 4304 18860 4326
rect 2317 4267 2375 4273
rect 2317 4264 2329 4267
rect 1688 4236 2329 4264
rect 1688 4182 1716 4236
rect 2317 4233 2329 4236
rect 2363 4264 2375 4267
rect 2498 4264 2504 4276
rect 2363 4236 2504 4264
rect 2363 4233 2375 4236
rect 2317 4227 2375 4233
rect 2498 4224 2504 4236
rect 2556 4224 2562 4276
rect 2958 4264 2964 4276
rect 2919 4236 2964 4264
rect 2958 4224 2964 4236
rect 3016 4224 3022 4276
rect 5534 4264 5540 4276
rect 4908 4236 5540 4264
rect 3421 4199 3479 4205
rect 3421 4165 3433 4199
rect 3467 4196 3479 4199
rect 3467 4168 4844 4196
rect 3467 4165 3479 4168
rect 3421 4159 3479 4165
rect 2590 4128 2596 4140
rect 2551 4100 2596 4128
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4097 2743 4131
rect 2685 4091 2743 4097
rect 290 4060 296 4072
rect 251 4032 296 4060
rect 290 4020 296 4032
rect 348 4020 354 4072
rect 661 4063 719 4069
rect 661 4029 673 4063
rect 707 4060 719 4063
rect 842 4060 848 4072
rect 707 4032 848 4060
rect 707 4029 719 4032
rect 661 4023 719 4029
rect 842 4020 848 4032
rect 900 4020 906 4072
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4029 2191 4063
rect 2700 4060 2728 4091
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 3973 4131 4031 4137
rect 2832 4100 2877 4128
rect 2832 4088 2838 4100
rect 3973 4097 3985 4131
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 2133 4023 2191 4029
rect 2608 4032 2728 4060
rect 3513 4063 3571 4069
rect 2148 3992 2176 4023
rect 2608 3992 2636 4032
rect 3513 4029 3525 4063
rect 3559 4029 3571 4063
rect 3513 4023 3571 4029
rect 2682 3992 2688 4004
rect 2148 3964 2688 3992
rect 2682 3952 2688 3964
rect 2740 3992 2746 4004
rect 3528 3992 3556 4023
rect 3602 4020 3608 4072
rect 3660 4060 3666 4072
rect 3660 4032 3705 4060
rect 3660 4020 3666 4032
rect 3881 3995 3939 4001
rect 3881 3992 3893 3995
rect 2740 3964 3372 3992
rect 3528 3964 3893 3992
rect 2740 3952 2746 3964
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 3053 3927 3111 3933
rect 3053 3924 3065 3927
rect 2372 3896 3065 3924
rect 2372 3884 2378 3896
rect 3053 3893 3065 3896
rect 3099 3893 3111 3927
rect 3344 3924 3372 3964
rect 3881 3961 3893 3964
rect 3927 3961 3939 3995
rect 3881 3955 3939 3961
rect 3988 3924 4016 4091
rect 3344 3896 4016 3924
rect 3053 3887 3111 3893
rect 4338 3884 4344 3936
rect 4396 3924 4402 3936
rect 4617 3927 4675 3933
rect 4617 3924 4629 3927
rect 4396 3896 4629 3924
rect 4396 3884 4402 3896
rect 4617 3893 4629 3896
rect 4663 3893 4675 3927
rect 4816 3924 4844 4168
rect 4908 4137 4936 4236
rect 5534 4224 5540 4236
rect 5592 4264 5598 4276
rect 5994 4264 6000 4276
rect 5592 4236 6000 4264
rect 5592 4224 5598 4236
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 7650 4264 7656 4276
rect 7611 4236 7656 4264
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 8573 4267 8631 4273
rect 8573 4233 8585 4267
rect 8619 4264 8631 4267
rect 8938 4264 8944 4276
rect 8619 4236 8944 4264
rect 8619 4233 8631 4236
rect 8573 4227 8631 4233
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 9125 4267 9183 4273
rect 9125 4233 9137 4267
rect 9171 4264 9183 4267
rect 9677 4267 9735 4273
rect 9677 4264 9689 4267
rect 9171 4236 9689 4264
rect 9171 4233 9183 4236
rect 9125 4227 9183 4233
rect 9677 4233 9689 4236
rect 9723 4233 9735 4267
rect 10042 4264 10048 4276
rect 10003 4236 10048 4264
rect 9677 4227 9735 4233
rect 10042 4224 10048 4236
rect 10100 4224 10106 4276
rect 11241 4267 11299 4273
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 11422 4264 11428 4276
rect 11287 4236 11428 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11422 4224 11428 4236
rect 11480 4224 11486 4276
rect 12158 4224 12164 4276
rect 12216 4264 12222 4276
rect 12713 4267 12771 4273
rect 12713 4264 12725 4267
rect 12216 4236 12725 4264
rect 12216 4224 12222 4236
rect 12713 4233 12725 4236
rect 12759 4233 12771 4267
rect 12713 4227 12771 4233
rect 13541 4267 13599 4273
rect 13541 4233 13553 4267
rect 13587 4264 13599 4267
rect 13722 4264 13728 4276
rect 13587 4236 13728 4264
rect 13587 4233 13599 4236
rect 13541 4227 13599 4233
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 14277 4267 14335 4273
rect 14277 4233 14289 4267
rect 14323 4264 14335 4267
rect 14642 4264 14648 4276
rect 14323 4236 14648 4264
rect 14323 4233 14335 4236
rect 14277 4227 14335 4233
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 14918 4224 14924 4276
rect 14976 4264 14982 4276
rect 15838 4264 15844 4276
rect 14976 4236 15844 4264
rect 14976 4224 14982 4236
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 5626 4156 5632 4208
rect 5684 4156 5690 4208
rect 14550 4196 14556 4208
rect 9140 4168 10640 4196
rect 4893 4131 4951 4137
rect 4893 4097 4905 4131
rect 4939 4097 4951 4131
rect 4893 4091 4951 4097
rect 6687 4131 6745 4137
rect 6687 4097 6699 4131
rect 6733 4128 6745 4131
rect 7006 4128 7012 4140
rect 6733 4100 7012 4128
rect 6733 4097 6745 4100
rect 6687 4091 6745 4097
rect 7006 4088 7012 4100
rect 7064 4128 7070 4140
rect 8202 4128 8208 4140
rect 7064 4100 8208 4128
rect 7064 4088 7070 4100
rect 8202 4088 8208 4100
rect 8260 4128 8266 4140
rect 8481 4131 8539 4137
rect 8481 4128 8493 4131
rect 8260 4100 8493 4128
rect 8260 4088 8266 4100
rect 8481 4097 8493 4100
rect 8527 4097 8539 4131
rect 8481 4091 8539 4097
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 5261 4063 5319 4069
rect 5261 4029 5273 4063
rect 5307 4060 5319 4063
rect 6086 4060 6092 4072
rect 5307 4032 6092 4060
rect 5307 4029 5319 4032
rect 5261 4023 5319 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 7745 4063 7803 4069
rect 7745 4029 7757 4063
rect 7791 4029 7803 4063
rect 7745 4023 7803 4029
rect 7929 4063 7987 4069
rect 7929 4029 7941 4063
rect 7975 4029 7987 4063
rect 7929 4023 7987 4029
rect 7760 3992 7788 4023
rect 6012 3964 7788 3992
rect 7944 3992 7972 4023
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 8680 4060 8708 4091
rect 8754 4088 8760 4140
rect 8812 4128 8818 4140
rect 9140 4128 9168 4168
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 8812 4100 9168 4128
rect 9232 4100 10149 4128
rect 8812 4088 8818 4100
rect 9232 4072 9260 4100
rect 10137 4097 10149 4100
rect 10183 4128 10195 4131
rect 10612 4128 10640 4168
rect 12406 4168 14556 4196
rect 11149 4131 11207 4137
rect 11149 4128 11161 4131
rect 10183 4100 10456 4128
rect 10612 4100 11161 4128
rect 10183 4097 10195 4100
rect 10137 4091 10195 4097
rect 9214 4060 9220 4072
rect 8352 4032 8708 4060
rect 9175 4032 9220 4060
rect 8352 4020 8358 4032
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 9401 4063 9459 4069
rect 9401 4029 9413 4063
rect 9447 4060 9459 4063
rect 9858 4060 9864 4072
rect 9447 4032 9864 4060
rect 9447 4029 9459 4032
rect 9401 4023 9459 4029
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 10226 4020 10232 4072
rect 10284 4060 10290 4072
rect 10284 4032 10329 4060
rect 10284 4020 10290 4032
rect 10244 3992 10272 4020
rect 7944 3964 10272 3992
rect 10428 3992 10456 4100
rect 11149 4097 11161 4100
rect 11195 4097 11207 4131
rect 11330 4128 11336 4140
rect 11291 4100 11336 4128
rect 11149 4091 11207 4097
rect 11164 4060 11192 4091
rect 11330 4088 11336 4100
rect 11388 4128 11394 4140
rect 12406 4128 12434 4168
rect 11388 4100 12434 4128
rect 12897 4131 12955 4137
rect 11388 4088 11394 4100
rect 12897 4097 12909 4131
rect 12943 4128 12955 4131
rect 13170 4128 13176 4140
rect 12943 4100 13176 4128
rect 12943 4097 12955 4100
rect 12897 4091 12955 4097
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 13372 4137 13400 4168
rect 13740 4140 13768 4168
rect 14550 4156 14556 4168
rect 14608 4156 14614 4208
rect 15746 4156 15752 4208
rect 15804 4156 15810 4208
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4097 13415 4131
rect 13357 4091 13415 4097
rect 12621 4063 12679 4069
rect 11164 4032 12434 4060
rect 11330 3992 11336 4004
rect 10428 3964 11336 3992
rect 6012 3936 6040 3964
rect 5994 3924 6000 3936
rect 4816 3896 6000 3924
rect 4617 3887 4675 3893
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 7282 3924 7288 3936
rect 7243 3896 7288 3924
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 7760 3924 7788 3964
rect 11330 3952 11336 3964
rect 11388 3952 11394 4004
rect 12406 3992 12434 4032
rect 12621 4029 12633 4063
rect 12667 4060 12679 4063
rect 12986 4060 12992 4072
rect 12667 4032 12992 4060
rect 12667 4029 12679 4032
rect 12621 4023 12679 4029
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4060 13139 4063
rect 13372 4060 13400 4091
rect 13722 4088 13728 4140
rect 13780 4088 13786 4140
rect 13817 4131 13875 4137
rect 13817 4097 13829 4131
rect 13863 4128 13875 4131
rect 15102 4128 15108 4140
rect 13863 4100 15108 4128
rect 13863 4097 13875 4100
rect 13817 4091 13875 4097
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 18233 4131 18291 4137
rect 18233 4097 18245 4131
rect 18279 4128 18291 4131
rect 18506 4128 18512 4140
rect 18279 4100 18512 4128
rect 18279 4097 18291 4100
rect 18233 4091 18291 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 13127 4032 13400 4060
rect 13127 4029 13139 4032
rect 13081 4023 13139 4029
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 13504 4032 14228 4060
rect 13504 4020 13510 4032
rect 14200 3992 14228 4032
rect 14366 4020 14372 4072
rect 14424 4060 14430 4072
rect 14645 4063 14703 4069
rect 14645 4060 14657 4063
rect 14424 4032 14657 4060
rect 14424 4020 14430 4032
rect 14645 4029 14657 4032
rect 14691 4029 14703 4063
rect 14826 4060 14832 4072
rect 14787 4032 14832 4060
rect 14645 4023 14703 4029
rect 14826 4020 14832 4032
rect 14884 4020 14890 4072
rect 15197 4063 15255 4069
rect 15197 4029 15209 4063
rect 15243 4060 15255 4063
rect 15243 4032 18368 4060
rect 15243 4029 15255 4032
rect 15197 4023 15255 4029
rect 14461 3995 14519 4001
rect 14461 3992 14473 3995
rect 12406 3964 14136 3992
rect 14200 3964 14473 3992
rect 14108 3936 14136 3964
rect 14461 3961 14473 3964
rect 14507 3992 14519 3995
rect 14550 3992 14556 4004
rect 14507 3964 14556 3992
rect 14507 3961 14519 3964
rect 14461 3955 14519 3961
rect 14550 3952 14556 3964
rect 14608 3952 14614 4004
rect 18340 4001 18368 4032
rect 18325 3995 18383 4001
rect 18325 3961 18337 3995
rect 18371 3961 18383 3995
rect 18325 3955 18383 3961
rect 8662 3924 8668 3936
rect 7760 3896 8668 3924
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 8754 3884 8760 3936
rect 8812 3924 8818 3936
rect 8812 3896 8857 3924
rect 8812 3884 8818 3896
rect 9122 3884 9128 3936
rect 9180 3924 9186 3936
rect 12621 3927 12679 3933
rect 12621 3924 12633 3927
rect 9180 3896 12633 3924
rect 9180 3884 9186 3896
rect 12621 3893 12633 3896
rect 12667 3893 12679 3927
rect 12621 3887 12679 3893
rect 12802 3884 12808 3936
rect 12860 3924 12866 3936
rect 13173 3927 13231 3933
rect 13173 3924 13185 3927
rect 12860 3896 13185 3924
rect 12860 3884 12866 3896
rect 13173 3893 13185 3896
rect 13219 3893 13231 3927
rect 14090 3924 14096 3936
rect 14051 3896 14096 3924
rect 13173 3887 13231 3893
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 16623 3927 16681 3933
rect 16623 3924 16635 3927
rect 16172 3896 16635 3924
rect 16172 3884 16178 3896
rect 16623 3893 16635 3896
rect 16669 3893 16681 3927
rect 16623 3887 16681 3893
rect 0 3834 18860 3856
rect 0 3782 3110 3834
rect 3162 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 6210 3834
rect 6262 3782 6274 3834
rect 6326 3782 6338 3834
rect 6390 3782 6402 3834
rect 6454 3782 6466 3834
rect 6518 3782 9310 3834
rect 9362 3782 9374 3834
rect 9426 3782 9438 3834
rect 9490 3782 9502 3834
rect 9554 3782 9566 3834
rect 9618 3782 12410 3834
rect 12462 3782 12474 3834
rect 12526 3782 12538 3834
rect 12590 3782 12602 3834
rect 12654 3782 12666 3834
rect 12718 3782 15510 3834
rect 15562 3782 15574 3834
rect 15626 3782 15638 3834
rect 15690 3782 15702 3834
rect 15754 3782 15766 3834
rect 15818 3782 18860 3834
rect 0 3760 18860 3782
rect 842 3720 848 3732
rect 803 3692 848 3720
rect 842 3680 848 3692
rect 900 3680 906 3732
rect 6273 3723 6331 3729
rect 6273 3689 6285 3723
rect 6319 3720 6331 3723
rect 6546 3720 6552 3732
rect 6319 3692 6552 3720
rect 6319 3689 6331 3692
rect 6273 3683 6331 3689
rect 6546 3680 6552 3692
rect 6604 3680 6610 3732
rect 6730 3680 6736 3732
rect 6788 3680 6794 3732
rect 8478 3720 8484 3732
rect 8439 3692 8484 3720
rect 8478 3680 8484 3692
rect 8536 3680 8542 3732
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 8628 3692 10701 3720
rect 8628 3680 8634 3692
rect 10689 3689 10701 3692
rect 10735 3689 10747 3723
rect 10689 3683 10747 3689
rect 13078 3680 13084 3732
rect 13136 3720 13142 3732
rect 13538 3720 13544 3732
rect 13136 3692 13544 3720
rect 13136 3680 13142 3692
rect 13538 3680 13544 3692
rect 13596 3720 13602 3732
rect 13633 3723 13691 3729
rect 13633 3720 13645 3723
rect 13596 3692 13645 3720
rect 13596 3680 13602 3692
rect 13633 3689 13645 3692
rect 13679 3689 13691 3723
rect 14458 3720 14464 3732
rect 13633 3683 13691 3689
rect 13832 3692 14464 3720
rect 2590 3652 2596 3664
rect 2240 3624 2596 3652
rect 2240 3596 2268 3624
rect 2590 3612 2596 3624
rect 2648 3652 2654 3664
rect 3513 3655 3571 3661
rect 3513 3652 3525 3655
rect 2648 3624 3525 3652
rect 2648 3612 2654 3624
rect 3513 3621 3525 3624
rect 3559 3621 3571 3655
rect 3513 3615 3571 3621
rect 5905 3655 5963 3661
rect 5905 3621 5917 3655
rect 5951 3652 5963 3655
rect 6748 3652 6776 3680
rect 5951 3624 6776 3652
rect 5951 3621 5963 3624
rect 5905 3615 5963 3621
rect 6822 3612 6828 3664
rect 6880 3612 6886 3664
rect 8202 3612 8208 3664
rect 8260 3652 8266 3664
rect 11238 3652 11244 3664
rect 8260 3624 9628 3652
rect 11199 3624 11244 3652
rect 8260 3612 8266 3624
rect 2222 3584 2228 3596
rect 2183 3556 2228 3584
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 2608 3556 3280 3584
rect 2608 3528 2636 3556
rect 1029 3519 1087 3525
rect 1029 3485 1041 3519
rect 1075 3516 1087 3519
rect 1949 3519 2007 3525
rect 1075 3488 1624 3516
rect 1075 3485 1087 3488
rect 1029 3479 1087 3485
rect 1596 3389 1624 3488
rect 1949 3485 1961 3519
rect 1995 3516 2007 3519
rect 2314 3516 2320 3528
rect 1995 3488 2320 3516
rect 1995 3485 2007 3488
rect 1949 3479 2007 3485
rect 2314 3476 2320 3488
rect 2372 3476 2378 3528
rect 2590 3476 2596 3528
rect 2648 3476 2654 3528
rect 2774 3476 2780 3528
rect 2832 3516 2838 3528
rect 3252 3525 3280 3556
rect 5994 3544 6000 3596
rect 6052 3584 6058 3596
rect 6733 3587 6791 3593
rect 6733 3584 6745 3587
rect 6052 3556 6745 3584
rect 6052 3544 6058 3556
rect 6733 3553 6745 3556
rect 6779 3553 6791 3587
rect 6840 3584 6868 3612
rect 6917 3587 6975 3593
rect 6917 3584 6929 3587
rect 6840 3556 6929 3584
rect 6733 3547 6791 3553
rect 6917 3553 6929 3556
rect 6963 3553 6975 3587
rect 8754 3584 8760 3596
rect 8715 3556 8760 3584
rect 6917 3547 6975 3553
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2832 3488 3065 3516
rect 2832 3476 2838 3488
rect 3053 3485 3065 3488
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3485 3295 3519
rect 5902 3516 5908 3528
rect 5863 3488 5908 3516
rect 3237 3479 3295 3485
rect 5902 3476 5908 3488
rect 5960 3476 5966 3528
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3516 6699 3519
rect 7282 3516 7288 3528
rect 6687 3488 7288 3516
rect 6687 3485 6699 3488
rect 6641 3479 6699 3485
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 8662 3516 8668 3528
rect 8623 3488 8668 3516
rect 8662 3476 8668 3488
rect 8720 3476 8726 3528
rect 8938 3476 8944 3528
rect 8996 3518 9002 3528
rect 9600 3525 9628 3624
rect 11238 3612 11244 3624
rect 11296 3612 11302 3664
rect 12158 3612 12164 3664
rect 12216 3652 12222 3664
rect 12437 3655 12495 3661
rect 12437 3652 12449 3655
rect 12216 3624 12449 3652
rect 12216 3612 12222 3624
rect 12437 3621 12449 3624
rect 12483 3621 12495 3655
rect 12437 3615 12495 3621
rect 12526 3612 12532 3664
rect 12584 3652 12590 3664
rect 12989 3655 13047 3661
rect 12989 3652 13001 3655
rect 12584 3624 13001 3652
rect 12584 3612 12590 3624
rect 12989 3621 13001 3624
rect 13035 3621 13047 3655
rect 12989 3615 13047 3621
rect 11790 3544 11796 3596
rect 11848 3584 11854 3596
rect 12253 3587 12311 3593
rect 12253 3584 12265 3587
rect 11848 3556 12265 3584
rect 11848 3544 11854 3556
rect 12253 3553 12265 3556
rect 12299 3553 12311 3587
rect 12253 3547 12311 3553
rect 12342 3544 12348 3596
rect 12400 3584 12406 3596
rect 13081 3587 13139 3593
rect 12400 3556 12848 3584
rect 12400 3544 12406 3556
rect 9217 3519 9275 3525
rect 8996 3516 9076 3518
rect 9217 3516 9229 3519
rect 8996 3490 9229 3516
rect 8996 3476 9002 3490
rect 9048 3488 9229 3490
rect 9217 3485 9229 3488
rect 9263 3485 9275 3519
rect 9217 3479 9275 3485
rect 9585 3519 9643 3525
rect 9585 3485 9597 3519
rect 9631 3485 9643 3519
rect 9766 3516 9772 3528
rect 9727 3488 9772 3516
rect 9585 3479 9643 3485
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 10229 3519 10287 3525
rect 10229 3485 10241 3519
rect 10275 3516 10287 3519
rect 10410 3516 10416 3528
rect 10275 3488 10416 3516
rect 10275 3485 10287 3488
rect 10229 3479 10287 3485
rect 10410 3476 10416 3488
rect 10468 3476 10474 3528
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 11238 3516 11244 3528
rect 10551 3488 11244 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 12529 3519 12587 3525
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 12710 3516 12716 3528
rect 12575 3488 12716 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 12820 3525 12848 3556
rect 13081 3553 13093 3587
rect 13127 3584 13139 3587
rect 13832 3584 13860 3692
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 15102 3680 15108 3732
rect 15160 3720 15166 3732
rect 15197 3723 15255 3729
rect 15197 3720 15209 3723
rect 15160 3692 15209 3720
rect 15160 3680 15166 3692
rect 15197 3689 15209 3692
rect 15243 3689 15255 3723
rect 15197 3683 15255 3689
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15381 3723 15439 3729
rect 15381 3720 15393 3723
rect 15344 3692 15393 3720
rect 15344 3680 15350 3692
rect 15381 3689 15393 3692
rect 15427 3689 15439 3723
rect 15381 3683 15439 3689
rect 16114 3584 16120 3596
rect 13127 3556 13860 3584
rect 16075 3556 16120 3584
rect 13127 3553 13139 3556
rect 13081 3547 13139 3553
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 17494 3584 17500 3596
rect 17455 3556 17500 3584
rect 17494 3544 17500 3556
rect 17552 3544 17558 3596
rect 12805 3519 12863 3525
rect 12805 3485 12817 3519
rect 12851 3485 12863 3519
rect 13446 3516 13452 3528
rect 13407 3488 13452 3516
rect 12805 3479 12863 3485
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 13722 3516 13728 3528
rect 13683 3488 13728 3516
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 15749 3519 15807 3525
rect 13872 3488 13917 3516
rect 13872 3476 13878 3488
rect 15749 3485 15761 3519
rect 15795 3516 15807 3519
rect 15838 3516 15844 3528
rect 15795 3488 15844 3516
rect 15795 3485 15807 3488
rect 15749 3479 15807 3485
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 17512 3516 17540 3544
rect 18233 3519 18291 3525
rect 18233 3516 18245 3519
rect 17512 3488 18245 3516
rect 18233 3485 18245 3488
rect 18279 3485 18291 3519
rect 18233 3479 18291 3485
rect 2041 3451 2099 3457
rect 2041 3417 2053 3451
rect 2087 3448 2099 3451
rect 2608 3448 2636 3476
rect 3602 3448 3608 3460
rect 2087 3420 2636 3448
rect 3160 3420 3608 3448
rect 2087 3417 2099 3420
rect 2041 3411 2099 3417
rect 3160 3392 3188 3420
rect 3602 3408 3608 3420
rect 3660 3408 3666 3460
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 5629 3451 5687 3457
rect 5629 3448 5641 3451
rect 5316 3420 5641 3448
rect 5316 3408 5322 3420
rect 5629 3417 5641 3420
rect 5675 3417 5687 3451
rect 5629 3411 5687 3417
rect 5813 3451 5871 3457
rect 5813 3417 5825 3451
rect 5859 3448 5871 3451
rect 7006 3448 7012 3460
rect 5859 3420 7012 3448
rect 5859 3417 5871 3420
rect 5813 3411 5871 3417
rect 7006 3408 7012 3420
rect 7064 3408 7070 3460
rect 8294 3448 8300 3460
rect 7208 3420 8300 3448
rect 1581 3383 1639 3389
rect 1581 3349 1593 3383
rect 1627 3349 1639 3383
rect 1581 3343 1639 3349
rect 2222 3340 2228 3392
rect 2280 3380 2286 3392
rect 2409 3383 2467 3389
rect 2409 3380 2421 3383
rect 2280 3352 2421 3380
rect 2280 3340 2286 3352
rect 2409 3349 2421 3352
rect 2455 3349 2467 3383
rect 3142 3380 3148 3392
rect 3103 3352 3148 3380
rect 2409 3343 2467 3349
rect 3142 3340 3148 3352
rect 3200 3340 3206 3392
rect 3421 3383 3479 3389
rect 3421 3349 3433 3383
rect 3467 3380 3479 3383
rect 3510 3380 3516 3392
rect 3467 3352 3516 3380
rect 3467 3349 3479 3352
rect 3421 3343 3479 3349
rect 3510 3340 3516 3352
rect 3568 3340 3574 3392
rect 5442 3340 5448 3392
rect 5500 3380 5506 3392
rect 7208 3380 7236 3420
rect 8294 3408 8300 3420
rect 8352 3408 8358 3460
rect 5500 3352 7236 3380
rect 7285 3383 7343 3389
rect 5500 3340 5506 3352
rect 7285 3349 7297 3383
rect 7331 3380 7343 3383
rect 7374 3380 7380 3392
rect 7331 3352 7380 3380
rect 7331 3349 7343 3352
rect 7285 3343 7343 3349
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 8680 3380 8708 3476
rect 9030 3408 9036 3460
rect 9088 3448 9094 3460
rect 9309 3451 9367 3457
rect 9309 3448 9321 3451
rect 9088 3420 9321 3448
rect 9088 3408 9094 3420
rect 9309 3417 9321 3420
rect 9355 3417 9367 3451
rect 9309 3411 9367 3417
rect 9493 3451 9551 3457
rect 9493 3417 9505 3451
rect 9539 3448 9551 3451
rect 9950 3448 9956 3460
rect 9539 3420 9956 3448
rect 9539 3417 9551 3420
rect 9493 3411 9551 3417
rect 9950 3408 9956 3420
rect 10008 3448 10014 3460
rect 10321 3451 10379 3457
rect 10321 3448 10333 3451
rect 10008 3420 10333 3448
rect 10008 3408 10014 3420
rect 10321 3417 10333 3420
rect 10367 3417 10379 3451
rect 10321 3411 10379 3417
rect 10689 3451 10747 3457
rect 10689 3417 10701 3451
rect 10735 3448 10747 3451
rect 10873 3451 10931 3457
rect 10873 3448 10885 3451
rect 10735 3420 10885 3448
rect 10735 3417 10747 3420
rect 10689 3411 10747 3417
rect 10873 3417 10885 3420
rect 10919 3448 10931 3451
rect 11514 3448 11520 3460
rect 10919 3420 11520 3448
rect 10919 3417 10931 3420
rect 10873 3411 10931 3417
rect 11514 3408 11520 3420
rect 11572 3408 11578 3460
rect 11790 3408 11796 3460
rect 11848 3448 11854 3460
rect 14090 3457 14096 3460
rect 13265 3451 13323 3457
rect 13265 3448 13277 3451
rect 11848 3420 13277 3448
rect 11848 3408 11854 3420
rect 13265 3417 13277 3420
rect 13311 3417 13323 3451
rect 14084 3448 14096 3457
rect 14003 3420 14096 3448
rect 13265 3411 13323 3417
rect 14084 3411 14096 3420
rect 14148 3448 14154 3460
rect 14148 3420 15516 3448
rect 14090 3408 14096 3411
rect 14148 3408 14154 3420
rect 7524 3352 8708 3380
rect 9125 3383 9183 3389
rect 7524 3340 7530 3352
rect 9125 3349 9137 3383
rect 9171 3380 9183 3383
rect 9217 3383 9275 3389
rect 9217 3380 9229 3383
rect 9171 3352 9229 3380
rect 9171 3349 9183 3352
rect 9125 3343 9183 3349
rect 9217 3349 9229 3352
rect 9263 3349 9275 3383
rect 9217 3343 9275 3349
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 9677 3383 9735 3389
rect 9677 3380 9689 3383
rect 9456 3352 9689 3380
rect 9456 3340 9462 3352
rect 9677 3349 9689 3352
rect 9723 3349 9735 3383
rect 9677 3343 9735 3349
rect 9766 3340 9772 3392
rect 9824 3380 9830 3392
rect 10229 3383 10287 3389
rect 10229 3380 10241 3383
rect 9824 3352 10241 3380
rect 9824 3340 9830 3352
rect 10229 3349 10241 3352
rect 10275 3349 10287 3383
rect 11330 3380 11336 3392
rect 11291 3352 11336 3380
rect 10229 3343 10287 3349
rect 11330 3340 11336 3352
rect 11388 3340 11394 3392
rect 12253 3383 12311 3389
rect 12253 3349 12265 3383
rect 12299 3380 12311 3383
rect 12526 3380 12532 3392
rect 12299 3352 12532 3380
rect 12299 3349 12311 3352
rect 12253 3343 12311 3349
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 15488 3380 15516 3420
rect 16574 3408 16580 3460
rect 16632 3408 16638 3460
rect 18049 3451 18107 3457
rect 18049 3448 18061 3451
rect 17236 3420 18061 3448
rect 17236 3380 17264 3420
rect 18049 3417 18061 3420
rect 18095 3417 18107 3451
rect 18049 3411 18107 3417
rect 12676 3352 12721 3380
rect 15488 3352 17264 3380
rect 12676 3340 12682 3352
rect 0 3290 18860 3312
rect 0 3238 4660 3290
rect 4712 3238 4724 3290
rect 4776 3238 4788 3290
rect 4840 3238 4852 3290
rect 4904 3238 4916 3290
rect 4968 3238 7760 3290
rect 7812 3238 7824 3290
rect 7876 3238 7888 3290
rect 7940 3238 7952 3290
rect 8004 3238 8016 3290
rect 8068 3238 10860 3290
rect 10912 3238 10924 3290
rect 10976 3238 10988 3290
rect 11040 3238 11052 3290
rect 11104 3238 11116 3290
rect 11168 3238 13960 3290
rect 14012 3238 14024 3290
rect 14076 3238 14088 3290
rect 14140 3238 14152 3290
rect 14204 3238 14216 3290
rect 14268 3238 17060 3290
rect 17112 3238 17124 3290
rect 17176 3238 17188 3290
rect 17240 3238 17252 3290
rect 17304 3238 17316 3290
rect 17368 3238 18860 3290
rect 0 3216 18860 3238
rect 1946 3176 1952 3188
rect 1780 3148 1952 3176
rect 1780 3094 1808 3148
rect 1946 3136 1952 3148
rect 2004 3176 2010 3188
rect 2225 3179 2283 3185
rect 2225 3176 2237 3179
rect 2004 3148 2237 3176
rect 2004 3136 2010 3148
rect 2225 3145 2237 3148
rect 2271 3176 2283 3179
rect 2498 3176 2504 3188
rect 2271 3148 2504 3176
rect 2271 3145 2283 3148
rect 2225 3139 2283 3145
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 3145 3179 3203 3185
rect 3145 3145 3157 3179
rect 3191 3176 3203 3179
rect 3697 3179 3755 3185
rect 3697 3176 3709 3179
rect 3191 3148 3709 3176
rect 3191 3145 3203 3148
rect 3145 3139 3203 3145
rect 3697 3145 3709 3148
rect 3743 3145 3755 3179
rect 3697 3139 3755 3145
rect 5537 3179 5595 3185
rect 5537 3145 5549 3179
rect 5583 3176 5595 3179
rect 5629 3179 5687 3185
rect 5629 3176 5641 3179
rect 5583 3148 5641 3176
rect 5583 3145 5595 3148
rect 5537 3139 5595 3145
rect 5629 3145 5641 3148
rect 5675 3145 5687 3179
rect 5629 3139 5687 3145
rect 5718 3136 5724 3188
rect 5776 3176 5782 3188
rect 6733 3179 6791 3185
rect 5776 3148 6132 3176
rect 5776 3136 5782 3148
rect 5258 3108 5264 3120
rect 5219 3080 5264 3108
rect 5258 3068 5264 3080
rect 5316 3068 5322 3120
rect 5442 3108 5448 3120
rect 5403 3080 5448 3108
rect 5442 3068 5448 3080
rect 5500 3068 5506 3120
rect 6104 3108 6132 3148
rect 6733 3145 6745 3179
rect 6779 3176 6791 3179
rect 7285 3179 7343 3185
rect 7285 3176 7297 3179
rect 6779 3148 7297 3176
rect 6779 3145 6791 3148
rect 6733 3139 6791 3145
rect 7285 3145 7297 3148
rect 7331 3145 7343 3179
rect 7285 3139 7343 3145
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7432 3148 7757 3176
rect 7432 3136 7438 3148
rect 7745 3145 7757 3148
rect 7791 3176 7803 3179
rect 8202 3176 8208 3188
rect 7791 3148 8208 3176
rect 7791 3145 7803 3148
rect 7745 3139 7803 3145
rect 8202 3136 8208 3148
rect 8260 3176 8266 3188
rect 8570 3176 8576 3188
rect 8260 3148 8576 3176
rect 8260 3136 8266 3148
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 9950 3176 9956 3188
rect 8812 3148 9956 3176
rect 8812 3136 8818 3148
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 10410 3176 10416 3188
rect 10371 3148 10416 3176
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 11790 3176 11796 3188
rect 10704 3148 11796 3176
rect 6825 3111 6883 3117
rect 6825 3108 6837 3111
rect 6104 3080 6837 3108
rect 6825 3077 6837 3080
rect 6871 3108 6883 3111
rect 6914 3108 6920 3120
rect 6871 3080 6920 3108
rect 6871 3077 6883 3080
rect 6825 3071 6883 3077
rect 6914 3068 6920 3080
rect 6972 3068 6978 3120
rect 7190 3068 7196 3120
rect 7248 3108 7254 3120
rect 8938 3108 8944 3120
rect 7248 3080 8944 3108
rect 7248 3068 7254 3080
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 10060 3080 10364 3108
rect 290 3040 296 3052
rect 251 3012 296 3040
rect 290 3000 296 3012
rect 348 3000 354 3052
rect 2038 3000 2044 3052
rect 2096 3040 2102 3052
rect 2777 3043 2835 3049
rect 2777 3040 2789 3043
rect 2096 3012 2789 3040
rect 2096 3000 2102 3012
rect 2777 3009 2789 3012
rect 2823 3009 2835 3043
rect 2777 3003 2835 3009
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3040 3663 3043
rect 5537 3043 5595 3049
rect 3651 3012 5488 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 566 2972 572 2984
rect 527 2944 572 2972
rect 566 2932 572 2944
rect 624 2932 630 2984
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 2685 2975 2743 2981
rect 2685 2972 2697 2975
rect 2648 2944 2697 2972
rect 2648 2932 2654 2944
rect 2685 2941 2697 2944
rect 2731 2941 2743 2975
rect 2685 2935 2743 2941
rect 3142 2932 3148 2984
rect 3200 2972 3206 2984
rect 3789 2975 3847 2981
rect 3789 2972 3801 2975
rect 3200 2944 3801 2972
rect 3200 2932 3206 2944
rect 3789 2941 3801 2944
rect 3835 2941 3847 2975
rect 5460 2972 5488 3012
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 5902 3040 5908 3052
rect 5583 3012 5908 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 5902 3000 5908 3012
rect 5960 3040 5966 3052
rect 7208 3040 7236 3068
rect 5960 3012 7236 3040
rect 7653 3043 7711 3049
rect 5960 3000 5966 3012
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 7699 3012 8125 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8294 3040 8300 3052
rect 8255 3012 8300 3040
rect 8113 3003 8171 3009
rect 8294 3000 8300 3012
rect 8352 3040 8358 3052
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 8352 3012 8861 3040
rect 8352 3000 8358 3012
rect 8849 3009 8861 3012
rect 8895 3009 8907 3043
rect 8849 3003 8907 3009
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9398 3040 9404 3052
rect 9079 3012 9404 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 10060 3049 10088 3080
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 9646 3012 10057 3040
rect 5997 2975 6055 2981
rect 5460 2944 5948 2972
rect 3789 2935 3847 2941
rect 5920 2916 5948 2944
rect 5997 2941 6009 2975
rect 6043 2941 6055 2975
rect 5997 2935 6055 2941
rect 2866 2864 2872 2916
rect 2924 2904 2930 2916
rect 3237 2907 3295 2913
rect 3237 2904 3249 2907
rect 2924 2876 3249 2904
rect 2924 2864 2930 2876
rect 3237 2873 3249 2876
rect 3283 2873 3295 2907
rect 3237 2867 3295 2873
rect 3510 2864 3516 2916
rect 3568 2904 3574 2916
rect 5718 2904 5724 2916
rect 3568 2876 5724 2904
rect 3568 2864 3574 2876
rect 5718 2864 5724 2876
rect 5776 2864 5782 2916
rect 5902 2864 5908 2916
rect 5960 2864 5966 2916
rect 6012 2904 6040 2935
rect 6086 2932 6092 2984
rect 6144 2972 6150 2984
rect 6144 2944 6776 2972
rect 6144 2932 6150 2944
rect 6365 2907 6423 2913
rect 6365 2904 6377 2907
rect 6012 2876 6377 2904
rect 6365 2873 6377 2876
rect 6411 2873 6423 2907
rect 6748 2904 6776 2944
rect 6822 2932 6828 2984
rect 6880 2972 6886 2984
rect 7009 2975 7067 2981
rect 7009 2972 7021 2975
rect 6880 2944 7021 2972
rect 6880 2932 6886 2944
rect 7009 2941 7021 2944
rect 7055 2972 7067 2975
rect 7929 2975 7987 2981
rect 7055 2944 7880 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 6748 2876 6868 2904
rect 6365 2867 6423 2873
rect 6840 2848 6868 2876
rect 2038 2836 2044 2848
rect 1999 2808 2044 2836
rect 2038 2796 2044 2808
rect 2096 2796 2102 2848
rect 5626 2796 5632 2848
rect 5684 2836 5690 2848
rect 6273 2839 6331 2845
rect 6273 2836 6285 2839
rect 5684 2808 6285 2836
rect 5684 2796 5690 2808
rect 6273 2805 6285 2808
rect 6319 2805 6331 2839
rect 6273 2799 6331 2805
rect 6822 2796 6828 2848
rect 6880 2836 6886 2848
rect 7466 2836 7472 2848
rect 6880 2808 7472 2836
rect 6880 2796 6886 2808
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 7852 2836 7880 2944
rect 7929 2941 7941 2975
rect 7975 2941 7987 2975
rect 7929 2935 7987 2941
rect 8941 2975 8999 2981
rect 8941 2941 8953 2975
rect 8987 2972 8999 2975
rect 9646 2972 9674 3012
rect 10045 3009 10057 3012
rect 10091 3009 10103 3043
rect 10226 3040 10232 3052
rect 10187 3012 10232 3040
rect 10045 3003 10103 3009
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 8987 2944 9674 2972
rect 8987 2941 8999 2944
rect 8941 2935 8999 2941
rect 7944 2904 7972 2935
rect 10244 2904 10272 3000
rect 7944 2876 10272 2904
rect 10336 2904 10364 3080
rect 10594 3040 10600 3052
rect 10555 3012 10600 3040
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 10704 3049 10732 3148
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 12069 3179 12127 3185
rect 12069 3176 12081 3179
rect 11940 3148 12081 3176
rect 11940 3136 11946 3148
rect 12069 3145 12081 3148
rect 12115 3145 12127 3179
rect 12069 3139 12127 3145
rect 13538 3136 13544 3188
rect 13596 3176 13602 3188
rect 13596 3148 15148 3176
rect 13596 3136 13602 3148
rect 11330 3068 11336 3120
rect 11388 3108 11394 3120
rect 12529 3111 12587 3117
rect 11388 3080 11928 3108
rect 11388 3068 11394 3080
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 10778 3000 10784 3052
rect 10836 3040 10842 3052
rect 11146 3040 11152 3052
rect 10836 3012 10881 3040
rect 11107 3012 11152 3040
rect 10836 3000 10842 3012
rect 11146 3000 11152 3012
rect 11204 3000 11210 3052
rect 11422 3040 11428 3052
rect 11383 3012 11428 3040
rect 11422 3000 11428 3012
rect 11480 3000 11486 3052
rect 11900 3049 11928 3080
rect 12529 3077 12541 3111
rect 12575 3108 12587 3111
rect 12618 3108 12624 3120
rect 12575 3080 12624 3108
rect 12575 3077 12587 3080
rect 12529 3071 12587 3077
rect 12618 3068 12624 3080
rect 12676 3068 12682 3120
rect 14550 3068 14556 3120
rect 14608 3108 14614 3120
rect 14706 3111 14764 3117
rect 14706 3108 14718 3111
rect 14608 3080 14718 3108
rect 14608 3068 14614 3080
rect 14706 3077 14718 3080
rect 14752 3077 14764 3111
rect 14706 3071 14764 3077
rect 11885 3043 11943 3049
rect 11885 3009 11897 3043
rect 11931 3009 11943 3043
rect 12250 3040 12256 3052
rect 12211 3012 12256 3040
rect 11885 3003 11943 3009
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 13630 3000 13636 3052
rect 13688 3000 13694 3052
rect 13814 3000 13820 3052
rect 13872 3040 13878 3052
rect 14458 3040 14464 3052
rect 13872 3012 14464 3040
rect 13872 3000 13878 3012
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 15120 3040 15148 3148
rect 15378 3136 15384 3188
rect 15436 3176 15442 3188
rect 15841 3179 15899 3185
rect 15841 3176 15853 3179
rect 15436 3148 15853 3176
rect 15436 3136 15442 3148
rect 15841 3145 15853 3148
rect 15887 3145 15899 3179
rect 15841 3139 15899 3145
rect 15930 3136 15936 3188
rect 15988 3176 15994 3188
rect 15988 3148 16033 3176
rect 15988 3136 15994 3148
rect 15194 3068 15200 3120
rect 15252 3108 15258 3120
rect 16482 3108 16488 3120
rect 15252 3080 16488 3108
rect 15252 3068 15258 3080
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 16393 3043 16451 3049
rect 16393 3040 16405 3043
rect 15120 3012 16405 3040
rect 16393 3009 16405 3012
rect 16439 3040 16451 3043
rect 17494 3040 17500 3052
rect 16439 3012 17500 3040
rect 16439 3009 16451 3012
rect 16393 3003 16451 3009
rect 17494 3000 17500 3012
rect 17552 3040 17558 3052
rect 17862 3040 17868 3052
rect 17552 3012 17868 3040
rect 17552 3000 17558 3012
rect 17862 3000 17868 3012
rect 17920 3000 17926 3052
rect 11698 2972 11704 2984
rect 11659 2944 11704 2972
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 10778 2904 10784 2916
rect 10336 2876 10784 2904
rect 10778 2864 10784 2876
rect 10836 2864 10842 2916
rect 9858 2836 9864 2848
rect 7852 2808 9864 2836
rect 9858 2796 9864 2808
rect 9916 2796 9922 2848
rect 12268 2836 12296 3000
rect 14274 2972 14280 2984
rect 14235 2944 14280 2972
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 13814 2836 13820 2848
rect 12268 2808 13820 2836
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 15102 2796 15108 2848
rect 15160 2836 15166 2848
rect 16117 2839 16175 2845
rect 16117 2836 16129 2839
rect 15160 2808 16129 2836
rect 15160 2796 15166 2808
rect 16117 2805 16129 2808
rect 16163 2805 16175 2839
rect 16117 2799 16175 2805
rect 0 2746 18860 2768
rect 0 2694 3110 2746
rect 3162 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 6210 2746
rect 6262 2694 6274 2746
rect 6326 2694 6338 2746
rect 6390 2694 6402 2746
rect 6454 2694 6466 2746
rect 6518 2694 9310 2746
rect 9362 2694 9374 2746
rect 9426 2694 9438 2746
rect 9490 2694 9502 2746
rect 9554 2694 9566 2746
rect 9618 2694 12410 2746
rect 12462 2694 12474 2746
rect 12526 2694 12538 2746
rect 12590 2694 12602 2746
rect 12654 2694 12666 2746
rect 12718 2694 15510 2746
rect 15562 2694 15574 2746
rect 15626 2694 15638 2746
rect 15690 2694 15702 2746
rect 15754 2694 15766 2746
rect 15818 2694 18860 2746
rect 0 2672 18860 2694
rect 566 2592 572 2644
rect 624 2632 630 2644
rect 753 2635 811 2641
rect 753 2632 765 2635
rect 624 2604 765 2632
rect 624 2592 630 2604
rect 753 2601 765 2604
rect 799 2601 811 2635
rect 753 2595 811 2601
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 3145 2635 3203 2641
rect 2832 2604 2877 2632
rect 2832 2592 2838 2604
rect 3145 2601 3157 2635
rect 3191 2632 3203 2635
rect 3329 2635 3387 2641
rect 3329 2632 3341 2635
rect 3191 2604 3341 2632
rect 3191 2601 3203 2604
rect 3145 2595 3203 2601
rect 3329 2601 3341 2604
rect 3375 2632 3387 2635
rect 3510 2632 3516 2644
rect 3375 2604 3516 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 5442 2632 5448 2644
rect 4203 2604 5448 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 7101 2635 7159 2641
rect 7101 2601 7113 2635
rect 7147 2632 7159 2635
rect 7190 2632 7196 2644
rect 7147 2604 7196 2632
rect 7147 2601 7159 2604
rect 7101 2595 7159 2601
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 11057 2635 11115 2641
rect 11057 2601 11069 2635
rect 11103 2632 11115 2635
rect 11238 2632 11244 2644
rect 11103 2604 11244 2632
rect 11103 2601 11115 2604
rect 11057 2595 11115 2601
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 2593 2567 2651 2573
rect 2593 2564 2605 2567
rect 2056 2536 2605 2564
rect 2056 2508 2084 2536
rect 2593 2533 2605 2536
rect 2639 2533 2651 2567
rect 8754 2564 8760 2576
rect 8715 2536 8760 2564
rect 2593 2527 2651 2533
rect 2038 2496 2044 2508
rect 1999 2468 2044 2496
rect 2038 2456 2044 2468
rect 2096 2456 2102 2508
rect 2222 2496 2228 2508
rect 2183 2468 2228 2496
rect 2222 2456 2228 2468
rect 2280 2496 2286 2508
rect 2409 2499 2467 2505
rect 2409 2496 2421 2499
rect 2280 2468 2421 2496
rect 2280 2456 2286 2468
rect 2409 2465 2421 2468
rect 2455 2465 2467 2499
rect 2608 2496 2636 2527
rect 8754 2524 8760 2536
rect 8812 2524 8818 2576
rect 10594 2524 10600 2576
rect 10652 2564 10658 2576
rect 11333 2567 11391 2573
rect 11333 2564 11345 2567
rect 10652 2536 11345 2564
rect 10652 2524 10658 2536
rect 11333 2533 11345 2536
rect 11379 2564 11391 2567
rect 11517 2567 11575 2573
rect 11517 2564 11529 2567
rect 11379 2536 11529 2564
rect 11379 2533 11391 2536
rect 11333 2527 11391 2533
rect 11517 2533 11529 2536
rect 11563 2533 11575 2567
rect 11517 2527 11575 2533
rect 15286 2524 15292 2576
rect 15344 2564 15350 2576
rect 15657 2567 15715 2573
rect 15657 2564 15669 2567
rect 15344 2536 15669 2564
rect 15344 2524 15350 2536
rect 15657 2533 15669 2536
rect 15703 2533 15715 2567
rect 15657 2527 15715 2533
rect 2608 2468 2820 2496
rect 2409 2459 2467 2465
rect 937 2431 995 2437
rect 937 2397 949 2431
rect 983 2428 995 2431
rect 983 2400 1624 2428
rect 983 2397 995 2400
rect 937 2391 995 2397
rect 1596 2301 1624 2400
rect 2590 2388 2596 2440
rect 2648 2428 2654 2440
rect 2792 2437 2820 2468
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 5905 2499 5963 2505
rect 5905 2496 5917 2499
rect 5592 2468 5917 2496
rect 5592 2456 5598 2468
rect 5905 2465 5917 2468
rect 5951 2465 5963 2499
rect 5905 2459 5963 2465
rect 8849 2499 8907 2505
rect 8849 2465 8861 2499
rect 8895 2496 8907 2499
rect 9674 2496 9680 2508
rect 8895 2468 9680 2496
rect 8895 2465 8907 2468
rect 8849 2459 8907 2465
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 10778 2456 10784 2508
rect 10836 2496 10842 2508
rect 10836 2468 11100 2496
rect 10836 2456 10842 2468
rect 2685 2431 2743 2437
rect 2685 2428 2697 2431
rect 2648 2400 2697 2428
rect 2648 2388 2654 2400
rect 2685 2397 2697 2400
rect 2731 2397 2743 2431
rect 2685 2391 2743 2397
rect 2777 2431 2835 2437
rect 2777 2397 2789 2431
rect 2823 2397 2835 2431
rect 2958 2428 2964 2440
rect 2919 2400 2964 2428
rect 2777 2391 2835 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 6086 2388 6092 2440
rect 6144 2428 6150 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 6144 2400 6377 2428
rect 6144 2388 6150 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 9217 2431 9275 2437
rect 9217 2428 9229 2431
rect 6365 2391 6423 2397
rect 8956 2400 9229 2428
rect 1949 2363 2007 2369
rect 1949 2329 1961 2363
rect 1995 2360 2007 2363
rect 2866 2360 2872 2372
rect 1995 2332 2872 2360
rect 1995 2329 2007 2332
rect 1949 2323 2007 2329
rect 2866 2320 2872 2332
rect 2924 2320 2930 2372
rect 3973 2363 4031 2369
rect 3973 2329 3985 2363
rect 4019 2360 4031 2363
rect 4338 2360 4344 2372
rect 4019 2332 4344 2360
rect 4019 2329 4031 2332
rect 3973 2323 4031 2329
rect 4338 2320 4344 2332
rect 4396 2360 4402 2372
rect 5626 2360 5632 2372
rect 4396 2332 4462 2360
rect 5587 2332 5632 2360
rect 4396 2320 4402 2332
rect 5626 2320 5632 2332
rect 5684 2320 5690 2372
rect 7193 2363 7251 2369
rect 7193 2329 7205 2363
rect 7239 2360 7251 2363
rect 7466 2360 7472 2372
rect 7239 2332 7472 2360
rect 7239 2329 7251 2332
rect 7193 2323 7251 2329
rect 7466 2320 7472 2332
rect 7524 2320 7530 2372
rect 8570 2360 8576 2372
rect 8531 2332 8576 2360
rect 8570 2320 8576 2332
rect 8628 2320 8634 2372
rect 1581 2295 1639 2301
rect 1581 2261 1593 2295
rect 1627 2261 1639 2295
rect 1581 2255 1639 2261
rect 2685 2295 2743 2301
rect 2685 2261 2697 2295
rect 2731 2292 2743 2295
rect 2774 2292 2780 2304
rect 2731 2264 2780 2292
rect 2731 2261 2743 2264
rect 2685 2255 2743 2261
rect 2774 2252 2780 2264
rect 2832 2252 2838 2304
rect 4982 2252 4988 2304
rect 5040 2292 5046 2304
rect 6181 2295 6239 2301
rect 6181 2292 6193 2295
rect 5040 2264 6193 2292
rect 5040 2252 5046 2264
rect 6181 2261 6193 2264
rect 6227 2261 6239 2295
rect 8294 2292 8300 2304
rect 8255 2264 8300 2292
rect 6181 2255 6239 2261
rect 8294 2252 8300 2264
rect 8352 2252 8358 2304
rect 8956 2292 8984 2400
rect 9217 2397 9229 2400
rect 9263 2397 9275 2431
rect 10870 2428 10876 2440
rect 10831 2400 10876 2428
rect 9217 2391 9275 2397
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 11072 2437 11100 2468
rect 12802 2456 12808 2508
rect 12860 2496 12866 2508
rect 14274 2496 14280 2508
rect 12860 2468 14280 2496
rect 12860 2456 12866 2468
rect 14274 2456 14280 2468
rect 14332 2496 14338 2508
rect 15197 2499 15255 2505
rect 15197 2496 15209 2499
rect 14332 2468 15209 2496
rect 14332 2456 14338 2468
rect 15197 2465 15209 2468
rect 15243 2496 15255 2499
rect 15562 2496 15568 2508
rect 15243 2468 15568 2496
rect 15243 2465 15255 2468
rect 15197 2459 15255 2465
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 15838 2496 15844 2508
rect 15799 2468 15844 2496
rect 15838 2456 15844 2468
rect 15896 2456 15902 2508
rect 16482 2456 16488 2508
rect 16540 2496 16546 2508
rect 17865 2499 17923 2505
rect 17865 2496 17877 2499
rect 16540 2468 17877 2496
rect 16540 2456 16546 2468
rect 17865 2465 17877 2468
rect 17911 2465 17923 2499
rect 17865 2459 17923 2465
rect 11057 2431 11115 2437
rect 11057 2397 11069 2431
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 11425 2431 11483 2437
rect 11425 2397 11437 2431
rect 11471 2397 11483 2431
rect 11425 2391 11483 2397
rect 10643 2363 10701 2369
rect 9766 2292 9772 2304
rect 8956 2264 9772 2292
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 10134 2252 10140 2304
rect 10192 2292 10198 2304
rect 10244 2292 10272 2346
rect 10643 2329 10655 2363
rect 10689 2360 10701 2363
rect 11238 2360 11244 2372
rect 10689 2332 11244 2360
rect 10689 2329 10701 2332
rect 10643 2323 10701 2329
rect 11238 2320 11244 2332
rect 11296 2360 11302 2372
rect 11440 2360 11468 2391
rect 14550 2388 14556 2440
rect 14608 2428 14614 2440
rect 15013 2431 15071 2437
rect 15013 2428 15025 2431
rect 14608 2400 15025 2428
rect 14608 2388 14614 2400
rect 15013 2397 15025 2400
rect 15059 2428 15071 2431
rect 15381 2431 15439 2437
rect 15381 2428 15393 2431
rect 15059 2400 15393 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 15212 2372 15240 2400
rect 15381 2397 15393 2400
rect 15427 2397 15439 2431
rect 15381 2391 15439 2397
rect 11296 2332 11468 2360
rect 11296 2320 11302 2332
rect 11698 2320 11704 2372
rect 11756 2360 11762 2372
rect 11756 2332 15056 2360
rect 11756 2320 11762 2332
rect 11882 2292 11888 2304
rect 10192 2264 11888 2292
rect 10192 2252 10198 2264
rect 11882 2252 11888 2264
rect 11940 2252 11946 2304
rect 12710 2252 12716 2304
rect 12768 2292 12774 2304
rect 13630 2292 13636 2304
rect 12768 2264 13636 2292
rect 12768 2252 12774 2264
rect 13630 2252 13636 2264
rect 13688 2252 13694 2304
rect 14366 2252 14372 2304
rect 14424 2292 14430 2304
rect 14553 2295 14611 2301
rect 14553 2292 14565 2295
rect 14424 2264 14565 2292
rect 14424 2252 14430 2264
rect 14553 2261 14565 2264
rect 14599 2261 14611 2295
rect 14918 2292 14924 2304
rect 14879 2264 14924 2292
rect 14553 2255 14611 2261
rect 14918 2252 14924 2264
rect 14976 2252 14982 2304
rect 15028 2292 15056 2332
rect 15194 2320 15200 2372
rect 15252 2320 15258 2372
rect 15286 2320 15292 2372
rect 15344 2360 15350 2372
rect 15856 2360 15884 2456
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 18506 2428 18512 2440
rect 18279 2400 18512 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 18506 2388 18512 2400
rect 18564 2388 18570 2440
rect 16114 2360 16120 2372
rect 15344 2332 15884 2360
rect 16075 2332 16120 2360
rect 15344 2320 15350 2332
rect 16114 2320 16120 2332
rect 16172 2320 16178 2372
rect 16666 2320 16672 2372
rect 16724 2320 16730 2372
rect 17972 2332 18368 2360
rect 15304 2292 15332 2320
rect 15028 2264 15332 2292
rect 15838 2252 15844 2304
rect 15896 2292 15902 2304
rect 17972 2292 18000 2332
rect 18340 2301 18368 2332
rect 15896 2264 18000 2292
rect 18325 2295 18383 2301
rect 15896 2252 15902 2264
rect 18325 2261 18337 2295
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 0 2202 18860 2224
rect 0 2150 4660 2202
rect 4712 2150 4724 2202
rect 4776 2150 4788 2202
rect 4840 2150 4852 2202
rect 4904 2150 4916 2202
rect 4968 2150 7760 2202
rect 7812 2150 7824 2202
rect 7876 2150 7888 2202
rect 7940 2150 7952 2202
rect 8004 2150 8016 2202
rect 8068 2150 10860 2202
rect 10912 2150 10924 2202
rect 10976 2150 10988 2202
rect 11040 2150 11052 2202
rect 11104 2150 11116 2202
rect 11168 2150 13960 2202
rect 14012 2150 14024 2202
rect 14076 2150 14088 2202
rect 14140 2150 14152 2202
rect 14204 2150 14216 2202
rect 14268 2150 17060 2202
rect 17112 2150 17124 2202
rect 17176 2150 17188 2202
rect 17240 2150 17252 2202
rect 17304 2150 17316 2202
rect 17368 2150 18860 2202
rect 0 2128 18860 2150
rect 2041 2091 2099 2097
rect 2041 2057 2053 2091
rect 2087 2057 2099 2091
rect 9125 2091 9183 2097
rect 9125 2088 9137 2091
rect 2041 2051 2099 2057
rect 5920 2060 9137 2088
rect 1946 2020 1952 2032
rect 1794 1992 1952 2020
rect 1946 1980 1952 1992
rect 2004 1980 2010 2032
rect 2056 1952 2084 2051
rect 5534 2020 5540 2032
rect 3528 1992 5540 2020
rect 2869 1955 2927 1961
rect 2869 1952 2881 1955
rect 2056 1924 2881 1952
rect 2869 1921 2881 1924
rect 2915 1952 2927 1955
rect 2958 1952 2964 1964
rect 2915 1924 2964 1952
rect 2915 1921 2927 1924
rect 2869 1915 2927 1921
rect 2958 1912 2964 1924
rect 3016 1912 3022 1964
rect 3528 1961 3556 1992
rect 5534 1980 5540 1992
rect 5592 1980 5598 2032
rect 3513 1955 3571 1961
rect 3513 1921 3525 1955
rect 3559 1921 3571 1955
rect 3513 1915 3571 1921
rect 3697 1955 3755 1961
rect 3697 1921 3709 1955
rect 3743 1952 3755 1955
rect 4338 1952 4344 1964
rect 3743 1924 4344 1952
rect 3743 1921 3755 1924
rect 3697 1915 3755 1921
rect 290 1884 296 1896
rect 203 1856 296 1884
rect 290 1844 296 1856
rect 348 1844 354 1896
rect 569 1887 627 1893
rect 569 1853 581 1887
rect 615 1884 627 1887
rect 2501 1887 2559 1893
rect 2501 1884 2513 1887
rect 615 1856 2513 1884
rect 615 1853 627 1856
rect 569 1847 627 1853
rect 2501 1853 2513 1856
rect 2547 1853 2559 1887
rect 2501 1847 2559 1853
rect 2774 1844 2780 1896
rect 2832 1884 2838 1896
rect 2832 1856 2877 1884
rect 2832 1844 2838 1856
rect 308 1748 336 1844
rect 1762 1776 1768 1828
rect 1820 1816 1826 1828
rect 3528 1816 3556 1915
rect 4338 1912 4344 1924
rect 4396 1912 4402 1964
rect 4709 1955 4767 1961
rect 4709 1921 4721 1955
rect 4755 1952 4767 1955
rect 4982 1952 4988 1964
rect 4755 1924 4988 1952
rect 4755 1921 4767 1924
rect 4709 1915 4767 1921
rect 3973 1887 4031 1893
rect 3973 1853 3985 1887
rect 4019 1884 4031 1887
rect 4062 1884 4068 1896
rect 4019 1856 4068 1884
rect 4019 1853 4031 1856
rect 3973 1847 4031 1853
rect 4062 1844 4068 1856
rect 4120 1844 4126 1896
rect 1820 1788 3556 1816
rect 4341 1819 4399 1825
rect 1820 1776 1826 1788
rect 4341 1785 4353 1819
rect 4387 1816 4399 1819
rect 4724 1816 4752 1915
rect 4982 1912 4988 1924
rect 5040 1912 5046 1964
rect 5074 1912 5080 1964
rect 5132 1952 5138 1964
rect 5261 1955 5319 1961
rect 5261 1952 5273 1955
rect 5132 1924 5273 1952
rect 5132 1912 5138 1924
rect 5261 1921 5273 1924
rect 5307 1921 5319 1955
rect 5261 1915 5319 1921
rect 5353 1955 5411 1961
rect 5353 1921 5365 1955
rect 5399 1921 5411 1955
rect 5353 1915 5411 1921
rect 5368 1884 5396 1915
rect 5442 1912 5448 1964
rect 5500 1952 5506 1964
rect 5920 1952 5948 2060
rect 6086 2020 6092 2032
rect 6047 1992 6092 2020
rect 6086 1980 6092 1992
rect 6144 1980 6150 2032
rect 7484 2020 7512 2060
rect 9125 2057 9137 2060
rect 9171 2088 9183 2091
rect 9950 2088 9956 2100
rect 9171 2060 9956 2088
rect 9171 2057 9183 2060
rect 9125 2051 9183 2057
rect 9950 2048 9956 2060
rect 10008 2048 10014 2100
rect 11422 2088 11428 2100
rect 11383 2060 11428 2088
rect 11422 2048 11428 2060
rect 11480 2048 11486 2100
rect 12069 2091 12127 2097
rect 12069 2057 12081 2091
rect 12115 2088 12127 2091
rect 12253 2091 12311 2097
rect 12253 2088 12265 2091
rect 12115 2060 12265 2088
rect 12115 2057 12127 2060
rect 12069 2051 12127 2057
rect 12253 2057 12265 2060
rect 12299 2057 12311 2091
rect 12253 2051 12311 2057
rect 12621 2091 12679 2097
rect 12621 2057 12633 2091
rect 12667 2088 12679 2091
rect 13081 2091 13139 2097
rect 13081 2088 13093 2091
rect 12667 2060 13093 2088
rect 12667 2057 12679 2060
rect 12621 2051 12679 2057
rect 13081 2057 13093 2060
rect 13127 2057 13139 2091
rect 13081 2051 13139 2057
rect 13541 2091 13599 2097
rect 13541 2057 13553 2091
rect 13587 2088 13599 2091
rect 13630 2088 13636 2100
rect 13587 2060 13636 2088
rect 13587 2057 13599 2060
rect 13541 2051 13599 2057
rect 13630 2048 13636 2060
rect 13688 2048 13694 2100
rect 15838 2088 15844 2100
rect 15212 2060 15844 2088
rect 9674 2020 9680 2032
rect 7484 1992 7604 2020
rect 5500 1924 5948 1952
rect 5500 1912 5506 1924
rect 6104 1884 6132 1980
rect 6549 1955 6607 1961
rect 6549 1921 6561 1955
rect 6595 1921 6607 1955
rect 6730 1952 6736 1964
rect 6691 1924 6736 1952
rect 6549 1915 6607 1921
rect 5368 1856 6132 1884
rect 6564 1884 6592 1915
rect 6730 1912 6736 1924
rect 6788 1912 6794 1964
rect 6822 1912 6828 1964
rect 6880 1952 6886 1964
rect 7285 1955 7343 1961
rect 7285 1952 7297 1955
rect 6880 1924 7297 1952
rect 6880 1912 6886 1924
rect 7285 1921 7297 1924
rect 7331 1921 7343 1955
rect 7466 1952 7472 1964
rect 7427 1924 7472 1952
rect 7285 1915 7343 1921
rect 7466 1912 7472 1924
rect 7524 1912 7530 1964
rect 7576 1961 7604 1992
rect 8956 1992 9680 2020
rect 8956 1961 8984 1992
rect 9674 1980 9680 1992
rect 9732 1980 9738 2032
rect 9766 1980 9772 2032
rect 9824 2020 9830 2032
rect 15212 2029 15240 2060
rect 15838 2048 15844 2060
rect 15896 2048 15902 2100
rect 16114 2048 16120 2100
rect 16172 2088 16178 2100
rect 16669 2091 16727 2097
rect 16669 2088 16681 2091
rect 16172 2060 16681 2088
rect 16172 2048 16178 2060
rect 16669 2057 16681 2060
rect 16715 2057 16727 2091
rect 16669 2051 16727 2057
rect 17313 2091 17371 2097
rect 17313 2057 17325 2091
rect 17359 2088 17371 2091
rect 17494 2088 17500 2100
rect 17359 2060 17500 2088
rect 17359 2057 17371 2060
rect 17313 2051 17371 2057
rect 17494 2048 17500 2060
rect 17552 2088 17558 2100
rect 17862 2088 17868 2100
rect 17552 2060 17868 2088
rect 17552 2048 17558 2060
rect 17862 2048 17868 2060
rect 17920 2048 17926 2100
rect 18138 2088 18144 2100
rect 18099 2060 18144 2088
rect 18138 2048 18144 2060
rect 18196 2048 18202 2100
rect 10045 2023 10103 2029
rect 9824 1992 9869 2020
rect 9824 1980 9830 1992
rect 10045 1989 10057 2023
rect 10091 2020 10103 2023
rect 15197 2023 15255 2029
rect 10091 1992 14136 2020
rect 10091 1989 10103 1992
rect 10045 1983 10103 1989
rect 7561 1955 7619 1961
rect 7561 1921 7573 1955
rect 7607 1921 7619 1955
rect 7561 1915 7619 1921
rect 8941 1955 8999 1961
rect 8941 1921 8953 1955
rect 8987 1921 8999 1955
rect 8941 1915 8999 1921
rect 9217 1955 9275 1961
rect 9217 1921 9229 1955
rect 9263 1952 9275 1955
rect 9263 1924 9674 1952
rect 9853 1945 9911 1951
rect 9853 1942 9865 1945
rect 9263 1921 9275 1924
rect 9217 1915 9275 1921
rect 7374 1884 7380 1896
rect 6564 1856 7380 1884
rect 7374 1844 7380 1856
rect 7432 1844 7438 1896
rect 8570 1844 8576 1896
rect 8628 1884 8634 1896
rect 9232 1884 9260 1915
rect 8628 1856 9260 1884
rect 9646 1896 9674 1924
rect 9784 1914 9865 1942
rect 9646 1856 9680 1896
rect 8628 1844 8634 1856
rect 9674 1844 9680 1856
rect 9732 1844 9738 1896
rect 4387 1788 4752 1816
rect 4387 1785 4399 1788
rect 4341 1779 4399 1785
rect 8294 1776 8300 1828
rect 8352 1816 8358 1828
rect 8389 1819 8447 1825
rect 8389 1816 8401 1819
rect 8352 1788 8401 1816
rect 8352 1776 8358 1788
rect 8389 1785 8401 1788
rect 8435 1816 8447 1819
rect 9784 1816 9812 1914
rect 9853 1911 9865 1914
rect 9899 1911 9911 1945
rect 9950 1912 9956 1964
rect 10008 1952 10014 1964
rect 10137 1955 10195 1961
rect 10008 1924 10053 1952
rect 10008 1912 10014 1924
rect 10137 1921 10149 1955
rect 10183 1952 10195 1955
rect 10226 1952 10232 1964
rect 10183 1924 10232 1952
rect 10183 1921 10195 1924
rect 10137 1915 10195 1921
rect 10226 1912 10232 1924
rect 10284 1912 10290 1964
rect 11057 1955 11115 1961
rect 11057 1921 11069 1955
rect 11103 1952 11115 1955
rect 11238 1952 11244 1964
rect 11103 1924 11244 1952
rect 11103 1921 11115 1924
rect 11057 1915 11115 1921
rect 11238 1912 11244 1924
rect 11296 1912 11302 1964
rect 11716 1961 11744 1992
rect 11701 1955 11759 1961
rect 11701 1921 11713 1955
rect 11747 1921 11759 1955
rect 11701 1915 11759 1921
rect 11885 1955 11943 1961
rect 11885 1921 11897 1955
rect 11931 1952 11943 1955
rect 12069 1955 12127 1961
rect 12069 1952 12081 1955
rect 11931 1924 12081 1952
rect 11931 1921 11943 1924
rect 11885 1915 11943 1921
rect 12069 1921 12081 1924
rect 12115 1921 12127 1955
rect 12710 1952 12716 1964
rect 12671 1924 12716 1952
rect 12069 1915 12127 1921
rect 12710 1912 12716 1924
rect 12768 1912 12774 1964
rect 12894 1912 12900 1964
rect 12952 1952 12958 1964
rect 13449 1955 13507 1961
rect 13449 1952 13461 1955
rect 12952 1924 13461 1952
rect 12952 1912 12958 1924
rect 13449 1921 13461 1924
rect 13495 1921 13507 1955
rect 13449 1915 13507 1921
rect 13538 1912 13544 1964
rect 13596 1952 13602 1964
rect 14108 1961 14136 1992
rect 15197 1989 15209 2023
rect 15243 1989 15255 2023
rect 15197 1983 15255 1989
rect 13909 1955 13967 1961
rect 13909 1952 13921 1955
rect 13596 1924 13921 1952
rect 13596 1912 13602 1924
rect 13909 1921 13921 1924
rect 13955 1921 13967 1955
rect 13909 1915 13967 1921
rect 14093 1955 14151 1961
rect 14093 1921 14105 1955
rect 14139 1921 14151 1955
rect 14093 1915 14151 1921
rect 14277 1955 14335 1961
rect 14277 1921 14289 1955
rect 14323 1952 14335 1955
rect 14366 1952 14372 1964
rect 14323 1924 14372 1952
rect 14323 1921 14335 1924
rect 14277 1915 14335 1921
rect 9853 1905 9911 1911
rect 10962 1884 10968 1896
rect 10923 1856 10968 1884
rect 10962 1844 10968 1856
rect 11020 1844 11026 1896
rect 12802 1884 12808 1896
rect 12763 1856 12808 1884
rect 12802 1844 12808 1856
rect 12860 1844 12866 1896
rect 13725 1887 13783 1893
rect 13725 1853 13737 1887
rect 13771 1884 13783 1887
rect 13814 1884 13820 1896
rect 13771 1856 13820 1884
rect 13771 1853 13783 1856
rect 13725 1847 13783 1853
rect 13814 1844 13820 1856
rect 13872 1844 13878 1896
rect 9858 1816 9864 1828
rect 8435 1788 8800 1816
rect 9771 1788 9864 1816
rect 8435 1785 8447 1788
rect 8389 1779 8447 1785
rect 1780 1748 1808 1776
rect 308 1720 1808 1748
rect 1946 1708 1952 1760
rect 2004 1748 2010 1760
rect 2222 1748 2228 1760
rect 2004 1720 2228 1748
rect 2004 1708 2010 1720
rect 2222 1708 2228 1720
rect 2280 1708 2286 1760
rect 2498 1708 2504 1760
rect 2556 1748 2562 1760
rect 3237 1751 3295 1757
rect 3237 1748 3249 1751
rect 2556 1720 3249 1748
rect 2556 1708 2562 1720
rect 3237 1717 3249 1720
rect 3283 1717 3295 1751
rect 4430 1748 4436 1760
rect 4391 1720 4436 1748
rect 3237 1711 3295 1717
rect 4430 1708 4436 1720
rect 4488 1708 4494 1760
rect 4522 1708 4528 1760
rect 4580 1748 4586 1760
rect 4617 1751 4675 1757
rect 4617 1748 4629 1751
rect 4580 1720 4629 1748
rect 4580 1708 4586 1720
rect 4617 1717 4629 1720
rect 4663 1717 4675 1751
rect 4617 1711 4675 1717
rect 5166 1708 5172 1760
rect 5224 1748 5230 1760
rect 5629 1751 5687 1757
rect 5629 1748 5641 1751
rect 5224 1720 5641 1748
rect 5224 1708 5230 1720
rect 5629 1717 5641 1720
rect 5675 1717 5687 1751
rect 8662 1748 8668 1760
rect 8623 1720 8668 1748
rect 5629 1711 5687 1717
rect 8662 1708 8668 1720
rect 8720 1708 8726 1760
rect 8772 1748 8800 1788
rect 9858 1776 9864 1788
rect 9916 1816 9922 1828
rect 12820 1816 12848 1844
rect 9916 1788 12848 1816
rect 9916 1776 9922 1788
rect 10134 1748 10140 1760
rect 8772 1720 10140 1748
rect 10134 1708 10140 1720
rect 10192 1708 10198 1760
rect 11793 1751 11851 1757
rect 11793 1717 11805 1751
rect 11839 1748 11851 1751
rect 12158 1748 12164 1760
rect 11839 1720 12164 1748
rect 11839 1717 11851 1720
rect 11793 1711 11851 1717
rect 12158 1708 12164 1720
rect 12216 1708 12222 1760
rect 14108 1748 14136 1915
rect 14366 1912 14372 1924
rect 14424 1912 14430 1964
rect 14642 1912 14648 1964
rect 14700 1952 14706 1964
rect 14829 1955 14887 1961
rect 14829 1952 14841 1955
rect 14700 1924 14841 1952
rect 14700 1912 14706 1924
rect 14829 1921 14841 1924
rect 14875 1921 14887 1955
rect 16666 1952 16672 1964
rect 16330 1924 16672 1952
rect 14829 1915 14887 1921
rect 16666 1912 16672 1924
rect 16724 1912 16730 1964
rect 16942 1912 16948 1964
rect 17000 1952 17006 1964
rect 17221 1955 17279 1961
rect 17221 1952 17233 1955
rect 17000 1924 17233 1952
rect 17000 1912 17006 1924
rect 17221 1921 17233 1924
rect 17267 1921 17279 1955
rect 18230 1952 18236 1964
rect 18191 1924 18236 1952
rect 17221 1915 17279 1921
rect 18230 1912 18236 1924
rect 18288 1912 18294 1964
rect 14185 1887 14243 1893
rect 14185 1853 14197 1887
rect 14231 1884 14243 1887
rect 14553 1887 14611 1893
rect 14553 1884 14565 1887
rect 14231 1856 14565 1884
rect 14231 1853 14243 1856
rect 14185 1847 14243 1853
rect 14553 1853 14565 1856
rect 14599 1853 14611 1887
rect 14553 1847 14611 1853
rect 14921 1887 14979 1893
rect 14921 1853 14933 1887
rect 14967 1884 14979 1887
rect 15286 1884 15292 1896
rect 14967 1856 15292 1884
rect 14967 1853 14979 1856
rect 14921 1847 14979 1853
rect 15286 1844 15292 1856
rect 15344 1844 15350 1896
rect 15562 1844 15568 1896
rect 15620 1884 15626 1896
rect 17405 1887 17463 1893
rect 17405 1884 17417 1887
rect 15620 1856 17417 1884
rect 15620 1844 15626 1856
rect 17405 1853 17417 1856
rect 17451 1853 17463 1887
rect 17405 1847 17463 1853
rect 14645 1819 14703 1825
rect 14645 1785 14657 1819
rect 14691 1816 14703 1819
rect 14826 1816 14832 1828
rect 14691 1788 14832 1816
rect 14691 1785 14703 1788
rect 14645 1779 14703 1785
rect 14826 1776 14832 1788
rect 14884 1776 14890 1828
rect 16853 1819 16911 1825
rect 16853 1816 16865 1819
rect 16546 1788 16865 1816
rect 14737 1751 14795 1757
rect 14737 1748 14749 1751
rect 14108 1720 14749 1748
rect 14737 1717 14749 1720
rect 14783 1748 14795 1751
rect 15378 1748 15384 1760
rect 14783 1720 15384 1748
rect 14783 1717 14795 1720
rect 14737 1711 14795 1717
rect 15378 1708 15384 1720
rect 15436 1708 15442 1760
rect 15930 1708 15936 1760
rect 15988 1748 15994 1760
rect 16546 1748 16574 1788
rect 16853 1785 16865 1788
rect 16899 1785 16911 1819
rect 16853 1779 16911 1785
rect 15988 1720 16574 1748
rect 15988 1708 15994 1720
rect 0 1658 18860 1680
rect 0 1606 3110 1658
rect 3162 1606 3174 1658
rect 3226 1606 3238 1658
rect 3290 1606 3302 1658
rect 3354 1606 3366 1658
rect 3418 1606 6210 1658
rect 6262 1606 6274 1658
rect 6326 1606 6338 1658
rect 6390 1606 6402 1658
rect 6454 1606 6466 1658
rect 6518 1606 9310 1658
rect 9362 1606 9374 1658
rect 9426 1606 9438 1658
rect 9490 1606 9502 1658
rect 9554 1606 9566 1658
rect 9618 1606 12410 1658
rect 12462 1606 12474 1658
rect 12526 1606 12538 1658
rect 12590 1606 12602 1658
rect 12654 1606 12666 1658
rect 12718 1606 15510 1658
rect 15562 1606 15574 1658
rect 15626 1606 15638 1658
rect 15690 1606 15702 1658
rect 15754 1606 15766 1658
rect 15818 1606 18860 1658
rect 0 1584 18860 1606
rect 10134 1504 10140 1556
rect 10192 1544 10198 1556
rect 10597 1547 10655 1553
rect 10597 1544 10609 1547
rect 10192 1516 10609 1544
rect 10192 1504 10198 1516
rect 10597 1513 10609 1516
rect 10643 1513 10655 1547
rect 10597 1507 10655 1513
rect 14553 1547 14611 1553
rect 14553 1513 14565 1547
rect 14599 1544 14611 1547
rect 14642 1544 14648 1556
rect 14599 1516 14648 1544
rect 14599 1513 14611 1516
rect 14553 1507 14611 1513
rect 3513 1479 3571 1485
rect 3513 1445 3525 1479
rect 3559 1476 3571 1479
rect 4062 1476 4068 1488
rect 3559 1448 4068 1476
rect 3559 1445 3571 1448
rect 3513 1439 3571 1445
rect 3896 1417 3924 1448
rect 4062 1436 4068 1448
rect 4120 1476 4126 1488
rect 5074 1476 5080 1488
rect 4120 1448 5080 1476
rect 4120 1436 4126 1448
rect 5074 1436 5080 1448
rect 5132 1436 5138 1488
rect 7193 1479 7251 1485
rect 7193 1445 7205 1479
rect 7239 1476 7251 1479
rect 7466 1476 7472 1488
rect 7239 1448 7472 1476
rect 7239 1445 7251 1448
rect 7193 1439 7251 1445
rect 7466 1436 7472 1448
rect 7524 1436 7530 1488
rect 7929 1479 7987 1485
rect 7929 1445 7941 1479
rect 7975 1445 7987 1479
rect 7929 1439 7987 1445
rect 2041 1411 2099 1417
rect 2041 1377 2053 1411
rect 2087 1408 2099 1411
rect 3697 1411 3755 1417
rect 3697 1408 3709 1411
rect 2087 1380 3709 1408
rect 2087 1377 2099 1380
rect 2041 1371 2099 1377
rect 3697 1377 3709 1380
rect 3743 1377 3755 1411
rect 3697 1371 3755 1377
rect 3881 1411 3939 1417
rect 3881 1377 3893 1411
rect 3927 1377 3939 1411
rect 3881 1371 3939 1377
rect 3973 1411 4031 1417
rect 3973 1377 3985 1411
rect 4019 1408 4031 1411
rect 4522 1408 4528 1420
rect 4019 1380 4528 1408
rect 4019 1377 4031 1380
rect 3973 1371 4031 1377
rect 4522 1368 4528 1380
rect 4580 1408 4586 1420
rect 5169 1411 5227 1417
rect 5169 1408 5181 1411
rect 4580 1380 5181 1408
rect 4580 1368 4586 1380
rect 5169 1377 5181 1380
rect 5215 1377 5227 1411
rect 6730 1408 6736 1420
rect 5169 1371 5227 1377
rect 5644 1380 6736 1408
rect 1762 1340 1768 1352
rect 1723 1312 1768 1340
rect 1762 1300 1768 1312
rect 1820 1300 1826 1352
rect 4338 1340 4344 1352
rect 3174 1312 4344 1340
rect 4338 1300 4344 1312
rect 4396 1300 4402 1352
rect 4893 1343 4951 1349
rect 4893 1309 4905 1343
rect 4939 1309 4951 1343
rect 4893 1303 4951 1309
rect 4522 1272 4528 1284
rect 4483 1244 4528 1272
rect 4522 1232 4528 1244
rect 4580 1232 4586 1284
rect 4908 1272 4936 1303
rect 4982 1300 4988 1352
rect 5040 1340 5046 1352
rect 5644 1349 5672 1380
rect 6730 1368 6736 1380
rect 6788 1368 6794 1420
rect 5445 1343 5503 1349
rect 5445 1340 5457 1343
rect 5040 1312 5457 1340
rect 5040 1300 5046 1312
rect 5445 1309 5457 1312
rect 5491 1309 5503 1343
rect 5445 1303 5503 1309
rect 5629 1343 5687 1349
rect 5629 1309 5641 1343
rect 5675 1309 5687 1343
rect 5902 1340 5908 1352
rect 5863 1312 5908 1340
rect 5629 1303 5687 1309
rect 5902 1300 5908 1312
rect 5960 1300 5966 1352
rect 5994 1300 6000 1352
rect 6052 1340 6058 1352
rect 7006 1340 7012 1352
rect 6052 1312 7012 1340
rect 6052 1300 6058 1312
rect 7006 1300 7012 1312
rect 7064 1300 7070 1352
rect 7193 1343 7251 1349
rect 7193 1309 7205 1343
rect 7239 1309 7251 1343
rect 7193 1303 7251 1309
rect 5258 1272 5264 1284
rect 4908 1244 5264 1272
rect 5258 1232 5264 1244
rect 5316 1232 5322 1284
rect 6825 1275 6883 1281
rect 6825 1241 6837 1275
rect 6871 1241 6883 1275
rect 7208 1272 7236 1303
rect 7374 1300 7380 1352
rect 7432 1340 7438 1352
rect 7469 1343 7527 1349
rect 7469 1340 7481 1343
rect 7432 1312 7481 1340
rect 7432 1300 7438 1312
rect 7469 1309 7481 1312
rect 7515 1309 7527 1343
rect 7944 1340 7972 1439
rect 8481 1411 8539 1417
rect 8481 1377 8493 1411
rect 8527 1408 8539 1411
rect 8662 1408 8668 1420
rect 8527 1380 8668 1408
rect 8527 1377 8539 1380
rect 8481 1371 8539 1377
rect 8662 1368 8668 1380
rect 8720 1368 8726 1420
rect 8754 1368 8760 1420
rect 8812 1408 8818 1420
rect 9030 1408 9036 1420
rect 8812 1380 9036 1408
rect 8812 1368 8818 1380
rect 9030 1368 9036 1380
rect 9088 1368 9094 1420
rect 10612 1408 10640 1507
rect 14642 1504 14648 1516
rect 14700 1504 14706 1556
rect 14737 1547 14795 1553
rect 14737 1513 14749 1547
rect 14783 1544 14795 1547
rect 14918 1544 14924 1556
rect 14783 1516 14924 1544
rect 14783 1513 14795 1516
rect 14737 1507 14795 1513
rect 14918 1504 14924 1516
rect 14976 1504 14982 1556
rect 14660 1476 14688 1504
rect 15102 1476 15108 1488
rect 14660 1448 15108 1476
rect 15102 1436 15108 1448
rect 15160 1436 15166 1488
rect 10612 1380 11284 1408
rect 8570 1340 8576 1352
rect 7944 1312 8576 1340
rect 7469 1303 7527 1309
rect 8570 1300 8576 1312
rect 8628 1300 8634 1352
rect 8846 1340 8852 1352
rect 8807 1312 8852 1340
rect 8846 1300 8852 1312
rect 8904 1300 8910 1352
rect 10275 1343 10333 1349
rect 10275 1309 10287 1343
rect 10321 1340 10333 1343
rect 10410 1340 10416 1352
rect 10321 1312 10416 1340
rect 10321 1309 10333 1312
rect 10275 1303 10333 1309
rect 10410 1300 10416 1312
rect 10468 1340 10474 1352
rect 10962 1340 10968 1352
rect 10468 1312 10968 1340
rect 10468 1300 10474 1312
rect 10962 1300 10968 1312
rect 11020 1300 11026 1352
rect 11256 1326 11284 1380
rect 13814 1368 13820 1420
rect 13872 1408 13878 1420
rect 15289 1411 15347 1417
rect 15289 1408 15301 1411
rect 13872 1380 15301 1408
rect 13872 1368 13878 1380
rect 15289 1377 15301 1380
rect 15335 1377 15347 1411
rect 15289 1371 15347 1377
rect 12621 1343 12679 1349
rect 12621 1309 12633 1343
rect 12667 1309 12679 1343
rect 12621 1303 12679 1309
rect 13357 1343 13415 1349
rect 13357 1309 13369 1343
rect 13403 1340 13415 1343
rect 13446 1340 13452 1352
rect 13403 1312 13452 1340
rect 13403 1309 13415 1312
rect 13357 1303 13415 1309
rect 7558 1272 7564 1284
rect 7208 1244 7564 1272
rect 6825 1235 6883 1241
rect 4341 1207 4399 1213
rect 4341 1173 4353 1207
rect 4387 1204 4399 1207
rect 5166 1204 5172 1216
rect 4387 1176 5172 1204
rect 4387 1173 4399 1176
rect 4341 1167 4399 1173
rect 5166 1164 5172 1176
rect 5224 1164 5230 1216
rect 5350 1204 5356 1216
rect 5311 1176 5356 1204
rect 5350 1164 5356 1176
rect 5408 1164 5414 1216
rect 5810 1204 5816 1216
rect 5771 1176 5816 1204
rect 5810 1164 5816 1176
rect 5868 1164 5874 1216
rect 6840 1204 6868 1235
rect 7558 1232 7564 1244
rect 7616 1232 7622 1284
rect 10134 1272 10140 1284
rect 9890 1244 10140 1272
rect 10134 1232 10140 1244
rect 10192 1232 10198 1284
rect 12342 1272 12348 1284
rect 12303 1244 12348 1272
rect 12342 1232 12348 1244
rect 12400 1232 12406 1284
rect 12636 1272 12664 1303
rect 13446 1300 13452 1312
rect 13504 1300 13510 1352
rect 13541 1343 13599 1349
rect 13541 1309 13553 1343
rect 13587 1340 13599 1343
rect 14458 1340 14464 1352
rect 13587 1312 14464 1340
rect 13587 1309 13599 1312
rect 13541 1303 13599 1309
rect 14458 1300 14464 1312
rect 14516 1300 14522 1352
rect 15102 1340 15108 1352
rect 15063 1312 15108 1340
rect 15102 1300 15108 1312
rect 15160 1300 15166 1352
rect 15194 1300 15200 1352
rect 15252 1340 15258 1352
rect 15252 1312 15297 1340
rect 15252 1300 15258 1312
rect 15378 1300 15384 1352
rect 15436 1340 15442 1352
rect 15749 1343 15807 1349
rect 15749 1340 15761 1343
rect 15436 1312 15761 1340
rect 15436 1300 15442 1312
rect 15749 1309 15761 1312
rect 15795 1309 15807 1343
rect 15930 1340 15936 1352
rect 15891 1312 15936 1340
rect 15749 1303 15807 1309
rect 15930 1300 15936 1312
rect 15988 1300 15994 1352
rect 16025 1343 16083 1349
rect 16025 1309 16037 1343
rect 16071 1340 16083 1343
rect 16114 1340 16120 1352
rect 16071 1312 16120 1340
rect 16071 1309 16083 1312
rect 16025 1303 16083 1309
rect 16114 1300 16120 1312
rect 16172 1300 16178 1352
rect 16390 1340 16396 1352
rect 16351 1312 16396 1340
rect 16390 1300 16396 1312
rect 16448 1300 16454 1352
rect 14550 1272 14556 1284
rect 12636 1244 14556 1272
rect 14550 1232 14556 1244
rect 14608 1232 14614 1284
rect 16666 1232 16672 1284
rect 16724 1272 16730 1284
rect 17862 1272 17868 1284
rect 16724 1244 16790 1272
rect 17823 1244 17868 1272
rect 16724 1232 16730 1244
rect 17862 1232 17868 1244
rect 17920 1232 17926 1284
rect 6914 1204 6920 1216
rect 6827 1176 6920 1204
rect 6914 1164 6920 1176
rect 6972 1204 6978 1216
rect 8202 1204 8208 1216
rect 6972 1176 8208 1204
rect 6972 1164 6978 1176
rect 8202 1164 8208 1176
rect 8260 1204 8266 1216
rect 9398 1204 9404 1216
rect 8260 1176 9404 1204
rect 8260 1164 8266 1176
rect 9398 1164 9404 1176
rect 9456 1164 9462 1216
rect 10873 1207 10931 1213
rect 10873 1173 10885 1207
rect 10919 1204 10931 1207
rect 11514 1204 11520 1216
rect 10919 1176 11520 1204
rect 10919 1173 10931 1176
rect 10873 1167 10931 1173
rect 11514 1164 11520 1176
rect 11572 1164 11578 1216
rect 13354 1204 13360 1216
rect 13315 1176 13360 1204
rect 13354 1164 13360 1176
rect 13412 1164 13418 1216
rect 15841 1207 15899 1213
rect 15841 1173 15853 1207
rect 15887 1204 15899 1207
rect 16022 1204 16028 1216
rect 15887 1176 16028 1204
rect 15887 1173 15899 1176
rect 15841 1167 15899 1173
rect 16022 1164 16028 1176
rect 16080 1164 16086 1216
rect 0 1114 18860 1136
rect 0 1062 4660 1114
rect 4712 1062 4724 1114
rect 4776 1062 4788 1114
rect 4840 1062 4852 1114
rect 4904 1062 4916 1114
rect 4968 1062 7760 1114
rect 7812 1062 7824 1114
rect 7876 1062 7888 1114
rect 7940 1062 7952 1114
rect 8004 1062 8016 1114
rect 8068 1062 10860 1114
rect 10912 1062 10924 1114
rect 10976 1062 10988 1114
rect 11040 1062 11052 1114
rect 11104 1062 11116 1114
rect 11168 1062 13960 1114
rect 14012 1062 14024 1114
rect 14076 1062 14088 1114
rect 14140 1062 14152 1114
rect 14204 1062 14216 1114
rect 14268 1062 17060 1114
rect 17112 1062 17124 1114
rect 17176 1062 17188 1114
rect 17240 1062 17252 1114
rect 17304 1062 17316 1114
rect 17368 1062 18860 1114
rect 0 1040 18860 1062
rect 4295 1003 4353 1009
rect 4295 969 4307 1003
rect 4341 1000 4353 1003
rect 4982 1000 4988 1012
rect 4341 972 4844 1000
rect 4943 972 4988 1000
rect 4341 969 4353 972
rect 4295 963 4353 969
rect 2498 864 2504 876
rect 2459 836 2504 864
rect 2498 824 2504 836
rect 2556 824 2562 876
rect 3896 864 3924 918
rect 4430 892 4436 944
rect 4488 932 4494 944
rect 4816 932 4844 972
rect 4982 960 4988 972
rect 5040 960 5046 1012
rect 5902 960 5908 1012
rect 5960 1000 5966 1012
rect 7101 1003 7159 1009
rect 7101 1000 7113 1003
rect 5960 972 7113 1000
rect 5960 960 5966 972
rect 7101 969 7113 972
rect 7147 969 7159 1003
rect 7374 1000 7380 1012
rect 7335 972 7380 1000
rect 7101 963 7159 969
rect 4488 904 4660 932
rect 4816 904 4936 932
rect 4488 892 4494 904
rect 4338 864 4344 876
rect 3896 836 4344 864
rect 4338 824 4344 836
rect 4396 824 4402 876
rect 4632 873 4660 904
rect 4908 876 4936 904
rect 5442 892 5448 944
rect 5500 892 5506 944
rect 7116 932 7144 963
rect 7374 960 7380 972
rect 7432 960 7438 1012
rect 7558 960 7564 1012
rect 7616 1000 7622 1012
rect 8938 1000 8944 1012
rect 7616 972 8944 1000
rect 7616 960 7622 972
rect 7116 904 7604 932
rect 4617 867 4675 873
rect 4617 833 4629 867
rect 4663 833 4675 867
rect 4617 827 4675 833
rect 4706 824 4712 876
rect 4764 864 4770 876
rect 4764 836 4809 864
rect 4764 824 4770 836
rect 4890 824 4896 876
rect 4948 864 4954 876
rect 5074 864 5080 876
rect 4948 836 4993 864
rect 5035 836 5080 864
rect 4948 824 4954 836
rect 5074 824 5080 836
rect 5132 824 5138 876
rect 5353 867 5411 873
rect 5353 833 5365 867
rect 5399 864 5411 867
rect 5460 864 5488 892
rect 7282 864 7288 876
rect 5399 836 5488 864
rect 5399 833 5411 836
rect 5353 827 5411 833
rect 2869 799 2927 805
rect 2869 765 2881 799
rect 2915 796 2927 799
rect 4433 799 4491 805
rect 2915 768 3740 796
rect 2915 765 2927 768
rect 2869 759 2927 765
rect 3712 728 3740 768
rect 4433 765 4445 799
rect 4479 796 4491 799
rect 5626 796 5632 808
rect 4479 768 5396 796
rect 5587 768 5632 796
rect 4479 765 4491 768
rect 4433 759 4491 765
rect 5368 740 5396 768
rect 5626 756 5632 768
rect 5684 756 5690 808
rect 6748 796 6776 850
rect 7243 836 7288 864
rect 7282 824 7288 836
rect 7340 824 7346 876
rect 7466 864 7472 876
rect 7427 836 7472 864
rect 7466 824 7472 836
rect 7524 824 7530 876
rect 7576 873 7604 904
rect 7561 867 7619 873
rect 7561 833 7573 867
rect 7607 833 7619 867
rect 7742 864 7748 876
rect 7703 836 7748 864
rect 7561 827 7619 833
rect 7742 824 7748 836
rect 7800 824 7806 876
rect 8202 864 8208 876
rect 8163 836 8208 864
rect 8202 824 8208 836
rect 8260 824 8266 876
rect 8496 873 8524 972
rect 8938 960 8944 972
rect 8996 960 9002 1012
rect 9398 1000 9404 1012
rect 9359 972 9404 1000
rect 9398 960 9404 972
rect 9456 960 9462 1012
rect 11793 1003 11851 1009
rect 11793 969 11805 1003
rect 11839 969 11851 1003
rect 11793 963 11851 969
rect 12253 1003 12311 1009
rect 12253 969 12265 1003
rect 12299 1000 12311 1003
rect 12342 1000 12348 1012
rect 12299 972 12348 1000
rect 12299 969 12311 972
rect 12253 963 12311 969
rect 8570 892 8576 944
rect 8628 932 8634 944
rect 9125 935 9183 941
rect 8628 904 9076 932
rect 8628 892 8634 904
rect 8481 867 8539 873
rect 8481 833 8493 867
rect 8527 833 8539 867
rect 8754 864 8760 876
rect 8715 836 8760 864
rect 8481 827 8539 833
rect 8754 824 8760 836
rect 8812 824 8818 876
rect 9048 873 9076 904
rect 9125 901 9137 935
rect 9171 932 9183 935
rect 9674 932 9680 944
rect 9171 904 9680 932
rect 9171 901 9183 904
rect 9125 895 9183 901
rect 9674 892 9680 904
rect 9732 892 9738 944
rect 11514 932 11520 944
rect 11475 904 11520 932
rect 11514 892 11520 904
rect 11572 892 11578 944
rect 11808 932 11836 963
rect 12342 960 12348 972
rect 12400 960 12406 1012
rect 13538 960 13544 1012
rect 13596 1000 13602 1012
rect 14553 1003 14611 1009
rect 14553 1000 14565 1003
rect 13596 972 14565 1000
rect 13596 960 13602 972
rect 14553 969 14565 972
rect 14599 969 14611 1003
rect 16666 1000 16672 1012
rect 14553 963 14611 969
rect 16224 972 16672 1000
rect 11808 904 12112 932
rect 9033 867 9091 873
rect 9033 833 9045 867
rect 9079 833 9091 867
rect 9306 864 9312 876
rect 9267 836 9312 864
rect 9033 827 9091 833
rect 9306 824 9312 836
rect 9364 824 9370 876
rect 9953 867 10011 873
rect 9953 833 9965 867
rect 9999 833 10011 867
rect 10134 864 10140 876
rect 10095 836 10140 864
rect 9953 827 10011 833
rect 8294 796 8300 808
rect 6748 768 8300 796
rect 4525 731 4583 737
rect 4525 728 4537 731
rect 3712 700 4537 728
rect 4525 697 4537 700
rect 4571 697 4583 731
rect 4525 691 4583 697
rect 5350 688 5356 740
rect 5408 688 5414 740
rect 2222 620 2228 672
rect 2280 660 2286 672
rect 2317 663 2375 669
rect 2317 660 2329 663
rect 2280 632 2329 660
rect 2280 620 2286 632
rect 2317 629 2329 632
rect 2363 660 2375 663
rect 4338 660 4344 672
rect 2363 632 4344 660
rect 2363 629 2375 632
rect 2317 623 2375 629
rect 4338 620 4344 632
rect 4396 660 4402 672
rect 5261 663 5319 669
rect 5261 660 5273 663
rect 4396 632 5273 660
rect 4396 620 4402 632
rect 5261 629 5273 632
rect 5307 660 5319 663
rect 6748 660 6776 768
rect 8294 756 8300 768
rect 8352 756 8358 808
rect 9968 796 9996 827
rect 10134 824 10140 836
rect 10192 824 10198 876
rect 10410 864 10416 876
rect 10371 836 10416 864
rect 10410 824 10416 836
rect 10468 824 10474 876
rect 10226 796 10232 808
rect 8588 768 10232 796
rect 8588 737 8616 768
rect 10226 756 10232 768
rect 10284 796 10290 808
rect 11532 796 11560 892
rect 11698 864 11704 876
rect 11659 836 11704 864
rect 11698 824 11704 836
rect 11756 824 11762 876
rect 11790 824 11796 876
rect 11848 864 11854 876
rect 12084 873 12112 904
rect 12544 904 13216 932
rect 12069 867 12127 873
rect 11848 836 11893 864
rect 11848 824 11854 836
rect 12069 833 12081 867
rect 12115 833 12127 867
rect 12069 827 12127 833
rect 12158 824 12164 876
rect 12216 864 12222 876
rect 12544 873 12572 904
rect 12253 867 12311 873
rect 12253 864 12265 867
rect 12216 836 12265 864
rect 12216 824 12222 836
rect 12253 833 12265 836
rect 12299 833 12311 867
rect 12253 827 12311 833
rect 12529 867 12587 873
rect 12529 833 12541 867
rect 12575 833 12587 867
rect 12986 864 12992 876
rect 12947 836 12992 864
rect 12529 827 12587 833
rect 12544 796 12572 827
rect 12986 824 12992 836
rect 13044 824 13050 876
rect 13188 873 13216 904
rect 14826 892 14832 944
rect 14884 932 14890 944
rect 15013 935 15071 941
rect 15013 932 15025 935
rect 14884 904 15025 932
rect 14884 892 14890 904
rect 15013 901 15025 904
rect 15059 901 15071 935
rect 16224 918 16252 972
rect 16666 960 16672 972
rect 16724 960 16730 1012
rect 16942 960 16948 1012
rect 17000 1000 17006 1012
rect 17037 1003 17095 1009
rect 17037 1000 17049 1003
rect 17000 972 17049 1000
rect 17000 960 17006 972
rect 17037 969 17049 972
rect 17083 969 17095 1003
rect 17494 1000 17500 1012
rect 17455 972 17500 1000
rect 17037 963 17095 969
rect 17494 960 17500 972
rect 17552 960 17558 1012
rect 18230 960 18236 1012
rect 18288 1000 18294 1012
rect 18325 1003 18383 1009
rect 18325 1000 18337 1003
rect 18288 972 18337 1000
rect 18288 960 18294 972
rect 18325 969 18337 972
rect 18371 969 18383 1003
rect 18325 963 18383 969
rect 15013 895 15071 901
rect 13173 867 13231 873
rect 13173 833 13185 867
rect 13219 864 13231 867
rect 13262 864 13268 876
rect 13219 836 13268 864
rect 13219 833 13231 836
rect 13173 827 13231 833
rect 13262 824 13268 836
rect 13320 824 13326 876
rect 13722 864 13728 876
rect 13683 836 13728 864
rect 13722 824 13728 836
rect 13780 824 13786 876
rect 17310 824 17316 876
rect 17368 864 17374 876
rect 17405 867 17463 873
rect 17405 864 17417 867
rect 17368 836 17417 864
rect 17368 824 17374 836
rect 17405 833 17417 836
rect 17451 833 17463 867
rect 17405 827 17463 833
rect 18233 867 18291 873
rect 18233 833 18245 867
rect 18279 864 18291 867
rect 18506 864 18512 876
rect 18279 836 18512 864
rect 18279 833 18291 836
rect 18233 827 18291 833
rect 18506 824 18512 836
rect 18564 824 18570 876
rect 10284 768 10456 796
rect 11532 768 12572 796
rect 12621 799 12679 805
rect 10284 756 10290 768
rect 7745 731 7803 737
rect 7745 697 7757 731
rect 7791 728 7803 731
rect 8021 731 8079 737
rect 8021 728 8033 731
rect 7791 700 8033 728
rect 7791 697 7803 700
rect 7745 691 7803 697
rect 8021 697 8033 700
rect 8067 697 8079 731
rect 8021 691 8079 697
rect 8573 731 8631 737
rect 8573 697 8585 731
rect 8619 697 8631 731
rect 9674 728 9680 740
rect 9587 700 9680 728
rect 8573 691 8631 697
rect 9674 688 9680 700
rect 9732 728 9738 740
rect 10321 731 10379 737
rect 10321 728 10333 731
rect 9732 700 10333 728
rect 9732 688 9738 700
rect 10321 697 10333 700
rect 10367 697 10379 731
rect 10428 728 10456 768
rect 12621 765 12633 799
rect 12667 796 12679 799
rect 13538 796 13544 808
rect 12667 768 13544 796
rect 12667 765 12679 768
rect 12621 759 12679 765
rect 13538 756 13544 768
rect 13596 756 13602 808
rect 14274 796 14280 808
rect 14235 768 14280 796
rect 14274 756 14280 768
rect 14332 756 14338 808
rect 14550 756 14556 808
rect 14608 796 14614 808
rect 14737 799 14795 805
rect 14737 796 14749 799
rect 14608 768 14749 796
rect 14608 756 14614 768
rect 14737 765 14749 768
rect 14783 796 14795 799
rect 16206 796 16212 808
rect 14783 768 16212 796
rect 14783 765 14795 768
rect 14737 759 14795 765
rect 16206 756 16212 768
rect 16264 756 16270 808
rect 17586 756 17592 808
rect 17644 796 17650 808
rect 17644 768 17689 796
rect 17644 756 17650 768
rect 11790 728 11796 740
rect 10428 700 11796 728
rect 10321 691 10379 697
rect 11790 688 11796 700
rect 11848 688 11854 740
rect 12894 728 12900 740
rect 12855 700 12900 728
rect 12894 688 12900 700
rect 12952 688 12958 740
rect 14458 688 14464 740
rect 14516 728 14522 740
rect 14516 700 14688 728
rect 14516 688 14522 700
rect 5307 632 6776 660
rect 5307 629 5319 632
rect 5261 623 5319 629
rect 9122 620 9128 672
rect 9180 660 9186 672
rect 9217 663 9275 669
rect 9217 660 9229 663
rect 9180 632 9229 660
rect 9180 620 9186 632
rect 9217 629 9229 632
rect 9263 629 9275 663
rect 9950 660 9956 672
rect 9911 632 9956 660
rect 9217 623 9275 629
rect 9950 620 9956 632
rect 10008 620 10014 672
rect 14660 660 14688 700
rect 16482 660 16488 672
rect 14660 632 16488 660
rect 16482 620 16488 632
rect 16540 620 16546 672
rect 0 570 18860 592
rect 0 518 3110 570
rect 3162 518 3174 570
rect 3226 518 3238 570
rect 3290 518 3302 570
rect 3354 518 3366 570
rect 3418 518 6210 570
rect 6262 518 6274 570
rect 6326 518 6338 570
rect 6390 518 6402 570
rect 6454 518 6466 570
rect 6518 518 9310 570
rect 9362 518 9374 570
rect 9426 518 9438 570
rect 9490 518 9502 570
rect 9554 518 9566 570
rect 9618 518 12410 570
rect 12462 518 12474 570
rect 12526 518 12538 570
rect 12590 518 12602 570
rect 12654 518 12666 570
rect 12718 518 15510 570
rect 15562 518 15574 570
rect 15626 518 15638 570
rect 15690 518 15702 570
rect 15754 518 15766 570
rect 15818 518 18860 570
rect 0 496 18860 518
rect 5537 459 5595 465
rect 5537 425 5549 459
rect 5583 456 5595 459
rect 5626 456 5632 468
rect 5583 428 5632 456
rect 5583 425 5595 428
rect 5537 419 5595 425
rect 5626 416 5632 428
rect 5684 416 5690 468
rect 6181 459 6239 465
rect 6181 425 6193 459
rect 6227 456 6239 459
rect 7282 456 7288 468
rect 6227 428 7288 456
rect 6227 425 6239 428
rect 6181 419 6239 425
rect 5445 391 5503 397
rect 5445 357 5457 391
rect 5491 388 5503 391
rect 6196 388 6224 419
rect 7282 416 7288 428
rect 7340 416 7346 468
rect 8846 416 8852 468
rect 8904 456 8910 468
rect 9125 459 9183 465
rect 9125 456 9137 459
rect 8904 428 9137 456
rect 8904 416 8910 428
rect 9125 425 9137 428
rect 9171 425 9183 459
rect 13446 456 13452 468
rect 13407 428 13452 456
rect 9125 419 9183 425
rect 13446 416 13452 428
rect 13504 416 13510 468
rect 13538 416 13544 468
rect 13596 456 13602 468
rect 13596 428 13641 456
rect 13596 416 13602 428
rect 15194 416 15200 468
rect 15252 456 15258 468
rect 15657 459 15715 465
rect 15657 456 15669 459
rect 15252 428 15669 456
rect 15252 416 15258 428
rect 15657 425 15669 428
rect 15703 425 15715 459
rect 15657 419 15715 425
rect 16114 416 16120 468
rect 16172 456 16178 468
rect 16209 459 16267 465
rect 16209 456 16221 459
rect 16172 428 16221 456
rect 16172 416 16178 428
rect 16209 425 16221 428
rect 16255 425 16267 459
rect 17310 456 17316 468
rect 17271 428 17316 456
rect 16209 419 16267 425
rect 17310 416 17316 428
rect 17368 416 17374 468
rect 12250 388 12256 400
rect 5491 360 6224 388
rect 12211 360 12256 388
rect 5491 357 5503 360
rect 5445 351 5503 357
rect 12250 348 12256 360
rect 12308 348 12314 400
rect 15933 391 15991 397
rect 15933 357 15945 391
rect 15979 388 15991 391
rect 16390 388 16396 400
rect 15979 360 16396 388
rect 15979 357 15991 360
rect 15933 351 15991 357
rect 16390 348 16396 360
rect 16448 348 16454 400
rect 5810 280 5816 332
rect 5868 320 5874 332
rect 5868 292 6316 320
rect 5868 280 5874 292
rect 5166 212 5172 264
rect 5224 252 5230 264
rect 5353 255 5411 261
rect 5353 252 5365 255
rect 5224 224 5365 252
rect 5224 212 5230 224
rect 5353 221 5365 224
rect 5399 221 5411 255
rect 5902 252 5908 264
rect 5863 224 5908 252
rect 5353 215 5411 221
rect 5902 212 5908 224
rect 5960 212 5966 264
rect 6288 261 6316 292
rect 12360 292 13768 320
rect 6089 255 6147 261
rect 6089 221 6101 255
rect 6135 221 6147 255
rect 6089 215 6147 221
rect 6273 255 6331 261
rect 6273 221 6285 255
rect 6319 221 6331 255
rect 9122 252 9128 264
rect 9083 224 9128 252
rect 6273 215 6331 221
rect 4706 144 4712 196
rect 4764 184 4770 196
rect 6104 184 6132 215
rect 9122 212 9128 224
rect 9180 212 9186 264
rect 9217 255 9275 261
rect 9217 221 9229 255
rect 9263 252 9275 255
rect 9950 252 9956 264
rect 9263 224 9956 252
rect 9263 221 9275 224
rect 9217 215 9275 221
rect 9950 212 9956 224
rect 10008 212 10014 264
rect 11790 212 11796 264
rect 11848 252 11854 264
rect 12360 261 12388 292
rect 12069 255 12127 261
rect 12069 252 12081 255
rect 11848 224 12081 252
rect 11848 212 11854 224
rect 12069 221 12081 224
rect 12115 221 12127 255
rect 12069 215 12127 221
rect 12345 255 12403 261
rect 12345 221 12357 255
rect 12391 221 12403 255
rect 13262 252 13268 264
rect 13223 224 13268 252
rect 12345 215 12403 221
rect 13262 212 13268 224
rect 13320 212 13326 264
rect 13464 261 13492 292
rect 13740 264 13768 292
rect 16482 280 16488 332
rect 16540 320 16546 332
rect 16945 323 17003 329
rect 16945 320 16957 323
rect 16540 292 16957 320
rect 16540 280 16546 292
rect 16945 289 16957 292
rect 16991 289 17003 323
rect 16945 283 17003 289
rect 13449 255 13507 261
rect 13449 221 13461 255
rect 13495 221 13507 255
rect 13449 215 13507 221
rect 13541 255 13599 261
rect 13541 221 13553 255
rect 13587 221 13599 255
rect 13722 252 13728 264
rect 13683 224 13728 252
rect 13541 215 13599 221
rect 4764 156 6132 184
rect 4764 144 4770 156
rect 9030 144 9036 196
rect 9088 184 9094 196
rect 9401 187 9459 193
rect 9401 184 9413 187
rect 9088 156 9413 184
rect 9088 144 9094 156
rect 9401 153 9413 156
rect 9447 153 9459 187
rect 9401 147 9459 153
rect 11698 144 11704 196
rect 11756 184 11762 196
rect 12161 187 12219 193
rect 12161 184 12173 187
rect 11756 156 12173 184
rect 11756 144 11762 156
rect 12161 153 12173 156
rect 12207 153 12219 187
rect 12161 147 12219 153
rect 12986 144 12992 196
rect 13044 184 13050 196
rect 13556 184 13584 215
rect 13722 212 13728 224
rect 13780 212 13786 264
rect 15838 252 15844 264
rect 15799 224 15844 252
rect 15838 212 15844 224
rect 15896 212 15902 264
rect 16022 252 16028 264
rect 15983 224 16028 252
rect 16022 212 16028 224
rect 16080 212 16086 264
rect 16206 252 16212 264
rect 16167 224 16212 252
rect 16206 212 16212 224
rect 16264 212 16270 264
rect 17037 255 17095 261
rect 17037 221 17049 255
rect 17083 252 17095 255
rect 17862 252 17868 264
rect 17083 224 17868 252
rect 17083 221 17095 224
rect 17037 215 17095 221
rect 17862 212 17868 224
rect 17920 212 17926 264
rect 14458 184 14464 196
rect 13044 156 14464 184
rect 13044 144 13050 156
rect 14458 144 14464 156
rect 14516 144 14522 196
rect 5350 76 5356 128
rect 5408 116 5414 128
rect 5813 119 5871 125
rect 5813 116 5825 119
rect 5408 88 5825 116
rect 5408 76 5414 88
rect 5813 85 5825 88
rect 5859 85 5871 119
rect 5813 79 5871 85
rect 0 26 18860 48
rect 0 -26 4660 26
rect 4712 -26 4724 26
rect 4776 -26 4788 26
rect 4840 -26 4852 26
rect 4904 -26 4916 26
rect 4968 -26 7760 26
rect 7812 -26 7824 26
rect 7876 -26 7888 26
rect 7940 -26 7952 26
rect 8004 -26 8016 26
rect 8068 -26 10860 26
rect 10912 -26 10924 26
rect 10976 -26 10988 26
rect 11040 -26 11052 26
rect 11104 -26 11116 26
rect 11168 -26 13960 26
rect 14012 -26 14024 26
rect 14076 -26 14088 26
rect 14140 -26 14152 26
rect 14204 -26 14216 26
rect 14268 -26 17060 26
rect 17112 -26 17124 26
rect 17176 -26 17188 26
rect 17240 -26 17252 26
rect 17304 -26 17316 26
rect 17368 -26 18860 26
rect 0 -48 18860 -26
<< via1 >>
rect 4660 10854 4712 10906
rect 4724 10854 4776 10906
rect 4788 10854 4840 10906
rect 4852 10854 4904 10906
rect 4916 10854 4968 10906
rect 7760 10854 7812 10906
rect 7824 10854 7876 10906
rect 7888 10854 7940 10906
rect 7952 10854 8004 10906
rect 8016 10854 8068 10906
rect 10860 10854 10912 10906
rect 10924 10854 10976 10906
rect 10988 10854 11040 10906
rect 11052 10854 11104 10906
rect 11116 10854 11168 10906
rect 13960 10854 14012 10906
rect 14024 10854 14076 10906
rect 14088 10854 14140 10906
rect 14152 10854 14204 10906
rect 14216 10854 14268 10906
rect 17060 10854 17112 10906
rect 17124 10854 17176 10906
rect 17188 10854 17240 10906
rect 17252 10854 17304 10906
rect 17316 10854 17368 10906
rect 7104 10752 7156 10804
rect 296 10616 348 10668
rect 4160 10616 4212 10668
rect 9956 10752 10008 10804
rect 7656 10659 7708 10668
rect 7656 10625 7665 10659
rect 7665 10625 7699 10659
rect 7699 10625 7708 10659
rect 7656 10616 7708 10625
rect 8944 10616 8996 10668
rect 11336 10684 11388 10736
rect 12808 10752 12860 10804
rect 11244 10659 11296 10668
rect 11244 10625 11253 10659
rect 11253 10625 11287 10659
rect 11287 10625 11296 10659
rect 11244 10616 11296 10625
rect 3516 10548 3568 10600
rect 2688 10480 2740 10532
rect 1308 10412 1360 10464
rect 7012 10480 7064 10532
rect 8760 10548 8812 10600
rect 11060 10591 11112 10600
rect 11060 10557 11069 10591
rect 11069 10557 11103 10591
rect 11103 10557 11112 10591
rect 11060 10548 11112 10557
rect 10692 10480 10744 10532
rect 4436 10412 4488 10464
rect 8668 10412 8720 10464
rect 9220 10412 9272 10464
rect 11520 10412 11572 10464
rect 12808 10548 12860 10600
rect 15200 10616 15252 10668
rect 18052 10659 18104 10668
rect 18052 10625 18061 10659
rect 18061 10625 18095 10659
rect 18095 10625 18104 10659
rect 18052 10616 18104 10625
rect 13176 10480 13228 10532
rect 14372 10480 14424 10532
rect 18788 10616 18840 10668
rect 13360 10412 13412 10464
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 14464 10412 14516 10421
rect 14832 10412 14884 10464
rect 15292 10412 15344 10464
rect 16948 10455 17000 10464
rect 16948 10421 16957 10455
rect 16957 10421 16991 10455
rect 16991 10421 17000 10455
rect 16948 10412 17000 10421
rect 3110 10310 3162 10362
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 6210 10310 6262 10362
rect 6274 10310 6326 10362
rect 6338 10310 6390 10362
rect 6402 10310 6454 10362
rect 6466 10310 6518 10362
rect 9310 10310 9362 10362
rect 9374 10310 9426 10362
rect 9438 10310 9490 10362
rect 9502 10310 9554 10362
rect 9566 10310 9618 10362
rect 12410 10310 12462 10362
rect 12474 10310 12526 10362
rect 12538 10310 12590 10362
rect 12602 10310 12654 10362
rect 12666 10310 12718 10362
rect 15510 10310 15562 10362
rect 15574 10310 15626 10362
rect 15638 10310 15690 10362
rect 15702 10310 15754 10362
rect 15766 10310 15818 10362
rect 3516 10251 3568 10260
rect 3516 10217 3525 10251
rect 3525 10217 3559 10251
rect 3559 10217 3568 10251
rect 3516 10208 3568 10217
rect 7656 10208 7708 10260
rect 1308 10115 1360 10124
rect 1308 10081 1317 10115
rect 1317 10081 1351 10115
rect 1351 10081 1360 10115
rect 1308 10072 1360 10081
rect 2596 10072 2648 10124
rect 4344 10140 4396 10192
rect 4896 10140 4948 10192
rect 8760 10183 8812 10192
rect 8760 10149 8769 10183
rect 8769 10149 8803 10183
rect 8803 10149 8812 10183
rect 8760 10140 8812 10149
rect 10692 10183 10744 10192
rect 10692 10149 10701 10183
rect 10701 10149 10735 10183
rect 10735 10149 10744 10183
rect 10692 10140 10744 10149
rect 11244 10208 11296 10260
rect 13176 10208 13228 10260
rect 14924 10208 14976 10260
rect 15200 10208 15252 10260
rect 18052 10208 18104 10260
rect 2688 9936 2740 9988
rect 2228 9868 2280 9920
rect 4160 10072 4212 10124
rect 4068 9936 4120 9988
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 5448 10072 5500 10124
rect 6368 10072 6420 10124
rect 4896 10004 4948 10013
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 6184 10004 6236 10056
rect 6460 10047 6512 10056
rect 6460 10013 6469 10047
rect 6469 10013 6503 10047
rect 6503 10013 6512 10047
rect 6460 10004 6512 10013
rect 8668 10047 8720 10056
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 8668 10004 8720 10013
rect 7012 9936 7064 9988
rect 4528 9868 4580 9920
rect 5724 9868 5776 9920
rect 7656 9868 7708 9920
rect 8484 9911 8536 9920
rect 8484 9877 8493 9911
rect 8493 9877 8527 9911
rect 8527 9877 8536 9911
rect 8484 9868 8536 9877
rect 9956 10072 10008 10124
rect 13360 10115 13412 10124
rect 13360 10081 13369 10115
rect 13369 10081 13403 10115
rect 13403 10081 13412 10115
rect 13360 10072 13412 10081
rect 14464 10072 14516 10124
rect 16948 10072 17000 10124
rect 16488 10004 16540 10056
rect 18604 10004 18656 10056
rect 9220 9979 9272 9988
rect 9220 9945 9229 9979
rect 9229 9945 9263 9979
rect 9263 9945 9272 9979
rect 9220 9936 9272 9945
rect 9680 9936 9732 9988
rect 9864 9868 9916 9920
rect 14372 9868 14424 9920
rect 18328 9911 18380 9920
rect 18328 9877 18337 9911
rect 18337 9877 18371 9911
rect 18371 9877 18380 9911
rect 18328 9868 18380 9877
rect 4660 9766 4712 9818
rect 4724 9766 4776 9818
rect 4788 9766 4840 9818
rect 4852 9766 4904 9818
rect 4916 9766 4968 9818
rect 7760 9766 7812 9818
rect 7824 9766 7876 9818
rect 7888 9766 7940 9818
rect 7952 9766 8004 9818
rect 8016 9766 8068 9818
rect 10860 9766 10912 9818
rect 10924 9766 10976 9818
rect 10988 9766 11040 9818
rect 11052 9766 11104 9818
rect 11116 9766 11168 9818
rect 13960 9766 14012 9818
rect 14024 9766 14076 9818
rect 14088 9766 14140 9818
rect 14152 9766 14204 9818
rect 14216 9766 14268 9818
rect 17060 9766 17112 9818
rect 17124 9766 17176 9818
rect 17188 9766 17240 9818
rect 17252 9766 17304 9818
rect 17316 9766 17368 9818
rect 1952 9596 2004 9648
rect 2688 9596 2740 9648
rect 4160 9664 4212 9716
rect 3056 9596 3108 9648
rect 4068 9596 4120 9648
rect 5356 9639 5408 9648
rect 2136 9571 2188 9580
rect 2136 9537 2145 9571
rect 2145 9537 2179 9571
rect 2179 9537 2188 9571
rect 2136 9528 2188 9537
rect 2504 9571 2556 9580
rect 296 9503 348 9512
rect 296 9469 305 9503
rect 305 9469 339 9503
rect 339 9469 348 9503
rect 296 9460 348 9469
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 5356 9605 5365 9639
rect 5365 9605 5399 9639
rect 5399 9605 5408 9639
rect 5356 9596 5408 9605
rect 2504 9528 2556 9537
rect 3056 9460 3108 9512
rect 2688 9324 2740 9376
rect 4528 9528 4580 9580
rect 5448 9571 5500 9580
rect 5448 9537 5457 9571
rect 5457 9537 5491 9571
rect 5491 9537 5500 9571
rect 5448 9528 5500 9537
rect 6460 9664 6512 9716
rect 8944 9664 8996 9716
rect 5724 9639 5776 9648
rect 5724 9605 5733 9639
rect 5733 9605 5767 9639
rect 5767 9605 5776 9639
rect 5724 9596 5776 9605
rect 6184 9639 6236 9648
rect 6184 9605 6193 9639
rect 6193 9605 6227 9639
rect 6227 9605 6236 9639
rect 6184 9596 6236 9605
rect 6368 9596 6420 9648
rect 8484 9596 8536 9648
rect 9680 9596 9732 9648
rect 10048 9639 10100 9648
rect 10048 9605 10057 9639
rect 10057 9605 10091 9639
rect 10091 9605 10100 9639
rect 10048 9596 10100 9605
rect 10692 9596 10744 9648
rect 6092 9528 6144 9580
rect 7656 9528 7708 9580
rect 4344 9460 4396 9512
rect 6000 9460 6052 9512
rect 3608 9435 3660 9444
rect 3608 9401 3617 9435
rect 3617 9401 3651 9435
rect 3651 9401 3660 9435
rect 3608 9392 3660 9401
rect 5264 9324 5316 9376
rect 7564 9460 7616 9512
rect 9956 9528 10008 9580
rect 11796 9528 11848 9580
rect 14372 9664 14424 9716
rect 14464 9664 14516 9716
rect 16580 9664 16632 9716
rect 9680 9392 9732 9444
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 11152 9460 11204 9512
rect 11612 9460 11664 9512
rect 12808 9460 12860 9512
rect 14832 9571 14884 9580
rect 14832 9537 14841 9571
rect 14841 9537 14875 9571
rect 14875 9537 14884 9571
rect 14832 9528 14884 9537
rect 15292 9528 15344 9580
rect 18328 9460 18380 9512
rect 11428 9324 11480 9376
rect 13360 9324 13412 9376
rect 13452 9324 13504 9376
rect 14464 9324 14516 9376
rect 16672 9324 16724 9376
rect 3110 9222 3162 9274
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 6210 9222 6262 9274
rect 6274 9222 6326 9274
rect 6338 9222 6390 9274
rect 6402 9222 6454 9274
rect 6466 9222 6518 9274
rect 9310 9222 9362 9274
rect 9374 9222 9426 9274
rect 9438 9222 9490 9274
rect 9502 9222 9554 9274
rect 9566 9222 9618 9274
rect 12410 9222 12462 9274
rect 12474 9222 12526 9274
rect 12538 9222 12590 9274
rect 12602 9222 12654 9274
rect 12666 9222 12718 9274
rect 15510 9222 15562 9274
rect 15574 9222 15626 9274
rect 15638 9222 15690 9274
rect 15702 9222 15754 9274
rect 15766 9222 15818 9274
rect 1400 9163 1452 9172
rect 1400 9129 1409 9163
rect 1409 9129 1443 9163
rect 1443 9129 1452 9163
rect 1400 9120 1452 9129
rect 2964 9120 3016 9172
rect 10692 9163 10744 9172
rect 10692 9129 10701 9163
rect 10701 9129 10735 9163
rect 10735 9129 10744 9163
rect 10692 9120 10744 9129
rect 11796 9120 11848 9172
rect 14188 9120 14240 9172
rect 14464 9120 14516 9172
rect 1952 9027 2004 9036
rect 1952 8993 1961 9027
rect 1961 8993 1995 9027
rect 1995 8993 2004 9027
rect 1952 8984 2004 8993
rect 4528 8984 4580 9036
rect 1400 8916 1452 8968
rect 2688 8916 2740 8968
rect 4436 8959 4488 8968
rect 4436 8925 4445 8959
rect 4445 8925 4479 8959
rect 4479 8925 4488 8959
rect 4436 8916 4488 8925
rect 4988 8916 5040 8968
rect 5264 8916 5316 8968
rect 6092 8916 6144 8968
rect 8392 8916 8444 8968
rect 8484 8916 8536 8968
rect 10692 8984 10744 9036
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 10784 8916 10836 8968
rect 11244 8959 11296 8968
rect 11244 8925 11253 8959
rect 11253 8925 11287 8959
rect 11287 8925 11296 8959
rect 11244 8916 11296 8925
rect 13360 8984 13412 9036
rect 14464 8984 14516 9036
rect 16672 8984 16724 9036
rect 13452 8959 13504 8968
rect 4344 8848 4396 8900
rect 8300 8848 8352 8900
rect 1952 8780 2004 8832
rect 2504 8780 2556 8832
rect 3608 8780 3660 8832
rect 4160 8780 4212 8832
rect 4436 8780 4488 8832
rect 5264 8780 5316 8832
rect 8576 8780 8628 8832
rect 9128 8848 9180 8900
rect 9496 8848 9548 8900
rect 11796 8848 11848 8900
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 15844 8916 15896 8968
rect 11980 8780 12032 8832
rect 14188 8848 14240 8900
rect 16488 8848 16540 8900
rect 14372 8780 14424 8832
rect 18052 8780 18104 8832
rect 4660 8678 4712 8730
rect 4724 8678 4776 8730
rect 4788 8678 4840 8730
rect 4852 8678 4904 8730
rect 4916 8678 4968 8730
rect 7760 8678 7812 8730
rect 7824 8678 7876 8730
rect 7888 8678 7940 8730
rect 7952 8678 8004 8730
rect 8016 8678 8068 8730
rect 10860 8678 10912 8730
rect 10924 8678 10976 8730
rect 10988 8678 11040 8730
rect 11052 8678 11104 8730
rect 11116 8678 11168 8730
rect 13960 8678 14012 8730
rect 14024 8678 14076 8730
rect 14088 8678 14140 8730
rect 14152 8678 14204 8730
rect 14216 8678 14268 8730
rect 17060 8678 17112 8730
rect 17124 8678 17176 8730
rect 17188 8678 17240 8730
rect 17252 8678 17304 8730
rect 17316 8678 17368 8730
rect 2136 8619 2188 8628
rect 2136 8585 2145 8619
rect 2145 8585 2179 8619
rect 2179 8585 2188 8619
rect 2136 8576 2188 8585
rect 4160 8619 4212 8628
rect 4160 8585 4169 8619
rect 4169 8585 4203 8619
rect 4203 8585 4212 8619
rect 4160 8576 4212 8585
rect 4344 8576 4396 8628
rect 5264 8619 5316 8628
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 9496 8619 9548 8628
rect 1952 8508 2004 8560
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 296 8415 348 8424
rect 296 8381 305 8415
rect 305 8381 339 8415
rect 339 8381 348 8415
rect 296 8372 348 8381
rect 4068 8508 4120 8560
rect 4436 8508 4488 8560
rect 5356 8508 5408 8560
rect 7472 8508 7524 8560
rect 9496 8585 9505 8619
rect 9505 8585 9539 8619
rect 9539 8585 9548 8619
rect 9496 8576 9548 8585
rect 9680 8576 9732 8628
rect 11244 8576 11296 8628
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 2688 8483 2740 8492
rect 2228 8304 2280 8356
rect 2688 8449 2697 8483
rect 2697 8449 2731 8483
rect 2731 8449 2740 8483
rect 2688 8440 2740 8449
rect 2780 8483 2832 8492
rect 2780 8449 2789 8483
rect 2789 8449 2823 8483
rect 2823 8449 2832 8483
rect 2780 8440 2832 8449
rect 2412 8372 2464 8424
rect 4528 8440 4580 8492
rect 4988 8372 5040 8424
rect 5172 8304 5224 8356
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 2964 8236 3016 8245
rect 7288 8440 7340 8492
rect 10140 8508 10192 8560
rect 10600 8508 10652 8560
rect 8392 8440 8444 8492
rect 8576 8440 8628 8492
rect 12900 8508 12952 8560
rect 14556 8576 14608 8628
rect 13452 8508 13504 8560
rect 15844 8576 15896 8628
rect 15108 8508 15160 8560
rect 8668 8372 8720 8424
rect 11980 8440 12032 8492
rect 12808 8440 12860 8492
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 11704 8372 11756 8424
rect 6092 8236 6144 8288
rect 7656 8236 7708 8288
rect 7932 8279 7984 8288
rect 7932 8245 7941 8279
rect 7941 8245 7975 8279
rect 7975 8245 7984 8279
rect 8576 8279 8628 8288
rect 7932 8236 7984 8245
rect 8576 8245 8585 8279
rect 8585 8245 8619 8279
rect 8619 8245 8628 8279
rect 8576 8236 8628 8245
rect 8668 8236 8720 8288
rect 10784 8236 10836 8288
rect 11336 8304 11388 8356
rect 12164 8372 12216 8424
rect 13268 8415 13320 8424
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 13268 8372 13320 8381
rect 14372 8440 14424 8492
rect 14464 8372 14516 8424
rect 16672 8415 16724 8424
rect 16672 8381 16681 8415
rect 16681 8381 16715 8415
rect 16715 8381 16724 8415
rect 16672 8372 16724 8381
rect 17868 8372 17920 8424
rect 18604 8440 18656 8492
rect 12716 8304 12768 8356
rect 11244 8236 11296 8288
rect 12256 8236 12308 8288
rect 14280 8236 14332 8288
rect 3110 8134 3162 8186
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 6210 8134 6262 8186
rect 6274 8134 6326 8186
rect 6338 8134 6390 8186
rect 6402 8134 6454 8186
rect 6466 8134 6518 8186
rect 9310 8134 9362 8186
rect 9374 8134 9426 8186
rect 9438 8134 9490 8186
rect 9502 8134 9554 8186
rect 9566 8134 9618 8186
rect 12410 8134 12462 8186
rect 12474 8134 12526 8186
rect 12538 8134 12590 8186
rect 12602 8134 12654 8186
rect 12666 8134 12718 8186
rect 15510 8134 15562 8186
rect 15574 8134 15626 8186
rect 15638 8134 15690 8186
rect 15702 8134 15754 8186
rect 15766 8134 15818 8186
rect 2136 8032 2188 8084
rect 2688 8032 2740 8084
rect 4252 8032 4304 8084
rect 9772 8032 9824 8084
rect 12900 8032 12952 8084
rect 13360 8032 13412 8084
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 16488 8032 16540 8084
rect 2780 7964 2832 8016
rect 5080 7964 5132 8016
rect 5356 7964 5408 8016
rect 7656 8007 7708 8016
rect 7656 7973 7665 8007
rect 7665 7973 7699 8007
rect 7699 7973 7708 8007
rect 7656 7964 7708 7973
rect 7932 8007 7984 8016
rect 7932 7973 7941 8007
rect 7941 7973 7975 8007
rect 7975 7973 7984 8007
rect 7932 7964 7984 7973
rect 2228 7896 2280 7948
rect 2504 7939 2556 7948
rect 2504 7905 2513 7939
rect 2513 7905 2547 7939
rect 2547 7905 2556 7939
rect 2504 7896 2556 7905
rect 3516 7896 3568 7948
rect 5264 7939 5316 7948
rect 5264 7905 5273 7939
rect 5273 7905 5307 7939
rect 5307 7905 5316 7939
rect 5264 7896 5316 7905
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 2320 7871 2372 7880
rect 2320 7837 2329 7871
rect 2329 7837 2363 7871
rect 2363 7837 2372 7871
rect 2320 7828 2372 7837
rect 2964 7871 3016 7880
rect 2964 7837 2973 7871
rect 2973 7837 3007 7871
rect 3007 7837 3016 7871
rect 2964 7828 3016 7837
rect 4988 7828 5040 7880
rect 6644 7896 6696 7948
rect 7288 7939 7340 7948
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 8300 7896 8352 7948
rect 8484 7939 8536 7948
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 8484 7896 8536 7905
rect 9128 7896 9180 7948
rect 11336 7964 11388 8016
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 12808 7964 12860 8016
rect 6092 7828 6144 7880
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 8116 7871 8168 7880
rect 8116 7837 8125 7871
rect 8125 7837 8159 7871
rect 8159 7837 8168 7871
rect 8116 7828 8168 7837
rect 11980 7828 12032 7880
rect 5356 7760 5408 7812
rect 6552 7760 6604 7812
rect 8392 7760 8444 7812
rect 2504 7692 2556 7744
rect 4160 7692 4212 7744
rect 10048 7760 10100 7812
rect 10140 7760 10192 7812
rect 11796 7760 11848 7812
rect 11244 7692 11296 7744
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 13728 7896 13780 7948
rect 14280 7939 14332 7948
rect 14280 7905 14289 7939
rect 14289 7905 14323 7939
rect 14323 7905 14332 7939
rect 14280 7896 14332 7905
rect 12256 7828 12308 7837
rect 13544 7828 13596 7880
rect 14556 7871 14608 7880
rect 14556 7837 14565 7871
rect 14565 7837 14599 7871
rect 14599 7837 14608 7871
rect 14556 7828 14608 7837
rect 16672 7896 16724 7948
rect 13268 7760 13320 7812
rect 13636 7760 13688 7812
rect 13820 7760 13872 7812
rect 14372 7760 14424 7812
rect 16120 7803 16172 7812
rect 16120 7769 16129 7803
rect 16129 7769 16163 7803
rect 16163 7769 16172 7803
rect 16120 7760 16172 7769
rect 16580 7760 16632 7812
rect 17500 7760 17552 7812
rect 13452 7692 13504 7744
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 15016 7735 15068 7744
rect 15016 7701 15025 7735
rect 15025 7701 15059 7735
rect 15059 7701 15068 7735
rect 15016 7692 15068 7701
rect 4660 7590 4712 7642
rect 4724 7590 4776 7642
rect 4788 7590 4840 7642
rect 4852 7590 4904 7642
rect 4916 7590 4968 7642
rect 7760 7590 7812 7642
rect 7824 7590 7876 7642
rect 7888 7590 7940 7642
rect 7952 7590 8004 7642
rect 8016 7590 8068 7642
rect 10860 7590 10912 7642
rect 10924 7590 10976 7642
rect 10988 7590 11040 7642
rect 11052 7590 11104 7642
rect 11116 7590 11168 7642
rect 13960 7590 14012 7642
rect 14024 7590 14076 7642
rect 14088 7590 14140 7642
rect 14152 7590 14204 7642
rect 14216 7590 14268 7642
rect 17060 7590 17112 7642
rect 17124 7590 17176 7642
rect 17188 7590 17240 7642
rect 17252 7590 17304 7642
rect 17316 7590 17368 7642
rect 2136 7488 2188 7540
rect 2412 7488 2464 7540
rect 5448 7488 5500 7540
rect 7196 7488 7248 7540
rect 9128 7488 9180 7540
rect 10692 7531 10744 7540
rect 10692 7497 10701 7531
rect 10701 7497 10735 7531
rect 10735 7497 10744 7531
rect 10692 7488 10744 7497
rect 11244 7488 11296 7540
rect 11704 7531 11756 7540
rect 11704 7497 11713 7531
rect 11713 7497 11747 7531
rect 11747 7497 11756 7531
rect 11704 7488 11756 7497
rect 13728 7531 13780 7540
rect 13728 7497 13737 7531
rect 13737 7497 13771 7531
rect 13771 7497 13780 7531
rect 13728 7488 13780 7497
rect 1952 7420 2004 7472
rect 2044 7352 2096 7404
rect 2504 7352 2556 7404
rect 2872 7420 2924 7472
rect 296 7327 348 7336
rect 296 7293 305 7327
rect 305 7293 339 7327
rect 339 7293 348 7327
rect 296 7284 348 7293
rect 572 7327 624 7336
rect 572 7293 581 7327
rect 581 7293 615 7327
rect 615 7293 624 7327
rect 572 7284 624 7293
rect 3516 7352 3568 7404
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 5264 7420 5316 7472
rect 8392 7420 8444 7472
rect 4896 7352 4948 7404
rect 4988 7352 5040 7404
rect 5356 7395 5408 7404
rect 5356 7361 5365 7395
rect 5365 7361 5399 7395
rect 5399 7361 5408 7395
rect 5356 7352 5408 7361
rect 5632 7284 5684 7336
rect 6920 7352 6972 7404
rect 7104 7352 7156 7404
rect 5908 7284 5960 7336
rect 6644 7284 6696 7336
rect 8668 7352 8720 7404
rect 8852 7395 8904 7404
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 9864 7352 9916 7404
rect 10508 7352 10560 7404
rect 8024 7327 8076 7336
rect 8024 7293 8033 7327
rect 8033 7293 8067 7327
rect 8067 7293 8076 7327
rect 8024 7284 8076 7293
rect 5816 7216 5868 7268
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 10876 7395 10928 7404
rect 10876 7361 10885 7395
rect 10885 7361 10919 7395
rect 10919 7361 10928 7395
rect 10876 7352 10928 7361
rect 11336 7352 11388 7404
rect 11060 7284 11112 7336
rect 11796 7352 11848 7404
rect 12256 7352 12308 7404
rect 13452 7395 13504 7404
rect 13452 7361 13461 7395
rect 13461 7361 13495 7395
rect 13495 7361 13504 7395
rect 13452 7352 13504 7361
rect 13636 7395 13688 7404
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 13636 7352 13688 7361
rect 13728 7417 13780 7438
rect 13728 7386 13735 7417
rect 13735 7386 13769 7417
rect 13769 7386 13780 7417
rect 14004 7420 14056 7472
rect 14372 7420 14424 7472
rect 14556 7420 14608 7472
rect 15108 7420 15160 7472
rect 13912 7352 13964 7404
rect 14648 7352 14700 7404
rect 12164 7284 12216 7336
rect 15016 7284 15068 7336
rect 16304 7327 16356 7336
rect 16304 7293 16313 7327
rect 16313 7293 16347 7327
rect 16347 7293 16356 7327
rect 16304 7284 16356 7293
rect 10048 7216 10100 7268
rect 10232 7216 10284 7268
rect 2964 7148 3016 7200
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 7380 7191 7432 7200
rect 7380 7157 7389 7191
rect 7389 7157 7423 7191
rect 7423 7157 7432 7191
rect 7380 7148 7432 7157
rect 8300 7191 8352 7200
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 8484 7191 8536 7200
rect 8484 7157 8493 7191
rect 8493 7157 8527 7191
rect 8527 7157 8536 7191
rect 8484 7148 8536 7157
rect 10968 7191 11020 7200
rect 10968 7157 10977 7191
rect 10977 7157 11011 7191
rect 11011 7157 11020 7191
rect 10968 7148 11020 7157
rect 13728 7148 13780 7200
rect 14004 7148 14056 7200
rect 14372 7148 14424 7200
rect 18512 7148 18564 7200
rect 3110 7046 3162 7098
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 6210 7046 6262 7098
rect 6274 7046 6326 7098
rect 6338 7046 6390 7098
rect 6402 7046 6454 7098
rect 6466 7046 6518 7098
rect 9310 7046 9362 7098
rect 9374 7046 9426 7098
rect 9438 7046 9490 7098
rect 9502 7046 9554 7098
rect 9566 7046 9618 7098
rect 12410 7046 12462 7098
rect 12474 7046 12526 7098
rect 12538 7046 12590 7098
rect 12602 7046 12654 7098
rect 12666 7046 12718 7098
rect 15510 7046 15562 7098
rect 15574 7046 15626 7098
rect 15638 7046 15690 7098
rect 15702 7046 15754 7098
rect 15766 7046 15818 7098
rect 1952 6944 2004 6996
rect 6920 6987 6972 6996
rect 6920 6953 6929 6987
rect 6929 6953 6963 6987
rect 6963 6953 6972 6987
rect 6920 6944 6972 6953
rect 7472 6944 7524 6996
rect 10048 6944 10100 6996
rect 10968 6944 11020 6996
rect 15108 6944 15160 6996
rect 15844 6944 15896 6996
rect 16120 6987 16172 6996
rect 16120 6953 16129 6987
rect 16129 6953 16163 6987
rect 16163 6953 16172 6987
rect 16120 6944 16172 6953
rect 2320 6876 2372 6928
rect 4252 6876 4304 6928
rect 4068 6808 4120 6860
rect 5264 6876 5316 6928
rect 5816 6876 5868 6928
rect 2872 6783 2924 6792
rect 2872 6749 2881 6783
rect 2881 6749 2915 6783
rect 2915 6749 2924 6783
rect 2872 6740 2924 6749
rect 2964 6740 3016 6792
rect 5356 6808 5408 6860
rect 572 6672 624 6724
rect 2780 6715 2832 6724
rect 2780 6681 2789 6715
rect 2789 6681 2823 6715
rect 2823 6681 2832 6715
rect 4896 6740 4948 6792
rect 5080 6783 5132 6792
rect 5080 6749 5089 6783
rect 5089 6749 5123 6783
rect 5123 6749 5132 6783
rect 5080 6740 5132 6749
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 5632 6740 5684 6749
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 8116 6876 8168 6928
rect 9036 6876 9088 6928
rect 7380 6808 7432 6860
rect 7472 6808 7524 6860
rect 8024 6808 8076 6860
rect 5724 6740 5776 6749
rect 2780 6672 2832 6681
rect 2596 6604 2648 6656
rect 7656 6740 7708 6792
rect 8392 6808 8444 6860
rect 10508 6808 10560 6860
rect 10692 6808 10744 6860
rect 10876 6808 10928 6860
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 10416 6740 10468 6792
rect 11060 6740 11112 6792
rect 11796 6783 11848 6792
rect 11796 6749 11805 6783
rect 11805 6749 11839 6783
rect 11839 6749 11848 6783
rect 11796 6740 11848 6749
rect 8484 6672 8536 6724
rect 9680 6672 9732 6724
rect 10784 6672 10836 6724
rect 10968 6672 11020 6724
rect 6828 6647 6880 6656
rect 6828 6613 6837 6647
rect 6837 6613 6871 6647
rect 6871 6613 6880 6647
rect 6828 6604 6880 6613
rect 7196 6604 7248 6656
rect 7472 6604 7524 6656
rect 10416 6647 10468 6656
rect 10416 6613 10425 6647
rect 10425 6613 10459 6647
rect 10459 6613 10468 6647
rect 10416 6604 10468 6613
rect 10600 6604 10652 6656
rect 11244 6647 11296 6656
rect 11244 6613 11253 6647
rect 11253 6613 11287 6647
rect 11287 6613 11296 6647
rect 11244 6604 11296 6613
rect 12348 6604 12400 6656
rect 13544 6740 13596 6792
rect 14464 6808 14516 6860
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 18328 6808 18380 6860
rect 17868 6783 17920 6792
rect 17868 6749 17877 6783
rect 17877 6749 17911 6783
rect 17911 6749 17920 6783
rect 17868 6740 17920 6749
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 13728 6647 13780 6656
rect 13728 6613 13737 6647
rect 13737 6613 13771 6647
rect 13771 6613 13780 6647
rect 13728 6604 13780 6613
rect 15844 6672 15896 6724
rect 15200 6647 15252 6656
rect 15200 6613 15209 6647
rect 15209 6613 15243 6647
rect 15243 6613 15252 6647
rect 15200 6604 15252 6613
rect 4660 6502 4712 6554
rect 4724 6502 4776 6554
rect 4788 6502 4840 6554
rect 4852 6502 4904 6554
rect 4916 6502 4968 6554
rect 7760 6502 7812 6554
rect 7824 6502 7876 6554
rect 7888 6502 7940 6554
rect 7952 6502 8004 6554
rect 8016 6502 8068 6554
rect 10860 6502 10912 6554
rect 10924 6502 10976 6554
rect 10988 6502 11040 6554
rect 11052 6502 11104 6554
rect 11116 6502 11168 6554
rect 13960 6502 14012 6554
rect 14024 6502 14076 6554
rect 14088 6502 14140 6554
rect 14152 6502 14204 6554
rect 14216 6502 14268 6554
rect 17060 6502 17112 6554
rect 17124 6502 17176 6554
rect 17188 6502 17240 6554
rect 17252 6502 17304 6554
rect 17316 6502 17368 6554
rect 1952 6400 2004 6452
rect 2504 6400 2556 6452
rect 2780 6400 2832 6452
rect 2964 6400 3016 6452
rect 3700 6443 3752 6452
rect 3700 6409 3709 6443
rect 3709 6409 3743 6443
rect 3743 6409 3752 6443
rect 3700 6400 3752 6409
rect 5264 6443 5316 6452
rect 5264 6409 5273 6443
rect 5273 6409 5307 6443
rect 5307 6409 5316 6443
rect 5264 6400 5316 6409
rect 5724 6400 5776 6452
rect 5908 6443 5960 6452
rect 5908 6409 5917 6443
rect 5917 6409 5951 6443
rect 5951 6409 5960 6443
rect 5908 6400 5960 6409
rect 6644 6443 6696 6452
rect 6644 6409 6653 6443
rect 6653 6409 6687 6443
rect 6687 6409 6696 6443
rect 6644 6400 6696 6409
rect 7472 6400 7524 6452
rect 2596 6307 2648 6316
rect 2596 6273 2605 6307
rect 2605 6273 2639 6307
rect 2639 6273 2648 6307
rect 2596 6264 2648 6273
rect 3516 6332 3568 6384
rect 296 6239 348 6248
rect 296 6205 305 6239
rect 305 6205 339 6239
rect 339 6205 348 6239
rect 296 6196 348 6205
rect 572 6239 624 6248
rect 572 6205 581 6239
rect 581 6205 615 6239
rect 615 6205 624 6239
rect 572 6196 624 6205
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 2964 6196 3016 6248
rect 5632 6264 5684 6316
rect 6000 6307 6052 6316
rect 5172 6196 5224 6248
rect 5448 6239 5500 6248
rect 5448 6205 5457 6239
rect 5457 6205 5491 6239
rect 5491 6205 5500 6239
rect 6000 6273 6009 6307
rect 6009 6273 6043 6307
rect 6043 6273 6052 6307
rect 6000 6264 6052 6273
rect 6552 6332 6604 6384
rect 10232 6400 10284 6452
rect 10600 6400 10652 6452
rect 11888 6443 11940 6452
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 9772 6332 9824 6384
rect 10416 6332 10468 6384
rect 9036 6264 9088 6316
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 5448 6196 5500 6205
rect 7380 6196 7432 6248
rect 7656 6196 7708 6248
rect 10600 6264 10652 6316
rect 10692 6264 10744 6316
rect 13820 6400 13872 6452
rect 14372 6400 14424 6452
rect 15200 6400 15252 6452
rect 18052 6443 18104 6452
rect 12348 6375 12400 6384
rect 12348 6341 12357 6375
rect 12357 6341 12391 6375
rect 12391 6341 12400 6375
rect 12348 6332 12400 6341
rect 13728 6332 13780 6384
rect 10140 6239 10192 6248
rect 10140 6205 10149 6239
rect 10149 6205 10183 6239
rect 10183 6205 10192 6239
rect 10140 6196 10192 6205
rect 7104 6171 7156 6180
rect 7104 6137 7113 6171
rect 7113 6137 7147 6171
rect 7147 6137 7156 6171
rect 7104 6128 7156 6137
rect 8116 6128 8168 6180
rect 9864 6171 9916 6180
rect 2872 6060 2924 6112
rect 9128 6060 9180 6112
rect 9864 6137 9873 6171
rect 9873 6137 9907 6171
rect 9907 6137 9916 6171
rect 9864 6128 9916 6137
rect 10048 6128 10100 6180
rect 11888 6196 11940 6248
rect 18052 6409 18061 6443
rect 18061 6409 18095 6443
rect 18095 6409 18104 6443
rect 18052 6400 18104 6409
rect 13544 6128 13596 6180
rect 14372 6196 14424 6248
rect 17316 6239 17368 6248
rect 17316 6205 17325 6239
rect 17325 6205 17359 6239
rect 17359 6205 17368 6239
rect 17316 6196 17368 6205
rect 17500 6239 17552 6248
rect 17500 6205 17509 6239
rect 17509 6205 17543 6239
rect 17543 6205 17552 6239
rect 17500 6196 17552 6205
rect 18144 6239 18196 6248
rect 18144 6205 18153 6239
rect 18153 6205 18187 6239
rect 18187 6205 18196 6239
rect 18144 6196 18196 6205
rect 18328 6239 18380 6248
rect 18328 6205 18337 6239
rect 18337 6205 18371 6239
rect 18371 6205 18380 6239
rect 18328 6196 18380 6205
rect 10416 6060 10468 6112
rect 14096 6103 14148 6112
rect 14096 6069 14105 6103
rect 14105 6069 14139 6103
rect 14139 6069 14148 6103
rect 14096 6060 14148 6069
rect 16396 6060 16448 6112
rect 3110 5958 3162 6010
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 6210 5958 6262 6010
rect 6274 5958 6326 6010
rect 6338 5958 6390 6010
rect 6402 5958 6454 6010
rect 6466 5958 6518 6010
rect 9310 5958 9362 6010
rect 9374 5958 9426 6010
rect 9438 5958 9490 6010
rect 9502 5958 9554 6010
rect 9566 5958 9618 6010
rect 12410 5958 12462 6010
rect 12474 5958 12526 6010
rect 12538 5958 12590 6010
rect 12602 5958 12654 6010
rect 12666 5958 12718 6010
rect 15510 5958 15562 6010
rect 15574 5958 15626 6010
rect 15638 5958 15690 6010
rect 15702 5958 15754 6010
rect 15766 5958 15818 6010
rect 572 5856 624 5908
rect 5540 5856 5592 5908
rect 6000 5856 6052 5908
rect 3424 5831 3476 5840
rect 3424 5797 3433 5831
rect 3433 5797 3467 5831
rect 3467 5797 3476 5831
rect 3424 5788 3476 5797
rect 296 5720 348 5772
rect 3700 5763 3752 5772
rect 3700 5729 3709 5763
rect 3709 5729 3743 5763
rect 3743 5729 3752 5763
rect 3700 5720 3752 5729
rect 6092 5763 6144 5772
rect 6092 5729 6101 5763
rect 6101 5729 6135 5763
rect 6135 5729 6144 5763
rect 6092 5720 6144 5729
rect 6828 5720 6880 5772
rect 7656 5856 7708 5908
rect 8852 5856 8904 5908
rect 9680 5856 9732 5908
rect 2780 5652 2832 5704
rect 2964 5652 3016 5704
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 5448 5652 5500 5704
rect 10048 5720 10100 5772
rect 10416 5763 10468 5772
rect 10416 5729 10425 5763
rect 10425 5729 10459 5763
rect 10459 5729 10468 5763
rect 10416 5720 10468 5729
rect 10692 5763 10744 5772
rect 10692 5729 10701 5763
rect 10701 5729 10735 5763
rect 10735 5729 10744 5763
rect 10692 5720 10744 5729
rect 11244 5856 11296 5908
rect 15844 5899 15896 5908
rect 15844 5865 15853 5899
rect 15853 5865 15887 5899
rect 15887 5865 15896 5899
rect 15844 5856 15896 5865
rect 17316 5856 17368 5908
rect 11244 5720 11296 5772
rect 14096 5720 14148 5772
rect 14740 5763 14792 5772
rect 14740 5729 14749 5763
rect 14749 5729 14783 5763
rect 14783 5729 14792 5763
rect 14740 5720 14792 5729
rect 16396 5763 16448 5772
rect 16396 5729 16405 5763
rect 16405 5729 16439 5763
rect 16439 5729 16448 5763
rect 16396 5720 16448 5729
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 572 5627 624 5636
rect 572 5593 581 5627
rect 581 5593 615 5627
rect 615 5593 624 5627
rect 572 5584 624 5593
rect 7012 5584 7064 5636
rect 11888 5584 11940 5636
rect 13820 5584 13872 5636
rect 15016 5584 15068 5636
rect 16304 5652 16356 5704
rect 18144 5856 18196 5908
rect 2872 5516 2924 5568
rect 3700 5559 3752 5568
rect 3700 5525 3709 5559
rect 3709 5525 3743 5559
rect 3743 5525 3752 5559
rect 3700 5516 3752 5525
rect 8116 5516 8168 5568
rect 9772 5516 9824 5568
rect 15384 5516 15436 5568
rect 15844 5516 15896 5568
rect 4660 5414 4712 5466
rect 4724 5414 4776 5466
rect 4788 5414 4840 5466
rect 4852 5414 4904 5466
rect 4916 5414 4968 5466
rect 7760 5414 7812 5466
rect 7824 5414 7876 5466
rect 7888 5414 7940 5466
rect 7952 5414 8004 5466
rect 8016 5414 8068 5466
rect 10860 5414 10912 5466
rect 10924 5414 10976 5466
rect 10988 5414 11040 5466
rect 11052 5414 11104 5466
rect 11116 5414 11168 5466
rect 13960 5414 14012 5466
rect 14024 5414 14076 5466
rect 14088 5414 14140 5466
rect 14152 5414 14204 5466
rect 14216 5414 14268 5466
rect 17060 5414 17112 5466
rect 17124 5414 17176 5466
rect 17188 5414 17240 5466
rect 17252 5414 17304 5466
rect 17316 5414 17368 5466
rect 2504 5355 2556 5364
rect 2504 5321 2513 5355
rect 2513 5321 2547 5355
rect 2547 5321 2556 5355
rect 2504 5312 2556 5321
rect 3976 5312 4028 5364
rect 9772 5355 9824 5364
rect 9772 5321 9781 5355
rect 9781 5321 9815 5355
rect 9815 5321 9824 5355
rect 9772 5312 9824 5321
rect 9956 5312 10008 5364
rect 11336 5312 11388 5364
rect 11612 5312 11664 5364
rect 7012 5244 7064 5296
rect 8116 5244 8168 5296
rect 9128 5244 9180 5296
rect 11244 5244 11296 5296
rect 11888 5287 11940 5296
rect 11888 5253 11897 5287
rect 11897 5253 11931 5287
rect 11931 5253 11940 5287
rect 18144 5312 18196 5364
rect 11888 5244 11940 5253
rect 14280 5244 14332 5296
rect 15292 5244 15344 5296
rect 15660 5244 15712 5296
rect 15844 5244 15896 5296
rect 572 5176 624 5228
rect 2596 5176 2648 5228
rect 6000 5176 6052 5228
rect 7564 5219 7616 5228
rect 7564 5185 7573 5219
rect 7573 5185 7607 5219
rect 7607 5185 7616 5219
rect 7564 5176 7616 5185
rect 10600 5219 10652 5228
rect 10600 5185 10609 5219
rect 10609 5185 10643 5219
rect 10643 5185 10652 5219
rect 10600 5176 10652 5185
rect 14924 5219 14976 5228
rect 3700 5108 3752 5160
rect 8484 5108 8536 5160
rect 10048 5108 10100 5160
rect 10508 5108 10560 5160
rect 14924 5185 14933 5219
rect 14933 5185 14967 5219
rect 14967 5185 14976 5219
rect 14924 5176 14976 5185
rect 18512 5219 18564 5228
rect 18512 5185 18521 5219
rect 18521 5185 18555 5219
rect 18555 5185 18564 5219
rect 18512 5176 18564 5185
rect 13820 5151 13872 5160
rect 13820 5117 13829 5151
rect 13829 5117 13863 5151
rect 13863 5117 13872 5151
rect 13820 5108 13872 5117
rect 2504 4972 2556 5024
rect 4436 4972 4488 5024
rect 5448 4972 5500 5024
rect 7012 4972 7064 5024
rect 9036 4972 9088 5024
rect 16672 5015 16724 5024
rect 16672 4981 16681 5015
rect 16681 4981 16715 5015
rect 16715 4981 16724 5015
rect 16672 4972 16724 4981
rect 3110 4870 3162 4922
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 6210 4870 6262 4922
rect 6274 4870 6326 4922
rect 6338 4870 6390 4922
rect 6402 4870 6454 4922
rect 6466 4870 6518 4922
rect 9310 4870 9362 4922
rect 9374 4870 9426 4922
rect 9438 4870 9490 4922
rect 9502 4870 9554 4922
rect 9566 4870 9618 4922
rect 12410 4870 12462 4922
rect 12474 4870 12526 4922
rect 12538 4870 12590 4922
rect 12602 4870 12654 4922
rect 12666 4870 12718 4922
rect 15510 4870 15562 4922
rect 15574 4870 15626 4922
rect 15638 4870 15690 4922
rect 15702 4870 15754 4922
rect 15766 4870 15818 4922
rect 14372 4768 14424 4820
rect 14556 4768 14608 4820
rect 2964 4675 3016 4684
rect 2964 4641 2973 4675
rect 2973 4641 3007 4675
rect 3007 4641 3016 4675
rect 2964 4632 3016 4641
rect 11244 4700 11296 4752
rect 15292 4700 15344 4752
rect 6000 4632 6052 4684
rect 8300 4632 8352 4684
rect 8944 4675 8996 4684
rect 8944 4641 8953 4675
rect 8953 4641 8987 4675
rect 8987 4641 8996 4675
rect 8944 4632 8996 4641
rect 10048 4632 10100 4684
rect 11336 4675 11388 4684
rect 11336 4641 11345 4675
rect 11345 4641 11379 4675
rect 11379 4641 11388 4675
rect 11336 4632 11388 4641
rect 11428 4675 11480 4684
rect 11428 4641 11437 4675
rect 11437 4641 11471 4675
rect 11471 4641 11480 4675
rect 14740 4675 14792 4684
rect 11428 4632 11480 4641
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 15016 4675 15068 4684
rect 15016 4641 15025 4675
rect 15025 4641 15059 4675
rect 15059 4641 15068 4675
rect 15016 4632 15068 4641
rect 6184 4564 6236 4616
rect 6552 4564 6604 4616
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 9036 4607 9088 4616
rect 9036 4573 9045 4607
rect 9045 4573 9079 4607
rect 9079 4573 9088 4607
rect 9036 4564 9088 4573
rect 12256 4564 12308 4616
rect 4436 4496 4488 4548
rect 11336 4496 11388 4548
rect 14280 4496 14332 4548
rect 14648 4496 14700 4548
rect 15384 4539 15436 4548
rect 6092 4471 6144 4480
rect 6092 4437 6101 4471
rect 6101 4437 6135 4471
rect 6135 4437 6144 4471
rect 6092 4428 6144 4437
rect 6736 4471 6788 4480
rect 6736 4437 6745 4471
rect 6745 4437 6779 4471
rect 6779 4437 6788 4471
rect 6736 4428 6788 4437
rect 7656 4428 7708 4480
rect 13176 4428 13228 4480
rect 13728 4428 13780 4480
rect 14464 4428 14516 4480
rect 15384 4505 15393 4539
rect 15393 4505 15427 4539
rect 15427 4505 15436 4539
rect 15384 4496 15436 4505
rect 16672 4632 16724 4684
rect 15844 4607 15896 4616
rect 15844 4573 15853 4607
rect 15853 4573 15887 4607
rect 15887 4573 15896 4607
rect 15844 4564 15896 4573
rect 15752 4496 15804 4548
rect 16580 4496 16632 4548
rect 15936 4428 15988 4480
rect 4660 4326 4712 4378
rect 4724 4326 4776 4378
rect 4788 4326 4840 4378
rect 4852 4326 4904 4378
rect 4916 4326 4968 4378
rect 7760 4326 7812 4378
rect 7824 4326 7876 4378
rect 7888 4326 7940 4378
rect 7952 4326 8004 4378
rect 8016 4326 8068 4378
rect 10860 4326 10912 4378
rect 10924 4326 10976 4378
rect 10988 4326 11040 4378
rect 11052 4326 11104 4378
rect 11116 4326 11168 4378
rect 13960 4326 14012 4378
rect 14024 4326 14076 4378
rect 14088 4326 14140 4378
rect 14152 4326 14204 4378
rect 14216 4326 14268 4378
rect 17060 4326 17112 4378
rect 17124 4326 17176 4378
rect 17188 4326 17240 4378
rect 17252 4326 17304 4378
rect 17316 4326 17368 4378
rect 2504 4224 2556 4276
rect 2964 4267 3016 4276
rect 2964 4233 2973 4267
rect 2973 4233 3007 4267
rect 3007 4233 3016 4267
rect 2964 4224 3016 4233
rect 2596 4131 2648 4140
rect 2596 4097 2605 4131
rect 2605 4097 2639 4131
rect 2639 4097 2648 4131
rect 2596 4088 2648 4097
rect 296 4063 348 4072
rect 296 4029 305 4063
rect 305 4029 339 4063
rect 339 4029 348 4063
rect 296 4020 348 4029
rect 848 4020 900 4072
rect 2780 4131 2832 4140
rect 2780 4097 2789 4131
rect 2789 4097 2823 4131
rect 2823 4097 2832 4131
rect 2780 4088 2832 4097
rect 2688 3952 2740 4004
rect 3608 4063 3660 4072
rect 3608 4029 3617 4063
rect 3617 4029 3651 4063
rect 3651 4029 3660 4063
rect 3608 4020 3660 4029
rect 2320 3884 2372 3936
rect 4344 3884 4396 3936
rect 5540 4224 5592 4276
rect 6000 4224 6052 4276
rect 7656 4267 7708 4276
rect 7656 4233 7665 4267
rect 7665 4233 7699 4267
rect 7699 4233 7708 4267
rect 7656 4224 7708 4233
rect 8944 4224 8996 4276
rect 10048 4267 10100 4276
rect 10048 4233 10057 4267
rect 10057 4233 10091 4267
rect 10091 4233 10100 4267
rect 10048 4224 10100 4233
rect 11428 4224 11480 4276
rect 12164 4224 12216 4276
rect 13728 4224 13780 4276
rect 14648 4224 14700 4276
rect 14924 4224 14976 4276
rect 15844 4224 15896 4276
rect 5632 4156 5684 4208
rect 7012 4088 7064 4140
rect 8208 4088 8260 4140
rect 6092 4020 6144 4072
rect 8300 4020 8352 4072
rect 8760 4088 8812 4140
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 9864 4020 9916 4072
rect 10232 4063 10284 4072
rect 10232 4029 10241 4063
rect 10241 4029 10275 4063
rect 10275 4029 10284 4063
rect 10232 4020 10284 4029
rect 11336 4131 11388 4140
rect 11336 4097 11345 4131
rect 11345 4097 11379 4131
rect 11379 4097 11388 4131
rect 11336 4088 11388 4097
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 14556 4156 14608 4208
rect 15752 4156 15804 4208
rect 6000 3884 6052 3936
rect 7288 3927 7340 3936
rect 7288 3893 7297 3927
rect 7297 3893 7331 3927
rect 7331 3893 7340 3927
rect 7288 3884 7340 3893
rect 11336 3952 11388 4004
rect 12992 4020 13044 4072
rect 13728 4088 13780 4140
rect 15108 4088 15160 4140
rect 18512 4131 18564 4140
rect 18512 4097 18521 4131
rect 18521 4097 18555 4131
rect 18555 4097 18564 4131
rect 18512 4088 18564 4097
rect 13452 4020 13504 4072
rect 14372 4020 14424 4072
rect 14832 4063 14884 4072
rect 14832 4029 14841 4063
rect 14841 4029 14875 4063
rect 14875 4029 14884 4063
rect 14832 4020 14884 4029
rect 14556 3952 14608 4004
rect 8668 3884 8720 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 9128 3884 9180 3936
rect 12808 3884 12860 3936
rect 14096 3927 14148 3936
rect 14096 3893 14105 3927
rect 14105 3893 14139 3927
rect 14139 3893 14148 3927
rect 14096 3884 14148 3893
rect 16120 3884 16172 3936
rect 3110 3782 3162 3834
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 6210 3782 6262 3834
rect 6274 3782 6326 3834
rect 6338 3782 6390 3834
rect 6402 3782 6454 3834
rect 6466 3782 6518 3834
rect 9310 3782 9362 3834
rect 9374 3782 9426 3834
rect 9438 3782 9490 3834
rect 9502 3782 9554 3834
rect 9566 3782 9618 3834
rect 12410 3782 12462 3834
rect 12474 3782 12526 3834
rect 12538 3782 12590 3834
rect 12602 3782 12654 3834
rect 12666 3782 12718 3834
rect 15510 3782 15562 3834
rect 15574 3782 15626 3834
rect 15638 3782 15690 3834
rect 15702 3782 15754 3834
rect 15766 3782 15818 3834
rect 848 3723 900 3732
rect 848 3689 857 3723
rect 857 3689 891 3723
rect 891 3689 900 3723
rect 848 3680 900 3689
rect 6552 3680 6604 3732
rect 6736 3680 6788 3732
rect 8484 3723 8536 3732
rect 8484 3689 8493 3723
rect 8493 3689 8527 3723
rect 8527 3689 8536 3723
rect 8484 3680 8536 3689
rect 8576 3680 8628 3732
rect 13084 3680 13136 3732
rect 13544 3680 13596 3732
rect 2596 3612 2648 3664
rect 6828 3612 6880 3664
rect 8208 3612 8260 3664
rect 11244 3655 11296 3664
rect 2228 3587 2280 3596
rect 2228 3553 2237 3587
rect 2237 3553 2271 3587
rect 2271 3553 2280 3587
rect 2228 3544 2280 3553
rect 2320 3476 2372 3528
rect 2596 3476 2648 3528
rect 2780 3476 2832 3528
rect 6000 3544 6052 3596
rect 8760 3587 8812 3596
rect 8760 3553 8769 3587
rect 8769 3553 8803 3587
rect 8803 3553 8812 3587
rect 8760 3544 8812 3553
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 7288 3476 7340 3528
rect 8668 3519 8720 3528
rect 8668 3485 8677 3519
rect 8677 3485 8711 3519
rect 8711 3485 8720 3519
rect 8668 3476 8720 3485
rect 8944 3476 8996 3528
rect 11244 3621 11253 3655
rect 11253 3621 11287 3655
rect 11287 3621 11296 3655
rect 11244 3612 11296 3621
rect 12164 3612 12216 3664
rect 12532 3612 12584 3664
rect 11796 3544 11848 3596
rect 12348 3544 12400 3596
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 10416 3476 10468 3528
rect 11244 3476 11296 3528
rect 12716 3476 12768 3528
rect 14464 3680 14516 3732
rect 15108 3680 15160 3732
rect 15292 3680 15344 3732
rect 16120 3587 16172 3596
rect 16120 3553 16129 3587
rect 16129 3553 16163 3587
rect 16163 3553 16172 3587
rect 16120 3544 16172 3553
rect 17500 3587 17552 3596
rect 17500 3553 17509 3587
rect 17509 3553 17543 3587
rect 17543 3553 17552 3587
rect 17500 3544 17552 3553
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 13728 3519 13780 3528
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 13820 3519 13872 3528
rect 13820 3485 13829 3519
rect 13829 3485 13863 3519
rect 13863 3485 13872 3519
rect 13820 3476 13872 3485
rect 15844 3476 15896 3528
rect 3608 3408 3660 3460
rect 5264 3408 5316 3460
rect 7012 3408 7064 3460
rect 2228 3340 2280 3392
rect 3148 3383 3200 3392
rect 3148 3349 3157 3383
rect 3157 3349 3191 3383
rect 3191 3349 3200 3383
rect 3148 3340 3200 3349
rect 3516 3383 3568 3392
rect 3516 3349 3525 3383
rect 3525 3349 3559 3383
rect 3559 3349 3568 3383
rect 3516 3340 3568 3349
rect 5448 3340 5500 3392
rect 8300 3408 8352 3460
rect 7380 3340 7432 3392
rect 7472 3340 7524 3392
rect 9036 3408 9088 3460
rect 9956 3408 10008 3460
rect 11520 3451 11572 3460
rect 11520 3417 11529 3451
rect 11529 3417 11563 3451
rect 11563 3417 11572 3451
rect 11520 3408 11572 3417
rect 11796 3408 11848 3460
rect 14096 3451 14148 3460
rect 14096 3417 14130 3451
rect 14130 3417 14148 3451
rect 14096 3408 14148 3417
rect 9404 3340 9456 3392
rect 9772 3340 9824 3392
rect 11336 3383 11388 3392
rect 11336 3349 11345 3383
rect 11345 3349 11379 3383
rect 11379 3349 11388 3383
rect 11336 3340 11388 3349
rect 12532 3340 12584 3392
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 16580 3408 16632 3460
rect 12624 3340 12676 3349
rect 4660 3238 4712 3290
rect 4724 3238 4776 3290
rect 4788 3238 4840 3290
rect 4852 3238 4904 3290
rect 4916 3238 4968 3290
rect 7760 3238 7812 3290
rect 7824 3238 7876 3290
rect 7888 3238 7940 3290
rect 7952 3238 8004 3290
rect 8016 3238 8068 3290
rect 10860 3238 10912 3290
rect 10924 3238 10976 3290
rect 10988 3238 11040 3290
rect 11052 3238 11104 3290
rect 11116 3238 11168 3290
rect 13960 3238 14012 3290
rect 14024 3238 14076 3290
rect 14088 3238 14140 3290
rect 14152 3238 14204 3290
rect 14216 3238 14268 3290
rect 17060 3238 17112 3290
rect 17124 3238 17176 3290
rect 17188 3238 17240 3290
rect 17252 3238 17304 3290
rect 17316 3238 17368 3290
rect 1952 3136 2004 3188
rect 2504 3136 2556 3188
rect 5724 3136 5776 3188
rect 5264 3111 5316 3120
rect 5264 3077 5273 3111
rect 5273 3077 5307 3111
rect 5307 3077 5316 3111
rect 5264 3068 5316 3077
rect 5448 3111 5500 3120
rect 5448 3077 5457 3111
rect 5457 3077 5491 3111
rect 5491 3077 5500 3111
rect 5448 3068 5500 3077
rect 7380 3136 7432 3188
rect 8208 3136 8260 3188
rect 8576 3179 8628 3188
rect 8576 3145 8585 3179
rect 8585 3145 8619 3179
rect 8619 3145 8628 3179
rect 8576 3136 8628 3145
rect 8760 3136 8812 3188
rect 9956 3136 10008 3188
rect 10416 3179 10468 3188
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 6920 3068 6972 3120
rect 7196 3068 7248 3120
rect 8944 3068 8996 3120
rect 296 3043 348 3052
rect 296 3009 305 3043
rect 305 3009 339 3043
rect 339 3009 348 3043
rect 296 3000 348 3009
rect 2044 3000 2096 3052
rect 572 2975 624 2984
rect 572 2941 581 2975
rect 581 2941 615 2975
rect 615 2941 624 2975
rect 572 2932 624 2941
rect 2596 2932 2648 2984
rect 3148 2932 3200 2984
rect 5908 3000 5960 3052
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 9404 3000 9456 3052
rect 2872 2864 2924 2916
rect 3516 2864 3568 2916
rect 5724 2864 5776 2916
rect 5908 2864 5960 2916
rect 6092 2975 6144 2984
rect 6092 2941 6101 2975
rect 6101 2941 6135 2975
rect 6135 2941 6144 2975
rect 6092 2932 6144 2941
rect 6828 2932 6880 2984
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 5632 2796 5684 2848
rect 6828 2796 6880 2848
rect 7472 2796 7524 2848
rect 10232 3043 10284 3052
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 10600 3043 10652 3052
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 11796 3136 11848 3188
rect 11888 3136 11940 3188
rect 13544 3136 13596 3188
rect 11336 3068 11388 3120
rect 10784 3043 10836 3052
rect 10784 3009 10793 3043
rect 10793 3009 10827 3043
rect 10827 3009 10836 3043
rect 11152 3043 11204 3052
rect 10784 3000 10836 3009
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 11428 3043 11480 3052
rect 11428 3009 11437 3043
rect 11437 3009 11471 3043
rect 11471 3009 11480 3043
rect 11428 3000 11480 3009
rect 12624 3068 12676 3120
rect 14556 3068 14608 3120
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 13636 3000 13688 3052
rect 13820 3000 13872 3052
rect 14464 3043 14516 3052
rect 14464 3009 14473 3043
rect 14473 3009 14507 3043
rect 14507 3009 14516 3043
rect 14464 3000 14516 3009
rect 15384 3136 15436 3188
rect 15936 3179 15988 3188
rect 15936 3145 15945 3179
rect 15945 3145 15979 3179
rect 15979 3145 15988 3179
rect 15936 3136 15988 3145
rect 15200 3068 15252 3120
rect 16488 3111 16540 3120
rect 16488 3077 16497 3111
rect 16497 3077 16531 3111
rect 16531 3077 16540 3111
rect 16488 3068 16540 3077
rect 17500 3000 17552 3052
rect 17868 3000 17920 3052
rect 11704 2975 11756 2984
rect 11704 2941 11713 2975
rect 11713 2941 11747 2975
rect 11747 2941 11756 2975
rect 11704 2932 11756 2941
rect 10784 2864 10836 2916
rect 9864 2796 9916 2848
rect 14280 2975 14332 2984
rect 14280 2941 14289 2975
rect 14289 2941 14323 2975
rect 14323 2941 14332 2975
rect 14280 2932 14332 2941
rect 13820 2796 13872 2848
rect 15108 2796 15160 2848
rect 3110 2694 3162 2746
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 6210 2694 6262 2746
rect 6274 2694 6326 2746
rect 6338 2694 6390 2746
rect 6402 2694 6454 2746
rect 6466 2694 6518 2746
rect 9310 2694 9362 2746
rect 9374 2694 9426 2746
rect 9438 2694 9490 2746
rect 9502 2694 9554 2746
rect 9566 2694 9618 2746
rect 12410 2694 12462 2746
rect 12474 2694 12526 2746
rect 12538 2694 12590 2746
rect 12602 2694 12654 2746
rect 12666 2694 12718 2746
rect 15510 2694 15562 2746
rect 15574 2694 15626 2746
rect 15638 2694 15690 2746
rect 15702 2694 15754 2746
rect 15766 2694 15818 2746
rect 572 2592 624 2644
rect 2780 2635 2832 2644
rect 2780 2601 2789 2635
rect 2789 2601 2823 2635
rect 2823 2601 2832 2635
rect 2780 2592 2832 2601
rect 3516 2592 3568 2644
rect 5448 2592 5500 2644
rect 7196 2592 7248 2644
rect 11244 2592 11296 2644
rect 8760 2567 8812 2576
rect 2044 2499 2096 2508
rect 2044 2465 2053 2499
rect 2053 2465 2087 2499
rect 2087 2465 2096 2499
rect 2044 2456 2096 2465
rect 2228 2499 2280 2508
rect 2228 2465 2237 2499
rect 2237 2465 2271 2499
rect 2271 2465 2280 2499
rect 2228 2456 2280 2465
rect 8760 2533 8769 2567
rect 8769 2533 8803 2567
rect 8803 2533 8812 2567
rect 8760 2524 8812 2533
rect 10600 2524 10652 2576
rect 15292 2524 15344 2576
rect 2596 2388 2648 2440
rect 5540 2456 5592 2508
rect 9680 2456 9732 2508
rect 10784 2456 10836 2508
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 6092 2388 6144 2440
rect 2872 2320 2924 2372
rect 4344 2320 4396 2372
rect 5632 2363 5684 2372
rect 5632 2329 5641 2363
rect 5641 2329 5675 2363
rect 5675 2329 5684 2363
rect 5632 2320 5684 2329
rect 7472 2320 7524 2372
rect 8576 2363 8628 2372
rect 8576 2329 8585 2363
rect 8585 2329 8619 2363
rect 8619 2329 8628 2363
rect 8576 2320 8628 2329
rect 2780 2252 2832 2304
rect 4988 2252 5040 2304
rect 8300 2295 8352 2304
rect 8300 2261 8309 2295
rect 8309 2261 8343 2295
rect 8343 2261 8352 2295
rect 8300 2252 8352 2261
rect 10876 2431 10928 2440
rect 10876 2397 10885 2431
rect 10885 2397 10919 2431
rect 10919 2397 10928 2431
rect 10876 2388 10928 2397
rect 12808 2456 12860 2508
rect 14280 2456 14332 2508
rect 15568 2456 15620 2508
rect 15844 2499 15896 2508
rect 15844 2465 15853 2499
rect 15853 2465 15887 2499
rect 15887 2465 15896 2499
rect 15844 2456 15896 2465
rect 16488 2456 16540 2508
rect 9772 2252 9824 2304
rect 10140 2252 10192 2304
rect 11244 2320 11296 2372
rect 14556 2388 14608 2440
rect 11704 2320 11756 2372
rect 11888 2252 11940 2304
rect 12716 2252 12768 2304
rect 13636 2252 13688 2304
rect 14372 2252 14424 2304
rect 14924 2295 14976 2304
rect 14924 2261 14933 2295
rect 14933 2261 14967 2295
rect 14967 2261 14976 2295
rect 14924 2252 14976 2261
rect 15200 2320 15252 2372
rect 15292 2320 15344 2372
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 16120 2363 16172 2372
rect 16120 2329 16129 2363
rect 16129 2329 16163 2363
rect 16163 2329 16172 2363
rect 16120 2320 16172 2329
rect 16672 2320 16724 2372
rect 15844 2252 15896 2304
rect 4660 2150 4712 2202
rect 4724 2150 4776 2202
rect 4788 2150 4840 2202
rect 4852 2150 4904 2202
rect 4916 2150 4968 2202
rect 7760 2150 7812 2202
rect 7824 2150 7876 2202
rect 7888 2150 7940 2202
rect 7952 2150 8004 2202
rect 8016 2150 8068 2202
rect 10860 2150 10912 2202
rect 10924 2150 10976 2202
rect 10988 2150 11040 2202
rect 11052 2150 11104 2202
rect 11116 2150 11168 2202
rect 13960 2150 14012 2202
rect 14024 2150 14076 2202
rect 14088 2150 14140 2202
rect 14152 2150 14204 2202
rect 14216 2150 14268 2202
rect 17060 2150 17112 2202
rect 17124 2150 17176 2202
rect 17188 2150 17240 2202
rect 17252 2150 17304 2202
rect 17316 2150 17368 2202
rect 1952 1980 2004 2032
rect 2964 1912 3016 1964
rect 5540 1980 5592 2032
rect 296 1887 348 1896
rect 296 1853 305 1887
rect 305 1853 339 1887
rect 339 1853 348 1887
rect 296 1844 348 1853
rect 2780 1887 2832 1896
rect 2780 1853 2789 1887
rect 2789 1853 2823 1887
rect 2823 1853 2832 1887
rect 2780 1844 2832 1853
rect 1768 1776 1820 1828
rect 4344 1912 4396 1964
rect 4068 1844 4120 1896
rect 4988 1912 5040 1964
rect 5080 1912 5132 1964
rect 5448 1955 5500 1964
rect 5448 1921 5457 1955
rect 5457 1921 5491 1955
rect 5491 1921 5500 1955
rect 6092 2023 6144 2032
rect 6092 1989 6101 2023
rect 6101 1989 6135 2023
rect 6135 1989 6144 2023
rect 6092 1980 6144 1989
rect 9956 2048 10008 2100
rect 11428 2091 11480 2100
rect 11428 2057 11437 2091
rect 11437 2057 11471 2091
rect 11471 2057 11480 2091
rect 11428 2048 11480 2057
rect 13636 2048 13688 2100
rect 5448 1912 5500 1921
rect 6736 1955 6788 1964
rect 6736 1921 6745 1955
rect 6745 1921 6779 1955
rect 6779 1921 6788 1955
rect 6736 1912 6788 1921
rect 6828 1955 6880 1964
rect 6828 1921 6837 1955
rect 6837 1921 6871 1955
rect 6871 1921 6880 1955
rect 6828 1912 6880 1921
rect 7472 1955 7524 1964
rect 7472 1921 7481 1955
rect 7481 1921 7515 1955
rect 7515 1921 7524 1955
rect 7472 1912 7524 1921
rect 9680 1980 9732 2032
rect 9772 2023 9824 2032
rect 9772 1989 9781 2023
rect 9781 1989 9815 2023
rect 9815 1989 9824 2023
rect 15844 2048 15896 2100
rect 16120 2048 16172 2100
rect 17500 2048 17552 2100
rect 17868 2048 17920 2100
rect 18144 2091 18196 2100
rect 18144 2057 18153 2091
rect 18153 2057 18187 2091
rect 18187 2057 18196 2091
rect 18144 2048 18196 2057
rect 9772 1980 9824 1989
rect 7380 1844 7432 1896
rect 8576 1844 8628 1896
rect 9680 1844 9732 1896
rect 8300 1776 8352 1828
rect 9956 1955 10008 1964
rect 9956 1921 9965 1955
rect 9965 1921 9999 1955
rect 9999 1921 10008 1955
rect 9956 1912 10008 1921
rect 10232 1912 10284 1964
rect 11244 1912 11296 1964
rect 12716 1955 12768 1964
rect 12716 1921 12725 1955
rect 12725 1921 12759 1955
rect 12759 1921 12768 1955
rect 12716 1912 12768 1921
rect 12900 1912 12952 1964
rect 13544 1912 13596 1964
rect 10968 1887 11020 1896
rect 10968 1853 10977 1887
rect 10977 1853 11011 1887
rect 11011 1853 11020 1887
rect 10968 1844 11020 1853
rect 12808 1887 12860 1896
rect 12808 1853 12817 1887
rect 12817 1853 12851 1887
rect 12851 1853 12860 1887
rect 12808 1844 12860 1853
rect 13820 1844 13872 1896
rect 1952 1708 2004 1760
rect 2228 1751 2280 1760
rect 2228 1717 2237 1751
rect 2237 1717 2271 1751
rect 2271 1717 2280 1751
rect 2228 1708 2280 1717
rect 2504 1708 2556 1760
rect 4436 1751 4488 1760
rect 4436 1717 4445 1751
rect 4445 1717 4479 1751
rect 4479 1717 4488 1751
rect 4436 1708 4488 1717
rect 4528 1708 4580 1760
rect 5172 1708 5224 1760
rect 8668 1751 8720 1760
rect 8668 1717 8677 1751
rect 8677 1717 8711 1751
rect 8711 1717 8720 1751
rect 8668 1708 8720 1717
rect 9864 1776 9916 1828
rect 10140 1708 10192 1760
rect 12164 1708 12216 1760
rect 14372 1912 14424 1964
rect 14648 1912 14700 1964
rect 16672 1912 16724 1964
rect 16948 1912 17000 1964
rect 18236 1955 18288 1964
rect 18236 1921 18245 1955
rect 18245 1921 18279 1955
rect 18279 1921 18288 1955
rect 18236 1912 18288 1921
rect 15292 1844 15344 1896
rect 15568 1844 15620 1896
rect 14832 1776 14884 1828
rect 15384 1708 15436 1760
rect 15936 1708 15988 1760
rect 3110 1606 3162 1658
rect 3174 1606 3226 1658
rect 3238 1606 3290 1658
rect 3302 1606 3354 1658
rect 3366 1606 3418 1658
rect 6210 1606 6262 1658
rect 6274 1606 6326 1658
rect 6338 1606 6390 1658
rect 6402 1606 6454 1658
rect 6466 1606 6518 1658
rect 9310 1606 9362 1658
rect 9374 1606 9426 1658
rect 9438 1606 9490 1658
rect 9502 1606 9554 1658
rect 9566 1606 9618 1658
rect 12410 1606 12462 1658
rect 12474 1606 12526 1658
rect 12538 1606 12590 1658
rect 12602 1606 12654 1658
rect 12666 1606 12718 1658
rect 15510 1606 15562 1658
rect 15574 1606 15626 1658
rect 15638 1606 15690 1658
rect 15702 1606 15754 1658
rect 15766 1606 15818 1658
rect 10140 1504 10192 1556
rect 4068 1436 4120 1488
rect 5080 1436 5132 1488
rect 7472 1436 7524 1488
rect 4528 1368 4580 1420
rect 1768 1343 1820 1352
rect 1768 1309 1777 1343
rect 1777 1309 1811 1343
rect 1811 1309 1820 1343
rect 1768 1300 1820 1309
rect 4344 1300 4396 1352
rect 4528 1275 4580 1284
rect 4528 1241 4537 1275
rect 4537 1241 4571 1275
rect 4571 1241 4580 1275
rect 4528 1232 4580 1241
rect 4988 1300 5040 1352
rect 6736 1368 6788 1420
rect 5908 1343 5960 1352
rect 5908 1309 5917 1343
rect 5917 1309 5951 1343
rect 5951 1309 5960 1343
rect 5908 1300 5960 1309
rect 6000 1300 6052 1352
rect 7012 1343 7064 1352
rect 7012 1309 7021 1343
rect 7021 1309 7055 1343
rect 7055 1309 7064 1343
rect 7012 1300 7064 1309
rect 5264 1232 5316 1284
rect 7380 1300 7432 1352
rect 8668 1368 8720 1420
rect 8760 1368 8812 1420
rect 9036 1368 9088 1420
rect 14648 1504 14700 1556
rect 14924 1504 14976 1556
rect 15108 1436 15160 1488
rect 8576 1300 8628 1352
rect 8852 1343 8904 1352
rect 8852 1309 8861 1343
rect 8861 1309 8895 1343
rect 8895 1309 8904 1343
rect 8852 1300 8904 1309
rect 10416 1300 10468 1352
rect 10968 1300 11020 1352
rect 13820 1368 13872 1420
rect 5172 1164 5224 1216
rect 5356 1207 5408 1216
rect 5356 1173 5365 1207
rect 5365 1173 5399 1207
rect 5399 1173 5408 1207
rect 5356 1164 5408 1173
rect 5816 1207 5868 1216
rect 5816 1173 5825 1207
rect 5825 1173 5859 1207
rect 5859 1173 5868 1207
rect 5816 1164 5868 1173
rect 7564 1232 7616 1284
rect 10140 1232 10192 1284
rect 12348 1275 12400 1284
rect 12348 1241 12357 1275
rect 12357 1241 12391 1275
rect 12391 1241 12400 1275
rect 12348 1232 12400 1241
rect 13452 1300 13504 1352
rect 14464 1343 14516 1352
rect 14464 1309 14473 1343
rect 14473 1309 14507 1343
rect 14507 1309 14516 1343
rect 14464 1300 14516 1309
rect 15108 1343 15160 1352
rect 15108 1309 15117 1343
rect 15117 1309 15151 1343
rect 15151 1309 15160 1343
rect 15108 1300 15160 1309
rect 15200 1343 15252 1352
rect 15200 1309 15209 1343
rect 15209 1309 15243 1343
rect 15243 1309 15252 1343
rect 15200 1300 15252 1309
rect 15384 1300 15436 1352
rect 15936 1343 15988 1352
rect 15936 1309 15945 1343
rect 15945 1309 15979 1343
rect 15979 1309 15988 1343
rect 15936 1300 15988 1309
rect 16120 1300 16172 1352
rect 16396 1343 16448 1352
rect 16396 1309 16405 1343
rect 16405 1309 16439 1343
rect 16439 1309 16448 1343
rect 16396 1300 16448 1309
rect 14556 1232 14608 1284
rect 16672 1232 16724 1284
rect 17868 1275 17920 1284
rect 17868 1241 17877 1275
rect 17877 1241 17911 1275
rect 17911 1241 17920 1275
rect 17868 1232 17920 1241
rect 6920 1164 6972 1216
rect 8208 1207 8260 1216
rect 8208 1173 8217 1207
rect 8217 1173 8251 1207
rect 8251 1173 8260 1207
rect 8208 1164 8260 1173
rect 9404 1164 9456 1216
rect 11520 1164 11572 1216
rect 13360 1207 13412 1216
rect 13360 1173 13369 1207
rect 13369 1173 13403 1207
rect 13403 1173 13412 1207
rect 13360 1164 13412 1173
rect 16028 1164 16080 1216
rect 4660 1062 4712 1114
rect 4724 1062 4776 1114
rect 4788 1062 4840 1114
rect 4852 1062 4904 1114
rect 4916 1062 4968 1114
rect 7760 1062 7812 1114
rect 7824 1062 7876 1114
rect 7888 1062 7940 1114
rect 7952 1062 8004 1114
rect 8016 1062 8068 1114
rect 10860 1062 10912 1114
rect 10924 1062 10976 1114
rect 10988 1062 11040 1114
rect 11052 1062 11104 1114
rect 11116 1062 11168 1114
rect 13960 1062 14012 1114
rect 14024 1062 14076 1114
rect 14088 1062 14140 1114
rect 14152 1062 14204 1114
rect 14216 1062 14268 1114
rect 17060 1062 17112 1114
rect 17124 1062 17176 1114
rect 17188 1062 17240 1114
rect 17252 1062 17304 1114
rect 17316 1062 17368 1114
rect 4988 1003 5040 1012
rect 2504 867 2556 876
rect 2504 833 2513 867
rect 2513 833 2547 867
rect 2547 833 2556 867
rect 2504 824 2556 833
rect 4436 892 4488 944
rect 4988 969 4997 1003
rect 4997 969 5031 1003
rect 5031 969 5040 1003
rect 4988 960 5040 969
rect 5908 960 5960 1012
rect 7380 1003 7432 1012
rect 4344 824 4396 876
rect 5448 892 5500 944
rect 7380 969 7389 1003
rect 7389 969 7423 1003
rect 7423 969 7432 1003
rect 7380 960 7432 969
rect 7564 960 7616 1012
rect 4712 867 4764 876
rect 4712 833 4721 867
rect 4721 833 4755 867
rect 4755 833 4764 867
rect 4712 824 4764 833
rect 4896 867 4948 876
rect 4896 833 4905 867
rect 4905 833 4939 867
rect 4939 833 4948 867
rect 5080 867 5132 876
rect 4896 824 4948 833
rect 5080 833 5089 867
rect 5089 833 5123 867
rect 5123 833 5132 867
rect 5080 824 5132 833
rect 7288 867 7340 876
rect 5632 799 5684 808
rect 5632 765 5641 799
rect 5641 765 5675 799
rect 5675 765 5684 799
rect 5632 756 5684 765
rect 7288 833 7297 867
rect 7297 833 7331 867
rect 7331 833 7340 867
rect 7288 824 7340 833
rect 7472 867 7524 876
rect 7472 833 7481 867
rect 7481 833 7515 867
rect 7515 833 7524 867
rect 7472 824 7524 833
rect 7748 867 7800 876
rect 7748 833 7757 867
rect 7757 833 7791 867
rect 7791 833 7800 867
rect 7748 824 7800 833
rect 8208 867 8260 876
rect 8208 833 8217 867
rect 8217 833 8251 867
rect 8251 833 8260 867
rect 8208 824 8260 833
rect 8944 960 8996 1012
rect 9404 1003 9456 1012
rect 9404 969 9413 1003
rect 9413 969 9447 1003
rect 9447 969 9456 1003
rect 9404 960 9456 969
rect 8576 892 8628 944
rect 8760 867 8812 876
rect 8760 833 8769 867
rect 8769 833 8803 867
rect 8803 833 8812 867
rect 8760 824 8812 833
rect 9680 892 9732 944
rect 11520 935 11572 944
rect 11520 901 11529 935
rect 11529 901 11563 935
rect 11563 901 11572 935
rect 11520 892 11572 901
rect 12348 960 12400 1012
rect 13544 960 13596 1012
rect 16672 1003 16724 1012
rect 9312 867 9364 876
rect 9312 833 9321 867
rect 9321 833 9355 867
rect 9355 833 9364 867
rect 9312 824 9364 833
rect 10140 867 10192 876
rect 5356 688 5408 740
rect 2228 620 2280 672
rect 4344 620 4396 672
rect 8300 756 8352 808
rect 10140 833 10149 867
rect 10149 833 10183 867
rect 10183 833 10192 867
rect 10140 824 10192 833
rect 10416 867 10468 876
rect 10416 833 10425 867
rect 10425 833 10459 867
rect 10459 833 10468 867
rect 10416 824 10468 833
rect 10232 756 10284 808
rect 11704 867 11756 876
rect 11704 833 11713 867
rect 11713 833 11747 867
rect 11747 833 11756 867
rect 11704 824 11756 833
rect 11796 867 11848 876
rect 11796 833 11805 867
rect 11805 833 11839 867
rect 11839 833 11848 867
rect 11796 824 11848 833
rect 12164 824 12216 876
rect 12992 867 13044 876
rect 12992 833 13001 867
rect 13001 833 13035 867
rect 13035 833 13044 867
rect 12992 824 13044 833
rect 14832 892 14884 944
rect 16672 969 16681 1003
rect 16681 969 16715 1003
rect 16715 969 16724 1003
rect 16672 960 16724 969
rect 16948 960 17000 1012
rect 17500 1003 17552 1012
rect 17500 969 17509 1003
rect 17509 969 17543 1003
rect 17543 969 17552 1003
rect 17500 960 17552 969
rect 18236 960 18288 1012
rect 13268 824 13320 876
rect 13728 867 13780 876
rect 13728 833 13737 867
rect 13737 833 13771 867
rect 13771 833 13780 867
rect 13728 824 13780 833
rect 17316 824 17368 876
rect 18512 867 18564 876
rect 18512 833 18521 867
rect 18521 833 18555 867
rect 18555 833 18564 867
rect 18512 824 18564 833
rect 9680 731 9732 740
rect 9680 697 9689 731
rect 9689 697 9723 731
rect 9723 697 9732 731
rect 9680 688 9732 697
rect 13544 756 13596 808
rect 14280 799 14332 808
rect 14280 765 14289 799
rect 14289 765 14323 799
rect 14323 765 14332 799
rect 14280 756 14332 765
rect 14556 756 14608 808
rect 16212 756 16264 808
rect 17592 799 17644 808
rect 17592 765 17601 799
rect 17601 765 17635 799
rect 17635 765 17644 799
rect 17592 756 17644 765
rect 11796 688 11848 740
rect 12900 731 12952 740
rect 12900 697 12909 731
rect 12909 697 12943 731
rect 12943 697 12952 731
rect 12900 688 12952 697
rect 14464 688 14516 740
rect 9128 620 9180 672
rect 9956 663 10008 672
rect 9956 629 9965 663
rect 9965 629 9999 663
rect 9999 629 10008 663
rect 9956 620 10008 629
rect 16488 663 16540 672
rect 16488 629 16497 663
rect 16497 629 16531 663
rect 16531 629 16540 663
rect 16488 620 16540 629
rect 3110 518 3162 570
rect 3174 518 3226 570
rect 3238 518 3290 570
rect 3302 518 3354 570
rect 3366 518 3418 570
rect 6210 518 6262 570
rect 6274 518 6326 570
rect 6338 518 6390 570
rect 6402 518 6454 570
rect 6466 518 6518 570
rect 9310 518 9362 570
rect 9374 518 9426 570
rect 9438 518 9490 570
rect 9502 518 9554 570
rect 9566 518 9618 570
rect 12410 518 12462 570
rect 12474 518 12526 570
rect 12538 518 12590 570
rect 12602 518 12654 570
rect 12666 518 12718 570
rect 15510 518 15562 570
rect 15574 518 15626 570
rect 15638 518 15690 570
rect 15702 518 15754 570
rect 15766 518 15818 570
rect 5632 416 5684 468
rect 7288 416 7340 468
rect 8852 416 8904 468
rect 13452 459 13504 468
rect 13452 425 13461 459
rect 13461 425 13495 459
rect 13495 425 13504 459
rect 13452 416 13504 425
rect 13544 459 13596 468
rect 13544 425 13553 459
rect 13553 425 13587 459
rect 13587 425 13596 459
rect 13544 416 13596 425
rect 15200 416 15252 468
rect 16120 416 16172 468
rect 17316 459 17368 468
rect 17316 425 17325 459
rect 17325 425 17359 459
rect 17359 425 17368 459
rect 17316 416 17368 425
rect 12256 391 12308 400
rect 12256 357 12265 391
rect 12265 357 12299 391
rect 12299 357 12308 391
rect 12256 348 12308 357
rect 16396 348 16448 400
rect 5816 280 5868 332
rect 5172 212 5224 264
rect 5908 255 5960 264
rect 5908 221 5917 255
rect 5917 221 5951 255
rect 5951 221 5960 255
rect 5908 212 5960 221
rect 9128 255 9180 264
rect 4712 144 4764 196
rect 9128 221 9137 255
rect 9137 221 9171 255
rect 9171 221 9180 255
rect 9128 212 9180 221
rect 9956 212 10008 264
rect 11796 212 11848 264
rect 13268 255 13320 264
rect 13268 221 13277 255
rect 13277 221 13311 255
rect 13311 221 13320 255
rect 13268 212 13320 221
rect 16488 280 16540 332
rect 13728 255 13780 264
rect 9036 144 9088 196
rect 11704 144 11756 196
rect 12992 144 13044 196
rect 13728 221 13737 255
rect 13737 221 13771 255
rect 13771 221 13780 255
rect 13728 212 13780 221
rect 15844 255 15896 264
rect 15844 221 15853 255
rect 15853 221 15887 255
rect 15887 221 15896 255
rect 15844 212 15896 221
rect 16028 255 16080 264
rect 16028 221 16037 255
rect 16037 221 16071 255
rect 16071 221 16080 255
rect 16028 212 16080 221
rect 16212 255 16264 264
rect 16212 221 16221 255
rect 16221 221 16255 255
rect 16255 221 16264 255
rect 16212 212 16264 221
rect 17868 212 17920 264
rect 14464 144 14516 196
rect 5356 76 5408 128
rect 4660 -26 4712 26
rect 4724 -26 4776 26
rect 4788 -26 4840 26
rect 4852 -26 4904 26
rect 4916 -26 4968 26
rect 7760 -26 7812 26
rect 7824 -26 7876 26
rect 7888 -26 7940 26
rect 7952 -26 8004 26
rect 8016 -26 8068 26
rect 10860 -26 10912 26
rect 10924 -26 10976 26
rect 10988 -26 11040 26
rect 11052 -26 11104 26
rect 11116 -26 11168 26
rect 13960 -26 14012 26
rect 14024 -26 14076 26
rect 14088 -26 14140 26
rect 14152 -26 14204 26
rect 14216 -26 14268 26
rect 17060 -26 17112 26
rect 17124 -26 17176 26
rect 17188 -26 17240 26
rect 17252 -26 17304 26
rect 17316 -26 17368 26
<< metal2 >>
rect 1398 11200 1454 12000
rect 4250 11200 4306 12000
rect 7102 11200 7158 12000
rect 9954 11200 10010 12000
rect 12806 11200 12862 12000
rect 15396 11206 15608 11234
rect 296 10668 348 10674
rect 296 10610 348 10616
rect 308 9518 336 10610
rect 1308 10464 1360 10470
rect 1308 10406 1360 10412
rect 1320 10130 1348 10406
rect 1308 10124 1360 10130
rect 1308 10066 1360 10072
rect 296 9512 348 9518
rect 296 9454 348 9460
rect 308 8430 336 9454
rect 1412 9178 1440 11200
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 1952 9648 2004 9654
rect 1952 9590 2004 9596
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1412 8974 1440 9114
rect 1964 9042 1992 9590
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1964 8838 1992 8978
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1964 8566 1992 8774
rect 2148 8634 2176 9522
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 1952 8560 2004 8566
rect 1952 8502 2004 8508
rect 296 8424 348 8430
rect 296 8366 348 8372
rect 308 7342 336 8366
rect 1964 7478 1992 8502
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2148 8090 2176 8434
rect 2240 8362 2268 9862
rect 2502 9616 2558 9625
rect 2332 9560 2502 9568
rect 2332 9540 2504 9560
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2148 7970 2176 8026
rect 2056 7942 2176 7970
rect 2240 7954 2268 8298
rect 2228 7948 2280 7954
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 296 7336 348 7342
rect 296 7278 348 7284
rect 572 7336 624 7342
rect 572 7278 624 7284
rect 308 6254 336 7278
rect 584 6730 612 7278
rect 1964 7002 1992 7414
rect 2056 7410 2084 7942
rect 2228 7890 2280 7896
rect 2332 7886 2360 9540
rect 2556 9551 2558 9560
rect 2504 9522 2556 9528
rect 2608 9330 2636 10066
rect 2700 9994 2728 10474
rect 3110 10364 3418 10384
rect 3110 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3276 10364
rect 3332 10362 3356 10364
rect 3412 10362 3418 10364
rect 3172 10310 3174 10362
rect 3354 10310 3356 10362
rect 3110 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3276 10310
rect 3332 10308 3356 10310
rect 3412 10308 3418 10310
rect 3110 10288 3418 10308
rect 3528 10266 3556 10542
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 4172 10130 4200 10610
rect 4160 10124 4212 10130
rect 4160 10066 4212 10072
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 4080 9654 4108 9930
rect 4172 9722 4200 10066
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 2688 9648 2740 9654
rect 3056 9648 3108 9654
rect 2740 9608 3056 9636
rect 2688 9590 2740 9596
rect 2688 9376 2740 9382
rect 2608 9324 2688 9330
rect 2608 9318 2740 9324
rect 2608 9302 2728 9318
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2412 8424 2464 8430
rect 2412 8366 2464 8372
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2148 7546 2176 7822
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 572 6724 624 6730
rect 572 6666 624 6672
rect 1964 6458 1992 6938
rect 2332 6934 2360 7822
rect 2424 7546 2452 8366
rect 2516 7954 2544 8774
rect 2700 8498 2728 8910
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2700 8090 2728 8434
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2792 8022 2820 8434
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2516 7410 2544 7686
rect 2884 7478 2912 9608
rect 4068 9648 4120 9654
rect 3108 9608 3188 9636
rect 3056 9590 3108 9596
rect 3056 9512 3108 9518
rect 2976 9472 3056 9500
rect 2976 9178 3004 9472
rect 3160 9489 3188 9608
rect 4068 9590 4120 9596
rect 3056 9454 3108 9460
rect 3146 9480 3202 9489
rect 3146 9415 3202 9424
rect 3608 9444 3660 9450
rect 3608 9386 3660 9392
rect 3110 9276 3418 9296
rect 3110 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3276 9276
rect 3332 9274 3356 9276
rect 3412 9274 3418 9276
rect 3172 9222 3174 9274
rect 3354 9222 3356 9274
rect 3110 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3276 9222
rect 3332 9220 3356 9222
rect 3412 9220 3418 9222
rect 3110 9200 3418 9220
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 3620 8838 3648 9386
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4172 8634 4200 8774
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4068 8560 4120 8566
rect 4068 8502 4120 8508
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 4080 8242 4108 8502
rect 2976 7886 3004 8230
rect 4080 8214 4200 8242
rect 3110 8188 3418 8208
rect 3110 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3276 8188
rect 3332 8186 3356 8188
rect 3412 8186 3418 8188
rect 3172 8134 3174 8186
rect 3354 8134 3356 8186
rect 3110 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3276 8134
rect 3332 8132 3356 8134
rect 3412 8132 3418 8134
rect 3110 8112 3418 8132
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 3528 7410 3556 7890
rect 4172 7750 4200 8214
rect 4264 8090 4292 11200
rect 4660 10908 4968 10928
rect 4660 10906 4666 10908
rect 4722 10906 4746 10908
rect 4802 10906 4826 10908
rect 4882 10906 4906 10908
rect 4962 10906 4968 10908
rect 4722 10854 4724 10906
rect 4904 10854 4906 10906
rect 4660 10852 4666 10854
rect 4722 10852 4746 10854
rect 4802 10852 4826 10854
rect 4882 10852 4906 10854
rect 4962 10852 4968 10854
rect 4660 10832 4968 10852
rect 7116 10810 7144 11200
rect 7760 10908 8068 10928
rect 7760 10906 7766 10908
rect 7822 10906 7846 10908
rect 7902 10906 7926 10908
rect 7982 10906 8006 10908
rect 8062 10906 8068 10908
rect 7822 10854 7824 10906
rect 8004 10854 8006 10906
rect 7760 10852 7766 10854
rect 7822 10852 7846 10854
rect 7902 10852 7926 10854
rect 7982 10852 8006 10854
rect 8062 10852 8068 10854
rect 7760 10832 8068 10852
rect 9968 10810 9996 11200
rect 10860 10908 11168 10928
rect 10860 10906 10866 10908
rect 10922 10906 10946 10908
rect 11002 10906 11026 10908
rect 11082 10906 11106 10908
rect 11162 10906 11168 10908
rect 10922 10854 10924 10906
rect 11104 10854 11106 10906
rect 10860 10852 10866 10854
rect 10922 10852 10946 10854
rect 11002 10852 11026 10854
rect 11082 10852 11106 10854
rect 11162 10852 11168 10854
rect 10860 10832 11168 10852
rect 12820 10810 12848 11200
rect 13960 10908 14268 10928
rect 13960 10906 13966 10908
rect 14022 10906 14046 10908
rect 14102 10906 14126 10908
rect 14182 10906 14206 10908
rect 14262 10906 14268 10908
rect 14022 10854 14024 10906
rect 14204 10854 14206 10906
rect 13960 10852 13966 10854
rect 14022 10852 14046 10854
rect 14102 10852 14126 10854
rect 14182 10852 14206 10854
rect 14262 10852 14268 10854
rect 13960 10832 14268 10852
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 11336 10736 11388 10742
rect 11336 10678 11388 10684
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4356 9518 4384 10134
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4448 8974 4476 10406
rect 6210 10364 6518 10384
rect 6210 10362 6216 10364
rect 6272 10362 6296 10364
rect 6352 10362 6376 10364
rect 6432 10362 6456 10364
rect 6512 10362 6518 10364
rect 6272 10310 6274 10362
rect 6454 10310 6456 10362
rect 6210 10308 6216 10310
rect 6272 10308 6296 10310
rect 6352 10308 6376 10310
rect 6432 10308 6456 10310
rect 6512 10308 6518 10310
rect 6210 10288 6518 10308
rect 4896 10192 4948 10198
rect 4896 10134 4948 10140
rect 4908 10062 4936 10134
rect 5448 10124 5500 10130
rect 5368 10084 5448 10112
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4540 9586 4568 9862
rect 4660 9820 4968 9840
rect 4660 9818 4666 9820
rect 4722 9818 4746 9820
rect 4802 9818 4826 9820
rect 4882 9818 4906 9820
rect 4962 9818 4968 9820
rect 4722 9766 4724 9818
rect 4904 9766 4906 9818
rect 4660 9764 4666 9766
rect 4722 9764 4746 9766
rect 4802 9764 4826 9766
rect 4882 9764 4906 9766
rect 4962 9764 4968 9766
rect 4660 9744 4968 9764
rect 5368 9654 5396 10084
rect 5448 10066 5500 10072
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 5356 9648 5408 9654
rect 5552 9625 5580 9998
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5736 9654 5764 9862
rect 6196 9654 6224 9998
rect 6380 9654 6408 10066
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6472 9722 6500 9998
rect 7024 9994 7052 10474
rect 7668 10266 7696 10610
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 8680 10062 8708 10406
rect 8772 10198 8800 10542
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 7012 9988 7064 9994
rect 7012 9930 7064 9936
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 6460 9716 6512 9722
rect 6460 9658 6512 9664
rect 5724 9648 5776 9654
rect 5356 9590 5408 9596
rect 5538 9616 5594 9625
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 5448 9580 5500 9586
rect 5724 9590 5776 9596
rect 6184 9648 6236 9654
rect 6184 9590 6236 9596
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 7668 9586 7696 9862
rect 7760 9820 8068 9840
rect 7760 9818 7766 9820
rect 7822 9818 7846 9820
rect 7902 9818 7926 9820
rect 7982 9818 8006 9820
rect 8062 9818 8068 9820
rect 7822 9766 7824 9818
rect 8004 9766 8006 9818
rect 7760 9764 7766 9766
rect 7822 9764 7846 9766
rect 7902 9764 7926 9766
rect 7982 9764 8006 9766
rect 8062 9764 8068 9766
rect 7760 9744 8068 9764
rect 8496 9654 8524 9862
rect 8956 9722 8984 10610
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9232 9994 9260 10406
rect 9310 10364 9618 10384
rect 9310 10362 9316 10364
rect 9372 10362 9396 10364
rect 9452 10362 9476 10364
rect 9532 10362 9556 10364
rect 9612 10362 9618 10364
rect 9372 10310 9374 10362
rect 9554 10310 9556 10362
rect 9310 10308 9316 10310
rect 9372 10308 9396 10310
rect 9452 10308 9476 10310
rect 9532 10308 9556 10310
rect 9612 10308 9618 10310
rect 9310 10288 9618 10308
rect 10704 10198 10732 10474
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 9692 9654 9720 9930
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 5538 9551 5594 9560
rect 6092 9580 6144 9586
rect 5448 9522 5500 9528
rect 6092 9522 6144 9528
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 4540 9042 4568 9522
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4356 8634 4384 8842
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4448 8566 4476 8774
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4540 8498 4568 8978
rect 5276 8974 5304 9318
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 4660 8732 4968 8752
rect 4660 8730 4666 8732
rect 4722 8730 4746 8732
rect 4802 8730 4826 8732
rect 4882 8730 4906 8732
rect 4962 8730 4968 8732
rect 4722 8678 4724 8730
rect 4904 8678 4906 8730
rect 4660 8676 4666 8678
rect 4722 8676 4746 8678
rect 4802 8676 4826 8678
rect 4882 8676 4906 8678
rect 4962 8676 4968 8678
rect 4660 8656 4968 8676
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 5000 8430 5028 8910
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5276 8634 5304 8774
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 5000 7886 5028 8366
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5080 8016 5132 8022
rect 5080 7958 5132 7964
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 4068 7404 4120 7410
rect 4172 7392 4200 7686
rect 4660 7644 4968 7664
rect 4660 7642 4666 7644
rect 4722 7642 4746 7644
rect 4802 7642 4826 7644
rect 4882 7642 4906 7644
rect 4962 7642 4968 7644
rect 4722 7590 4724 7642
rect 4904 7590 4906 7642
rect 4660 7588 4666 7590
rect 4722 7588 4746 7590
rect 4802 7588 4826 7590
rect 4882 7588 4906 7590
rect 4962 7588 4968 7590
rect 4660 7568 4968 7588
rect 5000 7528 5028 7822
rect 4908 7500 5028 7528
rect 4908 7410 4936 7500
rect 4252 7404 4304 7410
rect 4172 7364 4252 7392
rect 4068 7346 4120 7352
rect 4252 7346 4304 7352
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4988 7404 5040 7410
rect 5092 7392 5120 7958
rect 5040 7364 5120 7392
rect 4988 7346 5040 7352
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2320 6928 2372 6934
rect 2320 6870 2372 6876
rect 2976 6798 3004 7142
rect 3110 7100 3418 7120
rect 3110 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3276 7100
rect 3332 7098 3356 7100
rect 3412 7098 3418 7100
rect 3172 7046 3174 7098
rect 3354 7046 3356 7098
rect 3110 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3276 7046
rect 3332 7044 3356 7046
rect 3412 7044 3418 7046
rect 3110 7024 3418 7044
rect 3528 6984 3556 7346
rect 3436 6956 3556 6984
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 1952 6452 2004 6458
rect 1952 6394 2004 6400
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 296 6248 348 6254
rect 296 6190 348 6196
rect 572 6248 624 6254
rect 572 6190 624 6196
rect 308 5778 336 6190
rect 584 5914 612 6190
rect 572 5908 624 5914
rect 572 5850 624 5856
rect 296 5772 348 5778
rect 296 5714 348 5720
rect 572 5636 624 5642
rect 572 5578 624 5584
rect 584 5234 612 5578
rect 2516 5370 2544 6394
rect 2608 6322 2636 6598
rect 2792 6458 2820 6666
rect 2780 6452 2832 6458
rect 2884 6440 2912 6734
rect 2964 6452 3016 6458
rect 2884 6412 2964 6440
rect 2780 6394 2832 6400
rect 2964 6394 3016 6400
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 572 5228 624 5234
rect 572 5170 624 5176
rect 2516 5030 2544 5306
rect 2608 5234 2636 6258
rect 2792 5710 2820 6394
rect 3436 6361 3464 6956
rect 4080 6866 4108 7346
rect 4264 6934 4292 7346
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4908 6798 4936 7346
rect 5092 6798 5120 7364
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 4660 6556 4968 6576
rect 4660 6554 4666 6556
rect 4722 6554 4746 6556
rect 4802 6554 4826 6556
rect 4882 6554 4906 6556
rect 4962 6554 4968 6556
rect 4722 6502 4724 6554
rect 4904 6502 4906 6554
rect 4660 6500 4666 6502
rect 4722 6500 4746 6502
rect 4802 6500 4826 6502
rect 4882 6500 4906 6502
rect 4962 6500 4968 6502
rect 4660 6480 4968 6500
rect 3700 6452 3752 6458
rect 3700 6394 3752 6400
rect 3516 6384 3568 6390
rect 3422 6352 3478 6361
rect 3516 6326 3568 6332
rect 3422 6287 3424 6296
rect 3476 6287 3478 6296
rect 3424 6258 3476 6264
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2884 5574 2912 6054
rect 2976 5710 3004 6190
rect 3110 6012 3418 6032
rect 3110 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3276 6012
rect 3332 6010 3356 6012
rect 3412 6010 3418 6012
rect 3172 5958 3174 6010
rect 3354 5958 3356 6010
rect 3110 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3276 5958
rect 3332 5956 3356 5958
rect 3412 5956 3418 5958
rect 3110 5936 3418 5956
rect 3424 5840 3476 5846
rect 3528 5794 3556 6326
rect 3476 5788 3556 5794
rect 3424 5782 3556 5788
rect 3436 5766 3556 5782
rect 3712 5778 3740 6394
rect 5184 6361 5212 8298
rect 5368 8022 5396 8502
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5276 7478 5304 7890
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5276 7018 5304 7414
rect 5368 7410 5396 7754
rect 5460 7546 5488 9522
rect 6000 9512 6052 9518
rect 5998 9480 6000 9489
rect 6052 9480 6054 9489
rect 5998 9415 6054 9424
rect 6104 8974 6132 9522
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 6210 9276 6518 9296
rect 6210 9274 6216 9276
rect 6272 9274 6296 9276
rect 6352 9274 6376 9276
rect 6432 9274 6456 9276
rect 6512 9274 6518 9276
rect 6272 9222 6274 9274
rect 6454 9222 6456 9274
rect 6210 9220 6216 9222
rect 6272 9220 6296 9222
rect 6352 9220 6376 9222
rect 6432 9220 6456 9222
rect 6512 9220 6518 9222
rect 6210 9200 6518 9220
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6104 8294 6132 8910
rect 7472 8560 7524 8566
rect 7472 8502 7524 8508
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6104 7886 6132 8230
rect 6210 8188 6518 8208
rect 6210 8186 6216 8188
rect 6272 8186 6296 8188
rect 6352 8186 6376 8188
rect 6432 8186 6456 8188
rect 6512 8186 6518 8188
rect 6272 8134 6274 8186
rect 6454 8134 6456 8186
rect 6210 8132 6216 8134
rect 6272 8132 6296 8134
rect 6352 8132 6376 8134
rect 6432 8132 6456 8134
rect 6512 8132 6518 8134
rect 6210 8112 6518 8132
rect 7300 7954 7328 8434
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5276 6990 5396 7018
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5276 6458 5304 6870
rect 5368 6866 5396 6990
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5170 6352 5226 6361
rect 5170 6287 5226 6296
rect 5184 6254 5212 6287
rect 5460 6254 5488 7482
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 5552 5914 5580 7142
rect 5644 7018 5672 7278
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5644 6990 5764 7018
rect 5736 6798 5764 6990
rect 5828 6934 5856 7210
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5644 6322 5672 6734
rect 5736 6458 5764 6734
rect 5920 6458 5948 7278
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6012 5914 6040 6258
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6104 5778 6132 7822
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6210 7100 6518 7120
rect 6210 7098 6216 7100
rect 6272 7098 6296 7100
rect 6352 7098 6376 7100
rect 6432 7098 6456 7100
rect 6512 7098 6518 7100
rect 6272 7046 6274 7098
rect 6454 7046 6456 7098
rect 6210 7044 6216 7046
rect 6272 7044 6296 7046
rect 6352 7044 6376 7046
rect 6432 7044 6456 7046
rect 6512 7044 6518 7046
rect 6210 7024 6518 7044
rect 6564 6390 6592 7754
rect 6656 7342 6684 7890
rect 7484 7886 7512 8502
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6656 6458 6684 7278
rect 6932 7002 6960 7346
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6210 6012 6518 6032
rect 6210 6010 6216 6012
rect 6272 6010 6296 6012
rect 6352 6010 6376 6012
rect 6432 6010 6456 6012
rect 6512 6010 6518 6012
rect 6272 5958 6274 6010
rect 6454 5958 6456 6010
rect 6210 5956 6216 5958
rect 6272 5956 6296 5958
rect 6352 5956 6376 5958
rect 6432 5956 6456 5958
rect 6512 5956 6518 5958
rect 6210 5936 6518 5956
rect 6840 5778 6868 6598
rect 7116 6186 7144 7346
rect 7208 6662 7236 7482
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7392 6866 7420 7142
rect 7484 7002 7512 7822
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7484 6746 7512 6802
rect 7392 6718 7512 6746
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7392 6254 7420 6718
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7484 6458 7512 6598
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7104 6180 7156 6186
rect 7104 6122 7156 6128
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 3712 5166 3740 5510
rect 3988 5370 4016 5646
rect 4660 5468 4968 5488
rect 4660 5466 4666 5468
rect 4722 5466 4746 5468
rect 4802 5466 4826 5468
rect 4882 5466 4906 5468
rect 4962 5466 4968 5468
rect 4722 5414 4724 5466
rect 4904 5414 4906 5466
rect 4660 5412 4666 5414
rect 4722 5412 4746 5414
rect 4802 5412 4826 5414
rect 4882 5412 4906 5414
rect 4962 5412 4968 5414
rect 4660 5392 4968 5412
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 5460 5030 5488 5646
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 7024 5302 7052 5578
rect 7012 5296 7064 5302
rect 7012 5238 7064 5244
rect 6000 5228 6052 5234
rect 6000 5170 6052 5176
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 2516 4282 2544 4966
rect 3110 4924 3418 4944
rect 3110 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3276 4924
rect 3332 4922 3356 4924
rect 3412 4922 3418 4924
rect 3172 4870 3174 4922
rect 3354 4870 3356 4922
rect 3110 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3276 4870
rect 3332 4868 3356 4870
rect 3412 4868 3418 4870
rect 3110 4848 3418 4868
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2976 4282 3004 4626
rect 4448 4554 4476 4966
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 296 4072 348 4078
rect 296 4014 348 4020
rect 848 4072 900 4078
rect 848 4014 900 4020
rect 308 3058 336 4014
rect 860 3738 888 4014
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 848 3732 900 3738
rect 848 3674 900 3680
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2240 3398 2268 3538
rect 2332 3534 2360 3878
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 296 3052 348 3058
rect 296 2994 348 3000
rect 308 1902 336 2994
rect 572 2984 624 2990
rect 572 2926 624 2932
rect 584 2650 612 2926
rect 572 2644 624 2650
rect 572 2586 624 2592
rect 1964 2038 1992 3130
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 2056 2854 2084 2994
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 2056 2514 2084 2790
rect 2240 2514 2268 3334
rect 2516 3194 2544 4218
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2608 3670 2636 4082
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2596 3664 2648 3670
rect 2596 3606 2648 3612
rect 2596 3528 2648 3534
rect 2700 3516 2728 3946
rect 2792 3534 2820 4082
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 3110 3836 3418 3856
rect 3110 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3276 3836
rect 3332 3834 3356 3836
rect 3412 3834 3418 3836
rect 3172 3782 3174 3834
rect 3354 3782 3356 3834
rect 3110 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3276 3782
rect 3332 3780 3356 3782
rect 3412 3780 3418 3782
rect 3110 3760 3418 3780
rect 2648 3488 2728 3516
rect 2780 3528 2832 3534
rect 2596 3470 2648 3476
rect 2780 3470 2832 3476
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2608 2990 2636 3470
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2608 2446 2636 2926
rect 2792 2650 2820 3470
rect 3620 3466 3648 4014
rect 4344 3936 4396 3942
rect 4448 3924 4476 4490
rect 5460 4434 5488 4966
rect 6012 4690 6040 5170
rect 7024 5030 7052 5238
rect 7576 5234 7604 9454
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9310 9276 9618 9296
rect 9310 9274 9316 9276
rect 9372 9274 9396 9276
rect 9452 9274 9476 9276
rect 9532 9274 9556 9276
rect 9612 9274 9618 9276
rect 9372 9222 9374 9274
rect 9554 9222 9556 9274
rect 9310 9220 9316 9222
rect 9372 9220 9396 9222
rect 9452 9220 9476 9222
rect 9532 9220 9556 9222
rect 9612 9220 9618 9222
rect 9310 9200 9618 9220
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 7760 8732 8068 8752
rect 7760 8730 7766 8732
rect 7822 8730 7846 8732
rect 7902 8730 7926 8732
rect 7982 8730 8006 8732
rect 8062 8730 8068 8732
rect 7822 8678 7824 8730
rect 8004 8678 8006 8730
rect 7760 8676 7766 8678
rect 7822 8676 7846 8678
rect 7902 8676 7926 8678
rect 7982 8676 8006 8678
rect 8062 8676 8068 8678
rect 7760 8656 8068 8676
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7668 8022 7696 8230
rect 7944 8022 7972 8230
rect 7656 8016 7708 8022
rect 7656 7958 7708 7964
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 8312 7954 8340 8842
rect 8404 8498 8432 8910
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8496 7954 8524 8910
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8498 8616 8774
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8588 8294 8616 8434
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8680 8294 8708 8366
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 7760 7644 8068 7664
rect 7760 7642 7766 7644
rect 7822 7642 7846 7644
rect 7902 7642 7926 7644
rect 7982 7642 8006 7644
rect 8062 7642 8068 7644
rect 7822 7590 7824 7642
rect 8004 7590 8006 7642
rect 7760 7588 7766 7590
rect 7822 7588 7846 7590
rect 7902 7588 7926 7590
rect 7982 7588 8006 7590
rect 8062 7588 8068 7590
rect 7760 7568 8068 7588
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8036 6866 8064 7278
rect 8128 6934 8156 7822
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 8404 7478 8432 7754
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8300 7200 8352 7206
rect 8220 7148 8300 7154
rect 8220 7142 8352 7148
rect 8220 7126 8340 7142
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 6254 7696 6734
rect 7760 6556 8068 6576
rect 7760 6554 7766 6556
rect 7822 6554 7846 6556
rect 7902 6554 7926 6556
rect 7982 6554 8006 6556
rect 8062 6554 8068 6556
rect 7822 6502 7824 6554
rect 8004 6502 8006 6554
rect 7760 6500 7766 6502
rect 7822 6500 7846 6502
rect 7902 6500 7926 6502
rect 7982 6500 8006 6502
rect 8062 6500 8068 6502
rect 7760 6480 8068 6500
rect 7656 6248 7708 6254
rect 7656 6190 7708 6196
rect 7668 5914 7696 6190
rect 8128 6186 8156 6870
rect 8116 6180 8168 6186
rect 8116 6122 8168 6128
rect 8220 6066 8248 7126
rect 8404 6866 8432 7414
rect 8680 7410 8708 8230
rect 9140 7954 9168 8842
rect 9508 8634 9536 8842
rect 9692 8634 9720 9386
rect 9772 9376 9824 9382
rect 9876 9364 9904 9862
rect 9968 9586 9996 10066
rect 11072 9976 11100 10542
rect 11256 10266 11284 10610
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11072 9948 11284 9976
rect 10860 9820 11168 9840
rect 10860 9818 10866 9820
rect 10922 9818 10946 9820
rect 11002 9818 11026 9820
rect 11082 9818 11106 9820
rect 11162 9818 11168 9820
rect 10922 9766 10924 9818
rect 11104 9766 11106 9818
rect 10860 9764 10866 9766
rect 10922 9764 10946 9766
rect 11002 9764 11026 9766
rect 11082 9764 11106 9766
rect 11162 9764 11168 9766
rect 10860 9744 11168 9764
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 10692 9648 10744 9654
rect 10692 9590 10744 9596
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9824 9336 9904 9364
rect 9772 9318 9824 9324
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9310 8188 9618 8208
rect 9310 8186 9316 8188
rect 9372 8186 9396 8188
rect 9452 8186 9476 8188
rect 9532 8186 9556 8188
rect 9612 8186 9618 8188
rect 9372 8134 9374 8186
rect 9554 8134 9556 8186
rect 9310 8132 9316 8134
rect 9372 8132 9396 8134
rect 9452 8132 9476 8134
rect 9532 8132 9556 8134
rect 9612 8132 9618 8134
rect 9310 8112 9618 8132
rect 9784 8090 9812 9318
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9140 7546 9168 7890
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8496 6730 8524 7142
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8128 6038 8248 6066
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 8128 5574 8156 6038
rect 8864 5914 8892 7346
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 6934 9076 7278
rect 9310 7100 9618 7120
rect 9310 7098 9316 7100
rect 9372 7098 9396 7100
rect 9452 7098 9476 7100
rect 9532 7098 9556 7100
rect 9612 7098 9618 7100
rect 9372 7046 9374 7098
rect 9554 7046 9556 7098
rect 9310 7044 9316 7046
rect 9372 7044 9396 7046
rect 9452 7044 9476 7046
rect 9532 7044 9556 7046
rect 9612 7044 9618 7046
rect 9310 7024 9618 7044
rect 9036 6928 9088 6934
rect 9036 6870 9088 6876
rect 9048 6322 9076 6870
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9692 6322 9720 6666
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 7760 5468 8068 5488
rect 7760 5466 7766 5468
rect 7822 5466 7846 5468
rect 7902 5466 7926 5468
rect 7982 5466 8006 5468
rect 8062 5466 8068 5468
rect 7822 5414 7824 5466
rect 8004 5414 8006 5466
rect 7760 5412 7766 5414
rect 7822 5412 7846 5414
rect 7902 5412 7926 5414
rect 7982 5412 8006 5414
rect 8062 5412 8068 5414
rect 7760 5392 8068 5412
rect 8128 5302 8156 5510
rect 9140 5302 9168 6054
rect 9310 6012 9618 6032
rect 9310 6010 9316 6012
rect 9372 6010 9396 6012
rect 9452 6010 9476 6012
rect 9532 6010 9556 6012
rect 9612 6010 9618 6012
rect 9372 5958 9374 6010
rect 9554 5958 9556 6010
rect 9310 5956 9316 5958
rect 9372 5956 9396 5958
rect 9452 5956 9476 5958
rect 9532 5956 9556 5958
rect 9612 5956 9618 5958
rect 9310 5936 9618 5956
rect 9692 5914 9720 6258
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9784 5574 9812 6326
rect 9876 6186 9904 7346
rect 9864 6180 9916 6186
rect 9864 6122 9916 6128
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9784 5370 9812 5510
rect 9968 5370 9996 9522
rect 10060 7818 10088 9590
rect 10704 9178 10732 9590
rect 11152 9512 11204 9518
rect 11256 9500 11284 9948
rect 11204 9472 11284 9500
rect 11152 9454 11204 9460
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10152 8566 10180 8910
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10152 7290 10180 7754
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10060 7274 10180 7290
rect 10048 7268 10180 7274
rect 10100 7262 10180 7268
rect 10048 7210 10100 7216
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10060 6186 10088 6938
rect 10152 6254 10180 7262
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10244 6798 10272 7210
rect 10520 6866 10548 7346
rect 10612 6984 10640 8502
rect 10704 7546 10732 8978
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 10796 8294 10824 8910
rect 10860 8732 11168 8752
rect 10860 8730 10866 8732
rect 10922 8730 10946 8732
rect 11002 8730 11026 8732
rect 11082 8730 11106 8732
rect 11162 8730 11168 8732
rect 10922 8678 10924 8730
rect 11104 8678 11106 8730
rect 10860 8676 10866 8678
rect 10922 8676 10946 8678
rect 11002 8676 11026 8678
rect 11082 8676 11106 8678
rect 11162 8676 11168 8678
rect 10860 8656 11168 8676
rect 11256 8634 11284 8910
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11348 8362 11376 10678
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11428 9376 11480 9382
rect 11428 9318 11480 9324
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10704 7154 10732 7482
rect 10796 7392 10824 8230
rect 11256 7750 11284 8230
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 10860 7644 11168 7664
rect 10860 7642 10866 7644
rect 10922 7642 10946 7644
rect 11002 7642 11026 7644
rect 11082 7642 11106 7644
rect 11162 7642 11168 7644
rect 10922 7590 10924 7642
rect 11104 7590 11106 7642
rect 10860 7588 10866 7590
rect 10922 7588 10946 7590
rect 11002 7588 11026 7590
rect 11082 7588 11106 7590
rect 11162 7588 11168 7590
rect 10860 7568 11168 7588
rect 11256 7546 11284 7686
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11348 7410 11376 7958
rect 11440 7954 11468 9318
rect 11532 8634 11560 10406
rect 12410 10364 12718 10384
rect 12410 10362 12416 10364
rect 12472 10362 12496 10364
rect 12552 10362 12576 10364
rect 12632 10362 12656 10364
rect 12712 10362 12718 10364
rect 12472 10310 12474 10362
rect 12654 10310 12656 10362
rect 12410 10308 12416 10310
rect 12472 10308 12496 10310
rect 12552 10308 12576 10310
rect 12632 10308 12656 10310
rect 12712 10308 12718 10310
rect 12410 10288 12718 10308
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 10876 7404 10928 7410
rect 10796 7364 10876 7392
rect 10876 7346 10928 7352
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10968 7200 11020 7206
rect 10704 7126 10916 7154
rect 10968 7142 11020 7148
rect 10612 6956 10824 6984
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10232 6792 10284 6798
rect 10416 6792 10468 6798
rect 10232 6734 10284 6740
rect 10336 6740 10416 6746
rect 10336 6734 10468 6740
rect 10336 6718 10456 6734
rect 10232 6452 10284 6458
rect 10336 6440 10364 6718
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10284 6412 10364 6440
rect 10232 6394 10284 6400
rect 10428 6390 10456 6598
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10428 5778 10456 6054
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 9772 5364 9824 5370
rect 9956 5364 10008 5370
rect 9772 5306 9824 5312
rect 9876 5324 9956 5352
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 9128 5296 9180 5302
rect 9876 5250 9904 5324
rect 9956 5306 10008 5312
rect 9128 5238 9180 5244
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 9692 5222 9904 5250
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6210 4924 6518 4944
rect 6210 4922 6216 4924
rect 6272 4922 6296 4924
rect 6352 4922 6376 4924
rect 6432 4922 6456 4924
rect 6512 4922 6518 4924
rect 6272 4870 6274 4922
rect 6454 4870 6456 4922
rect 6210 4868 6216 4870
rect 6272 4868 6296 4870
rect 6352 4868 6376 4870
rect 6432 4868 6456 4870
rect 6512 4868 6518 4870
rect 6210 4848 6518 4868
rect 6000 4684 6052 4690
rect 6000 4626 6052 4632
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 5460 4406 5672 4434
rect 4660 4380 4968 4400
rect 4660 4378 4666 4380
rect 4722 4378 4746 4380
rect 4802 4378 4826 4380
rect 4882 4378 4906 4380
rect 4962 4378 4968 4380
rect 4722 4326 4724 4378
rect 4904 4326 4906 4378
rect 4660 4324 4666 4326
rect 4722 4324 4746 4326
rect 4802 4324 4826 4326
rect 4882 4324 4906 4326
rect 4962 4324 4968 4326
rect 4660 4304 4968 4324
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 4396 3896 4476 3924
rect 4344 3878 4396 3884
rect 3608 3460 3660 3466
rect 3608 3402 3660 3408
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3160 2990 3188 3334
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 3528 2922 3556 3334
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2884 2378 2912 2858
rect 3110 2748 3418 2768
rect 3110 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3276 2748
rect 3332 2746 3356 2748
rect 3412 2746 3418 2748
rect 3172 2694 3174 2746
rect 3354 2694 3356 2746
rect 3110 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3276 2694
rect 3332 2692 3356 2694
rect 3412 2692 3418 2694
rect 3110 2672 3418 2692
rect 3528 2650 3556 2858
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 1952 2032 2004 2038
rect 1952 1974 2004 1980
rect 296 1896 348 1902
rect 296 1838 348 1844
rect 1768 1828 1820 1834
rect 1768 1770 1820 1776
rect 1780 1358 1808 1770
rect 1964 1766 1992 1974
rect 2792 1902 2820 2246
rect 2976 1970 3004 2382
rect 4356 2378 4384 3878
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 4660 3292 4968 3312
rect 4660 3290 4666 3292
rect 4722 3290 4746 3292
rect 4802 3290 4826 3292
rect 4882 3290 4906 3292
rect 4962 3290 4968 3292
rect 4722 3238 4724 3290
rect 4904 3238 4906 3290
rect 4660 3236 4666 3238
rect 4722 3236 4746 3238
rect 4802 3236 4826 3238
rect 4882 3236 4906 3238
rect 4962 3236 4968 3238
rect 4660 3216 4968 3236
rect 5276 3126 5304 3402
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 3126 5488 3334
rect 5264 3120 5316 3126
rect 5264 3062 5316 3068
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5276 2774 5304 3062
rect 5276 2746 5396 2774
rect 4344 2372 4396 2378
rect 4344 2314 4396 2320
rect 4356 1970 4384 2314
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 4660 2204 4968 2224
rect 4660 2202 4666 2204
rect 4722 2202 4746 2204
rect 4802 2202 4826 2204
rect 4882 2202 4906 2204
rect 4962 2202 4968 2204
rect 4722 2150 4724 2202
rect 4904 2150 4906 2202
rect 4660 2148 4666 2150
rect 4722 2148 4746 2150
rect 4802 2148 4826 2150
rect 4882 2148 4906 2150
rect 4962 2148 4968 2150
rect 4660 2128 4968 2148
rect 5000 1970 5028 2246
rect 2964 1964 3016 1970
rect 2964 1906 3016 1912
rect 4344 1964 4396 1970
rect 4344 1906 4396 1912
rect 4988 1964 5040 1970
rect 4988 1906 5040 1912
rect 5080 1964 5132 1970
rect 5368 1952 5396 2746
rect 5460 2650 5488 3062
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5552 2514 5580 4218
rect 5644 4214 5672 4406
rect 6012 4282 6040 4626
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 6104 4078 6132 4422
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6000 3936 6052 3942
rect 6196 3924 6224 4558
rect 6000 3878 6052 3884
rect 6104 3896 6224 3924
rect 6012 3602 6040 3878
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5736 2922 5764 3130
rect 5920 3058 5948 3470
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6104 2990 6132 3896
rect 6210 3836 6518 3856
rect 6210 3834 6216 3836
rect 6272 3834 6296 3836
rect 6352 3834 6376 3836
rect 6432 3834 6456 3836
rect 6512 3834 6518 3836
rect 6272 3782 6274 3834
rect 6454 3782 6456 3834
rect 6210 3780 6216 3782
rect 6272 3780 6296 3782
rect 6352 3780 6376 3782
rect 6432 3780 6456 3782
rect 6512 3780 6518 3782
rect 6210 3760 6518 3780
rect 6564 3738 6592 4558
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6748 3738 6776 4422
rect 7024 4146 7052 4558
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7668 4282 7696 4422
rect 7760 4380 8068 4400
rect 7760 4378 7766 4380
rect 7822 4378 7846 4380
rect 7902 4378 7926 4380
rect 7982 4378 8006 4380
rect 8062 4378 8068 4380
rect 7822 4326 7824 4378
rect 8004 4326 8006 4378
rect 7760 4324 7766 4326
rect 7822 4324 7846 4326
rect 7902 4324 7926 4326
rect 7982 4324 8006 4326
rect 8062 4324 8068 4326
rect 7760 4304 8068 4324
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6840 2990 6868 3606
rect 7024 3466 7052 4082
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7300 3534 7328 3878
rect 8220 3670 8248 4082
rect 8312 4078 8340 4626
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 8312 3466 8340 4014
rect 8496 3738 8524 5102
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8956 4282 8984 4626
rect 9048 4622 9076 4966
rect 9310 4924 9618 4944
rect 9310 4922 9316 4924
rect 9372 4922 9396 4924
rect 9452 4922 9476 4924
rect 9532 4922 9556 4924
rect 9612 4922 9618 4924
rect 9372 4870 9374 4922
rect 9554 4870 9556 4922
rect 9310 4868 9316 4870
rect 9372 4868 9396 4870
rect 9452 4868 9476 4870
rect 9532 4868 9556 4870
rect 9612 4868 9618 4870
rect 9310 4848 9618 4868
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8760 4140 8812 4146
rect 8680 4100 8760 4128
rect 8680 3942 8708 4100
rect 8760 4082 8812 4088
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7392 3194 7420 3334
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 6092 2984 6144 2990
rect 6828 2984 6880 2990
rect 6092 2926 6144 2932
rect 6748 2944 6828 2972
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5908 2916 5960 2922
rect 5908 2858 5960 2864
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5552 2038 5580 2450
rect 5644 2378 5672 2790
rect 5920 2774 5948 2858
rect 5920 2746 6040 2774
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 5540 2032 5592 2038
rect 5540 1974 5592 1980
rect 5448 1964 5500 1970
rect 5368 1924 5448 1952
rect 5080 1906 5132 1912
rect 5448 1906 5500 1912
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 4068 1896 4120 1902
rect 4068 1838 4120 1844
rect 1952 1760 2004 1766
rect 1952 1702 2004 1708
rect 2228 1760 2280 1766
rect 2228 1702 2280 1708
rect 2504 1760 2556 1766
rect 2504 1702 2556 1708
rect 1768 1352 1820 1358
rect 1768 1294 1820 1300
rect 2240 678 2268 1702
rect 2516 882 2544 1702
rect 3110 1660 3418 1680
rect 3110 1658 3116 1660
rect 3172 1658 3196 1660
rect 3252 1658 3276 1660
rect 3332 1658 3356 1660
rect 3412 1658 3418 1660
rect 3172 1606 3174 1658
rect 3354 1606 3356 1658
rect 3110 1604 3116 1606
rect 3172 1604 3196 1606
rect 3252 1604 3276 1606
rect 3332 1604 3356 1606
rect 3412 1604 3418 1606
rect 3110 1584 3418 1604
rect 4080 1494 4108 1838
rect 4068 1488 4120 1494
rect 4068 1430 4120 1436
rect 4356 1358 4384 1906
rect 4436 1760 4488 1766
rect 4436 1702 4488 1708
rect 4528 1760 4580 1766
rect 4528 1702 4580 1708
rect 4344 1352 4396 1358
rect 4344 1294 4396 1300
rect 4356 882 4384 1294
rect 4448 950 4476 1702
rect 4540 1426 4568 1702
rect 5092 1494 5120 1906
rect 5172 1760 5224 1766
rect 5172 1702 5224 1708
rect 5080 1488 5132 1494
rect 5080 1430 5132 1436
rect 4528 1420 4580 1426
rect 4528 1362 4580 1368
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 4528 1284 4580 1290
rect 4528 1226 4580 1232
rect 4436 944 4488 950
rect 4436 886 4488 892
rect 2504 876 2556 882
rect 2504 818 2556 824
rect 4344 876 4396 882
rect 4540 864 4568 1226
rect 4660 1116 4968 1136
rect 4660 1114 4666 1116
rect 4722 1114 4746 1116
rect 4802 1114 4826 1116
rect 4882 1114 4906 1116
rect 4962 1114 4968 1116
rect 4722 1062 4724 1114
rect 4904 1062 4906 1114
rect 4660 1060 4666 1062
rect 4722 1060 4746 1062
rect 4802 1060 4826 1062
rect 4882 1060 4906 1062
rect 4962 1060 4968 1062
rect 4660 1040 4968 1060
rect 5000 1018 5028 1294
rect 4988 1012 5040 1018
rect 4988 954 5040 960
rect 4894 912 4950 921
rect 4712 876 4764 882
rect 4540 836 4712 864
rect 4344 818 4396 824
rect 5092 882 5120 1430
rect 5184 1222 5212 1702
rect 5264 1284 5316 1290
rect 5264 1226 5316 1232
rect 5172 1216 5224 1222
rect 5172 1158 5224 1164
rect 4894 847 4896 856
rect 4712 818 4764 824
rect 4948 847 4950 856
rect 5080 876 5132 882
rect 4896 818 4948 824
rect 5080 818 5132 824
rect 4356 678 4384 818
rect 2228 672 2280 678
rect 2228 614 2280 620
rect 4344 672 4396 678
rect 4344 614 4396 620
rect 3110 572 3418 592
rect 3110 570 3116 572
rect 3172 570 3196 572
rect 3252 570 3276 572
rect 3332 570 3356 572
rect 3412 570 3418 572
rect 3172 518 3174 570
rect 3354 518 3356 570
rect 3110 516 3116 518
rect 3172 516 3196 518
rect 3252 516 3276 518
rect 3332 516 3356 518
rect 3412 516 3418 518
rect 3110 496 3418 516
rect 4724 202 4752 818
rect 5184 270 5212 1158
rect 5276 921 5304 1226
rect 5356 1216 5408 1222
rect 5356 1158 5408 1164
rect 5262 912 5318 921
rect 5262 847 5318 856
rect 5368 746 5396 1158
rect 5552 1034 5580 1974
rect 6012 1358 6040 2746
rect 6210 2748 6518 2768
rect 6210 2746 6216 2748
rect 6272 2746 6296 2748
rect 6352 2746 6376 2748
rect 6432 2746 6456 2748
rect 6512 2746 6518 2748
rect 6272 2694 6274 2746
rect 6454 2694 6456 2746
rect 6210 2692 6216 2694
rect 6272 2692 6296 2694
rect 6352 2692 6376 2694
rect 6432 2692 6456 2694
rect 6512 2692 6518 2694
rect 6210 2672 6518 2692
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 6104 2038 6132 2382
rect 6092 2032 6144 2038
rect 6092 1974 6144 1980
rect 6748 1970 6776 2944
rect 6828 2926 6880 2932
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6840 1970 6868 2790
rect 6736 1964 6788 1970
rect 6736 1906 6788 1912
rect 6828 1964 6880 1970
rect 6828 1906 6880 1912
rect 6210 1660 6518 1680
rect 6210 1658 6216 1660
rect 6272 1658 6296 1660
rect 6352 1658 6376 1660
rect 6432 1658 6456 1660
rect 6512 1658 6518 1660
rect 6272 1606 6274 1658
rect 6454 1606 6456 1658
rect 6210 1604 6216 1606
rect 6272 1604 6296 1606
rect 6352 1604 6376 1606
rect 6432 1604 6456 1606
rect 6512 1604 6518 1606
rect 6210 1584 6518 1604
rect 6748 1426 6776 1906
rect 6736 1420 6788 1426
rect 6736 1362 6788 1368
rect 5908 1352 5960 1358
rect 5908 1294 5960 1300
rect 6000 1352 6052 1358
rect 6000 1294 6052 1300
rect 5816 1216 5868 1222
rect 5816 1158 5868 1164
rect 5460 1006 5580 1034
rect 5460 950 5488 1006
rect 5448 944 5500 950
rect 5448 886 5500 892
rect 5632 808 5684 814
rect 5632 750 5684 756
rect 5356 740 5408 746
rect 5356 682 5408 688
rect 5172 264 5224 270
rect 5172 206 5224 212
rect 4712 196 4764 202
rect 4712 138 4764 144
rect 5368 134 5396 682
rect 5644 474 5672 750
rect 5632 468 5684 474
rect 5632 410 5684 416
rect 5828 338 5856 1158
rect 5920 1018 5948 1294
rect 6932 1222 6960 3062
rect 7208 2650 7236 3062
rect 7484 2854 7512 3334
rect 7760 3292 8068 3312
rect 7760 3290 7766 3292
rect 7822 3290 7846 3292
rect 7902 3290 7926 3292
rect 7982 3290 8006 3292
rect 8062 3290 8068 3292
rect 7822 3238 7824 3290
rect 8004 3238 8006 3290
rect 7760 3236 7766 3238
rect 7822 3236 7846 3238
rect 7902 3236 7926 3238
rect 7982 3236 8006 3238
rect 8062 3236 8068 3238
rect 7760 3216 8068 3236
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7472 2372 7524 2378
rect 7472 2314 7524 2320
rect 7484 1970 7512 2314
rect 7760 2204 8068 2224
rect 7760 2202 7766 2204
rect 7822 2202 7846 2204
rect 7902 2202 7926 2204
rect 7982 2202 8006 2204
rect 8062 2202 8068 2204
rect 7822 2150 7824 2202
rect 8004 2150 8006 2202
rect 7760 2148 7766 2150
rect 7822 2148 7846 2150
rect 7902 2148 7926 2150
rect 7982 2148 8006 2150
rect 8062 2148 8068 2150
rect 7760 2128 8068 2148
rect 7472 1964 7524 1970
rect 7472 1906 7524 1912
rect 7380 1896 7432 1902
rect 7380 1838 7432 1844
rect 7392 1358 7420 1838
rect 7484 1494 7512 1906
rect 7472 1488 7524 1494
rect 7472 1430 7524 1436
rect 7012 1352 7064 1358
rect 7010 1320 7012 1329
rect 7380 1352 7432 1358
rect 7064 1320 7066 1329
rect 7380 1294 7432 1300
rect 7010 1255 7066 1264
rect 6920 1216 6972 1222
rect 6920 1158 6972 1164
rect 7392 1018 7420 1294
rect 5908 1012 5960 1018
rect 5908 954 5960 960
rect 7380 1012 7432 1018
rect 7380 954 7432 960
rect 5816 332 5868 338
rect 5816 274 5868 280
rect 5920 270 5948 954
rect 7484 882 7512 1430
rect 7564 1284 7616 1290
rect 7564 1226 7616 1232
rect 7576 1018 7604 1226
rect 8220 1222 8248 3130
rect 8312 3058 8340 3402
rect 8588 3194 8616 3674
rect 8666 3632 8722 3641
rect 8772 3602 8800 3878
rect 8666 3567 8722 3576
rect 8760 3596 8812 3602
rect 8680 3534 8708 3567
rect 8760 3538 8812 3544
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8944 3528 8996 3534
rect 9048 3505 9076 4558
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 8944 3470 8996 3476
rect 9034 3496 9090 3505
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8772 2582 8800 3130
rect 8956 3126 8984 3470
rect 9034 3431 9036 3440
rect 9088 3431 9090 3440
rect 9036 3402 9088 3408
rect 9048 3371 9076 3402
rect 8944 3120 8996 3126
rect 8942 3088 8944 3097
rect 8996 3088 8998 3097
rect 8942 3023 8998 3032
rect 9140 2774 9168 3878
rect 8956 2746 9168 2774
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 8312 1834 8340 2246
rect 8588 1902 8616 2314
rect 8576 1896 8628 1902
rect 8576 1838 8628 1844
rect 8300 1828 8352 1834
rect 8300 1770 8352 1776
rect 8208 1216 8260 1222
rect 8208 1158 8260 1164
rect 7760 1116 8068 1136
rect 7760 1114 7766 1116
rect 7822 1114 7846 1116
rect 7902 1114 7926 1116
rect 7982 1114 8006 1116
rect 8062 1114 8068 1116
rect 7822 1062 7824 1114
rect 8004 1062 8006 1114
rect 7760 1060 7766 1062
rect 7822 1060 7846 1062
rect 7902 1060 7926 1062
rect 7982 1060 8006 1062
rect 8062 1060 8068 1062
rect 7760 1040 8068 1060
rect 7564 1012 7616 1018
rect 7564 954 7616 960
rect 7746 912 7802 921
rect 7288 876 7340 882
rect 7288 818 7340 824
rect 7472 876 7524 882
rect 8220 882 8248 1158
rect 7746 847 7748 856
rect 7472 818 7524 824
rect 7800 847 7802 856
rect 8208 876 8260 882
rect 7748 818 7800 824
rect 8208 818 8260 824
rect 6210 572 6518 592
rect 6210 570 6216 572
rect 6272 570 6296 572
rect 6352 570 6376 572
rect 6432 570 6456 572
rect 6512 570 6518 572
rect 6272 518 6274 570
rect 6454 518 6456 570
rect 6210 516 6216 518
rect 6272 516 6296 518
rect 6352 516 6376 518
rect 6432 516 6456 518
rect 6512 516 6518 518
rect 6210 496 6518 516
rect 7300 474 7328 818
rect 8312 814 8340 1770
rect 8668 1760 8720 1766
rect 8668 1702 8720 1708
rect 8680 1426 8708 1702
rect 8772 1426 8800 2518
rect 8668 1420 8720 1426
rect 8668 1362 8720 1368
rect 8760 1420 8812 1426
rect 8760 1362 8812 1368
rect 8576 1352 8628 1358
rect 8852 1352 8904 1358
rect 8576 1294 8628 1300
rect 8758 1320 8814 1329
rect 8588 950 8616 1294
rect 8852 1294 8904 1300
rect 8758 1255 8814 1264
rect 8576 944 8628 950
rect 8576 886 8628 892
rect 8772 882 8800 1255
rect 8760 876 8812 882
rect 8760 818 8812 824
rect 8300 808 8352 814
rect 8300 750 8352 756
rect 8864 474 8892 1294
rect 8956 1018 8984 2746
rect 9036 1420 9088 1426
rect 9036 1362 9088 1368
rect 8944 1012 8996 1018
rect 8944 954 8996 960
rect 7288 468 7340 474
rect 7288 410 7340 416
rect 8852 468 8904 474
rect 8852 410 8904 416
rect 9048 377 9076 1362
rect 9232 1329 9260 4014
rect 9310 3836 9618 3856
rect 9310 3834 9316 3836
rect 9372 3834 9396 3836
rect 9452 3834 9476 3836
rect 9532 3834 9556 3836
rect 9612 3834 9618 3836
rect 9372 3782 9374 3834
rect 9554 3782 9556 3834
rect 9310 3780 9316 3782
rect 9372 3780 9396 3782
rect 9452 3780 9476 3782
rect 9532 3780 9556 3782
rect 9612 3780 9618 3782
rect 9310 3760 9618 3780
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9416 3058 9444 3334
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9310 2748 9618 2768
rect 9310 2746 9316 2748
rect 9372 2746 9396 2748
rect 9452 2746 9476 2748
rect 9532 2746 9556 2748
rect 9612 2746 9618 2748
rect 9372 2694 9374 2746
rect 9554 2694 9556 2746
rect 9310 2692 9316 2694
rect 9372 2692 9396 2694
rect 9452 2692 9476 2694
rect 9532 2692 9556 2694
rect 9612 2692 9618 2694
rect 9310 2672 9618 2692
rect 9692 2514 9720 5222
rect 10060 5166 10088 5714
rect 10520 5166 10548 6802
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 6458 10640 6598
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10704 6322 10732 6802
rect 10796 6730 10824 6956
rect 10888 6866 10916 7126
rect 10980 7002 11008 7142
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10980 6730 11008 6938
rect 11072 6798 11100 7278
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 10860 6556 11168 6576
rect 10860 6554 10866 6556
rect 10922 6554 10946 6556
rect 11002 6554 11026 6556
rect 11082 6554 11106 6556
rect 11162 6554 11168 6556
rect 10922 6502 10924 6554
rect 11104 6502 11106 6554
rect 10860 6500 10866 6502
rect 10922 6500 10946 6502
rect 11002 6500 11026 6502
rect 11082 6500 11106 6502
rect 11162 6500 11168 6502
rect 10860 6480 11168 6500
rect 10600 6316 10652 6322
rect 10600 6258 10652 6264
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10612 5234 10640 6258
rect 10704 5778 10732 6258
rect 11256 5914 11284 6598
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 10692 5772 10744 5778
rect 10692 5714 10744 5720
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 10860 5468 11168 5488
rect 10860 5466 10866 5468
rect 10922 5466 10946 5468
rect 11002 5466 11026 5468
rect 11082 5466 11106 5468
rect 11162 5466 11168 5468
rect 10922 5414 10924 5466
rect 11104 5414 11106 5466
rect 10860 5412 10866 5414
rect 10922 5412 10946 5414
rect 11002 5412 11026 5414
rect 11082 5412 11106 5414
rect 11162 5412 11168 5414
rect 10860 5392 11168 5412
rect 11256 5302 11284 5714
rect 11624 5370 11652 9454
rect 11808 9178 11836 9522
rect 12820 9518 12848 10542
rect 13176 10532 13228 10538
rect 13176 10474 13228 10480
rect 14372 10532 14424 10538
rect 14372 10474 14424 10480
rect 13188 10266 13216 10474
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13176 10260 13228 10266
rect 13176 10202 13228 10208
rect 13372 10130 13400 10406
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 14384 9926 14412 10474
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14476 10130 14504 10406
rect 14464 10124 14516 10130
rect 14464 10066 14516 10072
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 13960 9820 14268 9840
rect 13960 9818 13966 9820
rect 14022 9818 14046 9820
rect 14102 9818 14126 9820
rect 14182 9818 14206 9820
rect 14262 9818 14268 9820
rect 14022 9766 14024 9818
rect 14204 9766 14206 9818
rect 13960 9764 13966 9766
rect 14022 9764 14046 9766
rect 14102 9764 14126 9766
rect 14182 9764 14206 9766
rect 14262 9764 14268 9766
rect 13960 9744 14268 9764
rect 14384 9722 14412 9862
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12410 9276 12718 9296
rect 12410 9274 12416 9276
rect 12472 9274 12496 9276
rect 12552 9274 12576 9276
rect 12632 9274 12656 9276
rect 12712 9274 12718 9276
rect 12472 9222 12474 9274
rect 12654 9222 12656 9274
rect 12410 9220 12416 9222
rect 12472 9220 12496 9222
rect 12552 9220 12576 9222
rect 12632 9220 12656 9222
rect 12712 9220 12718 9222
rect 12410 9200 12718 9220
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11808 8906 11836 9114
rect 11796 8900 11848 8906
rect 11848 8860 11928 8888
rect 11796 8842 11848 8848
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11716 7546 11744 8366
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11808 7410 11836 7754
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11808 6798 11836 7346
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11900 6458 11928 8860
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8498 12020 8774
rect 12820 8650 12848 9454
rect 14476 9382 14504 9658
rect 14844 9586 14872 10406
rect 15212 10266 15240 10610
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 13372 9042 13400 9318
rect 13360 9036 13412 9042
rect 13360 8978 13412 8984
rect 13464 8974 13492 9318
rect 14476 9178 14504 9318
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14464 9172 14516 9178
rect 14516 9132 14596 9160
rect 14464 9114 14516 9120
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 12728 8622 12848 8650
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11992 7886 12020 8434
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 12176 7342 12204 8366
rect 12728 8362 12756 8622
rect 13464 8566 13492 8910
rect 14200 8906 14228 9114
rect 14464 9036 14516 9042
rect 14464 8978 14516 8984
rect 14188 8900 14240 8906
rect 14188 8842 14240 8848
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 13960 8732 14268 8752
rect 13960 8730 13966 8732
rect 14022 8730 14046 8732
rect 14102 8730 14126 8732
rect 14182 8730 14206 8732
rect 14262 8730 14268 8732
rect 14022 8678 14024 8730
rect 14204 8678 14206 8730
rect 13960 8676 13966 8678
rect 14022 8676 14046 8678
rect 14102 8676 14126 8678
rect 14182 8676 14206 8678
rect 14262 8676 14268 8678
rect 13960 8656 14268 8676
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12268 7886 12296 8230
rect 12410 8188 12718 8208
rect 12410 8186 12416 8188
rect 12472 8186 12496 8188
rect 12552 8186 12576 8188
rect 12632 8186 12656 8188
rect 12712 8186 12718 8188
rect 12472 8134 12474 8186
rect 12654 8134 12656 8186
rect 12410 8132 12416 8134
rect 12472 8132 12496 8134
rect 12552 8132 12576 8134
rect 12632 8132 12656 8134
rect 12712 8132 12718 8134
rect 12410 8112 12718 8132
rect 12820 8022 12848 8434
rect 12912 8090 12940 8502
rect 14384 8498 14412 8774
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7410 12296 7822
rect 13280 7818 13308 8366
rect 13372 8090 13400 8434
rect 14476 8430 14504 8978
rect 14568 8634 14596 9132
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 14292 7954 14320 8230
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7410 13492 7686
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12410 7100 12718 7120
rect 12410 7098 12416 7100
rect 12472 7098 12496 7100
rect 12552 7098 12576 7100
rect 12632 7098 12656 7100
rect 12712 7098 12718 7100
rect 12472 7046 12474 7098
rect 12654 7046 12656 7098
rect 12410 7044 12416 7046
rect 12472 7044 12496 7046
rect 12552 7044 12576 7046
rect 12632 7044 12656 7046
rect 12712 7044 12718 7046
rect 12410 7024 12718 7044
rect 13556 6798 13584 7822
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 13648 7449 13676 7754
rect 13740 7546 13768 7890
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13634 7440 13690 7449
rect 13634 7375 13636 7384
rect 13688 7375 13690 7384
rect 13728 7438 13780 7444
rect 13728 7380 13780 7386
rect 13636 7346 13688 7352
rect 13648 7315 13676 7346
rect 13740 7206 13768 7380
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11900 6254 11928 6394
rect 12360 6390 12388 6598
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11900 5642 11928 6190
rect 13556 6186 13584 6734
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13740 6390 13768 6598
rect 13832 6458 13860 7754
rect 13960 7644 14268 7664
rect 13960 7642 13966 7644
rect 14022 7642 14046 7644
rect 14102 7642 14126 7644
rect 14182 7642 14206 7644
rect 14262 7642 14268 7644
rect 14022 7590 14024 7642
rect 14204 7590 14206 7642
rect 13960 7588 13966 7590
rect 14022 7588 14046 7590
rect 14102 7588 14126 7590
rect 14182 7588 14206 7590
rect 14262 7588 14268 7590
rect 13960 7568 14268 7588
rect 14384 7478 14412 7754
rect 14004 7472 14056 7478
rect 13910 7440 13966 7449
rect 14004 7414 14056 7420
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 13910 7375 13912 7384
rect 13964 7375 13966 7384
rect 13912 7346 13964 7352
rect 14016 7206 14044 7414
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14384 6798 14412 7142
rect 14476 6866 14504 8366
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14568 7478 14596 7822
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14660 7410 14688 7686
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 13960 6556 14268 6576
rect 13960 6554 13966 6556
rect 14022 6554 14046 6556
rect 14102 6554 14126 6556
rect 14182 6554 14206 6556
rect 14262 6554 14268 6556
rect 14022 6502 14024 6554
rect 14204 6502 14206 6554
rect 13960 6500 13966 6502
rect 14022 6500 14046 6502
rect 14102 6500 14126 6502
rect 14182 6500 14206 6502
rect 14262 6500 14268 6502
rect 13960 6480 14268 6500
rect 14384 6458 14412 6734
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 12410 6012 12718 6032
rect 12410 6010 12416 6012
rect 12472 6010 12496 6012
rect 12552 6010 12576 6012
rect 12632 6010 12656 6012
rect 12712 6010 12718 6012
rect 12472 5958 12474 6010
rect 12654 5958 12656 6010
rect 12410 5956 12416 5958
rect 12472 5956 12496 5958
rect 12552 5956 12576 5958
rect 12632 5956 12656 5958
rect 12712 5956 12718 5958
rect 12410 5936 12718 5956
rect 13832 5642 13860 6394
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14096 6112 14148 6118
rect 14096 6054 14148 6060
rect 14108 5778 14136 6054
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 14384 5710 14412 6190
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 11888 5636 11940 5642
rect 11888 5578 11940 5584
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11244 5296 11296 5302
rect 11244 5238 11296 5244
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10060 4282 10088 4626
rect 10860 4380 11168 4400
rect 10860 4378 10866 4380
rect 10922 4378 10946 4380
rect 11002 4378 11026 4380
rect 11082 4378 11106 4380
rect 11162 4378 11168 4380
rect 10922 4326 10924 4378
rect 11104 4326 11106 4378
rect 10860 4324 10866 4326
rect 10922 4324 10946 4326
rect 11002 4324 11026 4326
rect 11082 4324 11106 4326
rect 11162 4324 11168 4326
rect 10860 4304 11168 4324
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 9772 3528 9824 3534
rect 9770 3496 9772 3505
rect 9824 3496 9826 3505
rect 9770 3431 9826 3440
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9692 2038 9720 2450
rect 9784 2310 9812 3334
rect 9876 2854 9904 4014
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 9968 3194 9996 3402
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10244 3058 10272 4014
rect 11256 3670 11284 4694
rect 11348 4690 11376 5306
rect 11900 5302 11928 5578
rect 13960 5468 14268 5488
rect 13960 5466 13966 5468
rect 14022 5466 14046 5468
rect 14102 5466 14126 5468
rect 14182 5466 14206 5468
rect 14262 5466 14268 5468
rect 14022 5414 14024 5466
rect 14204 5414 14206 5466
rect 13960 5412 13966 5414
rect 14022 5412 14046 5414
rect 14102 5412 14126 5414
rect 14182 5412 14206 5414
rect 14262 5412 14268 5414
rect 13960 5392 14268 5412
rect 11888 5296 11940 5302
rect 11888 5238 11940 5244
rect 14280 5296 14332 5302
rect 14280 5238 14332 5244
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11348 4146 11376 4490
rect 11440 4282 11468 4626
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11348 4010 11376 4082
rect 11336 4004 11388 4010
rect 11336 3946 11388 3952
rect 11244 3664 11296 3670
rect 11244 3606 11296 3612
rect 11796 3596 11848 3602
rect 11796 3538 11848 3544
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11518 3496 11574 3505
rect 10428 3194 10456 3470
rect 10860 3292 11168 3312
rect 10860 3290 10866 3292
rect 10922 3290 10946 3292
rect 11002 3290 11026 3292
rect 11082 3290 11106 3292
rect 11162 3290 11168 3292
rect 10922 3238 10924 3290
rect 11104 3238 11106 3290
rect 10860 3236 10866 3238
rect 10922 3236 10946 3238
rect 11002 3236 11026 3238
rect 11082 3236 11106 3238
rect 11162 3236 11168 3238
rect 10860 3216 11168 3236
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10874 3088 10930 3097
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10784 3052 10836 3058
rect 10874 3023 10930 3032
rect 11150 3088 11206 3097
rect 11150 3023 11152 3032
rect 10784 2994 10836 3000
rect 9864 2848 9916 2854
rect 9864 2790 9916 2796
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9680 2032 9732 2038
rect 9680 1974 9732 1980
rect 9772 2032 9824 2038
rect 9772 1974 9824 1980
rect 9680 1896 9732 1902
rect 9784 1884 9812 1974
rect 9732 1856 9812 1884
rect 9680 1838 9732 1844
rect 9876 1834 9904 2790
rect 10612 2582 10640 2994
rect 10796 2922 10824 2994
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10600 2576 10652 2582
rect 10600 2518 10652 2524
rect 10796 2514 10824 2858
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10888 2446 10916 3023
rect 11204 3023 11206 3032
rect 11152 2994 11204 3000
rect 11256 2650 11284 3470
rect 11808 3466 11836 3538
rect 11518 3431 11520 3440
rect 11572 3431 11574 3440
rect 11796 3460 11848 3466
rect 11520 3402 11572 3408
rect 11796 3402 11848 3408
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11348 3126 11376 3334
rect 11808 3194 11836 3402
rect 11900 3194 11928 5238
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 12410 4924 12718 4944
rect 12410 4922 12416 4924
rect 12472 4922 12496 4924
rect 12552 4922 12576 4924
rect 12632 4922 12656 4924
rect 12712 4922 12718 4924
rect 12472 4870 12474 4922
rect 12654 4870 12656 4922
rect 12410 4868 12416 4870
rect 12472 4868 12496 4870
rect 12552 4868 12576 4870
rect 12632 4868 12656 4870
rect 12712 4868 12718 4870
rect 12410 4848 12718 4868
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12176 3670 12204 4218
rect 12164 3664 12216 3670
rect 12164 3606 12216 3612
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 11428 3052 11480 3058
rect 11428 2994 11480 3000
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 9968 1970 9996 2042
rect 9956 1964 10008 1970
rect 9956 1906 10008 1912
rect 9864 1828 9916 1834
rect 9864 1770 9916 1776
rect 10152 1766 10180 2246
rect 10860 2204 11168 2224
rect 10860 2202 10866 2204
rect 10922 2202 10946 2204
rect 11002 2202 11026 2204
rect 11082 2202 11106 2204
rect 11162 2202 11168 2204
rect 10922 2150 10924 2202
rect 11104 2150 11106 2202
rect 10860 2148 10866 2150
rect 10922 2148 10946 2150
rect 11002 2148 11026 2150
rect 11082 2148 11106 2150
rect 11162 2148 11168 2150
rect 10860 2128 11168 2148
rect 11256 1970 11284 2314
rect 11440 2106 11468 2994
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11716 2378 11744 2926
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 11900 2310 11928 3130
rect 12268 3058 12296 4558
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13188 4146 13216 4422
rect 13740 4282 13768 4422
rect 13728 4276 13780 4282
rect 13648 4236 13728 4264
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12410 3836 12718 3856
rect 12410 3834 12416 3836
rect 12472 3834 12496 3836
rect 12552 3834 12576 3836
rect 12632 3834 12656 3836
rect 12712 3834 12718 3836
rect 12472 3782 12474 3834
rect 12654 3782 12656 3834
rect 12410 3780 12416 3782
rect 12472 3780 12496 3782
rect 12552 3780 12576 3782
rect 12632 3780 12656 3782
rect 12712 3780 12718 3782
rect 12410 3760 12718 3780
rect 12532 3664 12584 3670
rect 12346 3632 12402 3641
rect 12532 3606 12584 3612
rect 12346 3567 12348 3576
rect 12400 3567 12402 3576
rect 12348 3538 12400 3544
rect 12544 3398 12572 3606
rect 12716 3528 12768 3534
rect 12820 3516 12848 3878
rect 13004 3754 13032 4014
rect 13004 3738 13124 3754
rect 13004 3732 13136 3738
rect 13004 3726 13084 3732
rect 13084 3674 13136 3680
rect 13464 3534 13492 4014
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 12768 3488 12848 3516
rect 13452 3528 13504 3534
rect 13450 3496 13452 3505
rect 13504 3496 13506 3505
rect 12716 3470 12768 3476
rect 13450 3431 13506 3440
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12636 3126 12664 3334
rect 13556 3194 13584 3674
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 13648 3058 13676 4236
rect 13728 4218 13780 4224
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13740 3534 13768 4082
rect 13832 3534 13860 5102
rect 14292 4554 14320 5238
rect 14384 4826 14412 5646
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14280 4548 14332 4554
rect 14332 4508 14412 4536
rect 14280 4490 14332 4496
rect 13960 4380 14268 4400
rect 13960 4378 13966 4380
rect 14022 4378 14046 4380
rect 14102 4378 14126 4380
rect 14182 4378 14206 4380
rect 14262 4378 14268 4380
rect 14022 4326 14024 4378
rect 14204 4326 14206 4378
rect 13960 4324 13966 4326
rect 14022 4324 14046 4326
rect 14102 4324 14126 4326
rect 14182 4324 14206 4326
rect 14262 4324 14268 4326
rect 13960 4304 14268 4324
rect 14384 4078 14412 4508
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 12256 3052 12308 3058
rect 13636 3052 13688 3058
rect 12256 2994 12308 3000
rect 13556 3012 13636 3040
rect 12410 2748 12718 2768
rect 12410 2746 12416 2748
rect 12472 2746 12496 2748
rect 12552 2746 12576 2748
rect 12632 2746 12656 2748
rect 12712 2746 12718 2748
rect 12472 2694 12474 2746
rect 12654 2694 12656 2746
rect 12410 2692 12416 2694
rect 12472 2692 12496 2694
rect 12552 2692 12576 2694
rect 12632 2692 12656 2694
rect 12712 2692 12718 2694
rect 12410 2672 12718 2692
rect 12808 2508 12860 2514
rect 12808 2450 12860 2456
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 11428 2100 11480 2106
rect 11428 2042 11480 2048
rect 12728 1970 12756 2246
rect 10232 1964 10284 1970
rect 10232 1906 10284 1912
rect 11244 1964 11296 1970
rect 11244 1906 11296 1912
rect 12716 1964 12768 1970
rect 12716 1906 12768 1912
rect 10140 1760 10192 1766
rect 10140 1702 10192 1708
rect 9310 1660 9618 1680
rect 9310 1658 9316 1660
rect 9372 1658 9396 1660
rect 9452 1658 9476 1660
rect 9532 1658 9556 1660
rect 9612 1658 9618 1660
rect 9372 1606 9374 1658
rect 9554 1606 9556 1658
rect 9310 1604 9316 1606
rect 9372 1604 9396 1606
rect 9452 1604 9476 1606
rect 9532 1604 9556 1606
rect 9612 1604 9618 1606
rect 9310 1584 9618 1604
rect 10152 1562 10180 1702
rect 10140 1556 10192 1562
rect 10140 1498 10192 1504
rect 9218 1320 9274 1329
rect 10152 1290 10180 1498
rect 9218 1255 9274 1264
rect 10140 1284 10192 1290
rect 10140 1226 10192 1232
rect 9404 1216 9456 1222
rect 9404 1158 9456 1164
rect 9416 1018 9444 1158
rect 9404 1012 9456 1018
rect 9404 954 9456 960
rect 9680 944 9732 950
rect 9680 886 9732 892
rect 10138 912 10194 921
rect 9312 876 9364 882
rect 9312 818 9364 824
rect 9324 785 9352 818
rect 9310 776 9366 785
rect 9692 746 9720 886
rect 10138 847 10140 856
rect 10192 847 10194 856
rect 10140 818 10192 824
rect 10244 814 10272 1906
rect 12820 1902 12848 2450
rect 13556 1970 13584 3012
rect 13636 2994 13688 3000
rect 13740 2774 13768 3470
rect 13832 3058 13860 3470
rect 14108 3466 14136 3878
rect 14476 3738 14504 4422
rect 14568 4214 14596 4762
rect 14752 4690 14780 5714
rect 14936 5234 14964 10202
rect 15304 9586 15332 10406
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 15120 8090 15148 8502
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15028 7342 15056 7686
rect 15120 7478 15148 8026
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15120 7002 15148 7414
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15212 6458 15240 6598
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14648 4548 14700 4554
rect 14648 4490 14700 4496
rect 14660 4282 14688 4490
rect 14936 4282 14964 5170
rect 15028 4690 15056 5578
rect 15396 5574 15424 11206
rect 15580 11098 15608 11206
rect 15658 11200 15714 12000
rect 18510 11200 18566 12000
rect 18786 11248 18842 11257
rect 15672 11098 15700 11200
rect 15580 11070 15700 11098
rect 17060 10908 17368 10928
rect 17060 10906 17066 10908
rect 17122 10906 17146 10908
rect 17202 10906 17226 10908
rect 17282 10906 17306 10908
rect 17362 10906 17368 10908
rect 17122 10854 17124 10906
rect 17304 10854 17306 10906
rect 17060 10852 17066 10854
rect 17122 10852 17146 10854
rect 17202 10852 17226 10854
rect 17282 10852 17306 10854
rect 17362 10852 17368 10854
rect 17060 10832 17368 10852
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 15510 10364 15818 10384
rect 15510 10362 15516 10364
rect 15572 10362 15596 10364
rect 15652 10362 15676 10364
rect 15732 10362 15756 10364
rect 15812 10362 15818 10364
rect 15572 10310 15574 10362
rect 15754 10310 15756 10362
rect 15510 10308 15516 10310
rect 15572 10308 15596 10310
rect 15652 10308 15676 10310
rect 15732 10308 15756 10310
rect 15812 10308 15818 10310
rect 15510 10288 15818 10308
rect 16960 10130 16988 10406
rect 18064 10266 18092 10610
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16488 10056 16540 10062
rect 16540 10004 16620 10010
rect 16488 9998 16620 10004
rect 16500 9982 16620 9998
rect 16592 9722 16620 9982
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 17060 9820 17368 9840
rect 17060 9818 17066 9820
rect 17122 9818 17146 9820
rect 17202 9818 17226 9820
rect 17282 9818 17306 9820
rect 17362 9818 17368 9820
rect 17122 9766 17124 9818
rect 17304 9766 17306 9818
rect 17060 9764 17066 9766
rect 17122 9764 17146 9766
rect 17202 9764 17226 9766
rect 17282 9764 17306 9766
rect 17362 9764 17368 9766
rect 17060 9744 17368 9764
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 18340 9518 18368 9862
rect 18328 9512 18380 9518
rect 18328 9454 18380 9460
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 15510 9276 15818 9296
rect 15510 9274 15516 9276
rect 15572 9274 15596 9276
rect 15652 9274 15676 9276
rect 15732 9274 15756 9276
rect 15812 9274 15818 9276
rect 15572 9222 15574 9274
rect 15754 9222 15756 9274
rect 15510 9220 15516 9222
rect 15572 9220 15596 9222
rect 15652 9220 15676 9222
rect 15732 9220 15756 9222
rect 15812 9220 15818 9222
rect 15510 9200 15818 9220
rect 16684 9042 16712 9318
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8634 15884 8910
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15510 8188 15818 8208
rect 15510 8186 15516 8188
rect 15572 8186 15596 8188
rect 15652 8186 15676 8188
rect 15732 8186 15756 8188
rect 15812 8186 15818 8188
rect 15572 8134 15574 8186
rect 15754 8134 15756 8186
rect 15510 8132 15516 8134
rect 15572 8132 15596 8134
rect 15652 8132 15676 8134
rect 15732 8132 15756 8134
rect 15812 8132 15818 8134
rect 15510 8112 15818 8132
rect 16500 8090 16528 8842
rect 16684 8430 16712 8978
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 17060 8732 17368 8752
rect 17060 8730 17066 8732
rect 17122 8730 17146 8732
rect 17202 8730 17226 8732
rect 17282 8730 17306 8732
rect 17362 8730 17368 8732
rect 17122 8678 17124 8730
rect 17304 8678 17306 8730
rect 17060 8676 17066 8678
rect 17122 8676 17146 8678
rect 17202 8676 17226 8678
rect 17282 8676 17306 8678
rect 17362 8676 17368 8678
rect 17060 8656 17368 8676
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 16488 8084 16540 8090
rect 16540 8044 16620 8072
rect 16488 8026 16540 8032
rect 16592 7818 16620 8044
rect 16684 7954 16712 8366
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 16580 7812 16632 7818
rect 16580 7754 16632 7760
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 15510 7100 15818 7120
rect 15510 7098 15516 7100
rect 15572 7098 15596 7100
rect 15652 7098 15676 7100
rect 15732 7098 15756 7100
rect 15812 7098 15818 7100
rect 15572 7046 15574 7098
rect 15754 7046 15756 7098
rect 15510 7044 15516 7046
rect 15572 7044 15596 7046
rect 15652 7044 15676 7046
rect 15732 7044 15756 7046
rect 15812 7044 15818 7046
rect 15510 7024 15818 7044
rect 16132 7002 16160 7754
rect 17060 7644 17368 7664
rect 17060 7642 17066 7644
rect 17122 7642 17146 7644
rect 17202 7642 17226 7644
rect 17282 7642 17306 7644
rect 17362 7642 17368 7644
rect 17122 7590 17124 7642
rect 17304 7590 17306 7642
rect 17060 7588 17066 7590
rect 17122 7588 17146 7590
rect 17202 7588 17226 7590
rect 17282 7588 17306 7590
rect 17362 7588 17368 7590
rect 17060 7568 17368 7588
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 16120 6996 16172 7002
rect 16120 6938 16172 6944
rect 15856 6730 15884 6938
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 15510 6012 15818 6032
rect 15510 6010 15516 6012
rect 15572 6010 15596 6012
rect 15652 6010 15676 6012
rect 15732 6010 15756 6012
rect 15812 6010 15818 6012
rect 15572 5958 15574 6010
rect 15754 5958 15756 6010
rect 15510 5956 15516 5958
rect 15572 5956 15596 5958
rect 15652 5956 15676 5958
rect 15732 5956 15756 5958
rect 15812 5956 15818 5958
rect 15510 5936 15818 5956
rect 15856 5914 15884 6666
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15856 5574 15884 5850
rect 16316 5710 16344 7278
rect 17060 6556 17368 6576
rect 17060 6554 17066 6556
rect 17122 6554 17146 6556
rect 17202 6554 17226 6556
rect 17282 6554 17306 6556
rect 17362 6554 17368 6556
rect 17122 6502 17124 6554
rect 17304 6502 17306 6554
rect 17060 6500 17066 6502
rect 17122 6500 17146 6502
rect 17202 6500 17226 6502
rect 17282 6500 17306 6502
rect 17362 6500 17368 6502
rect 17060 6480 17368 6500
rect 17512 6254 17540 7754
rect 17880 6798 17908 8366
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 18064 6458 18092 8774
rect 18524 7206 18552 11200
rect 18786 11183 18842 11192
rect 18800 10674 18828 11183
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18616 9761 18644 9998
rect 18602 9752 18658 9761
rect 18602 9687 18658 9696
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18616 8265 18644 8434
rect 18602 8256 18658 8265
rect 18602 8191 18658 8200
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18328 6860 18380 6866
rect 18328 6802 18380 6808
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 18340 6254 18368 6802
rect 18512 6792 18564 6798
rect 18510 6760 18512 6769
rect 18564 6760 18566 6769
rect 18510 6695 18566 6704
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16408 5778 16436 6054
rect 17328 5914 17356 6190
rect 18156 5914 18184 6190
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15844 5568 15896 5574
rect 15844 5510 15896 5516
rect 15856 5302 15884 5510
rect 17060 5468 17368 5488
rect 17060 5466 17066 5468
rect 17122 5466 17146 5468
rect 17202 5466 17226 5468
rect 17282 5466 17306 5468
rect 17362 5466 17368 5468
rect 17122 5414 17124 5466
rect 17304 5414 17306 5466
rect 17060 5412 17066 5414
rect 17122 5412 17146 5414
rect 17202 5412 17226 5414
rect 17282 5412 17306 5414
rect 17362 5412 17368 5414
rect 17060 5392 17368 5412
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15660 5296 15712 5302
rect 15844 5296 15896 5302
rect 15712 5256 15844 5284
rect 15660 5238 15712 5244
rect 15844 5238 15896 5244
rect 15304 4758 15332 5238
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 15510 4924 15818 4944
rect 15510 4922 15516 4924
rect 15572 4922 15596 4924
rect 15652 4922 15676 4924
rect 15732 4922 15756 4924
rect 15812 4922 15818 4924
rect 15572 4870 15574 4922
rect 15754 4870 15756 4922
rect 15510 4868 15516 4870
rect 15572 4868 15596 4870
rect 15652 4868 15676 4870
rect 15732 4868 15756 4870
rect 15812 4868 15818 4870
rect 15510 4848 15818 4868
rect 15292 4752 15344 4758
rect 15292 4694 15344 4700
rect 15016 4684 15068 4690
rect 15016 4626 15068 4632
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 14556 4208 14608 4214
rect 14556 4150 14608 4156
rect 14832 4072 14884 4078
rect 14936 4060 14964 4218
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 14884 4032 14964 4060
rect 14832 4014 14884 4020
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14096 3460 14148 3466
rect 14096 3402 14148 3408
rect 13960 3292 14268 3312
rect 13960 3290 13966 3292
rect 14022 3290 14046 3292
rect 14102 3290 14126 3292
rect 14182 3290 14206 3292
rect 14262 3290 14268 3292
rect 14022 3238 14024 3290
rect 14204 3238 14206 3290
rect 13960 3236 13966 3238
rect 14022 3236 14046 3238
rect 14102 3236 14126 3238
rect 14182 3236 14206 3238
rect 14262 3236 14268 3238
rect 13960 3216 14268 3236
rect 14568 3126 14596 3946
rect 15120 3738 15148 4082
rect 15304 3738 15332 4694
rect 16684 4690 16712 4966
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 15844 4616 15896 4622
rect 15844 4558 15896 4564
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 14556 3120 14608 3126
rect 14556 3062 14608 3068
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 13832 2854 13860 2994
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13648 2746 13768 2774
rect 13648 2310 13676 2746
rect 14292 2514 14320 2926
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 14476 2258 14504 2994
rect 14568 2446 14596 3062
rect 15120 2854 15148 3674
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 15212 2378 15240 3062
rect 15304 2582 15332 3674
rect 15396 3194 15424 4490
rect 15764 4214 15792 4490
rect 15856 4282 15884 4558
rect 16580 4548 16632 4554
rect 16580 4490 16632 4496
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 15752 4208 15804 4214
rect 15752 4150 15804 4156
rect 15510 3836 15818 3856
rect 15510 3834 15516 3836
rect 15572 3834 15596 3836
rect 15652 3834 15676 3836
rect 15732 3834 15756 3836
rect 15812 3834 15818 3836
rect 15572 3782 15574 3834
rect 15754 3782 15756 3834
rect 15510 3780 15516 3782
rect 15572 3780 15596 3782
rect 15652 3780 15676 3782
rect 15732 3780 15756 3782
rect 15812 3780 15818 3782
rect 15510 3760 15818 3780
rect 15856 3534 15884 4218
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15510 2748 15818 2768
rect 15510 2746 15516 2748
rect 15572 2746 15596 2748
rect 15652 2746 15676 2748
rect 15732 2746 15756 2748
rect 15812 2746 15818 2748
rect 15572 2694 15574 2746
rect 15754 2694 15756 2746
rect 15510 2692 15516 2694
rect 15572 2692 15596 2694
rect 15652 2692 15676 2694
rect 15732 2692 15756 2694
rect 15812 2692 15818 2694
rect 15510 2672 15818 2692
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15856 2514 15884 3470
rect 15948 3194 15976 4422
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16132 3602 16160 3878
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 16592 3466 16620 4490
rect 17060 4380 17368 4400
rect 17060 4378 17066 4380
rect 17122 4378 17146 4380
rect 17202 4378 17226 4380
rect 17282 4378 17306 4380
rect 17362 4378 17368 4380
rect 17122 4326 17124 4378
rect 17304 4326 17306 4378
rect 17060 4324 17066 4326
rect 17122 4324 17146 4326
rect 17202 4324 17226 4326
rect 17282 4324 17306 4326
rect 17362 4324 17368 4326
rect 17060 4304 17368 4324
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 16580 3460 16632 3466
rect 16632 3420 16712 3448
rect 16580 3402 16632 3408
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 16500 2514 16528 3062
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15844 2508 15896 2514
rect 15844 2450 15896 2456
rect 16488 2508 16540 2514
rect 16488 2450 16540 2456
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 15292 2372 15344 2378
rect 15292 2314 15344 2320
rect 14924 2304 14976 2310
rect 13648 2106 13676 2246
rect 13960 2204 14268 2224
rect 13960 2202 13966 2204
rect 14022 2202 14046 2204
rect 14102 2202 14126 2204
rect 14182 2202 14206 2204
rect 14262 2202 14268 2204
rect 14022 2150 14024 2202
rect 14204 2150 14206 2202
rect 13960 2148 13966 2150
rect 14022 2148 14046 2150
rect 14102 2148 14126 2150
rect 14182 2148 14206 2150
rect 14262 2148 14268 2150
rect 13960 2128 14268 2148
rect 13636 2100 13688 2106
rect 13636 2042 13688 2048
rect 14384 1970 14412 2246
rect 14476 2230 14596 2258
rect 14924 2246 14976 2252
rect 12900 1964 12952 1970
rect 12900 1906 12952 1912
rect 13544 1964 13596 1970
rect 13544 1906 13596 1912
rect 14372 1964 14424 1970
rect 14372 1906 14424 1912
rect 10968 1896 11020 1902
rect 10968 1838 11020 1844
rect 12808 1896 12860 1902
rect 12808 1838 12860 1844
rect 10980 1358 11008 1838
rect 12164 1760 12216 1766
rect 12164 1702 12216 1708
rect 10416 1352 10468 1358
rect 10416 1294 10468 1300
rect 10968 1352 11020 1358
rect 10968 1294 11020 1300
rect 10428 882 10456 1294
rect 11520 1216 11572 1222
rect 11520 1158 11572 1164
rect 10860 1116 11168 1136
rect 10860 1114 10866 1116
rect 10922 1114 10946 1116
rect 11002 1114 11026 1116
rect 11082 1114 11106 1116
rect 11162 1114 11168 1116
rect 10922 1062 10924 1114
rect 11104 1062 11106 1114
rect 10860 1060 10866 1062
rect 10922 1060 10946 1062
rect 11002 1060 11026 1062
rect 11082 1060 11106 1062
rect 11162 1060 11168 1062
rect 10860 1040 11168 1060
rect 11532 950 11560 1158
rect 11520 944 11572 950
rect 11520 886 11572 892
rect 12176 882 12204 1702
rect 12410 1660 12718 1680
rect 12410 1658 12416 1660
rect 12472 1658 12496 1660
rect 12552 1658 12576 1660
rect 12632 1658 12656 1660
rect 12712 1658 12718 1660
rect 12472 1606 12474 1658
rect 12654 1606 12656 1658
rect 12410 1604 12416 1606
rect 12472 1604 12496 1606
rect 12552 1604 12576 1606
rect 12632 1604 12656 1606
rect 12712 1604 12718 1606
rect 12410 1584 12718 1604
rect 12348 1284 12400 1290
rect 12348 1226 12400 1232
rect 12360 1018 12388 1226
rect 12348 1012 12400 1018
rect 12348 954 12400 960
rect 10416 876 10468 882
rect 10416 818 10468 824
rect 11704 876 11756 882
rect 11704 818 11756 824
rect 11796 876 11848 882
rect 11796 818 11848 824
rect 12164 876 12216 882
rect 12164 818 12216 824
rect 10232 808 10284 814
rect 10232 750 10284 756
rect 9310 711 9366 720
rect 9680 740 9732 746
rect 9680 682 9732 688
rect 9128 672 9180 678
rect 9128 614 9180 620
rect 9956 672 10008 678
rect 9956 614 10008 620
rect 9034 368 9090 377
rect 9034 303 9090 312
rect 5908 264 5960 270
rect 5908 206 5960 212
rect 9048 202 9076 303
rect 9140 270 9168 614
rect 9310 572 9618 592
rect 9310 570 9316 572
rect 9372 570 9396 572
rect 9452 570 9476 572
rect 9532 570 9556 572
rect 9612 570 9618 572
rect 9372 518 9374 570
rect 9554 518 9556 570
rect 9310 516 9316 518
rect 9372 516 9396 518
rect 9452 516 9476 518
rect 9532 516 9556 518
rect 9612 516 9618 518
rect 9310 496 9618 516
rect 9968 270 9996 614
rect 11716 377 11744 818
rect 11808 746 11836 818
rect 12912 746 12940 1906
rect 13452 1352 13504 1358
rect 13452 1294 13504 1300
rect 13360 1216 13412 1222
rect 13360 1158 13412 1164
rect 13372 921 13400 1158
rect 13358 912 13414 921
rect 12992 876 13044 882
rect 12992 818 13044 824
rect 13268 876 13320 882
rect 13358 847 13414 856
rect 13268 818 13320 824
rect 11796 740 11848 746
rect 11796 682 11848 688
rect 12900 740 12952 746
rect 12900 682 12952 688
rect 11702 368 11758 377
rect 11702 303 11758 312
rect 9128 264 9180 270
rect 9128 206 9180 212
rect 9956 264 10008 270
rect 9956 206 10008 212
rect 11716 202 11744 303
rect 11808 270 11836 682
rect 12410 572 12718 592
rect 12410 570 12416 572
rect 12472 570 12496 572
rect 12552 570 12576 572
rect 12632 570 12656 572
rect 12712 570 12718 572
rect 12472 518 12474 570
rect 12654 518 12656 570
rect 12410 516 12416 518
rect 12472 516 12496 518
rect 12552 516 12576 518
rect 12632 516 12656 518
rect 12712 516 12718 518
rect 12410 496 12718 516
rect 12256 400 12308 406
rect 12254 368 12256 377
rect 12308 368 12310 377
rect 12254 303 12310 312
rect 11796 264 11848 270
rect 11796 206 11848 212
rect 13004 202 13032 818
rect 13280 270 13308 818
rect 13464 474 13492 1294
rect 13556 1018 13584 1906
rect 13820 1896 13872 1902
rect 13820 1838 13872 1844
rect 13832 1426 13860 1838
rect 13820 1420 13872 1426
rect 13820 1362 13872 1368
rect 13544 1012 13596 1018
rect 13544 954 13596 960
rect 13726 912 13782 921
rect 13726 847 13728 856
rect 13780 847 13782 856
rect 13728 818 13780 824
rect 13544 808 13596 814
rect 13544 750 13596 756
rect 13556 474 13584 750
rect 13452 468 13504 474
rect 13452 410 13504 416
rect 13544 468 13596 474
rect 13544 410 13596 416
rect 13740 270 13768 818
rect 13832 785 13860 1362
rect 14464 1352 14516 1358
rect 14464 1294 14516 1300
rect 13960 1116 14268 1136
rect 13960 1114 13966 1116
rect 14022 1114 14046 1116
rect 14102 1114 14126 1116
rect 14182 1114 14206 1116
rect 14262 1114 14268 1116
rect 14022 1062 14024 1114
rect 14204 1062 14206 1114
rect 13960 1060 13966 1062
rect 14022 1060 14046 1062
rect 14102 1060 14126 1062
rect 14182 1060 14206 1062
rect 14262 1060 14268 1062
rect 13960 1040 14268 1060
rect 14280 808 14332 814
rect 13818 776 13874 785
rect 13818 711 13874 720
rect 14278 776 14280 785
rect 14332 776 14334 785
rect 14476 746 14504 1294
rect 14568 1290 14596 2230
rect 14648 1964 14700 1970
rect 14648 1906 14700 1912
rect 14660 1562 14688 1906
rect 14832 1828 14884 1834
rect 14832 1770 14884 1776
rect 14648 1556 14700 1562
rect 14648 1498 14700 1504
rect 14556 1284 14608 1290
rect 14556 1226 14608 1232
rect 14568 814 14596 1226
rect 14844 950 14872 1770
rect 14936 1562 14964 2246
rect 14924 1556 14976 1562
rect 14924 1498 14976 1504
rect 15108 1488 15160 1494
rect 15108 1430 15160 1436
rect 15120 1358 15148 1430
rect 15212 1358 15240 2314
rect 15304 1902 15332 2314
rect 15580 1902 15608 2450
rect 16684 2378 16712 3420
rect 17060 3292 17368 3312
rect 17060 3290 17066 3292
rect 17122 3290 17146 3292
rect 17202 3290 17226 3292
rect 17282 3290 17306 3292
rect 17362 3290 17368 3292
rect 17122 3238 17124 3290
rect 17304 3238 17306 3290
rect 17060 3236 17066 3238
rect 17122 3236 17146 3238
rect 17202 3236 17226 3238
rect 17282 3236 17306 3238
rect 17362 3236 17368 3238
rect 17060 3216 17368 3236
rect 17512 3058 17540 3538
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 16120 2372 16172 2378
rect 16120 2314 16172 2320
rect 16672 2372 16724 2378
rect 16672 2314 16724 2320
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 15856 2106 15884 2246
rect 16132 2106 16160 2314
rect 15844 2100 15896 2106
rect 15844 2042 15896 2048
rect 16120 2100 16172 2106
rect 16120 2042 16172 2048
rect 16684 1970 16712 2314
rect 17060 2204 17368 2224
rect 17060 2202 17066 2204
rect 17122 2202 17146 2204
rect 17202 2202 17226 2204
rect 17282 2202 17306 2204
rect 17362 2202 17368 2204
rect 17122 2150 17124 2202
rect 17304 2150 17306 2202
rect 17060 2148 17066 2150
rect 17122 2148 17146 2150
rect 17202 2148 17226 2150
rect 17282 2148 17306 2150
rect 17362 2148 17368 2150
rect 17060 2128 17368 2148
rect 17880 2106 17908 2994
rect 18156 2106 18184 5306
rect 18510 5264 18566 5273
rect 18510 5199 18512 5208
rect 18564 5199 18566 5208
rect 18512 5170 18564 5176
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18524 3777 18552 4082
rect 18510 3768 18566 3777
rect 18510 3703 18566 3712
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18524 2281 18552 2382
rect 18510 2272 18566 2281
rect 18510 2207 18566 2216
rect 17500 2100 17552 2106
rect 17500 2042 17552 2048
rect 17868 2100 17920 2106
rect 17868 2042 17920 2048
rect 18144 2100 18196 2106
rect 18144 2042 18196 2048
rect 16672 1964 16724 1970
rect 16672 1906 16724 1912
rect 16948 1964 17000 1970
rect 16948 1906 17000 1912
rect 15292 1896 15344 1902
rect 15292 1838 15344 1844
rect 15568 1896 15620 1902
rect 15568 1838 15620 1844
rect 15384 1760 15436 1766
rect 15384 1702 15436 1708
rect 15936 1760 15988 1766
rect 15936 1702 15988 1708
rect 15396 1358 15424 1702
rect 15510 1660 15818 1680
rect 15510 1658 15516 1660
rect 15572 1658 15596 1660
rect 15652 1658 15676 1660
rect 15732 1658 15756 1660
rect 15812 1658 15818 1660
rect 15572 1606 15574 1658
rect 15754 1606 15756 1658
rect 15510 1604 15516 1606
rect 15572 1604 15596 1606
rect 15652 1604 15676 1606
rect 15732 1604 15756 1606
rect 15812 1604 15818 1606
rect 15510 1584 15818 1604
rect 15948 1358 15976 1702
rect 15108 1352 15160 1358
rect 15108 1294 15160 1300
rect 15200 1352 15252 1358
rect 15200 1294 15252 1300
rect 15384 1352 15436 1358
rect 15384 1294 15436 1300
rect 15936 1352 15988 1358
rect 15936 1294 15988 1300
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 16396 1352 16448 1358
rect 16396 1294 16448 1300
rect 14832 944 14884 950
rect 14832 886 14884 892
rect 14556 808 14608 814
rect 14556 750 14608 756
rect 14278 711 14334 720
rect 14464 740 14516 746
rect 14464 682 14516 688
rect 13268 264 13320 270
rect 13268 206 13320 212
rect 13728 264 13780 270
rect 13728 206 13780 212
rect 14476 202 14504 682
rect 15212 474 15240 1294
rect 16028 1216 16080 1222
rect 16028 1158 16080 1164
rect 15510 572 15818 592
rect 15510 570 15516 572
rect 15572 570 15596 572
rect 15652 570 15676 572
rect 15732 570 15756 572
rect 15812 570 15818 572
rect 15572 518 15574 570
rect 15754 518 15756 570
rect 15510 516 15516 518
rect 15572 516 15596 518
rect 15652 516 15676 518
rect 15732 516 15756 518
rect 15812 516 15818 518
rect 15510 496 15818 516
rect 15200 468 15252 474
rect 15200 410 15252 416
rect 15842 368 15898 377
rect 15842 303 15898 312
rect 15856 270 15884 303
rect 16040 270 16068 1158
rect 16132 474 16160 1294
rect 16212 808 16264 814
rect 16212 750 16264 756
rect 16120 468 16172 474
rect 16120 410 16172 416
rect 16224 270 16252 750
rect 16408 406 16436 1294
rect 16684 1290 16712 1906
rect 16672 1284 16724 1290
rect 16672 1226 16724 1232
rect 16684 1018 16712 1226
rect 16960 1018 16988 1906
rect 17060 1116 17368 1136
rect 17060 1114 17066 1116
rect 17122 1114 17146 1116
rect 17202 1114 17226 1116
rect 17282 1114 17306 1116
rect 17362 1114 17368 1116
rect 17122 1062 17124 1114
rect 17304 1062 17306 1114
rect 17060 1060 17066 1062
rect 17122 1060 17146 1062
rect 17202 1060 17226 1062
rect 17282 1060 17306 1062
rect 17362 1060 17368 1062
rect 17060 1040 17368 1060
rect 17512 1018 17540 2042
rect 18236 1964 18288 1970
rect 18236 1906 18288 1912
rect 17868 1284 17920 1290
rect 17868 1226 17920 1232
rect 16672 1012 16724 1018
rect 16672 954 16724 960
rect 16948 1012 17000 1018
rect 16948 954 17000 960
rect 17500 1012 17552 1018
rect 17500 954 17552 960
rect 17880 921 17908 1226
rect 18248 1018 18276 1906
rect 18236 1012 18288 1018
rect 18236 954 18288 960
rect 17866 912 17922 921
rect 17316 876 17368 882
rect 17866 847 17922 856
rect 18512 876 18564 882
rect 17316 818 17368 824
rect 16488 672 16540 678
rect 16488 614 16540 620
rect 16396 400 16448 406
rect 16396 342 16448 348
rect 16500 338 16528 614
rect 17328 474 17356 818
rect 17592 808 17644 814
rect 17590 776 17592 785
rect 17644 776 17646 785
rect 17590 711 17646 720
rect 17316 468 17368 474
rect 17316 410 17368 416
rect 16488 332 16540 338
rect 16488 274 16540 280
rect 17880 270 17908 847
rect 18512 818 18564 824
rect 18524 785 18552 818
rect 18510 776 18566 785
rect 18510 711 18566 720
rect 15844 264 15896 270
rect 15844 206 15896 212
rect 16028 264 16080 270
rect 16028 206 16080 212
rect 16212 264 16264 270
rect 16212 206 16264 212
rect 17868 264 17920 270
rect 17868 206 17920 212
rect 9036 196 9088 202
rect 9036 138 9088 144
rect 11704 196 11756 202
rect 11704 138 11756 144
rect 12992 196 13044 202
rect 12992 138 13044 144
rect 14464 196 14516 202
rect 14464 138 14516 144
rect 5356 128 5408 134
rect 5356 70 5408 76
rect 4660 28 4968 48
rect 4660 26 4666 28
rect 4722 26 4746 28
rect 4802 26 4826 28
rect 4882 26 4906 28
rect 4962 26 4968 28
rect 4722 -26 4724 26
rect 4904 -26 4906 26
rect 4660 -28 4666 -26
rect 4722 -28 4746 -26
rect 4802 -28 4826 -26
rect 4882 -28 4906 -26
rect 4962 -28 4968 -26
rect 4660 -48 4968 -28
rect 7760 28 8068 48
rect 7760 26 7766 28
rect 7822 26 7846 28
rect 7902 26 7926 28
rect 7982 26 8006 28
rect 8062 26 8068 28
rect 7822 -26 7824 26
rect 8004 -26 8006 26
rect 7760 -28 7766 -26
rect 7822 -28 7846 -26
rect 7902 -28 7926 -26
rect 7982 -28 8006 -26
rect 8062 -28 8068 -26
rect 7760 -48 8068 -28
rect 10860 28 11168 48
rect 10860 26 10866 28
rect 10922 26 10946 28
rect 11002 26 11026 28
rect 11082 26 11106 28
rect 11162 26 11168 28
rect 10922 -26 10924 26
rect 11104 -26 11106 26
rect 10860 -28 10866 -26
rect 10922 -28 10946 -26
rect 11002 -28 11026 -26
rect 11082 -28 11106 -26
rect 11162 -28 11168 -26
rect 10860 -48 11168 -28
rect 13960 28 14268 48
rect 13960 26 13966 28
rect 14022 26 14046 28
rect 14102 26 14126 28
rect 14182 26 14206 28
rect 14262 26 14268 28
rect 14022 -26 14024 26
rect 14204 -26 14206 26
rect 13960 -28 13966 -26
rect 14022 -28 14046 -26
rect 14102 -28 14126 -26
rect 14182 -28 14206 -26
rect 14262 -28 14268 -26
rect 13960 -48 14268 -28
rect 17060 28 17368 48
rect 17060 26 17066 28
rect 17122 26 17146 28
rect 17202 26 17226 28
rect 17282 26 17306 28
rect 17362 26 17368 28
rect 17122 -26 17124 26
rect 17304 -26 17306 26
rect 17060 -28 17066 -26
rect 17122 -28 17146 -26
rect 17202 -28 17226 -26
rect 17282 -28 17306 -26
rect 17362 -28 17368 -26
rect 17060 -48 17368 -28
<< via2 >>
rect 2502 9580 2558 9616
rect 2502 9560 2504 9580
rect 2504 9560 2556 9580
rect 2556 9560 2558 9580
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 3276 10362 3332 10364
rect 3356 10362 3412 10364
rect 3116 10310 3162 10362
rect 3162 10310 3172 10362
rect 3196 10310 3226 10362
rect 3226 10310 3238 10362
rect 3238 10310 3252 10362
rect 3276 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3332 10362
rect 3356 10310 3366 10362
rect 3366 10310 3412 10362
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 3276 10308 3332 10310
rect 3356 10308 3412 10310
rect 3146 9424 3202 9480
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 3276 9274 3332 9276
rect 3356 9274 3412 9276
rect 3116 9222 3162 9274
rect 3162 9222 3172 9274
rect 3196 9222 3226 9274
rect 3226 9222 3238 9274
rect 3238 9222 3252 9274
rect 3276 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3332 9274
rect 3356 9222 3366 9274
rect 3366 9222 3412 9274
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3276 9220 3332 9222
rect 3356 9220 3412 9222
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 3276 8186 3332 8188
rect 3356 8186 3412 8188
rect 3116 8134 3162 8186
rect 3162 8134 3172 8186
rect 3196 8134 3226 8186
rect 3226 8134 3238 8186
rect 3238 8134 3252 8186
rect 3276 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3332 8186
rect 3356 8134 3366 8186
rect 3366 8134 3412 8186
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 3276 8132 3332 8134
rect 3356 8132 3412 8134
rect 4666 10906 4722 10908
rect 4746 10906 4802 10908
rect 4826 10906 4882 10908
rect 4906 10906 4962 10908
rect 4666 10854 4712 10906
rect 4712 10854 4722 10906
rect 4746 10854 4776 10906
rect 4776 10854 4788 10906
rect 4788 10854 4802 10906
rect 4826 10854 4840 10906
rect 4840 10854 4852 10906
rect 4852 10854 4882 10906
rect 4906 10854 4916 10906
rect 4916 10854 4962 10906
rect 4666 10852 4722 10854
rect 4746 10852 4802 10854
rect 4826 10852 4882 10854
rect 4906 10852 4962 10854
rect 7766 10906 7822 10908
rect 7846 10906 7902 10908
rect 7926 10906 7982 10908
rect 8006 10906 8062 10908
rect 7766 10854 7812 10906
rect 7812 10854 7822 10906
rect 7846 10854 7876 10906
rect 7876 10854 7888 10906
rect 7888 10854 7902 10906
rect 7926 10854 7940 10906
rect 7940 10854 7952 10906
rect 7952 10854 7982 10906
rect 8006 10854 8016 10906
rect 8016 10854 8062 10906
rect 7766 10852 7822 10854
rect 7846 10852 7902 10854
rect 7926 10852 7982 10854
rect 8006 10852 8062 10854
rect 10866 10906 10922 10908
rect 10946 10906 11002 10908
rect 11026 10906 11082 10908
rect 11106 10906 11162 10908
rect 10866 10854 10912 10906
rect 10912 10854 10922 10906
rect 10946 10854 10976 10906
rect 10976 10854 10988 10906
rect 10988 10854 11002 10906
rect 11026 10854 11040 10906
rect 11040 10854 11052 10906
rect 11052 10854 11082 10906
rect 11106 10854 11116 10906
rect 11116 10854 11162 10906
rect 10866 10852 10922 10854
rect 10946 10852 11002 10854
rect 11026 10852 11082 10854
rect 11106 10852 11162 10854
rect 13966 10906 14022 10908
rect 14046 10906 14102 10908
rect 14126 10906 14182 10908
rect 14206 10906 14262 10908
rect 13966 10854 14012 10906
rect 14012 10854 14022 10906
rect 14046 10854 14076 10906
rect 14076 10854 14088 10906
rect 14088 10854 14102 10906
rect 14126 10854 14140 10906
rect 14140 10854 14152 10906
rect 14152 10854 14182 10906
rect 14206 10854 14216 10906
rect 14216 10854 14262 10906
rect 13966 10852 14022 10854
rect 14046 10852 14102 10854
rect 14126 10852 14182 10854
rect 14206 10852 14262 10854
rect 6216 10362 6272 10364
rect 6296 10362 6352 10364
rect 6376 10362 6432 10364
rect 6456 10362 6512 10364
rect 6216 10310 6262 10362
rect 6262 10310 6272 10362
rect 6296 10310 6326 10362
rect 6326 10310 6338 10362
rect 6338 10310 6352 10362
rect 6376 10310 6390 10362
rect 6390 10310 6402 10362
rect 6402 10310 6432 10362
rect 6456 10310 6466 10362
rect 6466 10310 6512 10362
rect 6216 10308 6272 10310
rect 6296 10308 6352 10310
rect 6376 10308 6432 10310
rect 6456 10308 6512 10310
rect 4666 9818 4722 9820
rect 4746 9818 4802 9820
rect 4826 9818 4882 9820
rect 4906 9818 4962 9820
rect 4666 9766 4712 9818
rect 4712 9766 4722 9818
rect 4746 9766 4776 9818
rect 4776 9766 4788 9818
rect 4788 9766 4802 9818
rect 4826 9766 4840 9818
rect 4840 9766 4852 9818
rect 4852 9766 4882 9818
rect 4906 9766 4916 9818
rect 4916 9766 4962 9818
rect 4666 9764 4722 9766
rect 4746 9764 4802 9766
rect 4826 9764 4882 9766
rect 4906 9764 4962 9766
rect 5538 9560 5594 9616
rect 7766 9818 7822 9820
rect 7846 9818 7902 9820
rect 7926 9818 7982 9820
rect 8006 9818 8062 9820
rect 7766 9766 7812 9818
rect 7812 9766 7822 9818
rect 7846 9766 7876 9818
rect 7876 9766 7888 9818
rect 7888 9766 7902 9818
rect 7926 9766 7940 9818
rect 7940 9766 7952 9818
rect 7952 9766 7982 9818
rect 8006 9766 8016 9818
rect 8016 9766 8062 9818
rect 7766 9764 7822 9766
rect 7846 9764 7902 9766
rect 7926 9764 7982 9766
rect 8006 9764 8062 9766
rect 9316 10362 9372 10364
rect 9396 10362 9452 10364
rect 9476 10362 9532 10364
rect 9556 10362 9612 10364
rect 9316 10310 9362 10362
rect 9362 10310 9372 10362
rect 9396 10310 9426 10362
rect 9426 10310 9438 10362
rect 9438 10310 9452 10362
rect 9476 10310 9490 10362
rect 9490 10310 9502 10362
rect 9502 10310 9532 10362
rect 9556 10310 9566 10362
rect 9566 10310 9612 10362
rect 9316 10308 9372 10310
rect 9396 10308 9452 10310
rect 9476 10308 9532 10310
rect 9556 10308 9612 10310
rect 4666 8730 4722 8732
rect 4746 8730 4802 8732
rect 4826 8730 4882 8732
rect 4906 8730 4962 8732
rect 4666 8678 4712 8730
rect 4712 8678 4722 8730
rect 4746 8678 4776 8730
rect 4776 8678 4788 8730
rect 4788 8678 4802 8730
rect 4826 8678 4840 8730
rect 4840 8678 4852 8730
rect 4852 8678 4882 8730
rect 4906 8678 4916 8730
rect 4916 8678 4962 8730
rect 4666 8676 4722 8678
rect 4746 8676 4802 8678
rect 4826 8676 4882 8678
rect 4906 8676 4962 8678
rect 4666 7642 4722 7644
rect 4746 7642 4802 7644
rect 4826 7642 4882 7644
rect 4906 7642 4962 7644
rect 4666 7590 4712 7642
rect 4712 7590 4722 7642
rect 4746 7590 4776 7642
rect 4776 7590 4788 7642
rect 4788 7590 4802 7642
rect 4826 7590 4840 7642
rect 4840 7590 4852 7642
rect 4852 7590 4882 7642
rect 4906 7590 4916 7642
rect 4916 7590 4962 7642
rect 4666 7588 4722 7590
rect 4746 7588 4802 7590
rect 4826 7588 4882 7590
rect 4906 7588 4962 7590
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 3276 7098 3332 7100
rect 3356 7098 3412 7100
rect 3116 7046 3162 7098
rect 3162 7046 3172 7098
rect 3196 7046 3226 7098
rect 3226 7046 3238 7098
rect 3238 7046 3252 7098
rect 3276 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3332 7098
rect 3356 7046 3366 7098
rect 3366 7046 3412 7098
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3276 7044 3332 7046
rect 3356 7044 3412 7046
rect 4666 6554 4722 6556
rect 4746 6554 4802 6556
rect 4826 6554 4882 6556
rect 4906 6554 4962 6556
rect 4666 6502 4712 6554
rect 4712 6502 4722 6554
rect 4746 6502 4776 6554
rect 4776 6502 4788 6554
rect 4788 6502 4802 6554
rect 4826 6502 4840 6554
rect 4840 6502 4852 6554
rect 4852 6502 4882 6554
rect 4906 6502 4916 6554
rect 4916 6502 4962 6554
rect 4666 6500 4722 6502
rect 4746 6500 4802 6502
rect 4826 6500 4882 6502
rect 4906 6500 4962 6502
rect 3422 6316 3478 6352
rect 3422 6296 3424 6316
rect 3424 6296 3476 6316
rect 3476 6296 3478 6316
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 3276 6010 3332 6012
rect 3356 6010 3412 6012
rect 3116 5958 3162 6010
rect 3162 5958 3172 6010
rect 3196 5958 3226 6010
rect 3226 5958 3238 6010
rect 3238 5958 3252 6010
rect 3276 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3332 6010
rect 3356 5958 3366 6010
rect 3366 5958 3412 6010
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 3276 5956 3332 5958
rect 3356 5956 3412 5958
rect 5998 9460 6000 9480
rect 6000 9460 6052 9480
rect 6052 9460 6054 9480
rect 5998 9424 6054 9460
rect 6216 9274 6272 9276
rect 6296 9274 6352 9276
rect 6376 9274 6432 9276
rect 6456 9274 6512 9276
rect 6216 9222 6262 9274
rect 6262 9222 6272 9274
rect 6296 9222 6326 9274
rect 6326 9222 6338 9274
rect 6338 9222 6352 9274
rect 6376 9222 6390 9274
rect 6390 9222 6402 9274
rect 6402 9222 6432 9274
rect 6456 9222 6466 9274
rect 6466 9222 6512 9274
rect 6216 9220 6272 9222
rect 6296 9220 6352 9222
rect 6376 9220 6432 9222
rect 6456 9220 6512 9222
rect 6216 8186 6272 8188
rect 6296 8186 6352 8188
rect 6376 8186 6432 8188
rect 6456 8186 6512 8188
rect 6216 8134 6262 8186
rect 6262 8134 6272 8186
rect 6296 8134 6326 8186
rect 6326 8134 6338 8186
rect 6338 8134 6352 8186
rect 6376 8134 6390 8186
rect 6390 8134 6402 8186
rect 6402 8134 6432 8186
rect 6456 8134 6466 8186
rect 6466 8134 6512 8186
rect 6216 8132 6272 8134
rect 6296 8132 6352 8134
rect 6376 8132 6432 8134
rect 6456 8132 6512 8134
rect 5170 6296 5226 6352
rect 6216 7098 6272 7100
rect 6296 7098 6352 7100
rect 6376 7098 6432 7100
rect 6456 7098 6512 7100
rect 6216 7046 6262 7098
rect 6262 7046 6272 7098
rect 6296 7046 6326 7098
rect 6326 7046 6338 7098
rect 6338 7046 6352 7098
rect 6376 7046 6390 7098
rect 6390 7046 6402 7098
rect 6402 7046 6432 7098
rect 6456 7046 6466 7098
rect 6466 7046 6512 7098
rect 6216 7044 6272 7046
rect 6296 7044 6352 7046
rect 6376 7044 6432 7046
rect 6456 7044 6512 7046
rect 6216 6010 6272 6012
rect 6296 6010 6352 6012
rect 6376 6010 6432 6012
rect 6456 6010 6512 6012
rect 6216 5958 6262 6010
rect 6262 5958 6272 6010
rect 6296 5958 6326 6010
rect 6326 5958 6338 6010
rect 6338 5958 6352 6010
rect 6376 5958 6390 6010
rect 6390 5958 6402 6010
rect 6402 5958 6432 6010
rect 6456 5958 6466 6010
rect 6466 5958 6512 6010
rect 6216 5956 6272 5958
rect 6296 5956 6352 5958
rect 6376 5956 6432 5958
rect 6456 5956 6512 5958
rect 4666 5466 4722 5468
rect 4746 5466 4802 5468
rect 4826 5466 4882 5468
rect 4906 5466 4962 5468
rect 4666 5414 4712 5466
rect 4712 5414 4722 5466
rect 4746 5414 4776 5466
rect 4776 5414 4788 5466
rect 4788 5414 4802 5466
rect 4826 5414 4840 5466
rect 4840 5414 4852 5466
rect 4852 5414 4882 5466
rect 4906 5414 4916 5466
rect 4916 5414 4962 5466
rect 4666 5412 4722 5414
rect 4746 5412 4802 5414
rect 4826 5412 4882 5414
rect 4906 5412 4962 5414
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 3276 4922 3332 4924
rect 3356 4922 3412 4924
rect 3116 4870 3162 4922
rect 3162 4870 3172 4922
rect 3196 4870 3226 4922
rect 3226 4870 3238 4922
rect 3238 4870 3252 4922
rect 3276 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3332 4922
rect 3356 4870 3366 4922
rect 3366 4870 3412 4922
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 3276 4868 3332 4870
rect 3356 4868 3412 4870
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 3276 3834 3332 3836
rect 3356 3834 3412 3836
rect 3116 3782 3162 3834
rect 3162 3782 3172 3834
rect 3196 3782 3226 3834
rect 3226 3782 3238 3834
rect 3238 3782 3252 3834
rect 3276 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3332 3834
rect 3356 3782 3366 3834
rect 3366 3782 3412 3834
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 3276 3780 3332 3782
rect 3356 3780 3412 3782
rect 9316 9274 9372 9276
rect 9396 9274 9452 9276
rect 9476 9274 9532 9276
rect 9556 9274 9612 9276
rect 9316 9222 9362 9274
rect 9362 9222 9372 9274
rect 9396 9222 9426 9274
rect 9426 9222 9438 9274
rect 9438 9222 9452 9274
rect 9476 9222 9490 9274
rect 9490 9222 9502 9274
rect 9502 9222 9532 9274
rect 9556 9222 9566 9274
rect 9566 9222 9612 9274
rect 9316 9220 9372 9222
rect 9396 9220 9452 9222
rect 9476 9220 9532 9222
rect 9556 9220 9612 9222
rect 7766 8730 7822 8732
rect 7846 8730 7902 8732
rect 7926 8730 7982 8732
rect 8006 8730 8062 8732
rect 7766 8678 7812 8730
rect 7812 8678 7822 8730
rect 7846 8678 7876 8730
rect 7876 8678 7888 8730
rect 7888 8678 7902 8730
rect 7926 8678 7940 8730
rect 7940 8678 7952 8730
rect 7952 8678 7982 8730
rect 8006 8678 8016 8730
rect 8016 8678 8062 8730
rect 7766 8676 7822 8678
rect 7846 8676 7902 8678
rect 7926 8676 7982 8678
rect 8006 8676 8062 8678
rect 7766 7642 7822 7644
rect 7846 7642 7902 7644
rect 7926 7642 7982 7644
rect 8006 7642 8062 7644
rect 7766 7590 7812 7642
rect 7812 7590 7822 7642
rect 7846 7590 7876 7642
rect 7876 7590 7888 7642
rect 7888 7590 7902 7642
rect 7926 7590 7940 7642
rect 7940 7590 7952 7642
rect 7952 7590 7982 7642
rect 8006 7590 8016 7642
rect 8016 7590 8062 7642
rect 7766 7588 7822 7590
rect 7846 7588 7902 7590
rect 7926 7588 7982 7590
rect 8006 7588 8062 7590
rect 7766 6554 7822 6556
rect 7846 6554 7902 6556
rect 7926 6554 7982 6556
rect 8006 6554 8062 6556
rect 7766 6502 7812 6554
rect 7812 6502 7822 6554
rect 7846 6502 7876 6554
rect 7876 6502 7888 6554
rect 7888 6502 7902 6554
rect 7926 6502 7940 6554
rect 7940 6502 7952 6554
rect 7952 6502 7982 6554
rect 8006 6502 8016 6554
rect 8016 6502 8062 6554
rect 7766 6500 7822 6502
rect 7846 6500 7902 6502
rect 7926 6500 7982 6502
rect 8006 6500 8062 6502
rect 10866 9818 10922 9820
rect 10946 9818 11002 9820
rect 11026 9818 11082 9820
rect 11106 9818 11162 9820
rect 10866 9766 10912 9818
rect 10912 9766 10922 9818
rect 10946 9766 10976 9818
rect 10976 9766 10988 9818
rect 10988 9766 11002 9818
rect 11026 9766 11040 9818
rect 11040 9766 11052 9818
rect 11052 9766 11082 9818
rect 11106 9766 11116 9818
rect 11116 9766 11162 9818
rect 10866 9764 10922 9766
rect 10946 9764 11002 9766
rect 11026 9764 11082 9766
rect 11106 9764 11162 9766
rect 9316 8186 9372 8188
rect 9396 8186 9452 8188
rect 9476 8186 9532 8188
rect 9556 8186 9612 8188
rect 9316 8134 9362 8186
rect 9362 8134 9372 8186
rect 9396 8134 9426 8186
rect 9426 8134 9438 8186
rect 9438 8134 9452 8186
rect 9476 8134 9490 8186
rect 9490 8134 9502 8186
rect 9502 8134 9532 8186
rect 9556 8134 9566 8186
rect 9566 8134 9612 8186
rect 9316 8132 9372 8134
rect 9396 8132 9452 8134
rect 9476 8132 9532 8134
rect 9556 8132 9612 8134
rect 9316 7098 9372 7100
rect 9396 7098 9452 7100
rect 9476 7098 9532 7100
rect 9556 7098 9612 7100
rect 9316 7046 9362 7098
rect 9362 7046 9372 7098
rect 9396 7046 9426 7098
rect 9426 7046 9438 7098
rect 9438 7046 9452 7098
rect 9476 7046 9490 7098
rect 9490 7046 9502 7098
rect 9502 7046 9532 7098
rect 9556 7046 9566 7098
rect 9566 7046 9612 7098
rect 9316 7044 9372 7046
rect 9396 7044 9452 7046
rect 9476 7044 9532 7046
rect 9556 7044 9612 7046
rect 7766 5466 7822 5468
rect 7846 5466 7902 5468
rect 7926 5466 7982 5468
rect 8006 5466 8062 5468
rect 7766 5414 7812 5466
rect 7812 5414 7822 5466
rect 7846 5414 7876 5466
rect 7876 5414 7888 5466
rect 7888 5414 7902 5466
rect 7926 5414 7940 5466
rect 7940 5414 7952 5466
rect 7952 5414 7982 5466
rect 8006 5414 8016 5466
rect 8016 5414 8062 5466
rect 7766 5412 7822 5414
rect 7846 5412 7902 5414
rect 7926 5412 7982 5414
rect 8006 5412 8062 5414
rect 9316 6010 9372 6012
rect 9396 6010 9452 6012
rect 9476 6010 9532 6012
rect 9556 6010 9612 6012
rect 9316 5958 9362 6010
rect 9362 5958 9372 6010
rect 9396 5958 9426 6010
rect 9426 5958 9438 6010
rect 9438 5958 9452 6010
rect 9476 5958 9490 6010
rect 9490 5958 9502 6010
rect 9502 5958 9532 6010
rect 9556 5958 9566 6010
rect 9566 5958 9612 6010
rect 9316 5956 9372 5958
rect 9396 5956 9452 5958
rect 9476 5956 9532 5958
rect 9556 5956 9612 5958
rect 10866 8730 10922 8732
rect 10946 8730 11002 8732
rect 11026 8730 11082 8732
rect 11106 8730 11162 8732
rect 10866 8678 10912 8730
rect 10912 8678 10922 8730
rect 10946 8678 10976 8730
rect 10976 8678 10988 8730
rect 10988 8678 11002 8730
rect 11026 8678 11040 8730
rect 11040 8678 11052 8730
rect 11052 8678 11082 8730
rect 11106 8678 11116 8730
rect 11116 8678 11162 8730
rect 10866 8676 10922 8678
rect 10946 8676 11002 8678
rect 11026 8676 11082 8678
rect 11106 8676 11162 8678
rect 10866 7642 10922 7644
rect 10946 7642 11002 7644
rect 11026 7642 11082 7644
rect 11106 7642 11162 7644
rect 10866 7590 10912 7642
rect 10912 7590 10922 7642
rect 10946 7590 10976 7642
rect 10976 7590 10988 7642
rect 10988 7590 11002 7642
rect 11026 7590 11040 7642
rect 11040 7590 11052 7642
rect 11052 7590 11082 7642
rect 11106 7590 11116 7642
rect 11116 7590 11162 7642
rect 10866 7588 10922 7590
rect 10946 7588 11002 7590
rect 11026 7588 11082 7590
rect 11106 7588 11162 7590
rect 12416 10362 12472 10364
rect 12496 10362 12552 10364
rect 12576 10362 12632 10364
rect 12656 10362 12712 10364
rect 12416 10310 12462 10362
rect 12462 10310 12472 10362
rect 12496 10310 12526 10362
rect 12526 10310 12538 10362
rect 12538 10310 12552 10362
rect 12576 10310 12590 10362
rect 12590 10310 12602 10362
rect 12602 10310 12632 10362
rect 12656 10310 12666 10362
rect 12666 10310 12712 10362
rect 12416 10308 12472 10310
rect 12496 10308 12552 10310
rect 12576 10308 12632 10310
rect 12656 10308 12712 10310
rect 6216 4922 6272 4924
rect 6296 4922 6352 4924
rect 6376 4922 6432 4924
rect 6456 4922 6512 4924
rect 6216 4870 6262 4922
rect 6262 4870 6272 4922
rect 6296 4870 6326 4922
rect 6326 4870 6338 4922
rect 6338 4870 6352 4922
rect 6376 4870 6390 4922
rect 6390 4870 6402 4922
rect 6402 4870 6432 4922
rect 6456 4870 6466 4922
rect 6466 4870 6512 4922
rect 6216 4868 6272 4870
rect 6296 4868 6352 4870
rect 6376 4868 6432 4870
rect 6456 4868 6512 4870
rect 4666 4378 4722 4380
rect 4746 4378 4802 4380
rect 4826 4378 4882 4380
rect 4906 4378 4962 4380
rect 4666 4326 4712 4378
rect 4712 4326 4722 4378
rect 4746 4326 4776 4378
rect 4776 4326 4788 4378
rect 4788 4326 4802 4378
rect 4826 4326 4840 4378
rect 4840 4326 4852 4378
rect 4852 4326 4882 4378
rect 4906 4326 4916 4378
rect 4916 4326 4962 4378
rect 4666 4324 4722 4326
rect 4746 4324 4802 4326
rect 4826 4324 4882 4326
rect 4906 4324 4962 4326
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 3276 2746 3332 2748
rect 3356 2746 3412 2748
rect 3116 2694 3162 2746
rect 3162 2694 3172 2746
rect 3196 2694 3226 2746
rect 3226 2694 3238 2746
rect 3238 2694 3252 2746
rect 3276 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3332 2746
rect 3356 2694 3366 2746
rect 3366 2694 3412 2746
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3276 2692 3332 2694
rect 3356 2692 3412 2694
rect 4666 3290 4722 3292
rect 4746 3290 4802 3292
rect 4826 3290 4882 3292
rect 4906 3290 4962 3292
rect 4666 3238 4712 3290
rect 4712 3238 4722 3290
rect 4746 3238 4776 3290
rect 4776 3238 4788 3290
rect 4788 3238 4802 3290
rect 4826 3238 4840 3290
rect 4840 3238 4852 3290
rect 4852 3238 4882 3290
rect 4906 3238 4916 3290
rect 4916 3238 4962 3290
rect 4666 3236 4722 3238
rect 4746 3236 4802 3238
rect 4826 3236 4882 3238
rect 4906 3236 4962 3238
rect 4666 2202 4722 2204
rect 4746 2202 4802 2204
rect 4826 2202 4882 2204
rect 4906 2202 4962 2204
rect 4666 2150 4712 2202
rect 4712 2150 4722 2202
rect 4746 2150 4776 2202
rect 4776 2150 4788 2202
rect 4788 2150 4802 2202
rect 4826 2150 4840 2202
rect 4840 2150 4852 2202
rect 4852 2150 4882 2202
rect 4906 2150 4916 2202
rect 4916 2150 4962 2202
rect 4666 2148 4722 2150
rect 4746 2148 4802 2150
rect 4826 2148 4882 2150
rect 4906 2148 4962 2150
rect 6216 3834 6272 3836
rect 6296 3834 6352 3836
rect 6376 3834 6432 3836
rect 6456 3834 6512 3836
rect 6216 3782 6262 3834
rect 6262 3782 6272 3834
rect 6296 3782 6326 3834
rect 6326 3782 6338 3834
rect 6338 3782 6352 3834
rect 6376 3782 6390 3834
rect 6390 3782 6402 3834
rect 6402 3782 6432 3834
rect 6456 3782 6466 3834
rect 6466 3782 6512 3834
rect 6216 3780 6272 3782
rect 6296 3780 6352 3782
rect 6376 3780 6432 3782
rect 6456 3780 6512 3782
rect 7766 4378 7822 4380
rect 7846 4378 7902 4380
rect 7926 4378 7982 4380
rect 8006 4378 8062 4380
rect 7766 4326 7812 4378
rect 7812 4326 7822 4378
rect 7846 4326 7876 4378
rect 7876 4326 7888 4378
rect 7888 4326 7902 4378
rect 7926 4326 7940 4378
rect 7940 4326 7952 4378
rect 7952 4326 7982 4378
rect 8006 4326 8016 4378
rect 8016 4326 8062 4378
rect 7766 4324 7822 4326
rect 7846 4324 7902 4326
rect 7926 4324 7982 4326
rect 8006 4324 8062 4326
rect 9316 4922 9372 4924
rect 9396 4922 9452 4924
rect 9476 4922 9532 4924
rect 9556 4922 9612 4924
rect 9316 4870 9362 4922
rect 9362 4870 9372 4922
rect 9396 4870 9426 4922
rect 9426 4870 9438 4922
rect 9438 4870 9452 4922
rect 9476 4870 9490 4922
rect 9490 4870 9502 4922
rect 9502 4870 9532 4922
rect 9556 4870 9566 4922
rect 9566 4870 9612 4922
rect 9316 4868 9372 4870
rect 9396 4868 9452 4870
rect 9476 4868 9532 4870
rect 9556 4868 9612 4870
rect 3116 1658 3172 1660
rect 3196 1658 3252 1660
rect 3276 1658 3332 1660
rect 3356 1658 3412 1660
rect 3116 1606 3162 1658
rect 3162 1606 3172 1658
rect 3196 1606 3226 1658
rect 3226 1606 3238 1658
rect 3238 1606 3252 1658
rect 3276 1606 3290 1658
rect 3290 1606 3302 1658
rect 3302 1606 3332 1658
rect 3356 1606 3366 1658
rect 3366 1606 3412 1658
rect 3116 1604 3172 1606
rect 3196 1604 3252 1606
rect 3276 1604 3332 1606
rect 3356 1604 3412 1606
rect 4666 1114 4722 1116
rect 4746 1114 4802 1116
rect 4826 1114 4882 1116
rect 4906 1114 4962 1116
rect 4666 1062 4712 1114
rect 4712 1062 4722 1114
rect 4746 1062 4776 1114
rect 4776 1062 4788 1114
rect 4788 1062 4802 1114
rect 4826 1062 4840 1114
rect 4840 1062 4852 1114
rect 4852 1062 4882 1114
rect 4906 1062 4916 1114
rect 4916 1062 4962 1114
rect 4666 1060 4722 1062
rect 4746 1060 4802 1062
rect 4826 1060 4882 1062
rect 4906 1060 4962 1062
rect 4894 876 4950 912
rect 4894 856 4896 876
rect 4896 856 4948 876
rect 4948 856 4950 876
rect 3116 570 3172 572
rect 3196 570 3252 572
rect 3276 570 3332 572
rect 3356 570 3412 572
rect 3116 518 3162 570
rect 3162 518 3172 570
rect 3196 518 3226 570
rect 3226 518 3238 570
rect 3238 518 3252 570
rect 3276 518 3290 570
rect 3290 518 3302 570
rect 3302 518 3332 570
rect 3356 518 3366 570
rect 3366 518 3412 570
rect 3116 516 3172 518
rect 3196 516 3252 518
rect 3276 516 3332 518
rect 3356 516 3412 518
rect 5262 856 5318 912
rect 6216 2746 6272 2748
rect 6296 2746 6352 2748
rect 6376 2746 6432 2748
rect 6456 2746 6512 2748
rect 6216 2694 6262 2746
rect 6262 2694 6272 2746
rect 6296 2694 6326 2746
rect 6326 2694 6338 2746
rect 6338 2694 6352 2746
rect 6376 2694 6390 2746
rect 6390 2694 6402 2746
rect 6402 2694 6432 2746
rect 6456 2694 6466 2746
rect 6466 2694 6512 2746
rect 6216 2692 6272 2694
rect 6296 2692 6352 2694
rect 6376 2692 6432 2694
rect 6456 2692 6512 2694
rect 6216 1658 6272 1660
rect 6296 1658 6352 1660
rect 6376 1658 6432 1660
rect 6456 1658 6512 1660
rect 6216 1606 6262 1658
rect 6262 1606 6272 1658
rect 6296 1606 6326 1658
rect 6326 1606 6338 1658
rect 6338 1606 6352 1658
rect 6376 1606 6390 1658
rect 6390 1606 6402 1658
rect 6402 1606 6432 1658
rect 6456 1606 6466 1658
rect 6466 1606 6512 1658
rect 6216 1604 6272 1606
rect 6296 1604 6352 1606
rect 6376 1604 6432 1606
rect 6456 1604 6512 1606
rect 7766 3290 7822 3292
rect 7846 3290 7902 3292
rect 7926 3290 7982 3292
rect 8006 3290 8062 3292
rect 7766 3238 7812 3290
rect 7812 3238 7822 3290
rect 7846 3238 7876 3290
rect 7876 3238 7888 3290
rect 7888 3238 7902 3290
rect 7926 3238 7940 3290
rect 7940 3238 7952 3290
rect 7952 3238 7982 3290
rect 8006 3238 8016 3290
rect 8016 3238 8062 3290
rect 7766 3236 7822 3238
rect 7846 3236 7902 3238
rect 7926 3236 7982 3238
rect 8006 3236 8062 3238
rect 7766 2202 7822 2204
rect 7846 2202 7902 2204
rect 7926 2202 7982 2204
rect 8006 2202 8062 2204
rect 7766 2150 7812 2202
rect 7812 2150 7822 2202
rect 7846 2150 7876 2202
rect 7876 2150 7888 2202
rect 7888 2150 7902 2202
rect 7926 2150 7940 2202
rect 7940 2150 7952 2202
rect 7952 2150 7982 2202
rect 8006 2150 8016 2202
rect 8016 2150 8062 2202
rect 7766 2148 7822 2150
rect 7846 2148 7902 2150
rect 7926 2148 7982 2150
rect 8006 2148 8062 2150
rect 7010 1300 7012 1320
rect 7012 1300 7064 1320
rect 7064 1300 7066 1320
rect 7010 1264 7066 1300
rect 8666 3576 8722 3632
rect 9034 3460 9090 3496
rect 9034 3440 9036 3460
rect 9036 3440 9088 3460
rect 9088 3440 9090 3460
rect 8942 3068 8944 3088
rect 8944 3068 8996 3088
rect 8996 3068 8998 3088
rect 8942 3032 8998 3068
rect 7766 1114 7822 1116
rect 7846 1114 7902 1116
rect 7926 1114 7982 1116
rect 8006 1114 8062 1116
rect 7766 1062 7812 1114
rect 7812 1062 7822 1114
rect 7846 1062 7876 1114
rect 7876 1062 7888 1114
rect 7888 1062 7902 1114
rect 7926 1062 7940 1114
rect 7940 1062 7952 1114
rect 7952 1062 7982 1114
rect 8006 1062 8016 1114
rect 8016 1062 8062 1114
rect 7766 1060 7822 1062
rect 7846 1060 7902 1062
rect 7926 1060 7982 1062
rect 8006 1060 8062 1062
rect 7746 876 7802 912
rect 7746 856 7748 876
rect 7748 856 7800 876
rect 7800 856 7802 876
rect 6216 570 6272 572
rect 6296 570 6352 572
rect 6376 570 6432 572
rect 6456 570 6512 572
rect 6216 518 6262 570
rect 6262 518 6272 570
rect 6296 518 6326 570
rect 6326 518 6338 570
rect 6338 518 6352 570
rect 6376 518 6390 570
rect 6390 518 6402 570
rect 6402 518 6432 570
rect 6456 518 6466 570
rect 6466 518 6512 570
rect 6216 516 6272 518
rect 6296 516 6352 518
rect 6376 516 6432 518
rect 6456 516 6512 518
rect 8758 1264 8814 1320
rect 9316 3834 9372 3836
rect 9396 3834 9452 3836
rect 9476 3834 9532 3836
rect 9556 3834 9612 3836
rect 9316 3782 9362 3834
rect 9362 3782 9372 3834
rect 9396 3782 9426 3834
rect 9426 3782 9438 3834
rect 9438 3782 9452 3834
rect 9476 3782 9490 3834
rect 9490 3782 9502 3834
rect 9502 3782 9532 3834
rect 9556 3782 9566 3834
rect 9566 3782 9612 3834
rect 9316 3780 9372 3782
rect 9396 3780 9452 3782
rect 9476 3780 9532 3782
rect 9556 3780 9612 3782
rect 9316 2746 9372 2748
rect 9396 2746 9452 2748
rect 9476 2746 9532 2748
rect 9556 2746 9612 2748
rect 9316 2694 9362 2746
rect 9362 2694 9372 2746
rect 9396 2694 9426 2746
rect 9426 2694 9438 2746
rect 9438 2694 9452 2746
rect 9476 2694 9490 2746
rect 9490 2694 9502 2746
rect 9502 2694 9532 2746
rect 9556 2694 9566 2746
rect 9566 2694 9612 2746
rect 9316 2692 9372 2694
rect 9396 2692 9452 2694
rect 9476 2692 9532 2694
rect 9556 2692 9612 2694
rect 10866 6554 10922 6556
rect 10946 6554 11002 6556
rect 11026 6554 11082 6556
rect 11106 6554 11162 6556
rect 10866 6502 10912 6554
rect 10912 6502 10922 6554
rect 10946 6502 10976 6554
rect 10976 6502 10988 6554
rect 10988 6502 11002 6554
rect 11026 6502 11040 6554
rect 11040 6502 11052 6554
rect 11052 6502 11082 6554
rect 11106 6502 11116 6554
rect 11116 6502 11162 6554
rect 10866 6500 10922 6502
rect 10946 6500 11002 6502
rect 11026 6500 11082 6502
rect 11106 6500 11162 6502
rect 10866 5466 10922 5468
rect 10946 5466 11002 5468
rect 11026 5466 11082 5468
rect 11106 5466 11162 5468
rect 10866 5414 10912 5466
rect 10912 5414 10922 5466
rect 10946 5414 10976 5466
rect 10976 5414 10988 5466
rect 10988 5414 11002 5466
rect 11026 5414 11040 5466
rect 11040 5414 11052 5466
rect 11052 5414 11082 5466
rect 11106 5414 11116 5466
rect 11116 5414 11162 5466
rect 10866 5412 10922 5414
rect 10946 5412 11002 5414
rect 11026 5412 11082 5414
rect 11106 5412 11162 5414
rect 13966 9818 14022 9820
rect 14046 9818 14102 9820
rect 14126 9818 14182 9820
rect 14206 9818 14262 9820
rect 13966 9766 14012 9818
rect 14012 9766 14022 9818
rect 14046 9766 14076 9818
rect 14076 9766 14088 9818
rect 14088 9766 14102 9818
rect 14126 9766 14140 9818
rect 14140 9766 14152 9818
rect 14152 9766 14182 9818
rect 14206 9766 14216 9818
rect 14216 9766 14262 9818
rect 13966 9764 14022 9766
rect 14046 9764 14102 9766
rect 14126 9764 14182 9766
rect 14206 9764 14262 9766
rect 12416 9274 12472 9276
rect 12496 9274 12552 9276
rect 12576 9274 12632 9276
rect 12656 9274 12712 9276
rect 12416 9222 12462 9274
rect 12462 9222 12472 9274
rect 12496 9222 12526 9274
rect 12526 9222 12538 9274
rect 12538 9222 12552 9274
rect 12576 9222 12590 9274
rect 12590 9222 12602 9274
rect 12602 9222 12632 9274
rect 12656 9222 12666 9274
rect 12666 9222 12712 9274
rect 12416 9220 12472 9222
rect 12496 9220 12552 9222
rect 12576 9220 12632 9222
rect 12656 9220 12712 9222
rect 13966 8730 14022 8732
rect 14046 8730 14102 8732
rect 14126 8730 14182 8732
rect 14206 8730 14262 8732
rect 13966 8678 14012 8730
rect 14012 8678 14022 8730
rect 14046 8678 14076 8730
rect 14076 8678 14088 8730
rect 14088 8678 14102 8730
rect 14126 8678 14140 8730
rect 14140 8678 14152 8730
rect 14152 8678 14182 8730
rect 14206 8678 14216 8730
rect 14216 8678 14262 8730
rect 13966 8676 14022 8678
rect 14046 8676 14102 8678
rect 14126 8676 14182 8678
rect 14206 8676 14262 8678
rect 12416 8186 12472 8188
rect 12496 8186 12552 8188
rect 12576 8186 12632 8188
rect 12656 8186 12712 8188
rect 12416 8134 12462 8186
rect 12462 8134 12472 8186
rect 12496 8134 12526 8186
rect 12526 8134 12538 8186
rect 12538 8134 12552 8186
rect 12576 8134 12590 8186
rect 12590 8134 12602 8186
rect 12602 8134 12632 8186
rect 12656 8134 12666 8186
rect 12666 8134 12712 8186
rect 12416 8132 12472 8134
rect 12496 8132 12552 8134
rect 12576 8132 12632 8134
rect 12656 8132 12712 8134
rect 12416 7098 12472 7100
rect 12496 7098 12552 7100
rect 12576 7098 12632 7100
rect 12656 7098 12712 7100
rect 12416 7046 12462 7098
rect 12462 7046 12472 7098
rect 12496 7046 12526 7098
rect 12526 7046 12538 7098
rect 12538 7046 12552 7098
rect 12576 7046 12590 7098
rect 12590 7046 12602 7098
rect 12602 7046 12632 7098
rect 12656 7046 12666 7098
rect 12666 7046 12712 7098
rect 12416 7044 12472 7046
rect 12496 7044 12552 7046
rect 12576 7044 12632 7046
rect 12656 7044 12712 7046
rect 13634 7404 13690 7440
rect 13634 7384 13636 7404
rect 13636 7384 13688 7404
rect 13688 7384 13690 7404
rect 13966 7642 14022 7644
rect 14046 7642 14102 7644
rect 14126 7642 14182 7644
rect 14206 7642 14262 7644
rect 13966 7590 14012 7642
rect 14012 7590 14022 7642
rect 14046 7590 14076 7642
rect 14076 7590 14088 7642
rect 14088 7590 14102 7642
rect 14126 7590 14140 7642
rect 14140 7590 14152 7642
rect 14152 7590 14182 7642
rect 14206 7590 14216 7642
rect 14216 7590 14262 7642
rect 13966 7588 14022 7590
rect 14046 7588 14102 7590
rect 14126 7588 14182 7590
rect 14206 7588 14262 7590
rect 13910 7404 13966 7440
rect 13910 7384 13912 7404
rect 13912 7384 13964 7404
rect 13964 7384 13966 7404
rect 13966 6554 14022 6556
rect 14046 6554 14102 6556
rect 14126 6554 14182 6556
rect 14206 6554 14262 6556
rect 13966 6502 14012 6554
rect 14012 6502 14022 6554
rect 14046 6502 14076 6554
rect 14076 6502 14088 6554
rect 14088 6502 14102 6554
rect 14126 6502 14140 6554
rect 14140 6502 14152 6554
rect 14152 6502 14182 6554
rect 14206 6502 14216 6554
rect 14216 6502 14262 6554
rect 13966 6500 14022 6502
rect 14046 6500 14102 6502
rect 14126 6500 14182 6502
rect 14206 6500 14262 6502
rect 12416 6010 12472 6012
rect 12496 6010 12552 6012
rect 12576 6010 12632 6012
rect 12656 6010 12712 6012
rect 12416 5958 12462 6010
rect 12462 5958 12472 6010
rect 12496 5958 12526 6010
rect 12526 5958 12538 6010
rect 12538 5958 12552 6010
rect 12576 5958 12590 6010
rect 12590 5958 12602 6010
rect 12602 5958 12632 6010
rect 12656 5958 12666 6010
rect 12666 5958 12712 6010
rect 12416 5956 12472 5958
rect 12496 5956 12552 5958
rect 12576 5956 12632 5958
rect 12656 5956 12712 5958
rect 10866 4378 10922 4380
rect 10946 4378 11002 4380
rect 11026 4378 11082 4380
rect 11106 4378 11162 4380
rect 10866 4326 10912 4378
rect 10912 4326 10922 4378
rect 10946 4326 10976 4378
rect 10976 4326 10988 4378
rect 10988 4326 11002 4378
rect 11026 4326 11040 4378
rect 11040 4326 11052 4378
rect 11052 4326 11082 4378
rect 11106 4326 11116 4378
rect 11116 4326 11162 4378
rect 10866 4324 10922 4326
rect 10946 4324 11002 4326
rect 11026 4324 11082 4326
rect 11106 4324 11162 4326
rect 9770 3476 9772 3496
rect 9772 3476 9824 3496
rect 9824 3476 9826 3496
rect 9770 3440 9826 3476
rect 13966 5466 14022 5468
rect 14046 5466 14102 5468
rect 14126 5466 14182 5468
rect 14206 5466 14262 5468
rect 13966 5414 14012 5466
rect 14012 5414 14022 5466
rect 14046 5414 14076 5466
rect 14076 5414 14088 5466
rect 14088 5414 14102 5466
rect 14126 5414 14140 5466
rect 14140 5414 14152 5466
rect 14152 5414 14182 5466
rect 14206 5414 14216 5466
rect 14216 5414 14262 5466
rect 13966 5412 14022 5414
rect 14046 5412 14102 5414
rect 14126 5412 14182 5414
rect 14206 5412 14262 5414
rect 10866 3290 10922 3292
rect 10946 3290 11002 3292
rect 11026 3290 11082 3292
rect 11106 3290 11162 3292
rect 10866 3238 10912 3290
rect 10912 3238 10922 3290
rect 10946 3238 10976 3290
rect 10976 3238 10988 3290
rect 10988 3238 11002 3290
rect 11026 3238 11040 3290
rect 11040 3238 11052 3290
rect 11052 3238 11082 3290
rect 11106 3238 11116 3290
rect 11116 3238 11162 3290
rect 10866 3236 10922 3238
rect 10946 3236 11002 3238
rect 11026 3236 11082 3238
rect 11106 3236 11162 3238
rect 10874 3032 10930 3088
rect 11150 3052 11206 3088
rect 11150 3032 11152 3052
rect 11152 3032 11204 3052
rect 11204 3032 11206 3052
rect 11518 3460 11574 3496
rect 11518 3440 11520 3460
rect 11520 3440 11572 3460
rect 11572 3440 11574 3460
rect 12416 4922 12472 4924
rect 12496 4922 12552 4924
rect 12576 4922 12632 4924
rect 12656 4922 12712 4924
rect 12416 4870 12462 4922
rect 12462 4870 12472 4922
rect 12496 4870 12526 4922
rect 12526 4870 12538 4922
rect 12538 4870 12552 4922
rect 12576 4870 12590 4922
rect 12590 4870 12602 4922
rect 12602 4870 12632 4922
rect 12656 4870 12666 4922
rect 12666 4870 12712 4922
rect 12416 4868 12472 4870
rect 12496 4868 12552 4870
rect 12576 4868 12632 4870
rect 12656 4868 12712 4870
rect 10866 2202 10922 2204
rect 10946 2202 11002 2204
rect 11026 2202 11082 2204
rect 11106 2202 11162 2204
rect 10866 2150 10912 2202
rect 10912 2150 10922 2202
rect 10946 2150 10976 2202
rect 10976 2150 10988 2202
rect 10988 2150 11002 2202
rect 11026 2150 11040 2202
rect 11040 2150 11052 2202
rect 11052 2150 11082 2202
rect 11106 2150 11116 2202
rect 11116 2150 11162 2202
rect 10866 2148 10922 2150
rect 10946 2148 11002 2150
rect 11026 2148 11082 2150
rect 11106 2148 11162 2150
rect 12416 3834 12472 3836
rect 12496 3834 12552 3836
rect 12576 3834 12632 3836
rect 12656 3834 12712 3836
rect 12416 3782 12462 3834
rect 12462 3782 12472 3834
rect 12496 3782 12526 3834
rect 12526 3782 12538 3834
rect 12538 3782 12552 3834
rect 12576 3782 12590 3834
rect 12590 3782 12602 3834
rect 12602 3782 12632 3834
rect 12656 3782 12666 3834
rect 12666 3782 12712 3834
rect 12416 3780 12472 3782
rect 12496 3780 12552 3782
rect 12576 3780 12632 3782
rect 12656 3780 12712 3782
rect 12346 3596 12402 3632
rect 12346 3576 12348 3596
rect 12348 3576 12400 3596
rect 12400 3576 12402 3596
rect 13450 3476 13452 3496
rect 13452 3476 13504 3496
rect 13504 3476 13506 3496
rect 13450 3440 13506 3476
rect 13966 4378 14022 4380
rect 14046 4378 14102 4380
rect 14126 4378 14182 4380
rect 14206 4378 14262 4380
rect 13966 4326 14012 4378
rect 14012 4326 14022 4378
rect 14046 4326 14076 4378
rect 14076 4326 14088 4378
rect 14088 4326 14102 4378
rect 14126 4326 14140 4378
rect 14140 4326 14152 4378
rect 14152 4326 14182 4378
rect 14206 4326 14216 4378
rect 14216 4326 14262 4378
rect 13966 4324 14022 4326
rect 14046 4324 14102 4326
rect 14126 4324 14182 4326
rect 14206 4324 14262 4326
rect 12416 2746 12472 2748
rect 12496 2746 12552 2748
rect 12576 2746 12632 2748
rect 12656 2746 12712 2748
rect 12416 2694 12462 2746
rect 12462 2694 12472 2746
rect 12496 2694 12526 2746
rect 12526 2694 12538 2746
rect 12538 2694 12552 2746
rect 12576 2694 12590 2746
rect 12590 2694 12602 2746
rect 12602 2694 12632 2746
rect 12656 2694 12666 2746
rect 12666 2694 12712 2746
rect 12416 2692 12472 2694
rect 12496 2692 12552 2694
rect 12576 2692 12632 2694
rect 12656 2692 12712 2694
rect 9316 1658 9372 1660
rect 9396 1658 9452 1660
rect 9476 1658 9532 1660
rect 9556 1658 9612 1660
rect 9316 1606 9362 1658
rect 9362 1606 9372 1658
rect 9396 1606 9426 1658
rect 9426 1606 9438 1658
rect 9438 1606 9452 1658
rect 9476 1606 9490 1658
rect 9490 1606 9502 1658
rect 9502 1606 9532 1658
rect 9556 1606 9566 1658
rect 9566 1606 9612 1658
rect 9316 1604 9372 1606
rect 9396 1604 9452 1606
rect 9476 1604 9532 1606
rect 9556 1604 9612 1606
rect 9218 1264 9274 1320
rect 9310 720 9366 776
rect 10138 876 10194 912
rect 10138 856 10140 876
rect 10140 856 10192 876
rect 10192 856 10194 876
rect 17066 10906 17122 10908
rect 17146 10906 17202 10908
rect 17226 10906 17282 10908
rect 17306 10906 17362 10908
rect 17066 10854 17112 10906
rect 17112 10854 17122 10906
rect 17146 10854 17176 10906
rect 17176 10854 17188 10906
rect 17188 10854 17202 10906
rect 17226 10854 17240 10906
rect 17240 10854 17252 10906
rect 17252 10854 17282 10906
rect 17306 10854 17316 10906
rect 17316 10854 17362 10906
rect 17066 10852 17122 10854
rect 17146 10852 17202 10854
rect 17226 10852 17282 10854
rect 17306 10852 17362 10854
rect 15516 10362 15572 10364
rect 15596 10362 15652 10364
rect 15676 10362 15732 10364
rect 15756 10362 15812 10364
rect 15516 10310 15562 10362
rect 15562 10310 15572 10362
rect 15596 10310 15626 10362
rect 15626 10310 15638 10362
rect 15638 10310 15652 10362
rect 15676 10310 15690 10362
rect 15690 10310 15702 10362
rect 15702 10310 15732 10362
rect 15756 10310 15766 10362
rect 15766 10310 15812 10362
rect 15516 10308 15572 10310
rect 15596 10308 15652 10310
rect 15676 10308 15732 10310
rect 15756 10308 15812 10310
rect 17066 9818 17122 9820
rect 17146 9818 17202 9820
rect 17226 9818 17282 9820
rect 17306 9818 17362 9820
rect 17066 9766 17112 9818
rect 17112 9766 17122 9818
rect 17146 9766 17176 9818
rect 17176 9766 17188 9818
rect 17188 9766 17202 9818
rect 17226 9766 17240 9818
rect 17240 9766 17252 9818
rect 17252 9766 17282 9818
rect 17306 9766 17316 9818
rect 17316 9766 17362 9818
rect 17066 9764 17122 9766
rect 17146 9764 17202 9766
rect 17226 9764 17282 9766
rect 17306 9764 17362 9766
rect 15516 9274 15572 9276
rect 15596 9274 15652 9276
rect 15676 9274 15732 9276
rect 15756 9274 15812 9276
rect 15516 9222 15562 9274
rect 15562 9222 15572 9274
rect 15596 9222 15626 9274
rect 15626 9222 15638 9274
rect 15638 9222 15652 9274
rect 15676 9222 15690 9274
rect 15690 9222 15702 9274
rect 15702 9222 15732 9274
rect 15756 9222 15766 9274
rect 15766 9222 15812 9274
rect 15516 9220 15572 9222
rect 15596 9220 15652 9222
rect 15676 9220 15732 9222
rect 15756 9220 15812 9222
rect 15516 8186 15572 8188
rect 15596 8186 15652 8188
rect 15676 8186 15732 8188
rect 15756 8186 15812 8188
rect 15516 8134 15562 8186
rect 15562 8134 15572 8186
rect 15596 8134 15626 8186
rect 15626 8134 15638 8186
rect 15638 8134 15652 8186
rect 15676 8134 15690 8186
rect 15690 8134 15702 8186
rect 15702 8134 15732 8186
rect 15756 8134 15766 8186
rect 15766 8134 15812 8186
rect 15516 8132 15572 8134
rect 15596 8132 15652 8134
rect 15676 8132 15732 8134
rect 15756 8132 15812 8134
rect 17066 8730 17122 8732
rect 17146 8730 17202 8732
rect 17226 8730 17282 8732
rect 17306 8730 17362 8732
rect 17066 8678 17112 8730
rect 17112 8678 17122 8730
rect 17146 8678 17176 8730
rect 17176 8678 17188 8730
rect 17188 8678 17202 8730
rect 17226 8678 17240 8730
rect 17240 8678 17252 8730
rect 17252 8678 17282 8730
rect 17306 8678 17316 8730
rect 17316 8678 17362 8730
rect 17066 8676 17122 8678
rect 17146 8676 17202 8678
rect 17226 8676 17282 8678
rect 17306 8676 17362 8678
rect 15516 7098 15572 7100
rect 15596 7098 15652 7100
rect 15676 7098 15732 7100
rect 15756 7098 15812 7100
rect 15516 7046 15562 7098
rect 15562 7046 15572 7098
rect 15596 7046 15626 7098
rect 15626 7046 15638 7098
rect 15638 7046 15652 7098
rect 15676 7046 15690 7098
rect 15690 7046 15702 7098
rect 15702 7046 15732 7098
rect 15756 7046 15766 7098
rect 15766 7046 15812 7098
rect 15516 7044 15572 7046
rect 15596 7044 15652 7046
rect 15676 7044 15732 7046
rect 15756 7044 15812 7046
rect 17066 7642 17122 7644
rect 17146 7642 17202 7644
rect 17226 7642 17282 7644
rect 17306 7642 17362 7644
rect 17066 7590 17112 7642
rect 17112 7590 17122 7642
rect 17146 7590 17176 7642
rect 17176 7590 17188 7642
rect 17188 7590 17202 7642
rect 17226 7590 17240 7642
rect 17240 7590 17252 7642
rect 17252 7590 17282 7642
rect 17306 7590 17316 7642
rect 17316 7590 17362 7642
rect 17066 7588 17122 7590
rect 17146 7588 17202 7590
rect 17226 7588 17282 7590
rect 17306 7588 17362 7590
rect 15516 6010 15572 6012
rect 15596 6010 15652 6012
rect 15676 6010 15732 6012
rect 15756 6010 15812 6012
rect 15516 5958 15562 6010
rect 15562 5958 15572 6010
rect 15596 5958 15626 6010
rect 15626 5958 15638 6010
rect 15638 5958 15652 6010
rect 15676 5958 15690 6010
rect 15690 5958 15702 6010
rect 15702 5958 15732 6010
rect 15756 5958 15766 6010
rect 15766 5958 15812 6010
rect 15516 5956 15572 5958
rect 15596 5956 15652 5958
rect 15676 5956 15732 5958
rect 15756 5956 15812 5958
rect 17066 6554 17122 6556
rect 17146 6554 17202 6556
rect 17226 6554 17282 6556
rect 17306 6554 17362 6556
rect 17066 6502 17112 6554
rect 17112 6502 17122 6554
rect 17146 6502 17176 6554
rect 17176 6502 17188 6554
rect 17188 6502 17202 6554
rect 17226 6502 17240 6554
rect 17240 6502 17252 6554
rect 17252 6502 17282 6554
rect 17306 6502 17316 6554
rect 17316 6502 17362 6554
rect 17066 6500 17122 6502
rect 17146 6500 17202 6502
rect 17226 6500 17282 6502
rect 17306 6500 17362 6502
rect 18786 11192 18842 11248
rect 18602 9696 18658 9752
rect 18602 8200 18658 8256
rect 18510 6740 18512 6760
rect 18512 6740 18564 6760
rect 18564 6740 18566 6760
rect 18510 6704 18566 6740
rect 17066 5466 17122 5468
rect 17146 5466 17202 5468
rect 17226 5466 17282 5468
rect 17306 5466 17362 5468
rect 17066 5414 17112 5466
rect 17112 5414 17122 5466
rect 17146 5414 17176 5466
rect 17176 5414 17188 5466
rect 17188 5414 17202 5466
rect 17226 5414 17240 5466
rect 17240 5414 17252 5466
rect 17252 5414 17282 5466
rect 17306 5414 17316 5466
rect 17316 5414 17362 5466
rect 17066 5412 17122 5414
rect 17146 5412 17202 5414
rect 17226 5412 17282 5414
rect 17306 5412 17362 5414
rect 15516 4922 15572 4924
rect 15596 4922 15652 4924
rect 15676 4922 15732 4924
rect 15756 4922 15812 4924
rect 15516 4870 15562 4922
rect 15562 4870 15572 4922
rect 15596 4870 15626 4922
rect 15626 4870 15638 4922
rect 15638 4870 15652 4922
rect 15676 4870 15690 4922
rect 15690 4870 15702 4922
rect 15702 4870 15732 4922
rect 15756 4870 15766 4922
rect 15766 4870 15812 4922
rect 15516 4868 15572 4870
rect 15596 4868 15652 4870
rect 15676 4868 15732 4870
rect 15756 4868 15812 4870
rect 13966 3290 14022 3292
rect 14046 3290 14102 3292
rect 14126 3290 14182 3292
rect 14206 3290 14262 3292
rect 13966 3238 14012 3290
rect 14012 3238 14022 3290
rect 14046 3238 14076 3290
rect 14076 3238 14088 3290
rect 14088 3238 14102 3290
rect 14126 3238 14140 3290
rect 14140 3238 14152 3290
rect 14152 3238 14182 3290
rect 14206 3238 14216 3290
rect 14216 3238 14262 3290
rect 13966 3236 14022 3238
rect 14046 3236 14102 3238
rect 14126 3236 14182 3238
rect 14206 3236 14262 3238
rect 15516 3834 15572 3836
rect 15596 3834 15652 3836
rect 15676 3834 15732 3836
rect 15756 3834 15812 3836
rect 15516 3782 15562 3834
rect 15562 3782 15572 3834
rect 15596 3782 15626 3834
rect 15626 3782 15638 3834
rect 15638 3782 15652 3834
rect 15676 3782 15690 3834
rect 15690 3782 15702 3834
rect 15702 3782 15732 3834
rect 15756 3782 15766 3834
rect 15766 3782 15812 3834
rect 15516 3780 15572 3782
rect 15596 3780 15652 3782
rect 15676 3780 15732 3782
rect 15756 3780 15812 3782
rect 15516 2746 15572 2748
rect 15596 2746 15652 2748
rect 15676 2746 15732 2748
rect 15756 2746 15812 2748
rect 15516 2694 15562 2746
rect 15562 2694 15572 2746
rect 15596 2694 15626 2746
rect 15626 2694 15638 2746
rect 15638 2694 15652 2746
rect 15676 2694 15690 2746
rect 15690 2694 15702 2746
rect 15702 2694 15732 2746
rect 15756 2694 15766 2746
rect 15766 2694 15812 2746
rect 15516 2692 15572 2694
rect 15596 2692 15652 2694
rect 15676 2692 15732 2694
rect 15756 2692 15812 2694
rect 17066 4378 17122 4380
rect 17146 4378 17202 4380
rect 17226 4378 17282 4380
rect 17306 4378 17362 4380
rect 17066 4326 17112 4378
rect 17112 4326 17122 4378
rect 17146 4326 17176 4378
rect 17176 4326 17188 4378
rect 17188 4326 17202 4378
rect 17226 4326 17240 4378
rect 17240 4326 17252 4378
rect 17252 4326 17282 4378
rect 17306 4326 17316 4378
rect 17316 4326 17362 4378
rect 17066 4324 17122 4326
rect 17146 4324 17202 4326
rect 17226 4324 17282 4326
rect 17306 4324 17362 4326
rect 13966 2202 14022 2204
rect 14046 2202 14102 2204
rect 14126 2202 14182 2204
rect 14206 2202 14262 2204
rect 13966 2150 14012 2202
rect 14012 2150 14022 2202
rect 14046 2150 14076 2202
rect 14076 2150 14088 2202
rect 14088 2150 14102 2202
rect 14126 2150 14140 2202
rect 14140 2150 14152 2202
rect 14152 2150 14182 2202
rect 14206 2150 14216 2202
rect 14216 2150 14262 2202
rect 13966 2148 14022 2150
rect 14046 2148 14102 2150
rect 14126 2148 14182 2150
rect 14206 2148 14262 2150
rect 10866 1114 10922 1116
rect 10946 1114 11002 1116
rect 11026 1114 11082 1116
rect 11106 1114 11162 1116
rect 10866 1062 10912 1114
rect 10912 1062 10922 1114
rect 10946 1062 10976 1114
rect 10976 1062 10988 1114
rect 10988 1062 11002 1114
rect 11026 1062 11040 1114
rect 11040 1062 11052 1114
rect 11052 1062 11082 1114
rect 11106 1062 11116 1114
rect 11116 1062 11162 1114
rect 10866 1060 10922 1062
rect 10946 1060 11002 1062
rect 11026 1060 11082 1062
rect 11106 1060 11162 1062
rect 12416 1658 12472 1660
rect 12496 1658 12552 1660
rect 12576 1658 12632 1660
rect 12656 1658 12712 1660
rect 12416 1606 12462 1658
rect 12462 1606 12472 1658
rect 12496 1606 12526 1658
rect 12526 1606 12538 1658
rect 12538 1606 12552 1658
rect 12576 1606 12590 1658
rect 12590 1606 12602 1658
rect 12602 1606 12632 1658
rect 12656 1606 12666 1658
rect 12666 1606 12712 1658
rect 12416 1604 12472 1606
rect 12496 1604 12552 1606
rect 12576 1604 12632 1606
rect 12656 1604 12712 1606
rect 9034 312 9090 368
rect 9316 570 9372 572
rect 9396 570 9452 572
rect 9476 570 9532 572
rect 9556 570 9612 572
rect 9316 518 9362 570
rect 9362 518 9372 570
rect 9396 518 9426 570
rect 9426 518 9438 570
rect 9438 518 9452 570
rect 9476 518 9490 570
rect 9490 518 9502 570
rect 9502 518 9532 570
rect 9556 518 9566 570
rect 9566 518 9612 570
rect 9316 516 9372 518
rect 9396 516 9452 518
rect 9476 516 9532 518
rect 9556 516 9612 518
rect 13358 856 13414 912
rect 11702 312 11758 368
rect 12416 570 12472 572
rect 12496 570 12552 572
rect 12576 570 12632 572
rect 12656 570 12712 572
rect 12416 518 12462 570
rect 12462 518 12472 570
rect 12496 518 12526 570
rect 12526 518 12538 570
rect 12538 518 12552 570
rect 12576 518 12590 570
rect 12590 518 12602 570
rect 12602 518 12632 570
rect 12656 518 12666 570
rect 12666 518 12712 570
rect 12416 516 12472 518
rect 12496 516 12552 518
rect 12576 516 12632 518
rect 12656 516 12712 518
rect 12254 348 12256 368
rect 12256 348 12308 368
rect 12308 348 12310 368
rect 12254 312 12310 348
rect 13726 876 13782 912
rect 13726 856 13728 876
rect 13728 856 13780 876
rect 13780 856 13782 876
rect 13966 1114 14022 1116
rect 14046 1114 14102 1116
rect 14126 1114 14182 1116
rect 14206 1114 14262 1116
rect 13966 1062 14012 1114
rect 14012 1062 14022 1114
rect 14046 1062 14076 1114
rect 14076 1062 14088 1114
rect 14088 1062 14102 1114
rect 14126 1062 14140 1114
rect 14140 1062 14152 1114
rect 14152 1062 14182 1114
rect 14206 1062 14216 1114
rect 14216 1062 14262 1114
rect 13966 1060 14022 1062
rect 14046 1060 14102 1062
rect 14126 1060 14182 1062
rect 14206 1060 14262 1062
rect 13818 720 13874 776
rect 14278 756 14280 776
rect 14280 756 14332 776
rect 14332 756 14334 776
rect 14278 720 14334 756
rect 17066 3290 17122 3292
rect 17146 3290 17202 3292
rect 17226 3290 17282 3292
rect 17306 3290 17362 3292
rect 17066 3238 17112 3290
rect 17112 3238 17122 3290
rect 17146 3238 17176 3290
rect 17176 3238 17188 3290
rect 17188 3238 17202 3290
rect 17226 3238 17240 3290
rect 17240 3238 17252 3290
rect 17252 3238 17282 3290
rect 17306 3238 17316 3290
rect 17316 3238 17362 3290
rect 17066 3236 17122 3238
rect 17146 3236 17202 3238
rect 17226 3236 17282 3238
rect 17306 3236 17362 3238
rect 17066 2202 17122 2204
rect 17146 2202 17202 2204
rect 17226 2202 17282 2204
rect 17306 2202 17362 2204
rect 17066 2150 17112 2202
rect 17112 2150 17122 2202
rect 17146 2150 17176 2202
rect 17176 2150 17188 2202
rect 17188 2150 17202 2202
rect 17226 2150 17240 2202
rect 17240 2150 17252 2202
rect 17252 2150 17282 2202
rect 17306 2150 17316 2202
rect 17316 2150 17362 2202
rect 17066 2148 17122 2150
rect 17146 2148 17202 2150
rect 17226 2148 17282 2150
rect 17306 2148 17362 2150
rect 18510 5228 18566 5264
rect 18510 5208 18512 5228
rect 18512 5208 18564 5228
rect 18564 5208 18566 5228
rect 18510 3712 18566 3768
rect 18510 2216 18566 2272
rect 15516 1658 15572 1660
rect 15596 1658 15652 1660
rect 15676 1658 15732 1660
rect 15756 1658 15812 1660
rect 15516 1606 15562 1658
rect 15562 1606 15572 1658
rect 15596 1606 15626 1658
rect 15626 1606 15638 1658
rect 15638 1606 15652 1658
rect 15676 1606 15690 1658
rect 15690 1606 15702 1658
rect 15702 1606 15732 1658
rect 15756 1606 15766 1658
rect 15766 1606 15812 1658
rect 15516 1604 15572 1606
rect 15596 1604 15652 1606
rect 15676 1604 15732 1606
rect 15756 1604 15812 1606
rect 15516 570 15572 572
rect 15596 570 15652 572
rect 15676 570 15732 572
rect 15756 570 15812 572
rect 15516 518 15562 570
rect 15562 518 15572 570
rect 15596 518 15626 570
rect 15626 518 15638 570
rect 15638 518 15652 570
rect 15676 518 15690 570
rect 15690 518 15702 570
rect 15702 518 15732 570
rect 15756 518 15766 570
rect 15766 518 15812 570
rect 15516 516 15572 518
rect 15596 516 15652 518
rect 15676 516 15732 518
rect 15756 516 15812 518
rect 15842 312 15898 368
rect 17066 1114 17122 1116
rect 17146 1114 17202 1116
rect 17226 1114 17282 1116
rect 17306 1114 17362 1116
rect 17066 1062 17112 1114
rect 17112 1062 17122 1114
rect 17146 1062 17176 1114
rect 17176 1062 17188 1114
rect 17188 1062 17202 1114
rect 17226 1062 17240 1114
rect 17240 1062 17252 1114
rect 17252 1062 17282 1114
rect 17306 1062 17316 1114
rect 17316 1062 17362 1114
rect 17066 1060 17122 1062
rect 17146 1060 17202 1062
rect 17226 1060 17282 1062
rect 17306 1060 17362 1062
rect 17866 856 17922 912
rect 17590 756 17592 776
rect 17592 756 17644 776
rect 17644 756 17646 776
rect 17590 720 17646 756
rect 18510 720 18566 776
rect 4666 26 4722 28
rect 4746 26 4802 28
rect 4826 26 4882 28
rect 4906 26 4962 28
rect 4666 -26 4712 26
rect 4712 -26 4722 26
rect 4746 -26 4776 26
rect 4776 -26 4788 26
rect 4788 -26 4802 26
rect 4826 -26 4840 26
rect 4840 -26 4852 26
rect 4852 -26 4882 26
rect 4906 -26 4916 26
rect 4916 -26 4962 26
rect 4666 -28 4722 -26
rect 4746 -28 4802 -26
rect 4826 -28 4882 -26
rect 4906 -28 4962 -26
rect 7766 26 7822 28
rect 7846 26 7902 28
rect 7926 26 7982 28
rect 8006 26 8062 28
rect 7766 -26 7812 26
rect 7812 -26 7822 26
rect 7846 -26 7876 26
rect 7876 -26 7888 26
rect 7888 -26 7902 26
rect 7926 -26 7940 26
rect 7940 -26 7952 26
rect 7952 -26 7982 26
rect 8006 -26 8016 26
rect 8016 -26 8062 26
rect 7766 -28 7822 -26
rect 7846 -28 7902 -26
rect 7926 -28 7982 -26
rect 8006 -28 8062 -26
rect 10866 26 10922 28
rect 10946 26 11002 28
rect 11026 26 11082 28
rect 11106 26 11162 28
rect 10866 -26 10912 26
rect 10912 -26 10922 26
rect 10946 -26 10976 26
rect 10976 -26 10988 26
rect 10988 -26 11002 26
rect 11026 -26 11040 26
rect 11040 -26 11052 26
rect 11052 -26 11082 26
rect 11106 -26 11116 26
rect 11116 -26 11162 26
rect 10866 -28 10922 -26
rect 10946 -28 11002 -26
rect 11026 -28 11082 -26
rect 11106 -28 11162 -26
rect 13966 26 14022 28
rect 14046 26 14102 28
rect 14126 26 14182 28
rect 14206 26 14262 28
rect 13966 -26 14012 26
rect 14012 -26 14022 26
rect 14046 -26 14076 26
rect 14076 -26 14088 26
rect 14088 -26 14102 26
rect 14126 -26 14140 26
rect 14140 -26 14152 26
rect 14152 -26 14182 26
rect 14206 -26 14216 26
rect 14216 -26 14262 26
rect 13966 -28 14022 -26
rect 14046 -28 14102 -26
rect 14126 -28 14182 -26
rect 14206 -28 14262 -26
rect 17066 26 17122 28
rect 17146 26 17202 28
rect 17226 26 17282 28
rect 17306 26 17362 28
rect 17066 -26 17112 26
rect 17112 -26 17122 26
rect 17146 -26 17176 26
rect 17176 -26 17188 26
rect 17188 -26 17202 26
rect 17226 -26 17240 26
rect 17240 -26 17252 26
rect 17252 -26 17282 26
rect 17306 -26 17316 26
rect 17316 -26 17362 26
rect 17066 -28 17122 -26
rect 17146 -28 17202 -26
rect 17226 -28 17282 -26
rect 17306 -28 17362 -26
<< metal3 >>
rect 18781 11250 18847 11253
rect 19200 11250 20000 11280
rect 18781 11248 20000 11250
rect 18781 11192 18786 11248
rect 18842 11192 20000 11248
rect 18781 11190 20000 11192
rect 18781 11187 18847 11190
rect 19200 11160 20000 11190
rect 4654 10912 4974 10913
rect 4654 10848 4662 10912
rect 4726 10848 4742 10912
rect 4806 10848 4822 10912
rect 4886 10848 4902 10912
rect 4966 10848 4974 10912
rect 4654 10847 4974 10848
rect 7754 10912 8074 10913
rect 7754 10848 7762 10912
rect 7826 10848 7842 10912
rect 7906 10848 7922 10912
rect 7986 10848 8002 10912
rect 8066 10848 8074 10912
rect 7754 10847 8074 10848
rect 10854 10912 11174 10913
rect 10854 10848 10862 10912
rect 10926 10848 10942 10912
rect 11006 10848 11022 10912
rect 11086 10848 11102 10912
rect 11166 10848 11174 10912
rect 10854 10847 11174 10848
rect 13954 10912 14274 10913
rect 13954 10848 13962 10912
rect 14026 10848 14042 10912
rect 14106 10848 14122 10912
rect 14186 10848 14202 10912
rect 14266 10848 14274 10912
rect 13954 10847 14274 10848
rect 17054 10912 17374 10913
rect 17054 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17222 10912
rect 17286 10848 17302 10912
rect 17366 10848 17374 10912
rect 17054 10847 17374 10848
rect 3104 10368 3424 10369
rect 3104 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3272 10368
rect 3336 10304 3352 10368
rect 3416 10304 3424 10368
rect 3104 10303 3424 10304
rect 6204 10368 6524 10369
rect 6204 10304 6212 10368
rect 6276 10304 6292 10368
rect 6356 10304 6372 10368
rect 6436 10304 6452 10368
rect 6516 10304 6524 10368
rect 6204 10303 6524 10304
rect 9304 10368 9624 10369
rect 9304 10304 9312 10368
rect 9376 10304 9392 10368
rect 9456 10304 9472 10368
rect 9536 10304 9552 10368
rect 9616 10304 9624 10368
rect 9304 10303 9624 10304
rect 12404 10368 12724 10369
rect 12404 10304 12412 10368
rect 12476 10304 12492 10368
rect 12556 10304 12572 10368
rect 12636 10304 12652 10368
rect 12716 10304 12724 10368
rect 12404 10303 12724 10304
rect 15504 10368 15824 10369
rect 15504 10304 15512 10368
rect 15576 10304 15592 10368
rect 15656 10304 15672 10368
rect 15736 10304 15752 10368
rect 15816 10304 15824 10368
rect 15504 10303 15824 10304
rect 4654 9824 4974 9825
rect 4654 9760 4662 9824
rect 4726 9760 4742 9824
rect 4806 9760 4822 9824
rect 4886 9760 4902 9824
rect 4966 9760 4974 9824
rect 4654 9759 4974 9760
rect 7754 9824 8074 9825
rect 7754 9760 7762 9824
rect 7826 9760 7842 9824
rect 7906 9760 7922 9824
rect 7986 9760 8002 9824
rect 8066 9760 8074 9824
rect 7754 9759 8074 9760
rect 10854 9824 11174 9825
rect 10854 9760 10862 9824
rect 10926 9760 10942 9824
rect 11006 9760 11022 9824
rect 11086 9760 11102 9824
rect 11166 9760 11174 9824
rect 10854 9759 11174 9760
rect 13954 9824 14274 9825
rect 13954 9760 13962 9824
rect 14026 9760 14042 9824
rect 14106 9760 14122 9824
rect 14186 9760 14202 9824
rect 14266 9760 14274 9824
rect 13954 9759 14274 9760
rect 17054 9824 17374 9825
rect 17054 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17222 9824
rect 17286 9760 17302 9824
rect 17366 9760 17374 9824
rect 17054 9759 17374 9760
rect 18597 9754 18663 9757
rect 19200 9754 20000 9784
rect 18597 9752 20000 9754
rect 18597 9696 18602 9752
rect 18658 9696 20000 9752
rect 18597 9694 20000 9696
rect 18597 9691 18663 9694
rect 19200 9664 20000 9694
rect 2497 9618 2563 9621
rect 5533 9618 5599 9621
rect 2497 9616 5599 9618
rect 2497 9560 2502 9616
rect 2558 9560 5538 9616
rect 5594 9560 5599 9616
rect 2497 9558 5599 9560
rect 2497 9555 2563 9558
rect 5533 9555 5599 9558
rect 3141 9482 3207 9485
rect 5993 9482 6059 9485
rect 3141 9480 6059 9482
rect 3141 9424 3146 9480
rect 3202 9424 5998 9480
rect 6054 9424 6059 9480
rect 3141 9422 6059 9424
rect 3141 9419 3207 9422
rect 5993 9419 6059 9422
rect 3104 9280 3424 9281
rect 3104 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3272 9280
rect 3336 9216 3352 9280
rect 3416 9216 3424 9280
rect 3104 9215 3424 9216
rect 6204 9280 6524 9281
rect 6204 9216 6212 9280
rect 6276 9216 6292 9280
rect 6356 9216 6372 9280
rect 6436 9216 6452 9280
rect 6516 9216 6524 9280
rect 6204 9215 6524 9216
rect 9304 9280 9624 9281
rect 9304 9216 9312 9280
rect 9376 9216 9392 9280
rect 9456 9216 9472 9280
rect 9536 9216 9552 9280
rect 9616 9216 9624 9280
rect 9304 9215 9624 9216
rect 12404 9280 12724 9281
rect 12404 9216 12412 9280
rect 12476 9216 12492 9280
rect 12556 9216 12572 9280
rect 12636 9216 12652 9280
rect 12716 9216 12724 9280
rect 12404 9215 12724 9216
rect 15504 9280 15824 9281
rect 15504 9216 15512 9280
rect 15576 9216 15592 9280
rect 15656 9216 15672 9280
rect 15736 9216 15752 9280
rect 15816 9216 15824 9280
rect 15504 9215 15824 9216
rect 4654 8736 4974 8737
rect 4654 8672 4662 8736
rect 4726 8672 4742 8736
rect 4806 8672 4822 8736
rect 4886 8672 4902 8736
rect 4966 8672 4974 8736
rect 4654 8671 4974 8672
rect 7754 8736 8074 8737
rect 7754 8672 7762 8736
rect 7826 8672 7842 8736
rect 7906 8672 7922 8736
rect 7986 8672 8002 8736
rect 8066 8672 8074 8736
rect 7754 8671 8074 8672
rect 10854 8736 11174 8737
rect 10854 8672 10862 8736
rect 10926 8672 10942 8736
rect 11006 8672 11022 8736
rect 11086 8672 11102 8736
rect 11166 8672 11174 8736
rect 10854 8671 11174 8672
rect 13954 8736 14274 8737
rect 13954 8672 13962 8736
rect 14026 8672 14042 8736
rect 14106 8672 14122 8736
rect 14186 8672 14202 8736
rect 14266 8672 14274 8736
rect 13954 8671 14274 8672
rect 17054 8736 17374 8737
rect 17054 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17222 8736
rect 17286 8672 17302 8736
rect 17366 8672 17374 8736
rect 17054 8671 17374 8672
rect 18597 8258 18663 8261
rect 19200 8258 20000 8288
rect 18597 8256 20000 8258
rect 18597 8200 18602 8256
rect 18658 8200 20000 8256
rect 18597 8198 20000 8200
rect 18597 8195 18663 8198
rect 3104 8192 3424 8193
rect 3104 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3272 8192
rect 3336 8128 3352 8192
rect 3416 8128 3424 8192
rect 3104 8127 3424 8128
rect 6204 8192 6524 8193
rect 6204 8128 6212 8192
rect 6276 8128 6292 8192
rect 6356 8128 6372 8192
rect 6436 8128 6452 8192
rect 6516 8128 6524 8192
rect 6204 8127 6524 8128
rect 9304 8192 9624 8193
rect 9304 8128 9312 8192
rect 9376 8128 9392 8192
rect 9456 8128 9472 8192
rect 9536 8128 9552 8192
rect 9616 8128 9624 8192
rect 9304 8127 9624 8128
rect 12404 8192 12724 8193
rect 12404 8128 12412 8192
rect 12476 8128 12492 8192
rect 12556 8128 12572 8192
rect 12636 8128 12652 8192
rect 12716 8128 12724 8192
rect 12404 8127 12724 8128
rect 15504 8192 15824 8193
rect 15504 8128 15512 8192
rect 15576 8128 15592 8192
rect 15656 8128 15672 8192
rect 15736 8128 15752 8192
rect 15816 8128 15824 8192
rect 19200 8168 20000 8198
rect 15504 8127 15824 8128
rect 4654 7648 4974 7649
rect 4654 7584 4662 7648
rect 4726 7584 4742 7648
rect 4806 7584 4822 7648
rect 4886 7584 4902 7648
rect 4966 7584 4974 7648
rect 4654 7583 4974 7584
rect 7754 7648 8074 7649
rect 7754 7584 7762 7648
rect 7826 7584 7842 7648
rect 7906 7584 7922 7648
rect 7986 7584 8002 7648
rect 8066 7584 8074 7648
rect 7754 7583 8074 7584
rect 10854 7648 11174 7649
rect 10854 7584 10862 7648
rect 10926 7584 10942 7648
rect 11006 7584 11022 7648
rect 11086 7584 11102 7648
rect 11166 7584 11174 7648
rect 10854 7583 11174 7584
rect 13954 7648 14274 7649
rect 13954 7584 13962 7648
rect 14026 7584 14042 7648
rect 14106 7584 14122 7648
rect 14186 7584 14202 7648
rect 14266 7584 14274 7648
rect 13954 7583 14274 7584
rect 17054 7648 17374 7649
rect 17054 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17222 7648
rect 17286 7584 17302 7648
rect 17366 7584 17374 7648
rect 17054 7583 17374 7584
rect 13629 7442 13695 7445
rect 13905 7442 13971 7445
rect 13629 7440 13971 7442
rect 13629 7384 13634 7440
rect 13690 7384 13910 7440
rect 13966 7384 13971 7440
rect 13629 7382 13971 7384
rect 13629 7379 13695 7382
rect 13905 7379 13971 7382
rect 3104 7104 3424 7105
rect 3104 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3272 7104
rect 3336 7040 3352 7104
rect 3416 7040 3424 7104
rect 3104 7039 3424 7040
rect 6204 7104 6524 7105
rect 6204 7040 6212 7104
rect 6276 7040 6292 7104
rect 6356 7040 6372 7104
rect 6436 7040 6452 7104
rect 6516 7040 6524 7104
rect 6204 7039 6524 7040
rect 9304 7104 9624 7105
rect 9304 7040 9312 7104
rect 9376 7040 9392 7104
rect 9456 7040 9472 7104
rect 9536 7040 9552 7104
rect 9616 7040 9624 7104
rect 9304 7039 9624 7040
rect 12404 7104 12724 7105
rect 12404 7040 12412 7104
rect 12476 7040 12492 7104
rect 12556 7040 12572 7104
rect 12636 7040 12652 7104
rect 12716 7040 12724 7104
rect 12404 7039 12724 7040
rect 15504 7104 15824 7105
rect 15504 7040 15512 7104
rect 15576 7040 15592 7104
rect 15656 7040 15672 7104
rect 15736 7040 15752 7104
rect 15816 7040 15824 7104
rect 15504 7039 15824 7040
rect 18505 6762 18571 6765
rect 19200 6762 20000 6792
rect 18505 6760 20000 6762
rect 18505 6704 18510 6760
rect 18566 6704 20000 6760
rect 18505 6702 20000 6704
rect 18505 6699 18571 6702
rect 19200 6672 20000 6702
rect 4654 6560 4974 6561
rect 4654 6496 4662 6560
rect 4726 6496 4742 6560
rect 4806 6496 4822 6560
rect 4886 6496 4902 6560
rect 4966 6496 4974 6560
rect 4654 6495 4974 6496
rect 7754 6560 8074 6561
rect 7754 6496 7762 6560
rect 7826 6496 7842 6560
rect 7906 6496 7922 6560
rect 7986 6496 8002 6560
rect 8066 6496 8074 6560
rect 7754 6495 8074 6496
rect 10854 6560 11174 6561
rect 10854 6496 10862 6560
rect 10926 6496 10942 6560
rect 11006 6496 11022 6560
rect 11086 6496 11102 6560
rect 11166 6496 11174 6560
rect 10854 6495 11174 6496
rect 13954 6560 14274 6561
rect 13954 6496 13962 6560
rect 14026 6496 14042 6560
rect 14106 6496 14122 6560
rect 14186 6496 14202 6560
rect 14266 6496 14274 6560
rect 13954 6495 14274 6496
rect 17054 6560 17374 6561
rect 17054 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17222 6560
rect 17286 6496 17302 6560
rect 17366 6496 17374 6560
rect 17054 6495 17374 6496
rect 3417 6354 3483 6357
rect 5165 6354 5231 6357
rect 3417 6352 5231 6354
rect 3417 6296 3422 6352
rect 3478 6296 5170 6352
rect 5226 6296 5231 6352
rect 3417 6294 5231 6296
rect 3417 6291 3483 6294
rect 5165 6291 5231 6294
rect 3104 6016 3424 6017
rect 3104 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3272 6016
rect 3336 5952 3352 6016
rect 3416 5952 3424 6016
rect 3104 5951 3424 5952
rect 6204 6016 6524 6017
rect 6204 5952 6212 6016
rect 6276 5952 6292 6016
rect 6356 5952 6372 6016
rect 6436 5952 6452 6016
rect 6516 5952 6524 6016
rect 6204 5951 6524 5952
rect 9304 6016 9624 6017
rect 9304 5952 9312 6016
rect 9376 5952 9392 6016
rect 9456 5952 9472 6016
rect 9536 5952 9552 6016
rect 9616 5952 9624 6016
rect 9304 5951 9624 5952
rect 12404 6016 12724 6017
rect 12404 5952 12412 6016
rect 12476 5952 12492 6016
rect 12556 5952 12572 6016
rect 12636 5952 12652 6016
rect 12716 5952 12724 6016
rect 12404 5951 12724 5952
rect 15504 6016 15824 6017
rect 15504 5952 15512 6016
rect 15576 5952 15592 6016
rect 15656 5952 15672 6016
rect 15736 5952 15752 6016
rect 15816 5952 15824 6016
rect 15504 5951 15824 5952
rect 4654 5472 4974 5473
rect 4654 5408 4662 5472
rect 4726 5408 4742 5472
rect 4806 5408 4822 5472
rect 4886 5408 4902 5472
rect 4966 5408 4974 5472
rect 4654 5407 4974 5408
rect 7754 5472 8074 5473
rect 7754 5408 7762 5472
rect 7826 5408 7842 5472
rect 7906 5408 7922 5472
rect 7986 5408 8002 5472
rect 8066 5408 8074 5472
rect 7754 5407 8074 5408
rect 10854 5472 11174 5473
rect 10854 5408 10862 5472
rect 10926 5408 10942 5472
rect 11006 5408 11022 5472
rect 11086 5408 11102 5472
rect 11166 5408 11174 5472
rect 10854 5407 11174 5408
rect 13954 5472 14274 5473
rect 13954 5408 13962 5472
rect 14026 5408 14042 5472
rect 14106 5408 14122 5472
rect 14186 5408 14202 5472
rect 14266 5408 14274 5472
rect 13954 5407 14274 5408
rect 17054 5472 17374 5473
rect 17054 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17222 5472
rect 17286 5408 17302 5472
rect 17366 5408 17374 5472
rect 17054 5407 17374 5408
rect 18505 5266 18571 5269
rect 19200 5266 20000 5296
rect 18505 5264 20000 5266
rect 18505 5208 18510 5264
rect 18566 5208 20000 5264
rect 18505 5206 20000 5208
rect 18505 5203 18571 5206
rect 19200 5176 20000 5206
rect 3104 4928 3424 4929
rect 3104 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3272 4928
rect 3336 4864 3352 4928
rect 3416 4864 3424 4928
rect 3104 4863 3424 4864
rect 6204 4928 6524 4929
rect 6204 4864 6212 4928
rect 6276 4864 6292 4928
rect 6356 4864 6372 4928
rect 6436 4864 6452 4928
rect 6516 4864 6524 4928
rect 6204 4863 6524 4864
rect 9304 4928 9624 4929
rect 9304 4864 9312 4928
rect 9376 4864 9392 4928
rect 9456 4864 9472 4928
rect 9536 4864 9552 4928
rect 9616 4864 9624 4928
rect 9304 4863 9624 4864
rect 12404 4928 12724 4929
rect 12404 4864 12412 4928
rect 12476 4864 12492 4928
rect 12556 4864 12572 4928
rect 12636 4864 12652 4928
rect 12716 4864 12724 4928
rect 12404 4863 12724 4864
rect 15504 4928 15824 4929
rect 15504 4864 15512 4928
rect 15576 4864 15592 4928
rect 15656 4864 15672 4928
rect 15736 4864 15752 4928
rect 15816 4864 15824 4928
rect 15504 4863 15824 4864
rect 4654 4384 4974 4385
rect 4654 4320 4662 4384
rect 4726 4320 4742 4384
rect 4806 4320 4822 4384
rect 4886 4320 4902 4384
rect 4966 4320 4974 4384
rect 4654 4319 4974 4320
rect 7754 4384 8074 4385
rect 7754 4320 7762 4384
rect 7826 4320 7842 4384
rect 7906 4320 7922 4384
rect 7986 4320 8002 4384
rect 8066 4320 8074 4384
rect 7754 4319 8074 4320
rect 10854 4384 11174 4385
rect 10854 4320 10862 4384
rect 10926 4320 10942 4384
rect 11006 4320 11022 4384
rect 11086 4320 11102 4384
rect 11166 4320 11174 4384
rect 10854 4319 11174 4320
rect 13954 4384 14274 4385
rect 13954 4320 13962 4384
rect 14026 4320 14042 4384
rect 14106 4320 14122 4384
rect 14186 4320 14202 4384
rect 14266 4320 14274 4384
rect 13954 4319 14274 4320
rect 17054 4384 17374 4385
rect 17054 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17222 4384
rect 17286 4320 17302 4384
rect 17366 4320 17374 4384
rect 17054 4319 17374 4320
rect 3104 3840 3424 3841
rect 3104 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3272 3840
rect 3336 3776 3352 3840
rect 3416 3776 3424 3840
rect 3104 3775 3424 3776
rect 6204 3840 6524 3841
rect 6204 3776 6212 3840
rect 6276 3776 6292 3840
rect 6356 3776 6372 3840
rect 6436 3776 6452 3840
rect 6516 3776 6524 3840
rect 6204 3775 6524 3776
rect 9304 3840 9624 3841
rect 9304 3776 9312 3840
rect 9376 3776 9392 3840
rect 9456 3776 9472 3840
rect 9536 3776 9552 3840
rect 9616 3776 9624 3840
rect 9304 3775 9624 3776
rect 12404 3840 12724 3841
rect 12404 3776 12412 3840
rect 12476 3776 12492 3840
rect 12556 3776 12572 3840
rect 12636 3776 12652 3840
rect 12716 3776 12724 3840
rect 12404 3775 12724 3776
rect 15504 3840 15824 3841
rect 15504 3776 15512 3840
rect 15576 3776 15592 3840
rect 15656 3776 15672 3840
rect 15736 3776 15752 3840
rect 15816 3776 15824 3840
rect 15504 3775 15824 3776
rect 18505 3770 18571 3773
rect 19200 3770 20000 3800
rect 18505 3768 20000 3770
rect 18505 3712 18510 3768
rect 18566 3712 20000 3768
rect 18505 3710 20000 3712
rect 18505 3707 18571 3710
rect 19200 3680 20000 3710
rect 8661 3634 8727 3637
rect 12341 3634 12407 3637
rect 8661 3632 12407 3634
rect 8661 3576 8666 3632
rect 8722 3576 12346 3632
rect 12402 3576 12407 3632
rect 8661 3574 12407 3576
rect 8661 3571 8727 3574
rect 12341 3571 12407 3574
rect 9029 3498 9095 3501
rect 9765 3498 9831 3501
rect 9029 3496 9831 3498
rect 9029 3440 9034 3496
rect 9090 3440 9770 3496
rect 9826 3440 9831 3496
rect 9029 3438 9831 3440
rect 9029 3435 9095 3438
rect 9765 3435 9831 3438
rect 11513 3498 11579 3501
rect 13445 3498 13511 3501
rect 11513 3496 13511 3498
rect 11513 3440 11518 3496
rect 11574 3440 13450 3496
rect 13506 3440 13511 3496
rect 11513 3438 13511 3440
rect 11513 3435 11579 3438
rect 13445 3435 13511 3438
rect 4654 3296 4974 3297
rect 4654 3232 4662 3296
rect 4726 3232 4742 3296
rect 4806 3232 4822 3296
rect 4886 3232 4902 3296
rect 4966 3232 4974 3296
rect 4654 3231 4974 3232
rect 7754 3296 8074 3297
rect 7754 3232 7762 3296
rect 7826 3232 7842 3296
rect 7906 3232 7922 3296
rect 7986 3232 8002 3296
rect 8066 3232 8074 3296
rect 7754 3231 8074 3232
rect 10854 3296 11174 3297
rect 10854 3232 10862 3296
rect 10926 3232 10942 3296
rect 11006 3232 11022 3296
rect 11086 3232 11102 3296
rect 11166 3232 11174 3296
rect 10854 3231 11174 3232
rect 13954 3296 14274 3297
rect 13954 3232 13962 3296
rect 14026 3232 14042 3296
rect 14106 3232 14122 3296
rect 14186 3232 14202 3296
rect 14266 3232 14274 3296
rect 13954 3231 14274 3232
rect 17054 3296 17374 3297
rect 17054 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17222 3296
rect 17286 3232 17302 3296
rect 17366 3232 17374 3296
rect 17054 3231 17374 3232
rect 8937 3090 9003 3093
rect 10869 3090 10935 3093
rect 11145 3090 11211 3093
rect 8937 3088 11211 3090
rect 8937 3032 8942 3088
rect 8998 3032 10874 3088
rect 10930 3032 11150 3088
rect 11206 3032 11211 3088
rect 8937 3030 11211 3032
rect 8937 3027 9003 3030
rect 10869 3027 10935 3030
rect 11145 3027 11211 3030
rect 3104 2752 3424 2753
rect 3104 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3272 2752
rect 3336 2688 3352 2752
rect 3416 2688 3424 2752
rect 3104 2687 3424 2688
rect 6204 2752 6524 2753
rect 6204 2688 6212 2752
rect 6276 2688 6292 2752
rect 6356 2688 6372 2752
rect 6436 2688 6452 2752
rect 6516 2688 6524 2752
rect 6204 2687 6524 2688
rect 9304 2752 9624 2753
rect 9304 2688 9312 2752
rect 9376 2688 9392 2752
rect 9456 2688 9472 2752
rect 9536 2688 9552 2752
rect 9616 2688 9624 2752
rect 9304 2687 9624 2688
rect 12404 2752 12724 2753
rect 12404 2688 12412 2752
rect 12476 2688 12492 2752
rect 12556 2688 12572 2752
rect 12636 2688 12652 2752
rect 12716 2688 12724 2752
rect 12404 2687 12724 2688
rect 15504 2752 15824 2753
rect 15504 2688 15512 2752
rect 15576 2688 15592 2752
rect 15656 2688 15672 2752
rect 15736 2688 15752 2752
rect 15816 2688 15824 2752
rect 15504 2687 15824 2688
rect 18505 2274 18571 2277
rect 19200 2274 20000 2304
rect 18505 2272 20000 2274
rect 18505 2216 18510 2272
rect 18566 2216 20000 2272
rect 18505 2214 20000 2216
rect 18505 2211 18571 2214
rect 4654 2208 4974 2209
rect 4654 2144 4662 2208
rect 4726 2144 4742 2208
rect 4806 2144 4822 2208
rect 4886 2144 4902 2208
rect 4966 2144 4974 2208
rect 4654 2143 4974 2144
rect 7754 2208 8074 2209
rect 7754 2144 7762 2208
rect 7826 2144 7842 2208
rect 7906 2144 7922 2208
rect 7986 2144 8002 2208
rect 8066 2144 8074 2208
rect 7754 2143 8074 2144
rect 10854 2208 11174 2209
rect 10854 2144 10862 2208
rect 10926 2144 10942 2208
rect 11006 2144 11022 2208
rect 11086 2144 11102 2208
rect 11166 2144 11174 2208
rect 10854 2143 11174 2144
rect 13954 2208 14274 2209
rect 13954 2144 13962 2208
rect 14026 2144 14042 2208
rect 14106 2144 14122 2208
rect 14186 2144 14202 2208
rect 14266 2144 14274 2208
rect 13954 2143 14274 2144
rect 17054 2208 17374 2209
rect 17054 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17222 2208
rect 17286 2144 17302 2208
rect 17366 2144 17374 2208
rect 19200 2184 20000 2214
rect 17054 2143 17374 2144
rect 3104 1664 3424 1665
rect 3104 1600 3112 1664
rect 3176 1600 3192 1664
rect 3256 1600 3272 1664
rect 3336 1600 3352 1664
rect 3416 1600 3424 1664
rect 3104 1599 3424 1600
rect 6204 1664 6524 1665
rect 6204 1600 6212 1664
rect 6276 1600 6292 1664
rect 6356 1600 6372 1664
rect 6436 1600 6452 1664
rect 6516 1600 6524 1664
rect 6204 1599 6524 1600
rect 9304 1664 9624 1665
rect 9304 1600 9312 1664
rect 9376 1600 9392 1664
rect 9456 1600 9472 1664
rect 9536 1600 9552 1664
rect 9616 1600 9624 1664
rect 9304 1599 9624 1600
rect 12404 1664 12724 1665
rect 12404 1600 12412 1664
rect 12476 1600 12492 1664
rect 12556 1600 12572 1664
rect 12636 1600 12652 1664
rect 12716 1600 12724 1664
rect 12404 1599 12724 1600
rect 15504 1664 15824 1665
rect 15504 1600 15512 1664
rect 15576 1600 15592 1664
rect 15656 1600 15672 1664
rect 15736 1600 15752 1664
rect 15816 1600 15824 1664
rect 15504 1599 15824 1600
rect 7005 1322 7071 1325
rect 8753 1322 8819 1325
rect 9213 1322 9279 1325
rect 7005 1320 9279 1322
rect 7005 1264 7010 1320
rect 7066 1264 8758 1320
rect 8814 1264 9218 1320
rect 9274 1264 9279 1320
rect 7005 1262 9279 1264
rect 7005 1259 7071 1262
rect 8753 1259 8819 1262
rect 9213 1259 9279 1262
rect 4654 1120 4974 1121
rect 4654 1056 4662 1120
rect 4726 1056 4742 1120
rect 4806 1056 4822 1120
rect 4886 1056 4902 1120
rect 4966 1056 4974 1120
rect 4654 1055 4974 1056
rect 7754 1120 8074 1121
rect 7754 1056 7762 1120
rect 7826 1056 7842 1120
rect 7906 1056 7922 1120
rect 7986 1056 8002 1120
rect 8066 1056 8074 1120
rect 7754 1055 8074 1056
rect 10854 1120 11174 1121
rect 10854 1056 10862 1120
rect 10926 1056 10942 1120
rect 11006 1056 11022 1120
rect 11086 1056 11102 1120
rect 11166 1056 11174 1120
rect 10854 1055 11174 1056
rect 13954 1120 14274 1121
rect 13954 1056 13962 1120
rect 14026 1056 14042 1120
rect 14106 1056 14122 1120
rect 14186 1056 14202 1120
rect 14266 1056 14274 1120
rect 13954 1055 14274 1056
rect 17054 1120 17374 1121
rect 17054 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17222 1120
rect 17286 1056 17302 1120
rect 17366 1056 17374 1120
rect 17054 1055 17374 1056
rect 4889 914 4955 917
rect 5257 914 5323 917
rect 7741 914 7807 917
rect 4889 912 7807 914
rect 4889 856 4894 912
rect 4950 856 5262 912
rect 5318 856 7746 912
rect 7802 856 7807 912
rect 4889 854 7807 856
rect 4889 851 4955 854
rect 5257 851 5323 854
rect 7741 851 7807 854
rect 10133 914 10199 917
rect 13353 914 13419 917
rect 10133 912 13419 914
rect 10133 856 10138 912
rect 10194 856 13358 912
rect 13414 856 13419 912
rect 10133 854 13419 856
rect 10133 851 10199 854
rect 13353 851 13419 854
rect 13721 914 13787 917
rect 17861 914 17927 917
rect 13721 912 17927 914
rect 13721 856 13726 912
rect 13782 856 17866 912
rect 17922 856 17927 912
rect 13721 854 17927 856
rect 13721 851 13787 854
rect 17861 851 17927 854
rect 9305 778 9371 781
rect 13813 778 13879 781
rect 14273 778 14339 781
rect 17585 778 17651 781
rect 9305 776 17651 778
rect 9305 720 9310 776
rect 9366 720 13818 776
rect 13874 720 14278 776
rect 14334 720 17590 776
rect 17646 720 17651 776
rect 9305 718 17651 720
rect 9305 715 9371 718
rect 13813 715 13879 718
rect 14273 715 14339 718
rect 17585 715 17651 718
rect 18505 778 18571 781
rect 19200 778 20000 808
rect 18505 776 20000 778
rect 18505 720 18510 776
rect 18566 720 20000 776
rect 18505 718 20000 720
rect 18505 715 18571 718
rect 19200 688 20000 718
rect 3104 576 3424 577
rect 3104 512 3112 576
rect 3176 512 3192 576
rect 3256 512 3272 576
rect 3336 512 3352 576
rect 3416 512 3424 576
rect 3104 511 3424 512
rect 6204 576 6524 577
rect 6204 512 6212 576
rect 6276 512 6292 576
rect 6356 512 6372 576
rect 6436 512 6452 576
rect 6516 512 6524 576
rect 6204 511 6524 512
rect 9304 576 9624 577
rect 9304 512 9312 576
rect 9376 512 9392 576
rect 9456 512 9472 576
rect 9536 512 9552 576
rect 9616 512 9624 576
rect 9304 511 9624 512
rect 12404 576 12724 577
rect 12404 512 12412 576
rect 12476 512 12492 576
rect 12556 512 12572 576
rect 12636 512 12652 576
rect 12716 512 12724 576
rect 12404 511 12724 512
rect 15504 576 15824 577
rect 15504 512 15512 576
rect 15576 512 15592 576
rect 15656 512 15672 576
rect 15736 512 15752 576
rect 15816 512 15824 576
rect 15504 511 15824 512
rect 9029 370 9095 373
rect 11697 370 11763 373
rect 9029 368 11763 370
rect 9029 312 9034 368
rect 9090 312 11702 368
rect 11758 312 11763 368
rect 9029 310 11763 312
rect 9029 307 9095 310
rect 11697 307 11763 310
rect 12249 370 12315 373
rect 15837 370 15903 373
rect 12249 368 15903 370
rect 12249 312 12254 368
rect 12310 312 15842 368
rect 15898 312 15903 368
rect 12249 310 15903 312
rect 12249 307 12315 310
rect 15837 307 15903 310
rect 4654 32 4974 33
rect 4654 -32 4662 32
rect 4726 -32 4742 32
rect 4806 -32 4822 32
rect 4886 -32 4902 32
rect 4966 -32 4974 32
rect 4654 -33 4974 -32
rect 7754 32 8074 33
rect 7754 -32 7762 32
rect 7826 -32 7842 32
rect 7906 -32 7922 32
rect 7986 -32 8002 32
rect 8066 -32 8074 32
rect 7754 -33 8074 -32
rect 10854 32 11174 33
rect 10854 -32 10862 32
rect 10926 -32 10942 32
rect 11006 -32 11022 32
rect 11086 -32 11102 32
rect 11166 -32 11174 32
rect 10854 -33 11174 -32
rect 13954 32 14274 33
rect 13954 -32 13962 32
rect 14026 -32 14042 32
rect 14106 -32 14122 32
rect 14186 -32 14202 32
rect 14266 -32 14274 32
rect 13954 -33 14274 -32
rect 17054 32 17374 33
rect 17054 -32 17062 32
rect 17126 -32 17142 32
rect 17206 -32 17222 32
rect 17286 -32 17302 32
rect 17366 -32 17374 32
rect 17054 -33 17374 -32
<< via3 >>
rect 4662 10908 4726 10912
rect 4662 10852 4666 10908
rect 4666 10852 4722 10908
rect 4722 10852 4726 10908
rect 4662 10848 4726 10852
rect 4742 10908 4806 10912
rect 4742 10852 4746 10908
rect 4746 10852 4802 10908
rect 4802 10852 4806 10908
rect 4742 10848 4806 10852
rect 4822 10908 4886 10912
rect 4822 10852 4826 10908
rect 4826 10852 4882 10908
rect 4882 10852 4886 10908
rect 4822 10848 4886 10852
rect 4902 10908 4966 10912
rect 4902 10852 4906 10908
rect 4906 10852 4962 10908
rect 4962 10852 4966 10908
rect 4902 10848 4966 10852
rect 7762 10908 7826 10912
rect 7762 10852 7766 10908
rect 7766 10852 7822 10908
rect 7822 10852 7826 10908
rect 7762 10848 7826 10852
rect 7842 10908 7906 10912
rect 7842 10852 7846 10908
rect 7846 10852 7902 10908
rect 7902 10852 7906 10908
rect 7842 10848 7906 10852
rect 7922 10908 7986 10912
rect 7922 10852 7926 10908
rect 7926 10852 7982 10908
rect 7982 10852 7986 10908
rect 7922 10848 7986 10852
rect 8002 10908 8066 10912
rect 8002 10852 8006 10908
rect 8006 10852 8062 10908
rect 8062 10852 8066 10908
rect 8002 10848 8066 10852
rect 10862 10908 10926 10912
rect 10862 10852 10866 10908
rect 10866 10852 10922 10908
rect 10922 10852 10926 10908
rect 10862 10848 10926 10852
rect 10942 10908 11006 10912
rect 10942 10852 10946 10908
rect 10946 10852 11002 10908
rect 11002 10852 11006 10908
rect 10942 10848 11006 10852
rect 11022 10908 11086 10912
rect 11022 10852 11026 10908
rect 11026 10852 11082 10908
rect 11082 10852 11086 10908
rect 11022 10848 11086 10852
rect 11102 10908 11166 10912
rect 11102 10852 11106 10908
rect 11106 10852 11162 10908
rect 11162 10852 11166 10908
rect 11102 10848 11166 10852
rect 13962 10908 14026 10912
rect 13962 10852 13966 10908
rect 13966 10852 14022 10908
rect 14022 10852 14026 10908
rect 13962 10848 14026 10852
rect 14042 10908 14106 10912
rect 14042 10852 14046 10908
rect 14046 10852 14102 10908
rect 14102 10852 14106 10908
rect 14042 10848 14106 10852
rect 14122 10908 14186 10912
rect 14122 10852 14126 10908
rect 14126 10852 14182 10908
rect 14182 10852 14186 10908
rect 14122 10848 14186 10852
rect 14202 10908 14266 10912
rect 14202 10852 14206 10908
rect 14206 10852 14262 10908
rect 14262 10852 14266 10908
rect 14202 10848 14266 10852
rect 17062 10908 17126 10912
rect 17062 10852 17066 10908
rect 17066 10852 17122 10908
rect 17122 10852 17126 10908
rect 17062 10848 17126 10852
rect 17142 10908 17206 10912
rect 17142 10852 17146 10908
rect 17146 10852 17202 10908
rect 17202 10852 17206 10908
rect 17142 10848 17206 10852
rect 17222 10908 17286 10912
rect 17222 10852 17226 10908
rect 17226 10852 17282 10908
rect 17282 10852 17286 10908
rect 17222 10848 17286 10852
rect 17302 10908 17366 10912
rect 17302 10852 17306 10908
rect 17306 10852 17362 10908
rect 17362 10852 17366 10908
rect 17302 10848 17366 10852
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 3272 10364 3336 10368
rect 3272 10308 3276 10364
rect 3276 10308 3332 10364
rect 3332 10308 3336 10364
rect 3272 10304 3336 10308
rect 3352 10364 3416 10368
rect 3352 10308 3356 10364
rect 3356 10308 3412 10364
rect 3412 10308 3416 10364
rect 3352 10304 3416 10308
rect 6212 10364 6276 10368
rect 6212 10308 6216 10364
rect 6216 10308 6272 10364
rect 6272 10308 6276 10364
rect 6212 10304 6276 10308
rect 6292 10364 6356 10368
rect 6292 10308 6296 10364
rect 6296 10308 6352 10364
rect 6352 10308 6356 10364
rect 6292 10304 6356 10308
rect 6372 10364 6436 10368
rect 6372 10308 6376 10364
rect 6376 10308 6432 10364
rect 6432 10308 6436 10364
rect 6372 10304 6436 10308
rect 6452 10364 6516 10368
rect 6452 10308 6456 10364
rect 6456 10308 6512 10364
rect 6512 10308 6516 10364
rect 6452 10304 6516 10308
rect 9312 10364 9376 10368
rect 9312 10308 9316 10364
rect 9316 10308 9372 10364
rect 9372 10308 9376 10364
rect 9312 10304 9376 10308
rect 9392 10364 9456 10368
rect 9392 10308 9396 10364
rect 9396 10308 9452 10364
rect 9452 10308 9456 10364
rect 9392 10304 9456 10308
rect 9472 10364 9536 10368
rect 9472 10308 9476 10364
rect 9476 10308 9532 10364
rect 9532 10308 9536 10364
rect 9472 10304 9536 10308
rect 9552 10364 9616 10368
rect 9552 10308 9556 10364
rect 9556 10308 9612 10364
rect 9612 10308 9616 10364
rect 9552 10304 9616 10308
rect 12412 10364 12476 10368
rect 12412 10308 12416 10364
rect 12416 10308 12472 10364
rect 12472 10308 12476 10364
rect 12412 10304 12476 10308
rect 12492 10364 12556 10368
rect 12492 10308 12496 10364
rect 12496 10308 12552 10364
rect 12552 10308 12556 10364
rect 12492 10304 12556 10308
rect 12572 10364 12636 10368
rect 12572 10308 12576 10364
rect 12576 10308 12632 10364
rect 12632 10308 12636 10364
rect 12572 10304 12636 10308
rect 12652 10364 12716 10368
rect 12652 10308 12656 10364
rect 12656 10308 12712 10364
rect 12712 10308 12716 10364
rect 12652 10304 12716 10308
rect 15512 10364 15576 10368
rect 15512 10308 15516 10364
rect 15516 10308 15572 10364
rect 15572 10308 15576 10364
rect 15512 10304 15576 10308
rect 15592 10364 15656 10368
rect 15592 10308 15596 10364
rect 15596 10308 15652 10364
rect 15652 10308 15656 10364
rect 15592 10304 15656 10308
rect 15672 10364 15736 10368
rect 15672 10308 15676 10364
rect 15676 10308 15732 10364
rect 15732 10308 15736 10364
rect 15672 10304 15736 10308
rect 15752 10364 15816 10368
rect 15752 10308 15756 10364
rect 15756 10308 15812 10364
rect 15812 10308 15816 10364
rect 15752 10304 15816 10308
rect 4662 9820 4726 9824
rect 4662 9764 4666 9820
rect 4666 9764 4722 9820
rect 4722 9764 4726 9820
rect 4662 9760 4726 9764
rect 4742 9820 4806 9824
rect 4742 9764 4746 9820
rect 4746 9764 4802 9820
rect 4802 9764 4806 9820
rect 4742 9760 4806 9764
rect 4822 9820 4886 9824
rect 4822 9764 4826 9820
rect 4826 9764 4882 9820
rect 4882 9764 4886 9820
rect 4822 9760 4886 9764
rect 4902 9820 4966 9824
rect 4902 9764 4906 9820
rect 4906 9764 4962 9820
rect 4962 9764 4966 9820
rect 4902 9760 4966 9764
rect 7762 9820 7826 9824
rect 7762 9764 7766 9820
rect 7766 9764 7822 9820
rect 7822 9764 7826 9820
rect 7762 9760 7826 9764
rect 7842 9820 7906 9824
rect 7842 9764 7846 9820
rect 7846 9764 7902 9820
rect 7902 9764 7906 9820
rect 7842 9760 7906 9764
rect 7922 9820 7986 9824
rect 7922 9764 7926 9820
rect 7926 9764 7982 9820
rect 7982 9764 7986 9820
rect 7922 9760 7986 9764
rect 8002 9820 8066 9824
rect 8002 9764 8006 9820
rect 8006 9764 8062 9820
rect 8062 9764 8066 9820
rect 8002 9760 8066 9764
rect 10862 9820 10926 9824
rect 10862 9764 10866 9820
rect 10866 9764 10922 9820
rect 10922 9764 10926 9820
rect 10862 9760 10926 9764
rect 10942 9820 11006 9824
rect 10942 9764 10946 9820
rect 10946 9764 11002 9820
rect 11002 9764 11006 9820
rect 10942 9760 11006 9764
rect 11022 9820 11086 9824
rect 11022 9764 11026 9820
rect 11026 9764 11082 9820
rect 11082 9764 11086 9820
rect 11022 9760 11086 9764
rect 11102 9820 11166 9824
rect 11102 9764 11106 9820
rect 11106 9764 11162 9820
rect 11162 9764 11166 9820
rect 11102 9760 11166 9764
rect 13962 9820 14026 9824
rect 13962 9764 13966 9820
rect 13966 9764 14022 9820
rect 14022 9764 14026 9820
rect 13962 9760 14026 9764
rect 14042 9820 14106 9824
rect 14042 9764 14046 9820
rect 14046 9764 14102 9820
rect 14102 9764 14106 9820
rect 14042 9760 14106 9764
rect 14122 9820 14186 9824
rect 14122 9764 14126 9820
rect 14126 9764 14182 9820
rect 14182 9764 14186 9820
rect 14122 9760 14186 9764
rect 14202 9820 14266 9824
rect 14202 9764 14206 9820
rect 14206 9764 14262 9820
rect 14262 9764 14266 9820
rect 14202 9760 14266 9764
rect 17062 9820 17126 9824
rect 17062 9764 17066 9820
rect 17066 9764 17122 9820
rect 17122 9764 17126 9820
rect 17062 9760 17126 9764
rect 17142 9820 17206 9824
rect 17142 9764 17146 9820
rect 17146 9764 17202 9820
rect 17202 9764 17206 9820
rect 17142 9760 17206 9764
rect 17222 9820 17286 9824
rect 17222 9764 17226 9820
rect 17226 9764 17282 9820
rect 17282 9764 17286 9820
rect 17222 9760 17286 9764
rect 17302 9820 17366 9824
rect 17302 9764 17306 9820
rect 17306 9764 17362 9820
rect 17362 9764 17366 9820
rect 17302 9760 17366 9764
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 3272 9276 3336 9280
rect 3272 9220 3276 9276
rect 3276 9220 3332 9276
rect 3332 9220 3336 9276
rect 3272 9216 3336 9220
rect 3352 9276 3416 9280
rect 3352 9220 3356 9276
rect 3356 9220 3412 9276
rect 3412 9220 3416 9276
rect 3352 9216 3416 9220
rect 6212 9276 6276 9280
rect 6212 9220 6216 9276
rect 6216 9220 6272 9276
rect 6272 9220 6276 9276
rect 6212 9216 6276 9220
rect 6292 9276 6356 9280
rect 6292 9220 6296 9276
rect 6296 9220 6352 9276
rect 6352 9220 6356 9276
rect 6292 9216 6356 9220
rect 6372 9276 6436 9280
rect 6372 9220 6376 9276
rect 6376 9220 6432 9276
rect 6432 9220 6436 9276
rect 6372 9216 6436 9220
rect 6452 9276 6516 9280
rect 6452 9220 6456 9276
rect 6456 9220 6512 9276
rect 6512 9220 6516 9276
rect 6452 9216 6516 9220
rect 9312 9276 9376 9280
rect 9312 9220 9316 9276
rect 9316 9220 9372 9276
rect 9372 9220 9376 9276
rect 9312 9216 9376 9220
rect 9392 9276 9456 9280
rect 9392 9220 9396 9276
rect 9396 9220 9452 9276
rect 9452 9220 9456 9276
rect 9392 9216 9456 9220
rect 9472 9276 9536 9280
rect 9472 9220 9476 9276
rect 9476 9220 9532 9276
rect 9532 9220 9536 9276
rect 9472 9216 9536 9220
rect 9552 9276 9616 9280
rect 9552 9220 9556 9276
rect 9556 9220 9612 9276
rect 9612 9220 9616 9276
rect 9552 9216 9616 9220
rect 12412 9276 12476 9280
rect 12412 9220 12416 9276
rect 12416 9220 12472 9276
rect 12472 9220 12476 9276
rect 12412 9216 12476 9220
rect 12492 9276 12556 9280
rect 12492 9220 12496 9276
rect 12496 9220 12552 9276
rect 12552 9220 12556 9276
rect 12492 9216 12556 9220
rect 12572 9276 12636 9280
rect 12572 9220 12576 9276
rect 12576 9220 12632 9276
rect 12632 9220 12636 9276
rect 12572 9216 12636 9220
rect 12652 9276 12716 9280
rect 12652 9220 12656 9276
rect 12656 9220 12712 9276
rect 12712 9220 12716 9276
rect 12652 9216 12716 9220
rect 15512 9276 15576 9280
rect 15512 9220 15516 9276
rect 15516 9220 15572 9276
rect 15572 9220 15576 9276
rect 15512 9216 15576 9220
rect 15592 9276 15656 9280
rect 15592 9220 15596 9276
rect 15596 9220 15652 9276
rect 15652 9220 15656 9276
rect 15592 9216 15656 9220
rect 15672 9276 15736 9280
rect 15672 9220 15676 9276
rect 15676 9220 15732 9276
rect 15732 9220 15736 9276
rect 15672 9216 15736 9220
rect 15752 9276 15816 9280
rect 15752 9220 15756 9276
rect 15756 9220 15812 9276
rect 15812 9220 15816 9276
rect 15752 9216 15816 9220
rect 4662 8732 4726 8736
rect 4662 8676 4666 8732
rect 4666 8676 4722 8732
rect 4722 8676 4726 8732
rect 4662 8672 4726 8676
rect 4742 8732 4806 8736
rect 4742 8676 4746 8732
rect 4746 8676 4802 8732
rect 4802 8676 4806 8732
rect 4742 8672 4806 8676
rect 4822 8732 4886 8736
rect 4822 8676 4826 8732
rect 4826 8676 4882 8732
rect 4882 8676 4886 8732
rect 4822 8672 4886 8676
rect 4902 8732 4966 8736
rect 4902 8676 4906 8732
rect 4906 8676 4962 8732
rect 4962 8676 4966 8732
rect 4902 8672 4966 8676
rect 7762 8732 7826 8736
rect 7762 8676 7766 8732
rect 7766 8676 7822 8732
rect 7822 8676 7826 8732
rect 7762 8672 7826 8676
rect 7842 8732 7906 8736
rect 7842 8676 7846 8732
rect 7846 8676 7902 8732
rect 7902 8676 7906 8732
rect 7842 8672 7906 8676
rect 7922 8732 7986 8736
rect 7922 8676 7926 8732
rect 7926 8676 7982 8732
rect 7982 8676 7986 8732
rect 7922 8672 7986 8676
rect 8002 8732 8066 8736
rect 8002 8676 8006 8732
rect 8006 8676 8062 8732
rect 8062 8676 8066 8732
rect 8002 8672 8066 8676
rect 10862 8732 10926 8736
rect 10862 8676 10866 8732
rect 10866 8676 10922 8732
rect 10922 8676 10926 8732
rect 10862 8672 10926 8676
rect 10942 8732 11006 8736
rect 10942 8676 10946 8732
rect 10946 8676 11002 8732
rect 11002 8676 11006 8732
rect 10942 8672 11006 8676
rect 11022 8732 11086 8736
rect 11022 8676 11026 8732
rect 11026 8676 11082 8732
rect 11082 8676 11086 8732
rect 11022 8672 11086 8676
rect 11102 8732 11166 8736
rect 11102 8676 11106 8732
rect 11106 8676 11162 8732
rect 11162 8676 11166 8732
rect 11102 8672 11166 8676
rect 13962 8732 14026 8736
rect 13962 8676 13966 8732
rect 13966 8676 14022 8732
rect 14022 8676 14026 8732
rect 13962 8672 14026 8676
rect 14042 8732 14106 8736
rect 14042 8676 14046 8732
rect 14046 8676 14102 8732
rect 14102 8676 14106 8732
rect 14042 8672 14106 8676
rect 14122 8732 14186 8736
rect 14122 8676 14126 8732
rect 14126 8676 14182 8732
rect 14182 8676 14186 8732
rect 14122 8672 14186 8676
rect 14202 8732 14266 8736
rect 14202 8676 14206 8732
rect 14206 8676 14262 8732
rect 14262 8676 14266 8732
rect 14202 8672 14266 8676
rect 17062 8732 17126 8736
rect 17062 8676 17066 8732
rect 17066 8676 17122 8732
rect 17122 8676 17126 8732
rect 17062 8672 17126 8676
rect 17142 8732 17206 8736
rect 17142 8676 17146 8732
rect 17146 8676 17202 8732
rect 17202 8676 17206 8732
rect 17142 8672 17206 8676
rect 17222 8732 17286 8736
rect 17222 8676 17226 8732
rect 17226 8676 17282 8732
rect 17282 8676 17286 8732
rect 17222 8672 17286 8676
rect 17302 8732 17366 8736
rect 17302 8676 17306 8732
rect 17306 8676 17362 8732
rect 17362 8676 17366 8732
rect 17302 8672 17366 8676
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 3272 8188 3336 8192
rect 3272 8132 3276 8188
rect 3276 8132 3332 8188
rect 3332 8132 3336 8188
rect 3272 8128 3336 8132
rect 3352 8188 3416 8192
rect 3352 8132 3356 8188
rect 3356 8132 3412 8188
rect 3412 8132 3416 8188
rect 3352 8128 3416 8132
rect 6212 8188 6276 8192
rect 6212 8132 6216 8188
rect 6216 8132 6272 8188
rect 6272 8132 6276 8188
rect 6212 8128 6276 8132
rect 6292 8188 6356 8192
rect 6292 8132 6296 8188
rect 6296 8132 6352 8188
rect 6352 8132 6356 8188
rect 6292 8128 6356 8132
rect 6372 8188 6436 8192
rect 6372 8132 6376 8188
rect 6376 8132 6432 8188
rect 6432 8132 6436 8188
rect 6372 8128 6436 8132
rect 6452 8188 6516 8192
rect 6452 8132 6456 8188
rect 6456 8132 6512 8188
rect 6512 8132 6516 8188
rect 6452 8128 6516 8132
rect 9312 8188 9376 8192
rect 9312 8132 9316 8188
rect 9316 8132 9372 8188
rect 9372 8132 9376 8188
rect 9312 8128 9376 8132
rect 9392 8188 9456 8192
rect 9392 8132 9396 8188
rect 9396 8132 9452 8188
rect 9452 8132 9456 8188
rect 9392 8128 9456 8132
rect 9472 8188 9536 8192
rect 9472 8132 9476 8188
rect 9476 8132 9532 8188
rect 9532 8132 9536 8188
rect 9472 8128 9536 8132
rect 9552 8188 9616 8192
rect 9552 8132 9556 8188
rect 9556 8132 9612 8188
rect 9612 8132 9616 8188
rect 9552 8128 9616 8132
rect 12412 8188 12476 8192
rect 12412 8132 12416 8188
rect 12416 8132 12472 8188
rect 12472 8132 12476 8188
rect 12412 8128 12476 8132
rect 12492 8188 12556 8192
rect 12492 8132 12496 8188
rect 12496 8132 12552 8188
rect 12552 8132 12556 8188
rect 12492 8128 12556 8132
rect 12572 8188 12636 8192
rect 12572 8132 12576 8188
rect 12576 8132 12632 8188
rect 12632 8132 12636 8188
rect 12572 8128 12636 8132
rect 12652 8188 12716 8192
rect 12652 8132 12656 8188
rect 12656 8132 12712 8188
rect 12712 8132 12716 8188
rect 12652 8128 12716 8132
rect 15512 8188 15576 8192
rect 15512 8132 15516 8188
rect 15516 8132 15572 8188
rect 15572 8132 15576 8188
rect 15512 8128 15576 8132
rect 15592 8188 15656 8192
rect 15592 8132 15596 8188
rect 15596 8132 15652 8188
rect 15652 8132 15656 8188
rect 15592 8128 15656 8132
rect 15672 8188 15736 8192
rect 15672 8132 15676 8188
rect 15676 8132 15732 8188
rect 15732 8132 15736 8188
rect 15672 8128 15736 8132
rect 15752 8188 15816 8192
rect 15752 8132 15756 8188
rect 15756 8132 15812 8188
rect 15812 8132 15816 8188
rect 15752 8128 15816 8132
rect 4662 7644 4726 7648
rect 4662 7588 4666 7644
rect 4666 7588 4722 7644
rect 4722 7588 4726 7644
rect 4662 7584 4726 7588
rect 4742 7644 4806 7648
rect 4742 7588 4746 7644
rect 4746 7588 4802 7644
rect 4802 7588 4806 7644
rect 4742 7584 4806 7588
rect 4822 7644 4886 7648
rect 4822 7588 4826 7644
rect 4826 7588 4882 7644
rect 4882 7588 4886 7644
rect 4822 7584 4886 7588
rect 4902 7644 4966 7648
rect 4902 7588 4906 7644
rect 4906 7588 4962 7644
rect 4962 7588 4966 7644
rect 4902 7584 4966 7588
rect 7762 7644 7826 7648
rect 7762 7588 7766 7644
rect 7766 7588 7822 7644
rect 7822 7588 7826 7644
rect 7762 7584 7826 7588
rect 7842 7644 7906 7648
rect 7842 7588 7846 7644
rect 7846 7588 7902 7644
rect 7902 7588 7906 7644
rect 7842 7584 7906 7588
rect 7922 7644 7986 7648
rect 7922 7588 7926 7644
rect 7926 7588 7982 7644
rect 7982 7588 7986 7644
rect 7922 7584 7986 7588
rect 8002 7644 8066 7648
rect 8002 7588 8006 7644
rect 8006 7588 8062 7644
rect 8062 7588 8066 7644
rect 8002 7584 8066 7588
rect 10862 7644 10926 7648
rect 10862 7588 10866 7644
rect 10866 7588 10922 7644
rect 10922 7588 10926 7644
rect 10862 7584 10926 7588
rect 10942 7644 11006 7648
rect 10942 7588 10946 7644
rect 10946 7588 11002 7644
rect 11002 7588 11006 7644
rect 10942 7584 11006 7588
rect 11022 7644 11086 7648
rect 11022 7588 11026 7644
rect 11026 7588 11082 7644
rect 11082 7588 11086 7644
rect 11022 7584 11086 7588
rect 11102 7644 11166 7648
rect 11102 7588 11106 7644
rect 11106 7588 11162 7644
rect 11162 7588 11166 7644
rect 11102 7584 11166 7588
rect 13962 7644 14026 7648
rect 13962 7588 13966 7644
rect 13966 7588 14022 7644
rect 14022 7588 14026 7644
rect 13962 7584 14026 7588
rect 14042 7644 14106 7648
rect 14042 7588 14046 7644
rect 14046 7588 14102 7644
rect 14102 7588 14106 7644
rect 14042 7584 14106 7588
rect 14122 7644 14186 7648
rect 14122 7588 14126 7644
rect 14126 7588 14182 7644
rect 14182 7588 14186 7644
rect 14122 7584 14186 7588
rect 14202 7644 14266 7648
rect 14202 7588 14206 7644
rect 14206 7588 14262 7644
rect 14262 7588 14266 7644
rect 14202 7584 14266 7588
rect 17062 7644 17126 7648
rect 17062 7588 17066 7644
rect 17066 7588 17122 7644
rect 17122 7588 17126 7644
rect 17062 7584 17126 7588
rect 17142 7644 17206 7648
rect 17142 7588 17146 7644
rect 17146 7588 17202 7644
rect 17202 7588 17206 7644
rect 17142 7584 17206 7588
rect 17222 7644 17286 7648
rect 17222 7588 17226 7644
rect 17226 7588 17282 7644
rect 17282 7588 17286 7644
rect 17222 7584 17286 7588
rect 17302 7644 17366 7648
rect 17302 7588 17306 7644
rect 17306 7588 17362 7644
rect 17362 7588 17366 7644
rect 17302 7584 17366 7588
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 3272 7100 3336 7104
rect 3272 7044 3276 7100
rect 3276 7044 3332 7100
rect 3332 7044 3336 7100
rect 3272 7040 3336 7044
rect 3352 7100 3416 7104
rect 3352 7044 3356 7100
rect 3356 7044 3412 7100
rect 3412 7044 3416 7100
rect 3352 7040 3416 7044
rect 6212 7100 6276 7104
rect 6212 7044 6216 7100
rect 6216 7044 6272 7100
rect 6272 7044 6276 7100
rect 6212 7040 6276 7044
rect 6292 7100 6356 7104
rect 6292 7044 6296 7100
rect 6296 7044 6352 7100
rect 6352 7044 6356 7100
rect 6292 7040 6356 7044
rect 6372 7100 6436 7104
rect 6372 7044 6376 7100
rect 6376 7044 6432 7100
rect 6432 7044 6436 7100
rect 6372 7040 6436 7044
rect 6452 7100 6516 7104
rect 6452 7044 6456 7100
rect 6456 7044 6512 7100
rect 6512 7044 6516 7100
rect 6452 7040 6516 7044
rect 9312 7100 9376 7104
rect 9312 7044 9316 7100
rect 9316 7044 9372 7100
rect 9372 7044 9376 7100
rect 9312 7040 9376 7044
rect 9392 7100 9456 7104
rect 9392 7044 9396 7100
rect 9396 7044 9452 7100
rect 9452 7044 9456 7100
rect 9392 7040 9456 7044
rect 9472 7100 9536 7104
rect 9472 7044 9476 7100
rect 9476 7044 9532 7100
rect 9532 7044 9536 7100
rect 9472 7040 9536 7044
rect 9552 7100 9616 7104
rect 9552 7044 9556 7100
rect 9556 7044 9612 7100
rect 9612 7044 9616 7100
rect 9552 7040 9616 7044
rect 12412 7100 12476 7104
rect 12412 7044 12416 7100
rect 12416 7044 12472 7100
rect 12472 7044 12476 7100
rect 12412 7040 12476 7044
rect 12492 7100 12556 7104
rect 12492 7044 12496 7100
rect 12496 7044 12552 7100
rect 12552 7044 12556 7100
rect 12492 7040 12556 7044
rect 12572 7100 12636 7104
rect 12572 7044 12576 7100
rect 12576 7044 12632 7100
rect 12632 7044 12636 7100
rect 12572 7040 12636 7044
rect 12652 7100 12716 7104
rect 12652 7044 12656 7100
rect 12656 7044 12712 7100
rect 12712 7044 12716 7100
rect 12652 7040 12716 7044
rect 15512 7100 15576 7104
rect 15512 7044 15516 7100
rect 15516 7044 15572 7100
rect 15572 7044 15576 7100
rect 15512 7040 15576 7044
rect 15592 7100 15656 7104
rect 15592 7044 15596 7100
rect 15596 7044 15652 7100
rect 15652 7044 15656 7100
rect 15592 7040 15656 7044
rect 15672 7100 15736 7104
rect 15672 7044 15676 7100
rect 15676 7044 15732 7100
rect 15732 7044 15736 7100
rect 15672 7040 15736 7044
rect 15752 7100 15816 7104
rect 15752 7044 15756 7100
rect 15756 7044 15812 7100
rect 15812 7044 15816 7100
rect 15752 7040 15816 7044
rect 4662 6556 4726 6560
rect 4662 6500 4666 6556
rect 4666 6500 4722 6556
rect 4722 6500 4726 6556
rect 4662 6496 4726 6500
rect 4742 6556 4806 6560
rect 4742 6500 4746 6556
rect 4746 6500 4802 6556
rect 4802 6500 4806 6556
rect 4742 6496 4806 6500
rect 4822 6556 4886 6560
rect 4822 6500 4826 6556
rect 4826 6500 4882 6556
rect 4882 6500 4886 6556
rect 4822 6496 4886 6500
rect 4902 6556 4966 6560
rect 4902 6500 4906 6556
rect 4906 6500 4962 6556
rect 4962 6500 4966 6556
rect 4902 6496 4966 6500
rect 7762 6556 7826 6560
rect 7762 6500 7766 6556
rect 7766 6500 7822 6556
rect 7822 6500 7826 6556
rect 7762 6496 7826 6500
rect 7842 6556 7906 6560
rect 7842 6500 7846 6556
rect 7846 6500 7902 6556
rect 7902 6500 7906 6556
rect 7842 6496 7906 6500
rect 7922 6556 7986 6560
rect 7922 6500 7926 6556
rect 7926 6500 7982 6556
rect 7982 6500 7986 6556
rect 7922 6496 7986 6500
rect 8002 6556 8066 6560
rect 8002 6500 8006 6556
rect 8006 6500 8062 6556
rect 8062 6500 8066 6556
rect 8002 6496 8066 6500
rect 10862 6556 10926 6560
rect 10862 6500 10866 6556
rect 10866 6500 10922 6556
rect 10922 6500 10926 6556
rect 10862 6496 10926 6500
rect 10942 6556 11006 6560
rect 10942 6500 10946 6556
rect 10946 6500 11002 6556
rect 11002 6500 11006 6556
rect 10942 6496 11006 6500
rect 11022 6556 11086 6560
rect 11022 6500 11026 6556
rect 11026 6500 11082 6556
rect 11082 6500 11086 6556
rect 11022 6496 11086 6500
rect 11102 6556 11166 6560
rect 11102 6500 11106 6556
rect 11106 6500 11162 6556
rect 11162 6500 11166 6556
rect 11102 6496 11166 6500
rect 13962 6556 14026 6560
rect 13962 6500 13966 6556
rect 13966 6500 14022 6556
rect 14022 6500 14026 6556
rect 13962 6496 14026 6500
rect 14042 6556 14106 6560
rect 14042 6500 14046 6556
rect 14046 6500 14102 6556
rect 14102 6500 14106 6556
rect 14042 6496 14106 6500
rect 14122 6556 14186 6560
rect 14122 6500 14126 6556
rect 14126 6500 14182 6556
rect 14182 6500 14186 6556
rect 14122 6496 14186 6500
rect 14202 6556 14266 6560
rect 14202 6500 14206 6556
rect 14206 6500 14262 6556
rect 14262 6500 14266 6556
rect 14202 6496 14266 6500
rect 17062 6556 17126 6560
rect 17062 6500 17066 6556
rect 17066 6500 17122 6556
rect 17122 6500 17126 6556
rect 17062 6496 17126 6500
rect 17142 6556 17206 6560
rect 17142 6500 17146 6556
rect 17146 6500 17202 6556
rect 17202 6500 17206 6556
rect 17142 6496 17206 6500
rect 17222 6556 17286 6560
rect 17222 6500 17226 6556
rect 17226 6500 17282 6556
rect 17282 6500 17286 6556
rect 17222 6496 17286 6500
rect 17302 6556 17366 6560
rect 17302 6500 17306 6556
rect 17306 6500 17362 6556
rect 17362 6500 17366 6556
rect 17302 6496 17366 6500
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 3272 6012 3336 6016
rect 3272 5956 3276 6012
rect 3276 5956 3332 6012
rect 3332 5956 3336 6012
rect 3272 5952 3336 5956
rect 3352 6012 3416 6016
rect 3352 5956 3356 6012
rect 3356 5956 3412 6012
rect 3412 5956 3416 6012
rect 3352 5952 3416 5956
rect 6212 6012 6276 6016
rect 6212 5956 6216 6012
rect 6216 5956 6272 6012
rect 6272 5956 6276 6012
rect 6212 5952 6276 5956
rect 6292 6012 6356 6016
rect 6292 5956 6296 6012
rect 6296 5956 6352 6012
rect 6352 5956 6356 6012
rect 6292 5952 6356 5956
rect 6372 6012 6436 6016
rect 6372 5956 6376 6012
rect 6376 5956 6432 6012
rect 6432 5956 6436 6012
rect 6372 5952 6436 5956
rect 6452 6012 6516 6016
rect 6452 5956 6456 6012
rect 6456 5956 6512 6012
rect 6512 5956 6516 6012
rect 6452 5952 6516 5956
rect 9312 6012 9376 6016
rect 9312 5956 9316 6012
rect 9316 5956 9372 6012
rect 9372 5956 9376 6012
rect 9312 5952 9376 5956
rect 9392 6012 9456 6016
rect 9392 5956 9396 6012
rect 9396 5956 9452 6012
rect 9452 5956 9456 6012
rect 9392 5952 9456 5956
rect 9472 6012 9536 6016
rect 9472 5956 9476 6012
rect 9476 5956 9532 6012
rect 9532 5956 9536 6012
rect 9472 5952 9536 5956
rect 9552 6012 9616 6016
rect 9552 5956 9556 6012
rect 9556 5956 9612 6012
rect 9612 5956 9616 6012
rect 9552 5952 9616 5956
rect 12412 6012 12476 6016
rect 12412 5956 12416 6012
rect 12416 5956 12472 6012
rect 12472 5956 12476 6012
rect 12412 5952 12476 5956
rect 12492 6012 12556 6016
rect 12492 5956 12496 6012
rect 12496 5956 12552 6012
rect 12552 5956 12556 6012
rect 12492 5952 12556 5956
rect 12572 6012 12636 6016
rect 12572 5956 12576 6012
rect 12576 5956 12632 6012
rect 12632 5956 12636 6012
rect 12572 5952 12636 5956
rect 12652 6012 12716 6016
rect 12652 5956 12656 6012
rect 12656 5956 12712 6012
rect 12712 5956 12716 6012
rect 12652 5952 12716 5956
rect 15512 6012 15576 6016
rect 15512 5956 15516 6012
rect 15516 5956 15572 6012
rect 15572 5956 15576 6012
rect 15512 5952 15576 5956
rect 15592 6012 15656 6016
rect 15592 5956 15596 6012
rect 15596 5956 15652 6012
rect 15652 5956 15656 6012
rect 15592 5952 15656 5956
rect 15672 6012 15736 6016
rect 15672 5956 15676 6012
rect 15676 5956 15732 6012
rect 15732 5956 15736 6012
rect 15672 5952 15736 5956
rect 15752 6012 15816 6016
rect 15752 5956 15756 6012
rect 15756 5956 15812 6012
rect 15812 5956 15816 6012
rect 15752 5952 15816 5956
rect 4662 5468 4726 5472
rect 4662 5412 4666 5468
rect 4666 5412 4722 5468
rect 4722 5412 4726 5468
rect 4662 5408 4726 5412
rect 4742 5468 4806 5472
rect 4742 5412 4746 5468
rect 4746 5412 4802 5468
rect 4802 5412 4806 5468
rect 4742 5408 4806 5412
rect 4822 5468 4886 5472
rect 4822 5412 4826 5468
rect 4826 5412 4882 5468
rect 4882 5412 4886 5468
rect 4822 5408 4886 5412
rect 4902 5468 4966 5472
rect 4902 5412 4906 5468
rect 4906 5412 4962 5468
rect 4962 5412 4966 5468
rect 4902 5408 4966 5412
rect 7762 5468 7826 5472
rect 7762 5412 7766 5468
rect 7766 5412 7822 5468
rect 7822 5412 7826 5468
rect 7762 5408 7826 5412
rect 7842 5468 7906 5472
rect 7842 5412 7846 5468
rect 7846 5412 7902 5468
rect 7902 5412 7906 5468
rect 7842 5408 7906 5412
rect 7922 5468 7986 5472
rect 7922 5412 7926 5468
rect 7926 5412 7982 5468
rect 7982 5412 7986 5468
rect 7922 5408 7986 5412
rect 8002 5468 8066 5472
rect 8002 5412 8006 5468
rect 8006 5412 8062 5468
rect 8062 5412 8066 5468
rect 8002 5408 8066 5412
rect 10862 5468 10926 5472
rect 10862 5412 10866 5468
rect 10866 5412 10922 5468
rect 10922 5412 10926 5468
rect 10862 5408 10926 5412
rect 10942 5468 11006 5472
rect 10942 5412 10946 5468
rect 10946 5412 11002 5468
rect 11002 5412 11006 5468
rect 10942 5408 11006 5412
rect 11022 5468 11086 5472
rect 11022 5412 11026 5468
rect 11026 5412 11082 5468
rect 11082 5412 11086 5468
rect 11022 5408 11086 5412
rect 11102 5468 11166 5472
rect 11102 5412 11106 5468
rect 11106 5412 11162 5468
rect 11162 5412 11166 5468
rect 11102 5408 11166 5412
rect 13962 5468 14026 5472
rect 13962 5412 13966 5468
rect 13966 5412 14022 5468
rect 14022 5412 14026 5468
rect 13962 5408 14026 5412
rect 14042 5468 14106 5472
rect 14042 5412 14046 5468
rect 14046 5412 14102 5468
rect 14102 5412 14106 5468
rect 14042 5408 14106 5412
rect 14122 5468 14186 5472
rect 14122 5412 14126 5468
rect 14126 5412 14182 5468
rect 14182 5412 14186 5468
rect 14122 5408 14186 5412
rect 14202 5468 14266 5472
rect 14202 5412 14206 5468
rect 14206 5412 14262 5468
rect 14262 5412 14266 5468
rect 14202 5408 14266 5412
rect 17062 5468 17126 5472
rect 17062 5412 17066 5468
rect 17066 5412 17122 5468
rect 17122 5412 17126 5468
rect 17062 5408 17126 5412
rect 17142 5468 17206 5472
rect 17142 5412 17146 5468
rect 17146 5412 17202 5468
rect 17202 5412 17206 5468
rect 17142 5408 17206 5412
rect 17222 5468 17286 5472
rect 17222 5412 17226 5468
rect 17226 5412 17282 5468
rect 17282 5412 17286 5468
rect 17222 5408 17286 5412
rect 17302 5468 17366 5472
rect 17302 5412 17306 5468
rect 17306 5412 17362 5468
rect 17362 5412 17366 5468
rect 17302 5408 17366 5412
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 3272 4924 3336 4928
rect 3272 4868 3276 4924
rect 3276 4868 3332 4924
rect 3332 4868 3336 4924
rect 3272 4864 3336 4868
rect 3352 4924 3416 4928
rect 3352 4868 3356 4924
rect 3356 4868 3412 4924
rect 3412 4868 3416 4924
rect 3352 4864 3416 4868
rect 6212 4924 6276 4928
rect 6212 4868 6216 4924
rect 6216 4868 6272 4924
rect 6272 4868 6276 4924
rect 6212 4864 6276 4868
rect 6292 4924 6356 4928
rect 6292 4868 6296 4924
rect 6296 4868 6352 4924
rect 6352 4868 6356 4924
rect 6292 4864 6356 4868
rect 6372 4924 6436 4928
rect 6372 4868 6376 4924
rect 6376 4868 6432 4924
rect 6432 4868 6436 4924
rect 6372 4864 6436 4868
rect 6452 4924 6516 4928
rect 6452 4868 6456 4924
rect 6456 4868 6512 4924
rect 6512 4868 6516 4924
rect 6452 4864 6516 4868
rect 9312 4924 9376 4928
rect 9312 4868 9316 4924
rect 9316 4868 9372 4924
rect 9372 4868 9376 4924
rect 9312 4864 9376 4868
rect 9392 4924 9456 4928
rect 9392 4868 9396 4924
rect 9396 4868 9452 4924
rect 9452 4868 9456 4924
rect 9392 4864 9456 4868
rect 9472 4924 9536 4928
rect 9472 4868 9476 4924
rect 9476 4868 9532 4924
rect 9532 4868 9536 4924
rect 9472 4864 9536 4868
rect 9552 4924 9616 4928
rect 9552 4868 9556 4924
rect 9556 4868 9612 4924
rect 9612 4868 9616 4924
rect 9552 4864 9616 4868
rect 12412 4924 12476 4928
rect 12412 4868 12416 4924
rect 12416 4868 12472 4924
rect 12472 4868 12476 4924
rect 12412 4864 12476 4868
rect 12492 4924 12556 4928
rect 12492 4868 12496 4924
rect 12496 4868 12552 4924
rect 12552 4868 12556 4924
rect 12492 4864 12556 4868
rect 12572 4924 12636 4928
rect 12572 4868 12576 4924
rect 12576 4868 12632 4924
rect 12632 4868 12636 4924
rect 12572 4864 12636 4868
rect 12652 4924 12716 4928
rect 12652 4868 12656 4924
rect 12656 4868 12712 4924
rect 12712 4868 12716 4924
rect 12652 4864 12716 4868
rect 15512 4924 15576 4928
rect 15512 4868 15516 4924
rect 15516 4868 15572 4924
rect 15572 4868 15576 4924
rect 15512 4864 15576 4868
rect 15592 4924 15656 4928
rect 15592 4868 15596 4924
rect 15596 4868 15652 4924
rect 15652 4868 15656 4924
rect 15592 4864 15656 4868
rect 15672 4924 15736 4928
rect 15672 4868 15676 4924
rect 15676 4868 15732 4924
rect 15732 4868 15736 4924
rect 15672 4864 15736 4868
rect 15752 4924 15816 4928
rect 15752 4868 15756 4924
rect 15756 4868 15812 4924
rect 15812 4868 15816 4924
rect 15752 4864 15816 4868
rect 4662 4380 4726 4384
rect 4662 4324 4666 4380
rect 4666 4324 4722 4380
rect 4722 4324 4726 4380
rect 4662 4320 4726 4324
rect 4742 4380 4806 4384
rect 4742 4324 4746 4380
rect 4746 4324 4802 4380
rect 4802 4324 4806 4380
rect 4742 4320 4806 4324
rect 4822 4380 4886 4384
rect 4822 4324 4826 4380
rect 4826 4324 4882 4380
rect 4882 4324 4886 4380
rect 4822 4320 4886 4324
rect 4902 4380 4966 4384
rect 4902 4324 4906 4380
rect 4906 4324 4962 4380
rect 4962 4324 4966 4380
rect 4902 4320 4966 4324
rect 7762 4380 7826 4384
rect 7762 4324 7766 4380
rect 7766 4324 7822 4380
rect 7822 4324 7826 4380
rect 7762 4320 7826 4324
rect 7842 4380 7906 4384
rect 7842 4324 7846 4380
rect 7846 4324 7902 4380
rect 7902 4324 7906 4380
rect 7842 4320 7906 4324
rect 7922 4380 7986 4384
rect 7922 4324 7926 4380
rect 7926 4324 7982 4380
rect 7982 4324 7986 4380
rect 7922 4320 7986 4324
rect 8002 4380 8066 4384
rect 8002 4324 8006 4380
rect 8006 4324 8062 4380
rect 8062 4324 8066 4380
rect 8002 4320 8066 4324
rect 10862 4380 10926 4384
rect 10862 4324 10866 4380
rect 10866 4324 10922 4380
rect 10922 4324 10926 4380
rect 10862 4320 10926 4324
rect 10942 4380 11006 4384
rect 10942 4324 10946 4380
rect 10946 4324 11002 4380
rect 11002 4324 11006 4380
rect 10942 4320 11006 4324
rect 11022 4380 11086 4384
rect 11022 4324 11026 4380
rect 11026 4324 11082 4380
rect 11082 4324 11086 4380
rect 11022 4320 11086 4324
rect 11102 4380 11166 4384
rect 11102 4324 11106 4380
rect 11106 4324 11162 4380
rect 11162 4324 11166 4380
rect 11102 4320 11166 4324
rect 13962 4380 14026 4384
rect 13962 4324 13966 4380
rect 13966 4324 14022 4380
rect 14022 4324 14026 4380
rect 13962 4320 14026 4324
rect 14042 4380 14106 4384
rect 14042 4324 14046 4380
rect 14046 4324 14102 4380
rect 14102 4324 14106 4380
rect 14042 4320 14106 4324
rect 14122 4380 14186 4384
rect 14122 4324 14126 4380
rect 14126 4324 14182 4380
rect 14182 4324 14186 4380
rect 14122 4320 14186 4324
rect 14202 4380 14266 4384
rect 14202 4324 14206 4380
rect 14206 4324 14262 4380
rect 14262 4324 14266 4380
rect 14202 4320 14266 4324
rect 17062 4380 17126 4384
rect 17062 4324 17066 4380
rect 17066 4324 17122 4380
rect 17122 4324 17126 4380
rect 17062 4320 17126 4324
rect 17142 4380 17206 4384
rect 17142 4324 17146 4380
rect 17146 4324 17202 4380
rect 17202 4324 17206 4380
rect 17142 4320 17206 4324
rect 17222 4380 17286 4384
rect 17222 4324 17226 4380
rect 17226 4324 17282 4380
rect 17282 4324 17286 4380
rect 17222 4320 17286 4324
rect 17302 4380 17366 4384
rect 17302 4324 17306 4380
rect 17306 4324 17362 4380
rect 17362 4324 17366 4380
rect 17302 4320 17366 4324
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 3272 3836 3336 3840
rect 3272 3780 3276 3836
rect 3276 3780 3332 3836
rect 3332 3780 3336 3836
rect 3272 3776 3336 3780
rect 3352 3836 3416 3840
rect 3352 3780 3356 3836
rect 3356 3780 3412 3836
rect 3412 3780 3416 3836
rect 3352 3776 3416 3780
rect 6212 3836 6276 3840
rect 6212 3780 6216 3836
rect 6216 3780 6272 3836
rect 6272 3780 6276 3836
rect 6212 3776 6276 3780
rect 6292 3836 6356 3840
rect 6292 3780 6296 3836
rect 6296 3780 6352 3836
rect 6352 3780 6356 3836
rect 6292 3776 6356 3780
rect 6372 3836 6436 3840
rect 6372 3780 6376 3836
rect 6376 3780 6432 3836
rect 6432 3780 6436 3836
rect 6372 3776 6436 3780
rect 6452 3836 6516 3840
rect 6452 3780 6456 3836
rect 6456 3780 6512 3836
rect 6512 3780 6516 3836
rect 6452 3776 6516 3780
rect 9312 3836 9376 3840
rect 9312 3780 9316 3836
rect 9316 3780 9372 3836
rect 9372 3780 9376 3836
rect 9312 3776 9376 3780
rect 9392 3836 9456 3840
rect 9392 3780 9396 3836
rect 9396 3780 9452 3836
rect 9452 3780 9456 3836
rect 9392 3776 9456 3780
rect 9472 3836 9536 3840
rect 9472 3780 9476 3836
rect 9476 3780 9532 3836
rect 9532 3780 9536 3836
rect 9472 3776 9536 3780
rect 9552 3836 9616 3840
rect 9552 3780 9556 3836
rect 9556 3780 9612 3836
rect 9612 3780 9616 3836
rect 9552 3776 9616 3780
rect 12412 3836 12476 3840
rect 12412 3780 12416 3836
rect 12416 3780 12472 3836
rect 12472 3780 12476 3836
rect 12412 3776 12476 3780
rect 12492 3836 12556 3840
rect 12492 3780 12496 3836
rect 12496 3780 12552 3836
rect 12552 3780 12556 3836
rect 12492 3776 12556 3780
rect 12572 3836 12636 3840
rect 12572 3780 12576 3836
rect 12576 3780 12632 3836
rect 12632 3780 12636 3836
rect 12572 3776 12636 3780
rect 12652 3836 12716 3840
rect 12652 3780 12656 3836
rect 12656 3780 12712 3836
rect 12712 3780 12716 3836
rect 12652 3776 12716 3780
rect 15512 3836 15576 3840
rect 15512 3780 15516 3836
rect 15516 3780 15572 3836
rect 15572 3780 15576 3836
rect 15512 3776 15576 3780
rect 15592 3836 15656 3840
rect 15592 3780 15596 3836
rect 15596 3780 15652 3836
rect 15652 3780 15656 3836
rect 15592 3776 15656 3780
rect 15672 3836 15736 3840
rect 15672 3780 15676 3836
rect 15676 3780 15732 3836
rect 15732 3780 15736 3836
rect 15672 3776 15736 3780
rect 15752 3836 15816 3840
rect 15752 3780 15756 3836
rect 15756 3780 15812 3836
rect 15812 3780 15816 3836
rect 15752 3776 15816 3780
rect 4662 3292 4726 3296
rect 4662 3236 4666 3292
rect 4666 3236 4722 3292
rect 4722 3236 4726 3292
rect 4662 3232 4726 3236
rect 4742 3292 4806 3296
rect 4742 3236 4746 3292
rect 4746 3236 4802 3292
rect 4802 3236 4806 3292
rect 4742 3232 4806 3236
rect 4822 3292 4886 3296
rect 4822 3236 4826 3292
rect 4826 3236 4882 3292
rect 4882 3236 4886 3292
rect 4822 3232 4886 3236
rect 4902 3292 4966 3296
rect 4902 3236 4906 3292
rect 4906 3236 4962 3292
rect 4962 3236 4966 3292
rect 4902 3232 4966 3236
rect 7762 3292 7826 3296
rect 7762 3236 7766 3292
rect 7766 3236 7822 3292
rect 7822 3236 7826 3292
rect 7762 3232 7826 3236
rect 7842 3292 7906 3296
rect 7842 3236 7846 3292
rect 7846 3236 7902 3292
rect 7902 3236 7906 3292
rect 7842 3232 7906 3236
rect 7922 3292 7986 3296
rect 7922 3236 7926 3292
rect 7926 3236 7982 3292
rect 7982 3236 7986 3292
rect 7922 3232 7986 3236
rect 8002 3292 8066 3296
rect 8002 3236 8006 3292
rect 8006 3236 8062 3292
rect 8062 3236 8066 3292
rect 8002 3232 8066 3236
rect 10862 3292 10926 3296
rect 10862 3236 10866 3292
rect 10866 3236 10922 3292
rect 10922 3236 10926 3292
rect 10862 3232 10926 3236
rect 10942 3292 11006 3296
rect 10942 3236 10946 3292
rect 10946 3236 11002 3292
rect 11002 3236 11006 3292
rect 10942 3232 11006 3236
rect 11022 3292 11086 3296
rect 11022 3236 11026 3292
rect 11026 3236 11082 3292
rect 11082 3236 11086 3292
rect 11022 3232 11086 3236
rect 11102 3292 11166 3296
rect 11102 3236 11106 3292
rect 11106 3236 11162 3292
rect 11162 3236 11166 3292
rect 11102 3232 11166 3236
rect 13962 3292 14026 3296
rect 13962 3236 13966 3292
rect 13966 3236 14022 3292
rect 14022 3236 14026 3292
rect 13962 3232 14026 3236
rect 14042 3292 14106 3296
rect 14042 3236 14046 3292
rect 14046 3236 14102 3292
rect 14102 3236 14106 3292
rect 14042 3232 14106 3236
rect 14122 3292 14186 3296
rect 14122 3236 14126 3292
rect 14126 3236 14182 3292
rect 14182 3236 14186 3292
rect 14122 3232 14186 3236
rect 14202 3292 14266 3296
rect 14202 3236 14206 3292
rect 14206 3236 14262 3292
rect 14262 3236 14266 3292
rect 14202 3232 14266 3236
rect 17062 3292 17126 3296
rect 17062 3236 17066 3292
rect 17066 3236 17122 3292
rect 17122 3236 17126 3292
rect 17062 3232 17126 3236
rect 17142 3292 17206 3296
rect 17142 3236 17146 3292
rect 17146 3236 17202 3292
rect 17202 3236 17206 3292
rect 17142 3232 17206 3236
rect 17222 3292 17286 3296
rect 17222 3236 17226 3292
rect 17226 3236 17282 3292
rect 17282 3236 17286 3292
rect 17222 3232 17286 3236
rect 17302 3292 17366 3296
rect 17302 3236 17306 3292
rect 17306 3236 17362 3292
rect 17362 3236 17366 3292
rect 17302 3232 17366 3236
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 3272 2748 3336 2752
rect 3272 2692 3276 2748
rect 3276 2692 3332 2748
rect 3332 2692 3336 2748
rect 3272 2688 3336 2692
rect 3352 2748 3416 2752
rect 3352 2692 3356 2748
rect 3356 2692 3412 2748
rect 3412 2692 3416 2748
rect 3352 2688 3416 2692
rect 6212 2748 6276 2752
rect 6212 2692 6216 2748
rect 6216 2692 6272 2748
rect 6272 2692 6276 2748
rect 6212 2688 6276 2692
rect 6292 2748 6356 2752
rect 6292 2692 6296 2748
rect 6296 2692 6352 2748
rect 6352 2692 6356 2748
rect 6292 2688 6356 2692
rect 6372 2748 6436 2752
rect 6372 2692 6376 2748
rect 6376 2692 6432 2748
rect 6432 2692 6436 2748
rect 6372 2688 6436 2692
rect 6452 2748 6516 2752
rect 6452 2692 6456 2748
rect 6456 2692 6512 2748
rect 6512 2692 6516 2748
rect 6452 2688 6516 2692
rect 9312 2748 9376 2752
rect 9312 2692 9316 2748
rect 9316 2692 9372 2748
rect 9372 2692 9376 2748
rect 9312 2688 9376 2692
rect 9392 2748 9456 2752
rect 9392 2692 9396 2748
rect 9396 2692 9452 2748
rect 9452 2692 9456 2748
rect 9392 2688 9456 2692
rect 9472 2748 9536 2752
rect 9472 2692 9476 2748
rect 9476 2692 9532 2748
rect 9532 2692 9536 2748
rect 9472 2688 9536 2692
rect 9552 2748 9616 2752
rect 9552 2692 9556 2748
rect 9556 2692 9612 2748
rect 9612 2692 9616 2748
rect 9552 2688 9616 2692
rect 12412 2748 12476 2752
rect 12412 2692 12416 2748
rect 12416 2692 12472 2748
rect 12472 2692 12476 2748
rect 12412 2688 12476 2692
rect 12492 2748 12556 2752
rect 12492 2692 12496 2748
rect 12496 2692 12552 2748
rect 12552 2692 12556 2748
rect 12492 2688 12556 2692
rect 12572 2748 12636 2752
rect 12572 2692 12576 2748
rect 12576 2692 12632 2748
rect 12632 2692 12636 2748
rect 12572 2688 12636 2692
rect 12652 2748 12716 2752
rect 12652 2692 12656 2748
rect 12656 2692 12712 2748
rect 12712 2692 12716 2748
rect 12652 2688 12716 2692
rect 15512 2748 15576 2752
rect 15512 2692 15516 2748
rect 15516 2692 15572 2748
rect 15572 2692 15576 2748
rect 15512 2688 15576 2692
rect 15592 2748 15656 2752
rect 15592 2692 15596 2748
rect 15596 2692 15652 2748
rect 15652 2692 15656 2748
rect 15592 2688 15656 2692
rect 15672 2748 15736 2752
rect 15672 2692 15676 2748
rect 15676 2692 15732 2748
rect 15732 2692 15736 2748
rect 15672 2688 15736 2692
rect 15752 2748 15816 2752
rect 15752 2692 15756 2748
rect 15756 2692 15812 2748
rect 15812 2692 15816 2748
rect 15752 2688 15816 2692
rect 4662 2204 4726 2208
rect 4662 2148 4666 2204
rect 4666 2148 4722 2204
rect 4722 2148 4726 2204
rect 4662 2144 4726 2148
rect 4742 2204 4806 2208
rect 4742 2148 4746 2204
rect 4746 2148 4802 2204
rect 4802 2148 4806 2204
rect 4742 2144 4806 2148
rect 4822 2204 4886 2208
rect 4822 2148 4826 2204
rect 4826 2148 4882 2204
rect 4882 2148 4886 2204
rect 4822 2144 4886 2148
rect 4902 2204 4966 2208
rect 4902 2148 4906 2204
rect 4906 2148 4962 2204
rect 4962 2148 4966 2204
rect 4902 2144 4966 2148
rect 7762 2204 7826 2208
rect 7762 2148 7766 2204
rect 7766 2148 7822 2204
rect 7822 2148 7826 2204
rect 7762 2144 7826 2148
rect 7842 2204 7906 2208
rect 7842 2148 7846 2204
rect 7846 2148 7902 2204
rect 7902 2148 7906 2204
rect 7842 2144 7906 2148
rect 7922 2204 7986 2208
rect 7922 2148 7926 2204
rect 7926 2148 7982 2204
rect 7982 2148 7986 2204
rect 7922 2144 7986 2148
rect 8002 2204 8066 2208
rect 8002 2148 8006 2204
rect 8006 2148 8062 2204
rect 8062 2148 8066 2204
rect 8002 2144 8066 2148
rect 10862 2204 10926 2208
rect 10862 2148 10866 2204
rect 10866 2148 10922 2204
rect 10922 2148 10926 2204
rect 10862 2144 10926 2148
rect 10942 2204 11006 2208
rect 10942 2148 10946 2204
rect 10946 2148 11002 2204
rect 11002 2148 11006 2204
rect 10942 2144 11006 2148
rect 11022 2204 11086 2208
rect 11022 2148 11026 2204
rect 11026 2148 11082 2204
rect 11082 2148 11086 2204
rect 11022 2144 11086 2148
rect 11102 2204 11166 2208
rect 11102 2148 11106 2204
rect 11106 2148 11162 2204
rect 11162 2148 11166 2204
rect 11102 2144 11166 2148
rect 13962 2204 14026 2208
rect 13962 2148 13966 2204
rect 13966 2148 14022 2204
rect 14022 2148 14026 2204
rect 13962 2144 14026 2148
rect 14042 2204 14106 2208
rect 14042 2148 14046 2204
rect 14046 2148 14102 2204
rect 14102 2148 14106 2204
rect 14042 2144 14106 2148
rect 14122 2204 14186 2208
rect 14122 2148 14126 2204
rect 14126 2148 14182 2204
rect 14182 2148 14186 2204
rect 14122 2144 14186 2148
rect 14202 2204 14266 2208
rect 14202 2148 14206 2204
rect 14206 2148 14262 2204
rect 14262 2148 14266 2204
rect 14202 2144 14266 2148
rect 17062 2204 17126 2208
rect 17062 2148 17066 2204
rect 17066 2148 17122 2204
rect 17122 2148 17126 2204
rect 17062 2144 17126 2148
rect 17142 2204 17206 2208
rect 17142 2148 17146 2204
rect 17146 2148 17202 2204
rect 17202 2148 17206 2204
rect 17142 2144 17206 2148
rect 17222 2204 17286 2208
rect 17222 2148 17226 2204
rect 17226 2148 17282 2204
rect 17282 2148 17286 2204
rect 17222 2144 17286 2148
rect 17302 2204 17366 2208
rect 17302 2148 17306 2204
rect 17306 2148 17362 2204
rect 17362 2148 17366 2204
rect 17302 2144 17366 2148
rect 3112 1660 3176 1664
rect 3112 1604 3116 1660
rect 3116 1604 3172 1660
rect 3172 1604 3176 1660
rect 3112 1600 3176 1604
rect 3192 1660 3256 1664
rect 3192 1604 3196 1660
rect 3196 1604 3252 1660
rect 3252 1604 3256 1660
rect 3192 1600 3256 1604
rect 3272 1660 3336 1664
rect 3272 1604 3276 1660
rect 3276 1604 3332 1660
rect 3332 1604 3336 1660
rect 3272 1600 3336 1604
rect 3352 1660 3416 1664
rect 3352 1604 3356 1660
rect 3356 1604 3412 1660
rect 3412 1604 3416 1660
rect 3352 1600 3416 1604
rect 6212 1660 6276 1664
rect 6212 1604 6216 1660
rect 6216 1604 6272 1660
rect 6272 1604 6276 1660
rect 6212 1600 6276 1604
rect 6292 1660 6356 1664
rect 6292 1604 6296 1660
rect 6296 1604 6352 1660
rect 6352 1604 6356 1660
rect 6292 1600 6356 1604
rect 6372 1660 6436 1664
rect 6372 1604 6376 1660
rect 6376 1604 6432 1660
rect 6432 1604 6436 1660
rect 6372 1600 6436 1604
rect 6452 1660 6516 1664
rect 6452 1604 6456 1660
rect 6456 1604 6512 1660
rect 6512 1604 6516 1660
rect 6452 1600 6516 1604
rect 9312 1660 9376 1664
rect 9312 1604 9316 1660
rect 9316 1604 9372 1660
rect 9372 1604 9376 1660
rect 9312 1600 9376 1604
rect 9392 1660 9456 1664
rect 9392 1604 9396 1660
rect 9396 1604 9452 1660
rect 9452 1604 9456 1660
rect 9392 1600 9456 1604
rect 9472 1660 9536 1664
rect 9472 1604 9476 1660
rect 9476 1604 9532 1660
rect 9532 1604 9536 1660
rect 9472 1600 9536 1604
rect 9552 1660 9616 1664
rect 9552 1604 9556 1660
rect 9556 1604 9612 1660
rect 9612 1604 9616 1660
rect 9552 1600 9616 1604
rect 12412 1660 12476 1664
rect 12412 1604 12416 1660
rect 12416 1604 12472 1660
rect 12472 1604 12476 1660
rect 12412 1600 12476 1604
rect 12492 1660 12556 1664
rect 12492 1604 12496 1660
rect 12496 1604 12552 1660
rect 12552 1604 12556 1660
rect 12492 1600 12556 1604
rect 12572 1660 12636 1664
rect 12572 1604 12576 1660
rect 12576 1604 12632 1660
rect 12632 1604 12636 1660
rect 12572 1600 12636 1604
rect 12652 1660 12716 1664
rect 12652 1604 12656 1660
rect 12656 1604 12712 1660
rect 12712 1604 12716 1660
rect 12652 1600 12716 1604
rect 15512 1660 15576 1664
rect 15512 1604 15516 1660
rect 15516 1604 15572 1660
rect 15572 1604 15576 1660
rect 15512 1600 15576 1604
rect 15592 1660 15656 1664
rect 15592 1604 15596 1660
rect 15596 1604 15652 1660
rect 15652 1604 15656 1660
rect 15592 1600 15656 1604
rect 15672 1660 15736 1664
rect 15672 1604 15676 1660
rect 15676 1604 15732 1660
rect 15732 1604 15736 1660
rect 15672 1600 15736 1604
rect 15752 1660 15816 1664
rect 15752 1604 15756 1660
rect 15756 1604 15812 1660
rect 15812 1604 15816 1660
rect 15752 1600 15816 1604
rect 4662 1116 4726 1120
rect 4662 1060 4666 1116
rect 4666 1060 4722 1116
rect 4722 1060 4726 1116
rect 4662 1056 4726 1060
rect 4742 1116 4806 1120
rect 4742 1060 4746 1116
rect 4746 1060 4802 1116
rect 4802 1060 4806 1116
rect 4742 1056 4806 1060
rect 4822 1116 4886 1120
rect 4822 1060 4826 1116
rect 4826 1060 4882 1116
rect 4882 1060 4886 1116
rect 4822 1056 4886 1060
rect 4902 1116 4966 1120
rect 4902 1060 4906 1116
rect 4906 1060 4962 1116
rect 4962 1060 4966 1116
rect 4902 1056 4966 1060
rect 7762 1116 7826 1120
rect 7762 1060 7766 1116
rect 7766 1060 7822 1116
rect 7822 1060 7826 1116
rect 7762 1056 7826 1060
rect 7842 1116 7906 1120
rect 7842 1060 7846 1116
rect 7846 1060 7902 1116
rect 7902 1060 7906 1116
rect 7842 1056 7906 1060
rect 7922 1116 7986 1120
rect 7922 1060 7926 1116
rect 7926 1060 7982 1116
rect 7982 1060 7986 1116
rect 7922 1056 7986 1060
rect 8002 1116 8066 1120
rect 8002 1060 8006 1116
rect 8006 1060 8062 1116
rect 8062 1060 8066 1116
rect 8002 1056 8066 1060
rect 10862 1116 10926 1120
rect 10862 1060 10866 1116
rect 10866 1060 10922 1116
rect 10922 1060 10926 1116
rect 10862 1056 10926 1060
rect 10942 1116 11006 1120
rect 10942 1060 10946 1116
rect 10946 1060 11002 1116
rect 11002 1060 11006 1116
rect 10942 1056 11006 1060
rect 11022 1116 11086 1120
rect 11022 1060 11026 1116
rect 11026 1060 11082 1116
rect 11082 1060 11086 1116
rect 11022 1056 11086 1060
rect 11102 1116 11166 1120
rect 11102 1060 11106 1116
rect 11106 1060 11162 1116
rect 11162 1060 11166 1116
rect 11102 1056 11166 1060
rect 13962 1116 14026 1120
rect 13962 1060 13966 1116
rect 13966 1060 14022 1116
rect 14022 1060 14026 1116
rect 13962 1056 14026 1060
rect 14042 1116 14106 1120
rect 14042 1060 14046 1116
rect 14046 1060 14102 1116
rect 14102 1060 14106 1116
rect 14042 1056 14106 1060
rect 14122 1116 14186 1120
rect 14122 1060 14126 1116
rect 14126 1060 14182 1116
rect 14182 1060 14186 1116
rect 14122 1056 14186 1060
rect 14202 1116 14266 1120
rect 14202 1060 14206 1116
rect 14206 1060 14262 1116
rect 14262 1060 14266 1116
rect 14202 1056 14266 1060
rect 17062 1116 17126 1120
rect 17062 1060 17066 1116
rect 17066 1060 17122 1116
rect 17122 1060 17126 1116
rect 17062 1056 17126 1060
rect 17142 1116 17206 1120
rect 17142 1060 17146 1116
rect 17146 1060 17202 1116
rect 17202 1060 17206 1116
rect 17142 1056 17206 1060
rect 17222 1116 17286 1120
rect 17222 1060 17226 1116
rect 17226 1060 17282 1116
rect 17282 1060 17286 1116
rect 17222 1056 17286 1060
rect 17302 1116 17366 1120
rect 17302 1060 17306 1116
rect 17306 1060 17362 1116
rect 17362 1060 17366 1116
rect 17302 1056 17366 1060
rect 3112 572 3176 576
rect 3112 516 3116 572
rect 3116 516 3172 572
rect 3172 516 3176 572
rect 3112 512 3176 516
rect 3192 572 3256 576
rect 3192 516 3196 572
rect 3196 516 3252 572
rect 3252 516 3256 572
rect 3192 512 3256 516
rect 3272 572 3336 576
rect 3272 516 3276 572
rect 3276 516 3332 572
rect 3332 516 3336 572
rect 3272 512 3336 516
rect 3352 572 3416 576
rect 3352 516 3356 572
rect 3356 516 3412 572
rect 3412 516 3416 572
rect 3352 512 3416 516
rect 6212 572 6276 576
rect 6212 516 6216 572
rect 6216 516 6272 572
rect 6272 516 6276 572
rect 6212 512 6276 516
rect 6292 572 6356 576
rect 6292 516 6296 572
rect 6296 516 6352 572
rect 6352 516 6356 572
rect 6292 512 6356 516
rect 6372 572 6436 576
rect 6372 516 6376 572
rect 6376 516 6432 572
rect 6432 516 6436 572
rect 6372 512 6436 516
rect 6452 572 6516 576
rect 6452 516 6456 572
rect 6456 516 6512 572
rect 6512 516 6516 572
rect 6452 512 6516 516
rect 9312 572 9376 576
rect 9312 516 9316 572
rect 9316 516 9372 572
rect 9372 516 9376 572
rect 9312 512 9376 516
rect 9392 572 9456 576
rect 9392 516 9396 572
rect 9396 516 9452 572
rect 9452 516 9456 572
rect 9392 512 9456 516
rect 9472 572 9536 576
rect 9472 516 9476 572
rect 9476 516 9532 572
rect 9532 516 9536 572
rect 9472 512 9536 516
rect 9552 572 9616 576
rect 9552 516 9556 572
rect 9556 516 9612 572
rect 9612 516 9616 572
rect 9552 512 9616 516
rect 12412 572 12476 576
rect 12412 516 12416 572
rect 12416 516 12472 572
rect 12472 516 12476 572
rect 12412 512 12476 516
rect 12492 572 12556 576
rect 12492 516 12496 572
rect 12496 516 12552 572
rect 12552 516 12556 572
rect 12492 512 12556 516
rect 12572 572 12636 576
rect 12572 516 12576 572
rect 12576 516 12632 572
rect 12632 516 12636 572
rect 12572 512 12636 516
rect 12652 572 12716 576
rect 12652 516 12656 572
rect 12656 516 12712 572
rect 12712 516 12716 572
rect 12652 512 12716 516
rect 15512 572 15576 576
rect 15512 516 15516 572
rect 15516 516 15572 572
rect 15572 516 15576 572
rect 15512 512 15576 516
rect 15592 572 15656 576
rect 15592 516 15596 572
rect 15596 516 15652 572
rect 15652 516 15656 572
rect 15592 512 15656 516
rect 15672 572 15736 576
rect 15672 516 15676 572
rect 15676 516 15732 572
rect 15732 516 15736 572
rect 15672 512 15736 516
rect 15752 572 15816 576
rect 15752 516 15756 572
rect 15756 516 15812 572
rect 15812 516 15816 572
rect 15752 512 15816 516
rect 4662 28 4726 32
rect 4662 -28 4666 28
rect 4666 -28 4722 28
rect 4722 -28 4726 28
rect 4662 -32 4726 -28
rect 4742 28 4806 32
rect 4742 -28 4746 28
rect 4746 -28 4802 28
rect 4802 -28 4806 28
rect 4742 -32 4806 -28
rect 4822 28 4886 32
rect 4822 -28 4826 28
rect 4826 -28 4882 28
rect 4882 -28 4886 28
rect 4822 -32 4886 -28
rect 4902 28 4966 32
rect 4902 -28 4906 28
rect 4906 -28 4962 28
rect 4962 -28 4966 28
rect 4902 -32 4966 -28
rect 7762 28 7826 32
rect 7762 -28 7766 28
rect 7766 -28 7822 28
rect 7822 -28 7826 28
rect 7762 -32 7826 -28
rect 7842 28 7906 32
rect 7842 -28 7846 28
rect 7846 -28 7902 28
rect 7902 -28 7906 28
rect 7842 -32 7906 -28
rect 7922 28 7986 32
rect 7922 -28 7926 28
rect 7926 -28 7982 28
rect 7982 -28 7986 28
rect 7922 -32 7986 -28
rect 8002 28 8066 32
rect 8002 -28 8006 28
rect 8006 -28 8062 28
rect 8062 -28 8066 28
rect 8002 -32 8066 -28
rect 10862 28 10926 32
rect 10862 -28 10866 28
rect 10866 -28 10922 28
rect 10922 -28 10926 28
rect 10862 -32 10926 -28
rect 10942 28 11006 32
rect 10942 -28 10946 28
rect 10946 -28 11002 28
rect 11002 -28 11006 28
rect 10942 -32 11006 -28
rect 11022 28 11086 32
rect 11022 -28 11026 28
rect 11026 -28 11082 28
rect 11082 -28 11086 28
rect 11022 -32 11086 -28
rect 11102 28 11166 32
rect 11102 -28 11106 28
rect 11106 -28 11162 28
rect 11162 -28 11166 28
rect 11102 -32 11166 -28
rect 13962 28 14026 32
rect 13962 -28 13966 28
rect 13966 -28 14022 28
rect 14022 -28 14026 28
rect 13962 -32 14026 -28
rect 14042 28 14106 32
rect 14042 -28 14046 28
rect 14046 -28 14102 28
rect 14102 -28 14106 28
rect 14042 -32 14106 -28
rect 14122 28 14186 32
rect 14122 -28 14126 28
rect 14126 -28 14182 28
rect 14182 -28 14186 28
rect 14122 -32 14186 -28
rect 14202 28 14266 32
rect 14202 -28 14206 28
rect 14206 -28 14262 28
rect 14262 -28 14266 28
rect 14202 -32 14266 -28
rect 17062 28 17126 32
rect 17062 -28 17066 28
rect 17066 -28 17122 28
rect 17122 -28 17126 28
rect 17062 -32 17126 -28
rect 17142 28 17206 32
rect 17142 -28 17146 28
rect 17146 -28 17202 28
rect 17202 -28 17206 28
rect 17142 -32 17206 -28
rect 17222 28 17286 32
rect 17222 -28 17226 28
rect 17226 -28 17282 28
rect 17282 -28 17286 28
rect 17222 -32 17286 -28
rect 17302 28 17366 32
rect 17302 -28 17306 28
rect 17306 -28 17362 28
rect 17362 -28 17366 28
rect 17302 -32 17366 -28
<< metal4 >>
rect 3104 10368 3424 10928
rect 3104 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3272 10368
rect 3336 10304 3352 10368
rect 3416 10304 3424 10368
rect 3104 10160 3424 10304
rect 3104 9924 3146 10160
rect 3382 9924 3424 10160
rect 3104 9280 3424 9924
rect 3104 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3272 9280
rect 3336 9216 3352 9280
rect 3416 9216 3424 9280
rect 3104 8192 3424 9216
rect 3104 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3272 8192
rect 3336 8128 3352 8192
rect 3416 8128 3424 8192
rect 3104 7104 3424 8128
rect 3104 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3272 7104
rect 3336 7040 3352 7104
rect 3416 7040 3424 7104
rect 3104 6780 3424 7040
rect 3104 6544 3146 6780
rect 3382 6544 3424 6780
rect 3104 6016 3424 6544
rect 3104 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3272 6016
rect 3336 5952 3352 6016
rect 3416 5952 3424 6016
rect 3104 4928 3424 5952
rect 3104 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3272 4928
rect 3336 4864 3352 4928
rect 3416 4864 3424 4928
rect 3104 3840 3424 4864
rect 3104 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3272 3840
rect 3336 3776 3352 3840
rect 3416 3776 3424 3840
rect 3104 3400 3424 3776
rect 3104 3164 3146 3400
rect 3382 3164 3424 3400
rect 3104 2752 3424 3164
rect 3104 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3272 2752
rect 3336 2688 3352 2752
rect 3416 2688 3424 2752
rect 3104 1664 3424 2688
rect 3104 1600 3112 1664
rect 3176 1600 3192 1664
rect 3256 1600 3272 1664
rect 3336 1600 3352 1664
rect 3416 1600 3424 1664
rect 3104 576 3424 1600
rect 3104 512 3112 576
rect 3176 512 3192 576
rect 3256 512 3272 576
rect 3336 512 3352 576
rect 3416 512 3424 576
rect 3104 -48 3424 512
rect 4654 10912 4974 10928
rect 4654 10848 4662 10912
rect 4726 10848 4742 10912
rect 4806 10848 4822 10912
rect 4886 10848 4902 10912
rect 4966 10848 4974 10912
rect 4654 9824 4974 10848
rect 4654 9760 4662 9824
rect 4726 9760 4742 9824
rect 4806 9760 4822 9824
rect 4886 9760 4902 9824
rect 4966 9760 4974 9824
rect 4654 8736 4974 9760
rect 4654 8672 4662 8736
rect 4726 8672 4742 8736
rect 4806 8672 4822 8736
rect 4886 8672 4902 8736
rect 4966 8672 4974 8736
rect 4654 8470 4974 8672
rect 4654 8234 4696 8470
rect 4932 8234 4974 8470
rect 4654 7648 4974 8234
rect 4654 7584 4662 7648
rect 4726 7584 4742 7648
rect 4806 7584 4822 7648
rect 4886 7584 4902 7648
rect 4966 7584 4974 7648
rect 4654 6560 4974 7584
rect 4654 6496 4662 6560
rect 4726 6496 4742 6560
rect 4806 6496 4822 6560
rect 4886 6496 4902 6560
rect 4966 6496 4974 6560
rect 4654 5472 4974 6496
rect 4654 5408 4662 5472
rect 4726 5408 4742 5472
rect 4806 5408 4822 5472
rect 4886 5408 4902 5472
rect 4966 5408 4974 5472
rect 4654 5090 4974 5408
rect 4654 4854 4696 5090
rect 4932 4854 4974 5090
rect 4654 4384 4974 4854
rect 4654 4320 4662 4384
rect 4726 4320 4742 4384
rect 4806 4320 4822 4384
rect 4886 4320 4902 4384
rect 4966 4320 4974 4384
rect 4654 3296 4974 4320
rect 4654 3232 4662 3296
rect 4726 3232 4742 3296
rect 4806 3232 4822 3296
rect 4886 3232 4902 3296
rect 4966 3232 4974 3296
rect 4654 2208 4974 3232
rect 4654 2144 4662 2208
rect 4726 2144 4742 2208
rect 4806 2144 4822 2208
rect 4886 2144 4902 2208
rect 4966 2144 4974 2208
rect 4654 1120 4974 2144
rect 4654 1056 4662 1120
rect 4726 1056 4742 1120
rect 4806 1056 4822 1120
rect 4886 1056 4902 1120
rect 4966 1056 4974 1120
rect 4654 32 4974 1056
rect 4654 -32 4662 32
rect 4726 -32 4742 32
rect 4806 -32 4822 32
rect 4886 -32 4902 32
rect 4966 -32 4974 32
rect 4654 -48 4974 -32
rect 6204 10368 6524 10928
rect 6204 10304 6212 10368
rect 6276 10304 6292 10368
rect 6356 10304 6372 10368
rect 6436 10304 6452 10368
rect 6516 10304 6524 10368
rect 6204 10160 6524 10304
rect 6204 9924 6246 10160
rect 6482 9924 6524 10160
rect 6204 9280 6524 9924
rect 6204 9216 6212 9280
rect 6276 9216 6292 9280
rect 6356 9216 6372 9280
rect 6436 9216 6452 9280
rect 6516 9216 6524 9280
rect 6204 8192 6524 9216
rect 6204 8128 6212 8192
rect 6276 8128 6292 8192
rect 6356 8128 6372 8192
rect 6436 8128 6452 8192
rect 6516 8128 6524 8192
rect 6204 7104 6524 8128
rect 6204 7040 6212 7104
rect 6276 7040 6292 7104
rect 6356 7040 6372 7104
rect 6436 7040 6452 7104
rect 6516 7040 6524 7104
rect 6204 6780 6524 7040
rect 6204 6544 6246 6780
rect 6482 6544 6524 6780
rect 6204 6016 6524 6544
rect 6204 5952 6212 6016
rect 6276 5952 6292 6016
rect 6356 5952 6372 6016
rect 6436 5952 6452 6016
rect 6516 5952 6524 6016
rect 6204 4928 6524 5952
rect 6204 4864 6212 4928
rect 6276 4864 6292 4928
rect 6356 4864 6372 4928
rect 6436 4864 6452 4928
rect 6516 4864 6524 4928
rect 6204 3840 6524 4864
rect 6204 3776 6212 3840
rect 6276 3776 6292 3840
rect 6356 3776 6372 3840
rect 6436 3776 6452 3840
rect 6516 3776 6524 3840
rect 6204 3400 6524 3776
rect 6204 3164 6246 3400
rect 6482 3164 6524 3400
rect 6204 2752 6524 3164
rect 6204 2688 6212 2752
rect 6276 2688 6292 2752
rect 6356 2688 6372 2752
rect 6436 2688 6452 2752
rect 6516 2688 6524 2752
rect 6204 1664 6524 2688
rect 6204 1600 6212 1664
rect 6276 1600 6292 1664
rect 6356 1600 6372 1664
rect 6436 1600 6452 1664
rect 6516 1600 6524 1664
rect 6204 576 6524 1600
rect 6204 512 6212 576
rect 6276 512 6292 576
rect 6356 512 6372 576
rect 6436 512 6452 576
rect 6516 512 6524 576
rect 6204 -48 6524 512
rect 7754 10912 8074 10928
rect 7754 10848 7762 10912
rect 7826 10848 7842 10912
rect 7906 10848 7922 10912
rect 7986 10848 8002 10912
rect 8066 10848 8074 10912
rect 7754 9824 8074 10848
rect 7754 9760 7762 9824
rect 7826 9760 7842 9824
rect 7906 9760 7922 9824
rect 7986 9760 8002 9824
rect 8066 9760 8074 9824
rect 7754 8736 8074 9760
rect 7754 8672 7762 8736
rect 7826 8672 7842 8736
rect 7906 8672 7922 8736
rect 7986 8672 8002 8736
rect 8066 8672 8074 8736
rect 7754 8470 8074 8672
rect 7754 8234 7796 8470
rect 8032 8234 8074 8470
rect 7754 7648 8074 8234
rect 7754 7584 7762 7648
rect 7826 7584 7842 7648
rect 7906 7584 7922 7648
rect 7986 7584 8002 7648
rect 8066 7584 8074 7648
rect 7754 6560 8074 7584
rect 7754 6496 7762 6560
rect 7826 6496 7842 6560
rect 7906 6496 7922 6560
rect 7986 6496 8002 6560
rect 8066 6496 8074 6560
rect 7754 5472 8074 6496
rect 7754 5408 7762 5472
rect 7826 5408 7842 5472
rect 7906 5408 7922 5472
rect 7986 5408 8002 5472
rect 8066 5408 8074 5472
rect 7754 5090 8074 5408
rect 7754 4854 7796 5090
rect 8032 4854 8074 5090
rect 7754 4384 8074 4854
rect 7754 4320 7762 4384
rect 7826 4320 7842 4384
rect 7906 4320 7922 4384
rect 7986 4320 8002 4384
rect 8066 4320 8074 4384
rect 7754 3296 8074 4320
rect 7754 3232 7762 3296
rect 7826 3232 7842 3296
rect 7906 3232 7922 3296
rect 7986 3232 8002 3296
rect 8066 3232 8074 3296
rect 7754 2208 8074 3232
rect 7754 2144 7762 2208
rect 7826 2144 7842 2208
rect 7906 2144 7922 2208
rect 7986 2144 8002 2208
rect 8066 2144 8074 2208
rect 7754 1120 8074 2144
rect 7754 1056 7762 1120
rect 7826 1056 7842 1120
rect 7906 1056 7922 1120
rect 7986 1056 8002 1120
rect 8066 1056 8074 1120
rect 7754 32 8074 1056
rect 7754 -32 7762 32
rect 7826 -32 7842 32
rect 7906 -32 7922 32
rect 7986 -32 8002 32
rect 8066 -32 8074 32
rect 7754 -48 8074 -32
rect 9304 10368 9624 10928
rect 9304 10304 9312 10368
rect 9376 10304 9392 10368
rect 9456 10304 9472 10368
rect 9536 10304 9552 10368
rect 9616 10304 9624 10368
rect 9304 10160 9624 10304
rect 9304 9924 9346 10160
rect 9582 9924 9624 10160
rect 9304 9280 9624 9924
rect 9304 9216 9312 9280
rect 9376 9216 9392 9280
rect 9456 9216 9472 9280
rect 9536 9216 9552 9280
rect 9616 9216 9624 9280
rect 9304 8192 9624 9216
rect 9304 8128 9312 8192
rect 9376 8128 9392 8192
rect 9456 8128 9472 8192
rect 9536 8128 9552 8192
rect 9616 8128 9624 8192
rect 9304 7104 9624 8128
rect 9304 7040 9312 7104
rect 9376 7040 9392 7104
rect 9456 7040 9472 7104
rect 9536 7040 9552 7104
rect 9616 7040 9624 7104
rect 9304 6780 9624 7040
rect 9304 6544 9346 6780
rect 9582 6544 9624 6780
rect 9304 6016 9624 6544
rect 9304 5952 9312 6016
rect 9376 5952 9392 6016
rect 9456 5952 9472 6016
rect 9536 5952 9552 6016
rect 9616 5952 9624 6016
rect 9304 4928 9624 5952
rect 9304 4864 9312 4928
rect 9376 4864 9392 4928
rect 9456 4864 9472 4928
rect 9536 4864 9552 4928
rect 9616 4864 9624 4928
rect 9304 3840 9624 4864
rect 9304 3776 9312 3840
rect 9376 3776 9392 3840
rect 9456 3776 9472 3840
rect 9536 3776 9552 3840
rect 9616 3776 9624 3840
rect 9304 3400 9624 3776
rect 9304 3164 9346 3400
rect 9582 3164 9624 3400
rect 9304 2752 9624 3164
rect 9304 2688 9312 2752
rect 9376 2688 9392 2752
rect 9456 2688 9472 2752
rect 9536 2688 9552 2752
rect 9616 2688 9624 2752
rect 9304 1664 9624 2688
rect 9304 1600 9312 1664
rect 9376 1600 9392 1664
rect 9456 1600 9472 1664
rect 9536 1600 9552 1664
rect 9616 1600 9624 1664
rect 9304 576 9624 1600
rect 9304 512 9312 576
rect 9376 512 9392 576
rect 9456 512 9472 576
rect 9536 512 9552 576
rect 9616 512 9624 576
rect 9304 -48 9624 512
rect 10854 10912 11174 10928
rect 10854 10848 10862 10912
rect 10926 10848 10942 10912
rect 11006 10848 11022 10912
rect 11086 10848 11102 10912
rect 11166 10848 11174 10912
rect 10854 9824 11174 10848
rect 10854 9760 10862 9824
rect 10926 9760 10942 9824
rect 11006 9760 11022 9824
rect 11086 9760 11102 9824
rect 11166 9760 11174 9824
rect 10854 8736 11174 9760
rect 10854 8672 10862 8736
rect 10926 8672 10942 8736
rect 11006 8672 11022 8736
rect 11086 8672 11102 8736
rect 11166 8672 11174 8736
rect 10854 8470 11174 8672
rect 10854 8234 10896 8470
rect 11132 8234 11174 8470
rect 10854 7648 11174 8234
rect 10854 7584 10862 7648
rect 10926 7584 10942 7648
rect 11006 7584 11022 7648
rect 11086 7584 11102 7648
rect 11166 7584 11174 7648
rect 10854 6560 11174 7584
rect 10854 6496 10862 6560
rect 10926 6496 10942 6560
rect 11006 6496 11022 6560
rect 11086 6496 11102 6560
rect 11166 6496 11174 6560
rect 10854 5472 11174 6496
rect 10854 5408 10862 5472
rect 10926 5408 10942 5472
rect 11006 5408 11022 5472
rect 11086 5408 11102 5472
rect 11166 5408 11174 5472
rect 10854 5090 11174 5408
rect 10854 4854 10896 5090
rect 11132 4854 11174 5090
rect 10854 4384 11174 4854
rect 10854 4320 10862 4384
rect 10926 4320 10942 4384
rect 11006 4320 11022 4384
rect 11086 4320 11102 4384
rect 11166 4320 11174 4384
rect 10854 3296 11174 4320
rect 10854 3232 10862 3296
rect 10926 3232 10942 3296
rect 11006 3232 11022 3296
rect 11086 3232 11102 3296
rect 11166 3232 11174 3296
rect 10854 2208 11174 3232
rect 10854 2144 10862 2208
rect 10926 2144 10942 2208
rect 11006 2144 11022 2208
rect 11086 2144 11102 2208
rect 11166 2144 11174 2208
rect 10854 1120 11174 2144
rect 10854 1056 10862 1120
rect 10926 1056 10942 1120
rect 11006 1056 11022 1120
rect 11086 1056 11102 1120
rect 11166 1056 11174 1120
rect 10854 32 11174 1056
rect 10854 -32 10862 32
rect 10926 -32 10942 32
rect 11006 -32 11022 32
rect 11086 -32 11102 32
rect 11166 -32 11174 32
rect 10854 -48 11174 -32
rect 12404 10368 12724 10928
rect 12404 10304 12412 10368
rect 12476 10304 12492 10368
rect 12556 10304 12572 10368
rect 12636 10304 12652 10368
rect 12716 10304 12724 10368
rect 12404 10160 12724 10304
rect 12404 9924 12446 10160
rect 12682 9924 12724 10160
rect 12404 9280 12724 9924
rect 12404 9216 12412 9280
rect 12476 9216 12492 9280
rect 12556 9216 12572 9280
rect 12636 9216 12652 9280
rect 12716 9216 12724 9280
rect 12404 8192 12724 9216
rect 12404 8128 12412 8192
rect 12476 8128 12492 8192
rect 12556 8128 12572 8192
rect 12636 8128 12652 8192
rect 12716 8128 12724 8192
rect 12404 7104 12724 8128
rect 12404 7040 12412 7104
rect 12476 7040 12492 7104
rect 12556 7040 12572 7104
rect 12636 7040 12652 7104
rect 12716 7040 12724 7104
rect 12404 6780 12724 7040
rect 12404 6544 12446 6780
rect 12682 6544 12724 6780
rect 12404 6016 12724 6544
rect 12404 5952 12412 6016
rect 12476 5952 12492 6016
rect 12556 5952 12572 6016
rect 12636 5952 12652 6016
rect 12716 5952 12724 6016
rect 12404 4928 12724 5952
rect 12404 4864 12412 4928
rect 12476 4864 12492 4928
rect 12556 4864 12572 4928
rect 12636 4864 12652 4928
rect 12716 4864 12724 4928
rect 12404 3840 12724 4864
rect 12404 3776 12412 3840
rect 12476 3776 12492 3840
rect 12556 3776 12572 3840
rect 12636 3776 12652 3840
rect 12716 3776 12724 3840
rect 12404 3400 12724 3776
rect 12404 3164 12446 3400
rect 12682 3164 12724 3400
rect 12404 2752 12724 3164
rect 12404 2688 12412 2752
rect 12476 2688 12492 2752
rect 12556 2688 12572 2752
rect 12636 2688 12652 2752
rect 12716 2688 12724 2752
rect 12404 1664 12724 2688
rect 12404 1600 12412 1664
rect 12476 1600 12492 1664
rect 12556 1600 12572 1664
rect 12636 1600 12652 1664
rect 12716 1600 12724 1664
rect 12404 576 12724 1600
rect 12404 512 12412 576
rect 12476 512 12492 576
rect 12556 512 12572 576
rect 12636 512 12652 576
rect 12716 512 12724 576
rect 12404 -48 12724 512
rect 13954 10912 14274 10928
rect 13954 10848 13962 10912
rect 14026 10848 14042 10912
rect 14106 10848 14122 10912
rect 14186 10848 14202 10912
rect 14266 10848 14274 10912
rect 13954 9824 14274 10848
rect 13954 9760 13962 9824
rect 14026 9760 14042 9824
rect 14106 9760 14122 9824
rect 14186 9760 14202 9824
rect 14266 9760 14274 9824
rect 13954 8736 14274 9760
rect 13954 8672 13962 8736
rect 14026 8672 14042 8736
rect 14106 8672 14122 8736
rect 14186 8672 14202 8736
rect 14266 8672 14274 8736
rect 13954 8470 14274 8672
rect 13954 8234 13996 8470
rect 14232 8234 14274 8470
rect 13954 7648 14274 8234
rect 13954 7584 13962 7648
rect 14026 7584 14042 7648
rect 14106 7584 14122 7648
rect 14186 7584 14202 7648
rect 14266 7584 14274 7648
rect 13954 6560 14274 7584
rect 13954 6496 13962 6560
rect 14026 6496 14042 6560
rect 14106 6496 14122 6560
rect 14186 6496 14202 6560
rect 14266 6496 14274 6560
rect 13954 5472 14274 6496
rect 13954 5408 13962 5472
rect 14026 5408 14042 5472
rect 14106 5408 14122 5472
rect 14186 5408 14202 5472
rect 14266 5408 14274 5472
rect 13954 5090 14274 5408
rect 13954 4854 13996 5090
rect 14232 4854 14274 5090
rect 13954 4384 14274 4854
rect 13954 4320 13962 4384
rect 14026 4320 14042 4384
rect 14106 4320 14122 4384
rect 14186 4320 14202 4384
rect 14266 4320 14274 4384
rect 13954 3296 14274 4320
rect 13954 3232 13962 3296
rect 14026 3232 14042 3296
rect 14106 3232 14122 3296
rect 14186 3232 14202 3296
rect 14266 3232 14274 3296
rect 13954 2208 14274 3232
rect 13954 2144 13962 2208
rect 14026 2144 14042 2208
rect 14106 2144 14122 2208
rect 14186 2144 14202 2208
rect 14266 2144 14274 2208
rect 13954 1120 14274 2144
rect 13954 1056 13962 1120
rect 14026 1056 14042 1120
rect 14106 1056 14122 1120
rect 14186 1056 14202 1120
rect 14266 1056 14274 1120
rect 13954 32 14274 1056
rect 13954 -32 13962 32
rect 14026 -32 14042 32
rect 14106 -32 14122 32
rect 14186 -32 14202 32
rect 14266 -32 14274 32
rect 13954 -48 14274 -32
rect 15504 10368 15824 10928
rect 15504 10304 15512 10368
rect 15576 10304 15592 10368
rect 15656 10304 15672 10368
rect 15736 10304 15752 10368
rect 15816 10304 15824 10368
rect 15504 10160 15824 10304
rect 15504 9924 15546 10160
rect 15782 9924 15824 10160
rect 15504 9280 15824 9924
rect 15504 9216 15512 9280
rect 15576 9216 15592 9280
rect 15656 9216 15672 9280
rect 15736 9216 15752 9280
rect 15816 9216 15824 9280
rect 15504 8192 15824 9216
rect 15504 8128 15512 8192
rect 15576 8128 15592 8192
rect 15656 8128 15672 8192
rect 15736 8128 15752 8192
rect 15816 8128 15824 8192
rect 15504 7104 15824 8128
rect 15504 7040 15512 7104
rect 15576 7040 15592 7104
rect 15656 7040 15672 7104
rect 15736 7040 15752 7104
rect 15816 7040 15824 7104
rect 15504 6780 15824 7040
rect 15504 6544 15546 6780
rect 15782 6544 15824 6780
rect 15504 6016 15824 6544
rect 15504 5952 15512 6016
rect 15576 5952 15592 6016
rect 15656 5952 15672 6016
rect 15736 5952 15752 6016
rect 15816 5952 15824 6016
rect 15504 4928 15824 5952
rect 15504 4864 15512 4928
rect 15576 4864 15592 4928
rect 15656 4864 15672 4928
rect 15736 4864 15752 4928
rect 15816 4864 15824 4928
rect 15504 3840 15824 4864
rect 15504 3776 15512 3840
rect 15576 3776 15592 3840
rect 15656 3776 15672 3840
rect 15736 3776 15752 3840
rect 15816 3776 15824 3840
rect 15504 3400 15824 3776
rect 15504 3164 15546 3400
rect 15782 3164 15824 3400
rect 15504 2752 15824 3164
rect 15504 2688 15512 2752
rect 15576 2688 15592 2752
rect 15656 2688 15672 2752
rect 15736 2688 15752 2752
rect 15816 2688 15824 2752
rect 15504 1664 15824 2688
rect 15504 1600 15512 1664
rect 15576 1600 15592 1664
rect 15656 1600 15672 1664
rect 15736 1600 15752 1664
rect 15816 1600 15824 1664
rect 15504 576 15824 1600
rect 15504 512 15512 576
rect 15576 512 15592 576
rect 15656 512 15672 576
rect 15736 512 15752 576
rect 15816 512 15824 576
rect 15504 -48 15824 512
rect 17054 10912 17374 10928
rect 17054 10848 17062 10912
rect 17126 10848 17142 10912
rect 17206 10848 17222 10912
rect 17286 10848 17302 10912
rect 17366 10848 17374 10912
rect 17054 9824 17374 10848
rect 17054 9760 17062 9824
rect 17126 9760 17142 9824
rect 17206 9760 17222 9824
rect 17286 9760 17302 9824
rect 17366 9760 17374 9824
rect 17054 8736 17374 9760
rect 17054 8672 17062 8736
rect 17126 8672 17142 8736
rect 17206 8672 17222 8736
rect 17286 8672 17302 8736
rect 17366 8672 17374 8736
rect 17054 8470 17374 8672
rect 17054 8234 17096 8470
rect 17332 8234 17374 8470
rect 17054 7648 17374 8234
rect 17054 7584 17062 7648
rect 17126 7584 17142 7648
rect 17206 7584 17222 7648
rect 17286 7584 17302 7648
rect 17366 7584 17374 7648
rect 17054 6560 17374 7584
rect 17054 6496 17062 6560
rect 17126 6496 17142 6560
rect 17206 6496 17222 6560
rect 17286 6496 17302 6560
rect 17366 6496 17374 6560
rect 17054 5472 17374 6496
rect 17054 5408 17062 5472
rect 17126 5408 17142 5472
rect 17206 5408 17222 5472
rect 17286 5408 17302 5472
rect 17366 5408 17374 5472
rect 17054 5090 17374 5408
rect 17054 4854 17096 5090
rect 17332 4854 17374 5090
rect 17054 4384 17374 4854
rect 17054 4320 17062 4384
rect 17126 4320 17142 4384
rect 17206 4320 17222 4384
rect 17286 4320 17302 4384
rect 17366 4320 17374 4384
rect 17054 3296 17374 4320
rect 17054 3232 17062 3296
rect 17126 3232 17142 3296
rect 17206 3232 17222 3296
rect 17286 3232 17302 3296
rect 17366 3232 17374 3296
rect 17054 2208 17374 3232
rect 17054 2144 17062 2208
rect 17126 2144 17142 2208
rect 17206 2144 17222 2208
rect 17286 2144 17302 2208
rect 17366 2144 17374 2208
rect 17054 1120 17374 2144
rect 17054 1056 17062 1120
rect 17126 1056 17142 1120
rect 17206 1056 17222 1120
rect 17286 1056 17302 1120
rect 17366 1056 17374 1120
rect 17054 32 17374 1056
rect 17054 -32 17062 32
rect 17126 -32 17142 32
rect 17206 -32 17222 32
rect 17286 -32 17302 32
rect 17366 -32 17374 32
rect 17054 -48 17374 -32
<< via4 >>
rect 3146 9924 3382 10160
rect 3146 6544 3382 6780
rect 3146 3164 3382 3400
rect 4696 8234 4932 8470
rect 4696 4854 4932 5090
rect 6246 9924 6482 10160
rect 6246 6544 6482 6780
rect 6246 3164 6482 3400
rect 7796 8234 8032 8470
rect 7796 4854 8032 5090
rect 9346 9924 9582 10160
rect 9346 6544 9582 6780
rect 9346 3164 9582 3400
rect 10896 8234 11132 8470
rect 10896 4854 11132 5090
rect 12446 9924 12682 10160
rect 12446 6544 12682 6780
rect 12446 3164 12682 3400
rect 13996 8234 14232 8470
rect 13996 4854 14232 5090
rect 15546 9924 15782 10160
rect 15546 6544 15782 6780
rect 15546 3164 15782 3400
rect 17096 8234 17332 8470
rect 17096 4854 17332 5090
<< metal5 >>
rect 0 10160 18860 10202
rect 0 9924 3146 10160
rect 3382 9924 6246 10160
rect 6482 9924 9346 10160
rect 9582 9924 12446 10160
rect 12682 9924 15546 10160
rect 15782 9924 18860 10160
rect 0 9882 18860 9924
rect 0 8470 18860 8512
rect 0 8234 4696 8470
rect 4932 8234 7796 8470
rect 8032 8234 10896 8470
rect 11132 8234 13996 8470
rect 14232 8234 17096 8470
rect 17332 8234 18860 8470
rect 0 8192 18860 8234
rect 0 6780 18860 6822
rect 0 6544 3146 6780
rect 3382 6544 6246 6780
rect 6482 6544 9346 6780
rect 9582 6544 12446 6780
rect 12682 6544 15546 6780
rect 15782 6544 18860 6780
rect 0 6502 18860 6544
rect 0 5090 18860 5132
rect 0 4854 4696 5090
rect 4932 4854 7796 5090
rect 8032 4854 10896 5090
rect 11132 4854 13996 5090
rect 14232 4854 17096 5090
rect 17332 4854 18860 5090
rect 0 4812 18860 4854
rect 0 3400 18860 3442
rect 0 3164 3146 3400
rect 3382 3164 6246 3400
rect 6482 3164 9346 3400
rect 9582 3164 12446 3400
rect 12682 3164 15546 3400
rect 15782 3164 18860 3400
rect 0 3122 18860 3164
use sky130_fd_sc_hd__decap_3  PHY_2 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 0 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1636915332
transform 1 0 0 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 276 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1012 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1196 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_23 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2116 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 1636915332
transform 1 0 1380 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__449__SET_B OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 2392 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 276 0 -1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_14
timestamp 1636915332
transform 1 0 1288 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_27
timestamp 1636915332
transform 1 0 2484 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_40
timestamp 1636915332
transform 1 0 3680 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1636915332
transform 1 0 2392 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1636915332
transform 1 0 3588 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1636915332
transform 1 0 2392 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _300_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4784 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _449_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2484 0 -1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__o2bb2ai_1  _297_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5980 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _290_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5152 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1636915332
transform 1 0 4784 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1636915332
transform 1 0 4784 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1636915332
transform 1 0 5244 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 4876 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__450__RESET_B
timestamp 1636915332
transform -1 0 5336 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _296_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 6072 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1636915332
transform 1 0 5980 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69
timestamp 1636915332
transform 1 0 6348 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtn_1  _450_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5336 0 -1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__nor2_1  _309_
timestamp 1636915332
transform -1 0 7820 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _303_
timestamp 1636915332
transform 1 0 7268 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1636915332
transform 1 0 7176 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1636915332
transform 1 0 7176 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_85
timestamp 1636915332
transform 1 0 7820 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77
timestamp 1636915332
transform 1 0 7084 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _312_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9476 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_2  _310_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8004 0 -1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_1  _306_
timestamp 1636915332
transform -1 0 9384 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1636915332
transform 1 0 8372 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_97
timestamp 1636915332
transform 1 0 8924 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98
timestamp 1636915332
transform 1 0 9016 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8464 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_79
timestamp 1636915332
transform 1 0 7268 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__o21bai_1  _311_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 9660 0 -1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _304_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 10488 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1636915332
transform 1 0 9568 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1636915332
transform 1 0 9568 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_103
timestamp 1636915332
transform 1 0 9476 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__310__B1
timestamp 1636915332
transform 1 0 9384 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1636915332
transform 1 0 10764 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_122
timestamp 1636915332
transform 1 0 11224 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_114
timestamp 1636915332
transform 1 0 10488 0 -1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_118
timestamp 1636915332
transform 1 0 10856 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_105
timestamp 1636915332
transform 1 0 9660 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_1  _357_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12328 0 -1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _332_
timestamp 1636915332
transform -1 0 12420 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _329_
timestamp 1636915332
transform 1 0 12052 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _328_
timestamp 1636915332
transform 1 0 11500 0 -1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1636915332
transform 1 0 11960 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1636915332
transform 1 0 11960 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_129
timestamp 1636915332
transform 1 0 11868 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_135
timestamp 1636915332
transform 1 0 12420 0 1 0
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _356_
timestamp 1636915332
transform 1 0 13524 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _307_
timestamp 1636915332
transform -1 0 13524 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1636915332
transform 1 0 13156 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_4  _305_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12972 0 -1 1088
box -38 -48 1418 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1636915332
transform 1 0 14352 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1636915332
transform 1 0 14352 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_157
timestamp 1636915332
transform 1 0 14444 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_150
timestamp 1636915332
transform 1 0 13800 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__440__RESET_B
timestamp 1636915332
transform -1 0 14720 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _333_
timestamp 1636915332
transform 1 0 15824 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1636915332
transform 1 0 15548 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__385__A1
timestamp 1636915332
transform -1 0 15824 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtn_1  _440_
timestamp 1636915332
transform 1 0 14720 0 -1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_12  FILLER_0_157
timestamp 1636915332
transform 1 0 14444 0 1 0
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_1  _355_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 16836 0 1 0
box -38 -48 682 592
use sky130_fd_sc_hd__inv_4  _330__6 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 16560 0 1 0
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1636915332
transform 1 0 16744 0 -1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1636915332
transform 1 0 16744 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_183
timestamp 1636915332
transform 1 0 16836 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_180
timestamp 1636915332
transform 1 0 16560 0 1 0
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__441__SET_B
timestamp 1636915332
transform -1 0 16744 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _381_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 17020 0 -1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_190
timestamp 1636915332
transform 1 0 17480 0 1 0
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1636915332
transform 1 0 17940 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_194
timestamp 1636915332
transform 1 0 17848 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_196
timestamp 1636915332
transform 1 0 18032 0 1 0
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_194
timestamp 1636915332
transform 1 0 17848 0 1 0
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1636915332
transform -1 0 18308 0 -1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1636915332
transform -1 0 18860 0 1 0
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1636915332
transform -1 0 18860 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 18308 0 -1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_11
timestamp 1636915332
transform 1 0 1012 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1636915332
transform 1 0 1288 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_18
timestamp 1636915332
transform 1 0 1656 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1636915332
transform 1 0 276 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1636915332
transform 1 0 0 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1636915332
transform 1 0 1196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtn_1  _448_
timestamp 1636915332
transform 1 0 1748 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_2_48
timestamp 1636915332
transform 1 0 4416 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1636915332
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _295_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5152 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _301_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4416 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_66
timestamp 1636915332
transform 1 0 6072 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1636915332
transform 1 0 5980 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_2  _278_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 7452 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _292_
timestamp 1636915332
transform 1 0 5152 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _294_
timestamp 1636915332
transform -1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__B1
timestamp 1636915332
transform 1 0 8096 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_90
timestamp 1636915332
transform 1 0 8280 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1636915332
transform 1 0 8372 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _447_
timestamp 1636915332
transform 1 0 8464 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer5 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 7452 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__RESET_B
timestamp 1636915332
transform 1 0 10580 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_113
timestamp 1636915332
transform 1 0 10396 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1636915332
transform 1 0 10764 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtn_1  _442_
timestamp 1636915332
transform -1 0 12696 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_2_138
timestamp 1636915332
transform 1 0 12696 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_142
timestamp 1636915332
transform 1 0 13064 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_144
timestamp 1636915332
transform 1 0 13248 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_148
timestamp 1636915332
transform 1 0 13616 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1636915332
transform 1 0 13156 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _308_
timestamp 1636915332
transform -1 0 13616 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_156
timestamp 1636915332
transform 1 0 14352 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_170
timestamp 1636915332
transform 1 0 15640 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1636915332
transform 1 0 15548 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _331_
timestamp 1636915332
transform -1 0 16008 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _334_
timestamp 1636915332
transform 1 0 14444 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _385_
timestamp 1636915332
transform 1 0 14720 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_2_196
timestamp 1636915332
transform 1 0 18032 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1636915332
transform 1 0 17940 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_2  _441_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 16008 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1636915332
transform -1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__446__RESET_B
timestamp 1636915332
transform 1 0 2116 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1636915332
transform 1 0 0 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _446_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 276 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__448__RESET_B
timestamp 1636915332
transform 1 0 3588 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_25
timestamp 1636915332
transform 1 0 2300 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_41
timestamp 1636915332
transform 1 0 3772 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1636915332
transform 1 0 2392 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _291_
timestamp 1636915332
transform -1 0 4784 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _298__4
timestamp 1636915332
transform -1 0 3588 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _299_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3956 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _314_
timestamp 1636915332
transform -1 0 3128 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1636915332
transform 1 0 4876 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1636915332
transform 1 0 5704 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1636915332
transform 1 0 4784 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _293_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 5152 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _397_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 7176 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__447__SET_B
timestamp 1636915332
transform 1 0 8280 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_84
timestamp 1636915332
transform 1 0 7728 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_92
timestamp 1636915332
transform 1 0 8464 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1636915332
transform 1 0 7176 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _282_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9384 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _283_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 7728 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  _302__5
timestamp 1636915332
transform -1 0 9016 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__fill_2  FILLER_3_102
timestamp 1636915332
transform 1 0 9384 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_111
timestamp 1636915332
transform 1 0 10212 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_117
timestamp 1636915332
transform 1 0 10764 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1636915332
transform 1 0 9568 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1636915332
transform -1 0 9936 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _326_
timestamp 1636915332
transform 1 0 9936 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _349_
timestamp 1636915332
transform 1 0 10856 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_3_125
timestamp 1636915332
transform 1 0 11500 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_131
timestamp 1636915332
transform 1 0 12052 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1636915332
transform 1 0 11960 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _327_
timestamp 1636915332
transform -1 0 11960 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1636915332
transform 1 0 13064 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _407_
timestamp 1636915332
transform 1 0 12236 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__427__RESET_B
timestamp 1636915332
transform 1 0 13892 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_157
timestamp 1636915332
transform 1 0 14444 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1636915332
transform 1 0 14352 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _335_
timestamp 1636915332
transform -1 0 14352 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _336_
timestamp 1636915332
transform -1 0 14904 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _427_
timestamp 1636915332
transform 1 0 14904 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_3_192
timestamp 1636915332
transform 1 0 17664 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1636915332
transform 1 0 16744 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _374_
timestamp 1636915332
transform -1 0 18400 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _382_
timestamp 1636915332
transform 1 0 16836 0 -1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1636915332
transform 1 0 18400 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1636915332
transform -1 0 18860 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1636915332
transform 1 0 1012 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_14
timestamp 1636915332
transform 1 0 1288 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1636915332
transform 1 0 276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1636915332
transform 1 0 644 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1636915332
transform 1 0 0 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1636915332
transform 1 0 1196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _315_
timestamp 1636915332
transform 1 0 1564 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _316_
timestamp 1636915332
transform 1 0 736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__313__A
timestamp 1636915332
transform 1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__315__S
timestamp 1636915332
transform 1 0 3220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__451__RESET_B
timestamp 1636915332
transform 1 0 3864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_37
timestamp 1636915332
transform 1 0 3404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_40
timestamp 1636915332
transform 1 0 3680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1636915332
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__nor3_1  _313_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _337_
timestamp 1636915332
transform 1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _451_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5980 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_4_70
timestamp 1636915332
transform 1 0 6440 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1636915332
transform 1 0 5980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  rebuffer6 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 6440 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__454__SET_B
timestamp 1636915332
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_80
timestamp 1636915332
transform 1 0 7360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_88
timestamp 1636915332
transform 1 0 8096 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1636915332
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _277_
timestamp 1636915332
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _279_
timestamp 1636915332
transform -1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _454_
timestamp 1636915332
transform 1 0 8832 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1636915332
transform 1 0 10764 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1636915332
transform 1 0 11408 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _280_
timestamp 1636915332
transform -1 0 11408 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_127
timestamp 1636915332
transform 1 0 11684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_139
timestamp 1636915332
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1636915332
transform 1 0 13248 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1636915332
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__386__A1
timestamp 1636915332
transform 1 0 15364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__430__RESET_B
timestamp 1636915332
transform 1 0 15640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_156
timestamp 1636915332
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1636915332
transform 1 0 15548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp 1636915332
transform 1 0 14536 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _430_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 15824 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1636915332
transform -1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_196
timestamp 1636915332
transform 1 0 18032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1636915332
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1636915332
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1636915332
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__445__RESET_B
timestamp 1636915332
transform 1 0 2116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1636915332
transform 1 0 0 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _445_
timestamp 1636915332
transform 1 0 276 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_5_25
timestamp 1636915332
transform 1 0 2300 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_27
timestamp 1636915332
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_44
timestamp 1636915332
transform 1 0 4048 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1636915332
transform 1 0 2392 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _363_
timestamp 1636915332
transform 1 0 2576 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _403_
timestamp 1636915332
transform 1 0 3220 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_53
timestamp 1636915332
transform 1 0 4876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1636915332
transform 1 0 4784 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _288_
timestamp 1636915332
transform 1 0 5244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _289_
timestamp 1636915332
transform 1 0 5612 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _405_
timestamp 1636915332
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__404__A1
timestamp 1636915332
transform 1 0 8464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_94
timestamp 1636915332
transform 1 0 8648 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_99
timestamp 1636915332
transform 1 0 9108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1636915332
transform 1 0 7176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _272_
timestamp 1636915332
transform 1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _358_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1636915332
transform 1 0 7268 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_103
timestamp 1636915332
transform 1 0 9476 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_112
timestamp 1636915332
transform 1 0 10304 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_119
timestamp 1636915332
transform 1 0 10948 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1636915332
transform 1 0 9568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__nand3b_1  _275_
timestamp 1636915332
transform -1 0 10948 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  _345_
timestamp 1636915332
transform 1 0 9660 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_2  _351_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 11960 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__443__RESET_B
timestamp 1636915332
transform 1 0 12052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1636915332
transform 1 0 11960 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _443_
timestamp 1636915332
transform 1 0 12236 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1636915332
transform 1 0 14352 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _320_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 16468 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _414_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 14444 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__414__D
timestamp 1636915332
transform 1 0 16468 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_181
timestamp 1636915332
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_183
timestamp 1636915332
transform 1 0 16836 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_195
timestamp 1636915332
transform 1 0 17940 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1636915332
transform 1 0 16744 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_201
timestamp 1636915332
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1636915332
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _318_
timestamp 1636915332
transform 1 0 828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1636915332
transform 1 0 0 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1636915332
transform 1 0 0 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1636915332
transform 1 0 276 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_12
timestamp 1636915332
transform 1 0 1104 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _317_
timestamp 1636915332
transform 1 0 1564 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1636915332
transform 1 0 1196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_14
timestamp 1636915332
transform 1 0 1288 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__444__SET_B
timestamp 1636915332
transform 1 0 2208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_2  _444_
timestamp 1636915332
transform 1 0 276 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1636915332
transform 1 0 3036 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _364_
timestamp 1636915332
transform -1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _338_
timestamp 1636915332
transform 1 0 2484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1636915332
transform 1 0 2392 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_32
timestamp 1636915332
transform 1 0 2944 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_28
timestamp 1636915332
transform 1 0 2576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__338__A_N
timestamp 1636915332
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__317__S
timestamp 1636915332
transform 1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__clkinv_2  _362_
timestamp 1636915332
transform 1 0 3864 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1636915332
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_46
timestamp 1636915332
transform 1 0 4232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_38
timestamp 1636915332
transform 1 0 3496 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_40
timestamp 1636915332
transform 1 0 3680 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_1  _286_
timestamp 1636915332
transform 1 0 5612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1636915332
transform 1 0 4784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_60
timestamp 1636915332
transform 1 0 5520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_52
timestamp 1636915332
transform 1 0 4784 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__452__SET_B
timestamp 1636915332
transform 1 0 4600 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1636915332
transform 1 0 6256 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1636915332
transform 1 0 5980 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_74
timestamp 1636915332
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_66
timestamp 1636915332
transform 1 0 6072 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_1  _452_
timestamp 1636915332
transform 1 0 4876 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _401_
timestamp 1636915332
transform 1 0 7268 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1636915332
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_80
timestamp 1636915332
transform 1 0 7360 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_77
timestamp 1636915332
transform 1 0 7084 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__405__A1
timestamp 1636915332
transform 1 0 7176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _360_
timestamp 1636915332
transform -1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _285_
timestamp 1636915332
transform -1 0 9200 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1636915332
transform 1 0 8372 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_88
timestamp 1636915332
transform 1 0 8096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_88
timestamp 1636915332
transform 1 0 8096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _399_
timestamp 1636915332
transform 1 0 8740 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1636915332
transform 1 0 9660 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_1  _284_
timestamp 1636915332
transform -1 0 9568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _271_
timestamp 1636915332
transform 1 0 9568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1636915332
transform 1 0 9568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_107
timestamp 1636915332
transform 1 0 9844 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_2  _350_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 10856 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _281_
timestamp 1636915332
transform -1 0 10580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1636915332
transform 1 0 10764 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_114
timestamp 1636915332
transform 1 0 10488 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_115
timestamp 1636915332
transform 1 0 10580 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _348_
timestamp 1636915332
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_124
timestamp 1636915332
transform 1 0 11408 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_120
timestamp 1636915332
transform 1 0 11040 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1636915332
transform 1 0 11960 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_131
timestamp 1636915332
transform 1 0 12052 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_127
timestamp 1636915332
transform 1 0 11684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__350__A_N
timestamp 1636915332
transform 1 0 11500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_1  _325_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 12604 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _324_
timestamp 1636915332
transform -1 0 12604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_137
timestamp 1636915332
transform 1 0 12604 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__and2_1  _323_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 13156 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _322_
timestamp 1636915332
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _274_
timestamp 1636915332
transform 1 0 13248 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1636915332
transform 1 0 13156 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_148
timestamp 1636915332
transform 1 0 13616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__470__RESET_B
timestamp 1636915332
transform 1 0 13432 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__or2b_1  _319_
timestamp 1636915332
transform 1 0 13800 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1636915332
transform 1 0 14352 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__428__SET_B
timestamp 1636915332
transform 1 0 14628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__B1
timestamp 1636915332
transform 1 0 14444 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1636915332
transform 1 0 15548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_170
timestamp 1636915332
transform 1 0 15640 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_166
timestamp 1636915332
transform 1 0 15272 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__431__SET_B
timestamp 1636915332
transform 1 0 15364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_4  _431_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 15732 0 1 3264
box -38 -48 2246 592
use sky130_fd_sc_hd__dfstp_1  _428_
timestamp 1636915332
transform 1 0 14812 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _415_
timestamp 1636915332
transform 1 0 13800 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1636915332
transform -1 0 18308 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_183
timestamp 1636915332
transform 1 0 16836 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_195
timestamp 1636915332
transform 1 0 17940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1636915332
transform 1 0 16744 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1636915332
transform 1 0 17940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  split4
timestamp 1636915332
transform -1 0 18400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_200
timestamp 1636915332
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1636915332
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1636915332
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1636915332
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1636915332
transform 1 0 1012 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_14
timestamp 1636915332
transform 1 0 1288 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_3
timestamp 1636915332
transform 1 0 276 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1636915332
transform 1 0 0 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1636915332
transform 1 0 1196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_26
timestamp 1636915332
transform 1 0 2392 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1636915332
transform 1 0 2760 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_38
timestamp 1636915332
transform 1 0 3496 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1636915332
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _339_
timestamp 1636915332
transform 1 0 2852 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dfstp_1  _439_
timestamp 1636915332
transform 1 0 3680 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_8_61
timestamp 1636915332
transform 1 0 5612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1636915332
transform 1 0 5980 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_1  _287_
timestamp 1636915332
transform -1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _359_
timestamp 1636915332
transform 1 0 6808 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_8_81
timestamp 1636915332
transform 1 0 7452 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_89
timestamp 1636915332
transform 1 0 8188 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_92
timestamp 1636915332
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1636915332
transform 1 0 8372 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _361_
timestamp 1636915332
transform 1 0 8832 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_8_103
timestamp 1636915332
transform 1 0 9476 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_115
timestamp 1636915332
transform 1 0 10580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1636915332
transform 1 0 10764 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _411_
timestamp 1636915332
transform 1 0 10856 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1636915332
transform 1 0 13156 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _416_
timestamp 1636915332
transform 1 0 11684 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _470_
timestamp 1636915332
transform -1 0 15088 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__432__RESET_B
timestamp 1636915332
transform 1 0 15640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_168
timestamp 1636915332
transform 1 0 15456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1636915332
transform 1 0 15548 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _321_
timestamp 1636915332
transform -1 0 15456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _432_
timestamp 1636915332
transform 1 0 15824 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_8_196
timestamp 1636915332
transform 1 0 18032 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1636915332
transform 1 0 17940 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1636915332
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1636915332
transform 1 0 276 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1636915332
transform 1 0 0 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _461_
timestamp 1636915332
transform 1 0 460 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 1636915332
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1636915332
transform 1 0 2392 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_33
timestamp 1636915332
transform 1 0 3036 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_29
timestamp 1636915332
transform 1 0 2668 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__461__SET_B
timestamp 1636915332
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1636915332
transform 1 0 3680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_37
timestamp 1636915332
transform 1 0 3404 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__463__RESET_B
timestamp 1636915332
transform 1 0 3864 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__SET_B
timestamp 1636915332
transform 1 0 3496 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_44
timestamp 1636915332
transform 1 0 4048 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__464__SET_B
timestamp 1636915332
transform 1 0 5888 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_53
timestamp 1636915332
transform 1 0 4876 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_61
timestamp 1636915332
transform 1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_66
timestamp 1636915332
transform 1 0 6072 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_74
timestamp 1636915332
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1636915332
transform 1 0 4784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk
timestamp 1636915332
transform -1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__453__RESET_B
timestamp 1636915332
transform 1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_79
timestamp 1636915332
transform 1 0 7268 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1636915332
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _453_
timestamp 1636915332
transform 1 0 7544 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk_A
timestamp 1636915332
transform -1 0 9844 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_102
timestamp 1636915332
transform 1 0 9384 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1636915332
transform 1 0 9844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_118
timestamp 1636915332
transform 1 0 10856 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1636915332
transform 1 0 9568 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _370_
timestamp 1636915332
transform -1 0 10856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk
timestamp 1636915332
transform 1 0 10212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__424__RESET_B
timestamp 1636915332
transform 1 0 11776 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_126
timestamp 1636915332
transform 1 0 11592 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1636915332
transform 1 0 11960 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _424_
timestamp 1636915332
transform -1 0 13892 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__RESET_B
timestamp 1636915332
transform 1 0 14720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_151
timestamp 1636915332
transform 1 0 13892 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_155
timestamp 1636915332
transform 1 0 14260 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_157
timestamp 1636915332
transform 1 0 14444 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1636915332
transform 1 0 14352 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _429_
timestamp 1636915332
transform 1 0 14904 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1636915332
transform -1 0 18308 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_183
timestamp 1636915332
transform 1 0 16836 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_195
timestamp 1636915332
transform 1 0 17940 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1636915332
transform 1 0 16744 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1636915332
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1636915332
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1636915332
transform 1 0 1012 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_14
timestamp 1636915332
transform 1 0 1288 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1636915332
transform 1 0 276 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1636915332
transform 1 0 0 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1636915332
transform 1 0 1196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _239__1
timestamp 1636915332
transform -1 0 1012 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 1636915332
transform 1 0 2944 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1636915332
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__and2b_1  _241_
timestamp 1636915332
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _242_
timestamp 1636915332
transform -1 0 4048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _243_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2392 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_2  _463_
timestamp 1636915332
transform 1 0 4048 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1636915332
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _464_
timestamp 1636915332
transform 1 0 6072 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__RESET_B
timestamp 1636915332
transform 1 0 8740 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_92
timestamp 1636915332
transform 1 0 8464 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1636915332
transform 1 0 8372 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _368_
timestamp 1636915332
transform 1 0 8004 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_1  _465_
timestamp 1636915332
transform -1 0 10764 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1636915332
transform 1 0 10764 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _371_
timestamp 1636915332
transform 1 0 10856 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_10_125
timestamp 1636915332
transform 1 0 11500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_137
timestamp 1636915332
transform 1 0 12604 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_144
timestamp 1636915332
transform 1 0 13248 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1636915332
transform 1 0 13156 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__468__SET_B
timestamp 1636915332
transform 1 0 15824 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_152
timestamp 1636915332
transform 1 0 13984 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_161
timestamp 1636915332
transform 1 0 14812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_170
timestamp 1636915332
transform 1 0 15640 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1636915332
transform 1 0 15548 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _377_
timestamp 1636915332
transform 1 0 14168 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1636915332
transform 1 0 17940 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _372_
timestamp 1636915332
transform 1 0 18032 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _468_
timestamp 1636915332
transform 1 0 16008 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_10_200
timestamp 1636915332
transform 1 0 18400 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1636915332
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__460__RESET_B
timestamp 1636915332
transform 1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1636915332
transform 1 0 0 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _460_
timestamp 1636915332
transform 1 0 276 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_11_25
timestamp 1636915332
transform 1 0 2300 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp 1636915332
transform 1 0 2484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_46
timestamp 1636915332
transform 1 0 4232 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1636915332
transform 1 0 2392 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_1  _233_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 2852 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _235_
timestamp 1636915332
transform -1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1636915332
transform -1 0 4232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _237_
timestamp 1636915332
transform -1 0 3956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_11_66
timestamp 1636915332
transform 1 0 6072 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1636915332
transform 1 0 4784 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _231_
timestamp 1636915332
transform -1 0 6072 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1636915332
transform 1 0 4876 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _391_
timestamp 1636915332
transform -1 0 7176 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1636915332
transform 1 0 7268 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_83
timestamp 1636915332
transform 1 0 7636 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1636915332
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 9568 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1636915332
transform 1 0 9568 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _219_
timestamp 1636915332
transform -1 0 9936 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _228_
timestamp 1636915332
transform -1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _389_
timestamp 1636915332
transform -1 0 10764 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__469__RESET_B
timestamp 1636915332
transform 1 0 11776 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_125
timestamp 1636915332
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1636915332
transform 1 0 11960 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _469_
timestamp 1636915332
transform 1 0 12052 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_11_151
timestamp 1636915332
transform 1 0 13892 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1636915332
transform 1 0 14352 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_2  _265_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 14444 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _373_
timestamp 1636915332
transform -1 0 16008 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _376_
timestamp 1636915332
transform -1 0 14352 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_174
timestamp 1636915332
transform 1 0 16008 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_178
timestamp 1636915332
transform 1 0 16376 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1636915332
transform 1 0 16744 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 1636915332
transform 1 0 16836 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp 1636915332
transform 1 0 16468 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _387_
timestamp 1636915332
transform 1 0 17664 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_201
timestamp 1636915332
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1636915332
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__462__RESET_B
timestamp 1636915332
transform 1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1636915332
transform 1 0 1012 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_14
timestamp 1636915332
transform 1 0 1288 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_22
timestamp 1636915332
transform 1 0 2024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1636915332
transform 1 0 276 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1636915332
transform 1 0 0 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1636915332
transform 1 0 1196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_25
timestamp 1636915332
transform 1 0 2300 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_40
timestamp 1636915332
transform 1 0 3680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1636915332
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _234_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 3128 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _238_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 3128 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _251_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 5520 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_1  FILLER_12_60
timestamp 1636915332
transform 1 0 5520 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_66
timestamp 1636915332
transform 1 0 6072 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1636915332
transform 1 0 5980 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _229_
timestamp 1636915332
transform -1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _230_
timestamp 1636915332
transform 1 0 6164 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1636915332
transform 1 0 8372 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__xnor2_1  _369_
timestamp 1636915332
transform -1 0 8372 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1636915332
transform 1 0 6900 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_pll_clk90
timestamp 1636915332
transform -1 0 10304 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_12_116
timestamp 1636915332
transform 1 0 10672 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1636915332
transform 1 0 10764 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _227_
timestamp 1636915332
transform 1 0 10304 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _388_
timestamp 1636915332
transform 1 0 10856 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_134
timestamp 1636915332
transform 1 0 12328 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_139
timestamp 1636915332
transform 1 0 12788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1636915332
transform 1 0 13156 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _204_
timestamp 1636915332
transform 1 0 13248 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1636915332
transform 1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_4  _347_
timestamp 1636915332
transform 1 0 11684 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__433__RESET_B
timestamp 1636915332
transform 1 0 15916 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_170
timestamp 1636915332
transform 1 0 15640 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1636915332
transform 1 0 15548 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _346_
timestamp 1636915332
transform -1 0 14720 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1636915332
transform 1 0 14720 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1636915332
transform -1 0 18308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_196
timestamp 1636915332
transform 1 0 18032 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1636915332
transform 1 0 17940 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _433_
timestamp 1636915332
transform -1 0 17940 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1636915332
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1636915332
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1636915332
transform 1 0 0 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1636915332
transform 1 0 0 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1636915332
transform 1 0 276 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_11
timestamp 1636915332
transform 1 0 1012 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_1  _263_
timestamp 1636915332
transform -1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1636915332
transform -1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _254_
timestamp 1636915332
transform 1 0 2116 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1636915332
transform 1 0 1196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_22
timestamp 1636915332
transform 1 0 2024 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_18
timestamp 1636915332
transform 1 0 1656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1636915332
transform 1 0 1288 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtn_1  _462_
timestamp 1636915332
transform 1 0 276 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  _384_
timestamp 1636915332
transform 1 0 2576 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _223_
timestamp 1636915332
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  _216_
timestamp 1636915332
transform 1 0 2944 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1636915332
transform 1 0 2392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_37
timestamp 1636915332
transform 1 0 3404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_31
timestamp 1636915332
transform 1 0 2852 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__456__RESET_B
timestamp 1636915332
transform 1 0 2392 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__o211a_1  _245_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 4784 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1636915332
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_43
timestamp 1636915332
transform 1 0 3956 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_39
timestamp 1636915332
transform 1 0 3588 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_40
timestamp 1636915332
transform 1 0 3680 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _217_
timestamp 1636915332
transform 1 0 5060 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _215_
timestamp 1636915332
transform -1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1636915332
transform 1 0 4784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_56
timestamp 1636915332
transform 1 0 5152 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_52
timestamp 1636915332
transform 1 0 4784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1636915332
transform 1 0 4876 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_1  _232_
timestamp 1636915332
transform -1 0 6256 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _224_
timestamp 1636915332
transform 1 0 6072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1636915332
transform 1 0 5980 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_61
timestamp 1636915332
transform 1 0 5612 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_pll_clk90
timestamp 1636915332
transform -1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_74
timestamp 1636915332
transform 1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_68
timestamp 1636915332
transform 1 0 6256 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1636915332
transform 1 0 7360 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _218_
timestamp 1636915332
transform -1 0 8372 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _212_
timestamp 1636915332
transform 1 0 7268 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1636915332
transform 1 0 7176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_84
timestamp 1636915332
transform 1 0 7728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_78
timestamp 1636915332
transform 1 0 7176 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_79
timestamp 1636915332
transform 1 0 7268 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_76
timestamp 1636915332
transform 1 0 6992 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _379_
timestamp 1636915332
transform 1 0 8464 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1636915332
transform 1 0 8372 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_89
timestamp 1636915332
transform 1 0 8188 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__467__RESET_B
timestamp 1636915332
transform 1 0 8280 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  _467_
timestamp 1636915332
transform 1 0 8464 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1636915332
transform 1 0 9568 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_105
timestamp 1636915332
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_101
timestamp 1636915332
transform 1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_pll_clk90
timestamp 1636915332
transform 1 0 10488 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _220_
timestamp 1636915332
transform -1 0 10488 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_115
timestamp 1636915332
transform 1 0 10580 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_pll_clk90_A
timestamp 1636915332
transform 1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_1  _213_
timestamp 1636915332
transform -1 0 11408 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1636915332
transform 1 0 10764 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_122
timestamp 1636915332
transform 1 0 11224 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_118
timestamp 1636915332
transform 1 0 10856 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _353_
timestamp 1636915332
transform 1 0 11316 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _225_
timestamp 1636915332
transform -1 0 11960 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_4  _266_
timestamp 1636915332
transform 1 0 12512 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _222_
timestamp 1636915332
transform 1 0 11960 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1636915332
transform 1 0 11960 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _413_
timestamp 1636915332
transform 1 0 13708 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_1  _269_
timestamp 1636915332
transform 1 0 13432 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1636915332
transform 1 0 13156 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_148
timestamp 1636915332
transform 1 0 13616 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_144
timestamp 1636915332
transform 1 0 13248 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_143
timestamp 1636915332
transform 1 0 13156 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_131
timestamp 1636915332
transform 1 0 12052 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _270_
timestamp 1636915332
transform 1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _268_
timestamp 1636915332
transform -1 0 14352 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1636915332
transform 1 0 14536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1636915332
transform 1 0 14352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1636915332
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_166
timestamp 1636915332
transform 1 0 15272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__455__SET_B
timestamp 1636915332
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__436__RESET_B
timestamp 1636915332
transform 1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfstp_1  _455_
timestamp 1636915332
transform -1 0 16376 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _436_
timestamp 1636915332
transform 1 0 15824 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_13_178
timestamp 1636915332
transform 1 0 16376 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_183
timestamp 1636915332
transform 1 0 16836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_195
timestamp 1636915332
transform 1 0 17940 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_196
timestamp 1636915332
transform 1 0 18032 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1636915332
transform 1 0 16744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1636915332
transform 1 0 17940 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_201
timestamp 1636915332
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1636915332
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1636915332
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1636915332
transform 1 0 0 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _255_
timestamp 1636915332
transform -1 0 2392 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _456_
timestamp 1636915332
transform 1 0 276 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_15_31
timestamp 1636915332
transform 1 0 2852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1636915332
transform 1 0 2392 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_1  _264_
timestamp 1636915332
transform -1 0 2852 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _383_
timestamp 1636915332
transform 1 0 2944 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1636915332
transform 1 0 3772 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_50
timestamp 1636915332
transform 1 0 4600 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1636915332
transform 1 0 4784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _409_
timestamp 1636915332
transform 1 0 4876 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _419_
timestamp 1636915332
transform 1 0 5704 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_79
timestamp 1636915332
transform 1 0 7268 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_83
timestamp 1636915332
transform 1 0 7636 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_88
timestamp 1636915332
transform 1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1636915332
transform 1 0 7176 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_1  _208_
timestamp 1636915332
transform 1 0 8464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _209_
timestamp 1636915332
transform 1 0 9016 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _211_
timestamp 1636915332
transform -1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _214_
timestamp 1636915332
transform 1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_105
timestamp 1636915332
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1636915332
transform 1 0 9568 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _226_
timestamp 1636915332
transform 1 0 10764 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _394_
timestamp 1636915332
transform 1 0 11132 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_134
timestamp 1636915332
transform 1 0 12328 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_148
timestamp 1636915332
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1636915332
transform 1 0 11960 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 1636915332
transform -1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2ai_2  _354_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 13616 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__434__SET_B
timestamp 1636915332
transform 1 0 14628 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_155
timestamp 1636915332
transform 1 0 14260 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1636915332
transform 1 0 14444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1636915332
transform 1 0 14352 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _352_
timestamp 1636915332
transform 1 0 13984 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _434_
timestamp 1636915332
transform -1 0 16744 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1636915332
transform -1 0 18308 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_183
timestamp 1636915332
transform 1 0 16836 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_195
timestamp 1636915332
transform 1 0 17940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1636915332
transform 1 0 16744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1636915332
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1636915332
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1636915332
transform -1 0 1472 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1636915332
transform 1 0 1012 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1636915332
transform 1 0 276 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1636915332
transform 1 0 0 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1636915332
transform 1 0 1196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_12  input3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 1472 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_35
timestamp 1636915332
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_40
timestamp 1636915332
transform 1 0 3680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1636915332
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  _259_
timestamp 1636915332
transform -1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _395_
timestamp 1636915332
transform 1 0 4048 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_53
timestamp 1636915332
transform 1 0 4876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_63
timestamp 1636915332
transform 1 0 5796 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_66
timestamp 1636915332
transform 1 0 6072 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1636915332
transform 1 0 5980 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1636915332
transform 1 0 4968 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _418_
timestamp 1636915332
transform 1 0 6808 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_90
timestamp 1636915332
transform 1 0 8280 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_92
timestamp 1636915332
transform 1 0 8464 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1636915332
transform 1 0 8372 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  _417_
timestamp 1636915332
transform 1 0 8648 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__466__SET_B
timestamp 1636915332
transform 1 0 10580 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_114
timestamp 1636915332
transform 1 0 10488 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1636915332
transform 1 0 10764 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _210_
timestamp 1636915332
transform -1 0 10488 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _466_
timestamp 1636915332
transform 1 0 10856 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__438__RESET_B
timestamp 1636915332
transform 1 0 13248 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_139
timestamp 1636915332
transform 1 0 12788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1636915332
transform 1 0 13156 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _438_
timestamp 1636915332
transform 1 0 13432 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_16_170
timestamp 1636915332
transform 1 0 15640 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1636915332
transform 1 0 15548 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_4  _437_
timestamp 1636915332
transform 1 0 15732 0 1 8704
box -38 -48 2246 592
use sky130_fd_sc_hd__decap_6  FILLER_16_196
timestamp 1636915332
transform 1 0 18032 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1636915332
transform 1 0 17940 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1636915332
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1636915332
transform 1 0 0 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _257_
timestamp 1636915332
transform -1 0 2392 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtn_1  _458_
timestamp 1636915332
transform 1 0 276 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__458__RESET_B
timestamp 1636915332
transform 1 0 3496 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_40
timestamp 1636915332
transform 1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1636915332
transform 1 0 2392 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nand3_1  _256_
timestamp 1636915332
transform -1 0 2852 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _260_
timestamp 1636915332
transform -1 0 3220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _261_
timestamp 1636915332
transform -1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _365_
timestamp 1636915332
transform 1 0 3956 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__459__SET_B
timestamp 1636915332
transform 1 0 5980 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_50
timestamp 1636915332
transform 1 0 4600 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1636915332
transform 1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1636915332
transform 1 0 5520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_72
timestamp 1636915332
transform 1 0 6624 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1636915332
transform 1 0 4784 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _244__2
timestamp 1636915332
transform -1 0 6624 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _248_
timestamp 1636915332
transform 1 0 5152 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _253_
timestamp 1636915332
transform -1 0 5980 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1636915332
transform 1 0 7176 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _246_
timestamp 1636915332
transform -1 0 7912 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _420_
timestamp 1636915332
transform 1 0 7912 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__425__RESET_B
timestamp 1636915332
transform 1 0 9936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_ext_clk_A
timestamp 1636915332
transform -1 0 9936 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_102
timestamp 1636915332
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_105
timestamp 1636915332
transform 1 0 9660 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1636915332
transform 1 0 9568 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _425_
timestamp 1636915332
transform 1 0 10120 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__435__RESET_B
timestamp 1636915332
transform 1 0 12328 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_131
timestamp 1636915332
transform 1 0 12052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1636915332
transform 1 0 11960 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_1  _435_
timestamp 1636915332
transform -1 0 14352 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__422__SET_B
timestamp 1636915332
transform 1 0 14628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 1636915332
transform 1 0 14444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1636915332
transform 1 0 14352 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _422_
timestamp 1636915332
transform 1 0 14812 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_8  FILLER_17_191
timestamp 1636915332
transform 1 0 17572 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1636915332
transform 1 0 16744 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 16836 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_199
timestamp 1636915332
transform 1 0 18308 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1636915332
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_11
timestamp 1636915332
transform 1 0 1012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_3
timestamp 1636915332
transform 1 0 276 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1636915332
transform 1 0 0 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1636915332
transform 1 0 1196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _457_
timestamp 1636915332
transform 1 0 1288 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_18_35
timestamp 1636915332
transform 1 0 3220 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1636915332
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor3b_2  _247_
timestamp 1636915332
transform -1 0 4600 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _366_
timestamp 1636915332
transform -1 0 3588 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_56
timestamp 1636915332
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_64
timestamp 1636915332
transform 1 0 5888 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1636915332
transform 1 0 5980 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _249_
timestamp 1636915332
transform -1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _250_
timestamp 1636915332
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _252_
timestamp 1636915332
transform -1 0 5888 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dfstp_1  _459_
timestamp 1636915332
transform 1 0 6072 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__426__RESET_B
timestamp 1636915332
transform 1 0 8740 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1636915332
transform 1 0 8004 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1636915332
transform 1 0 8372 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _344_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 8740 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _426_
timestamp 1636915332
transform 1 0 8924 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1636915332
transform 1 0 10764 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ext_clk
timestamp 1636915332
transform 1 0 10856 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  FILLER_18_142
timestamp 1636915332
transform 1 0 13064 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_144
timestamp 1636915332
transform 1 0 13248 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1636915332
transform 1 0 13156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _423_
timestamp 1636915332
transform 1 0 13340 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_ext_clk
timestamp 1636915332
transform -1 0 13064 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__421__SET_B
timestamp 1636915332
transform 1 0 15824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__437__SET_B
timestamp 1636915332
transform 1 0 15640 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_166
timestamp 1636915332
transform 1 0 15272 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1636915332
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1636915332
transform -1 0 18308 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_196
timestamp 1636915332
transform 1 0 18032 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1636915332
transform 1 0 17940 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dfstp_1  _421_
timestamp 1636915332
transform 1 0 16008 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1636915332
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1636915332
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1636915332
transform 1 0 1012 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_14
timestamp 1636915332
transform 1 0 1288 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_20
timestamp 1636915332
transform 1 0 1840 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1636915332
transform 1 0 276 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1636915332
transform 1 0 0 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1636915332
transform 1 0 1196 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _258__3
timestamp 1636915332
transform -1 0 1840 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__457__SET_B
timestamp 1636915332
transform 1 0 3220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_27
timestamp 1636915332
transform 1 0 2484 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1636915332
transform 1 0 3404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_47
timestamp 1636915332
transform 1 0 4324 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1636915332
transform 1 0 2392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1636915332
transform 1 0 3588 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  _367_
timestamp 1636915332
transform 1 0 3680 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_19_51
timestamp 1636915332
transform 1 0 4692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_53
timestamp 1636915332
transform 1 0 4876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_66
timestamp 1636915332
transform 1 0 6072 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1636915332
transform 1 0 4784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1636915332
transform 1 0 5980 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__343__S
timestamp 1636915332
transform 1 0 8188 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_86
timestamp 1636915332
transform 1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1636915332
transform 1 0 7176 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1636915332
transform 1 0 8372 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _343_ OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform 1 0 8464 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_ext_clk
timestamp 1636915332
transform 1 0 7544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output10
timestamp 1636915332
transform 1 0 7268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_101
timestamp 1636915332
transform 1 0 9292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_116
timestamp 1636915332
transform 1 0 10672 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1636915332
transform 1 0 9568 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1636915332
transform 1 0 10764 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _412_
timestamp 1636915332
transform -1 0 11684 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1
timestamp 1636915332
transform 1 0 9660 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  output12
timestamp 1636915332
transform 1 0 10396 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__423__SET_B
timestamp 1636915332
transform 1 0 13248 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_127
timestamp 1636915332
transform 1 0 11684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_140
timestamp 1636915332
transform 1 0 12880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1636915332
transform 1 0 11960 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1636915332
transform 1 0 13156 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _340__9
timestamp 1636915332
transform -1 0 13892 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _393_
timestamp 1636915332
transform 1 0 12052 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_155
timestamp 1636915332
transform 1 0 14260 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1636915332
transform 1 0 14720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_167
timestamp 1636915332
transform 1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1636915332
transform 1 0 14352 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1636915332
transform 1 0 15548 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _341__8
timestamp 1636915332
transform -1 0 15364 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__conb_1  _378__13 OpenLane/pdks//sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1636915332
transform -1 0 14720 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1636915332
transform 1 0 15640 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1636915332
transform -1 0 14260 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1636915332
transform -1 0 17940 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1636915332
transform 1 0 16376 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_188
timestamp 1636915332
transform 1 0 17296 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_192
timestamp 1636915332
transform 1 0 17664 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1636915332
transform 1 0 16744 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1636915332
transform 1 0 17940 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_4  _342__7
timestamp 1636915332
transform -1 0 17296 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _375_
timestamp 1636915332
transform 1 0 18032 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1636915332
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1636915332
transform 1 0 18308 0 -1 10880
box -38 -48 314 592
<< labels >>
rlabel metal5 s 0 4812 18860 5132 6 VGND
port 0 nsew ground input
rlabel metal5 s 0 8192 18860 8512 6 VGND
port 0 nsew ground input
rlabel metal4 s 4654 -48 4974 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 7754 -48 8074 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 10854 -48 11174 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 13954 -48 14274 10928 6 VGND
port 0 nsew ground input
rlabel metal4 s 17054 -48 17374 10928 6 VGND
port 0 nsew ground input
rlabel metal5 s 0 3122 18860 3442 6 VPWR
port 1 nsew power input
rlabel metal5 s 0 6502 18860 6822 6 VPWR
port 1 nsew power input
rlabel metal5 s 0 9882 18860 10202 6 VPWR
port 1 nsew power input
rlabel metal4 s 3104 -48 3424 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 6204 -48 6524 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 9304 -48 9624 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 12404 -48 12724 10928 6 VPWR
port 1 nsew power input
rlabel metal4 s 15504 -48 15824 10928 6 VPWR
port 1 nsew power input
rlabel metal2 s 7102 11200 7158 12000 6 core_clk
port 2 nsew signal tristate
rlabel metal2 s 4250 11200 4306 12000 6 ext_clk
port 3 nsew signal input
rlabel metal3 s 19200 688 20000 808 6 ext_clk_sel
port 4 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 ext_reset
port 5 nsew signal input
rlabel metal2 s 15658 11200 15714 12000 6 pll_clk
port 6 nsew signal input
rlabel metal2 s 18510 11200 18566 12000 6 pll_clk90
port 7 nsew signal input
rlabel metal2 s 1398 11200 1454 12000 6 resetb
port 8 nsew signal input
rlabel metal2 s 12806 11200 12862 12000 6 resetb_sync
port 9 nsew signal tristate
rlabel metal3 s 19200 6672 20000 6792 6 sel2[0]
port 10 nsew signal input
rlabel metal3 s 19200 8168 20000 8288 6 sel2[1]
port 11 nsew signal input
rlabel metal3 s 19200 9664 20000 9784 6 sel2[2]
port 12 nsew signal input
rlabel metal3 s 19200 2184 20000 2304 6 sel[0]
port 13 nsew signal input
rlabel metal3 s 19200 3680 20000 3800 6 sel[1]
port 14 nsew signal input
rlabel metal3 s 19200 5176 20000 5296 6 sel[2]
port 15 nsew signal input
rlabel metal2 s 9954 11200 10010 12000 6 user_clk
port 16 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 12000
<< end >>
