magic
tech sky130A
magscale 1 2
timestamp 1686151263
<< checkpaint >>
rect -1260 996747 718860 1038860
rect -1260 996340 42060 996747
rect -1260 971594 40853 996340
rect 68429 995258 93594 996747
rect 68429 994534 73601 995258
rect 74797 994147 93594 995258
rect 119629 995258 144994 996747
rect 119629 994534 124801 995258
rect 126197 994147 144994 995258
rect 170829 995258 196394 996747
rect 170829 994534 176001 995258
rect 177597 994147 196394 995258
rect 222029 995258 247794 996747
rect 222029 994534 227201 995258
rect 228997 994147 247794 995258
rect 273229 995258 299394 996747
rect 332140 996340 349660 996747
rect 273229 994534 278401 995258
rect 280597 994147 299394 995258
rect 377629 994534 401194 996747
rect 466629 994534 490194 996747
rect 517829 994534 541594 996747
rect 574340 996340 591860 996747
rect 617229 995258 643394 996747
rect 676340 995540 718860 996747
rect 617229 994534 622401 995258
rect 382397 994147 401194 994534
rect 471397 994147 490194 994534
rect 522797 994147 541594 994534
rect 624597 994147 643394 995258
rect 88689 994059 91412 994147
rect 140092 994068 142815 994147
rect 191496 994050 194219 994147
rect 242902 994086 245625 994147
rect 294504 994038 297227 994147
rect 396305 994083 399028 994147
rect 485285 994047 488008 994147
rect 536713 994008 539436 994147
rect 638473 993970 641185 994147
rect 676747 972411 718860 995540
rect -1260 971564 43453 971594
rect -1260 969399 43454 971564
rect 674545 970312 718860 972411
rect -1260 966701 43595 969399
rect -1260 964260 43457 966701
rect -1260 951488 43454 964260
rect 674146 957540 718860 970312
rect 674143 955127 718860 957540
rect 674053 952395 718860 955127
rect -1260 950747 42152 951488
rect -1260 945575 43062 950747
rect 674146 950236 718860 952395
rect 674147 950206 718860 950236
rect -1260 930447 40853 945575
rect -1260 910740 43030 930447
rect 676747 923860 718860 950206
rect -1260 886060 40853 910740
rect 674570 904153 718860 923860
rect -1260 868540 41260 886060
rect 676747 882411 718860 904153
rect 674545 881112 718860 882411
rect -1260 843860 40853 868540
rect 674146 868340 718860 881112
rect 674143 865952 718860 868340
rect 674079 863220 718860 865952
rect 674146 861036 718860 863220
rect 674147 861006 718860 861036
rect -1260 826340 41260 843860
rect 676747 834660 718860 861006
rect -1260 801794 40853 826340
rect 676340 817140 718860 834660
rect -1260 801764 43453 801794
rect -1260 799604 43454 801764
rect -1260 796906 43574 799604
rect -1260 794460 43457 796906
rect -1260 781688 43454 794460
rect 676747 793411 718860 817140
rect 674545 791912 718860 793411
rect -1260 780747 42152 781688
rect -1260 775575 43062 780747
rect 674146 779140 718860 791912
rect 674143 776750 718860 779140
rect -1260 758594 40853 775575
rect 674041 774018 718860 776750
rect 674146 771836 718860 774018
rect 674147 771806 718860 771836
rect -1260 758564 43453 758594
rect -1260 756407 43454 758564
rect -1260 753709 43568 756407
rect -1260 751260 43457 753709
rect -1260 738488 43454 751260
rect 676747 748411 718860 771806
rect 674545 746912 718860 748411
rect -1260 737747 42152 738488
rect -1260 732575 43062 737747
rect 674146 734140 718860 746912
rect -1260 715394 40853 732575
rect 674143 731756 718860 734140
rect 674050 729024 718860 731756
rect 674146 726836 718860 729024
rect 674147 726806 718860 726836
rect -1260 715364 43453 715394
rect -1260 713205 43454 715364
rect -1260 710504 43503 713205
rect -1260 708060 43457 710504
rect -1260 695288 43454 708060
rect 676747 703411 718860 726806
rect 674545 701912 718860 703411
rect -1260 694747 42152 695288
rect -1260 689575 43062 694747
rect -1260 672194 40853 689575
rect 674146 689140 718860 701912
rect 674143 686729 718860 689140
rect 674061 683997 718860 686729
rect 674146 681836 718860 683997
rect 674147 681806 718860 681836
rect -1260 672164 43453 672194
rect -1260 669996 43454 672164
rect -1260 667295 43521 669996
rect -1260 664860 43457 667295
rect -1260 652088 43454 664860
rect 676747 658411 718860 681806
rect 674545 656712 718860 658411
rect -1260 651747 42152 652088
rect -1260 646575 43062 651747
rect -1260 628994 40853 646575
rect 674146 643940 718860 656712
rect 674143 641546 718860 643940
rect 674058 638814 718860 641546
rect 674146 636636 718860 638814
rect 674147 636606 718860 636636
rect -1260 628964 43453 628994
rect -1260 626775 43454 628964
rect -1260 624074 43560 626775
rect -1260 621660 43457 624074
rect -1260 608888 43454 621660
rect 676747 613411 718860 636606
rect 674545 611712 718860 613411
rect -1260 608747 42152 608888
rect -1260 603575 43062 608747
rect -1260 585794 40853 603575
rect 674146 598940 718860 611712
rect 674143 596526 718860 598940
rect 674038 593794 718860 596526
rect 674146 591636 718860 593794
rect 674147 591606 718860 591636
rect -1260 585764 43453 585794
rect -1260 583599 43454 585764
rect -1260 580898 43557 583599
rect -1260 578460 43457 580898
rect -1260 565688 43454 578460
rect 676747 568411 718860 591606
rect 674545 566512 718860 568411
rect -1260 560575 43062 565688
rect -1260 542594 40853 560575
rect 674146 553740 718860 566512
rect 674143 551322 718860 553740
rect 673985 548590 718860 551322
rect 674146 546436 718860 548590
rect 674147 546406 718860 546436
rect -1260 542564 43453 542594
rect -1260 540417 43454 542564
rect -1260 537716 43524 540417
rect -1260 535260 43457 537716
rect -1260 522488 43454 535260
rect -1260 517575 43062 522488
rect 676747 520060 718860 546406
rect -1260 499260 40853 517575
rect 676340 502540 718860 520060
rect -1260 481740 41260 499260
rect -1260 459247 40853 481740
rect 676747 476060 718860 502540
rect -1260 439540 43030 459247
rect 674570 456353 718860 476060
rect -1260 414994 40853 439540
rect 676747 431860 718860 456353
rect -1260 414964 43453 414994
rect -1260 412794 43454 414964
rect 676340 414340 718860 431860
rect -1260 410093 43578 412794
rect -1260 407660 43457 410093
rect -1260 394888 43454 407660
rect -1260 393747 42152 394888
rect -1260 388575 43062 393747
rect 676747 391411 718860 414340
rect 674545 389312 718860 391411
rect -1260 371794 40853 388575
rect 674146 376540 718860 389312
rect 674143 374089 718860 376540
rect -1260 371764 43453 371794
rect -1260 369576 43454 371764
rect 674082 371404 718860 374089
rect -1260 366875 43563 369576
rect 674146 369236 718860 371404
rect 674147 369206 718860 369236
rect -1260 364460 43457 366875
rect -1260 351688 43454 364460
rect -1260 350747 42152 351688
rect -1260 345575 43062 350747
rect 676747 346411 718860 369206
rect -1260 328594 40853 345575
rect 674545 344112 718860 346411
rect 674146 331340 718860 344112
rect 674143 328891 718860 331340
rect -1260 328564 43453 328594
rect -1260 326398 43454 328564
rect -1260 323697 43581 326398
rect 674088 326206 718860 328891
rect 674104 325013 718860 326206
rect 674146 324036 718860 325013
rect 674147 324006 718860 324036
rect -1260 321260 43457 323697
rect -1260 308488 43454 321260
rect -1260 307747 42152 308488
rect -1260 302575 43062 307747
rect -1260 285394 40853 302575
rect 676747 301411 718860 324006
rect 674545 299112 718860 301411
rect 674146 286340 718860 299112
rect -1260 285364 43453 285394
rect -1260 283181 43454 285364
rect 674143 283987 718860 286340
rect -1260 280512 43530 283181
rect 674061 281197 718860 283987
rect -1260 278060 43457 280512
rect 674146 279036 718860 281197
rect 674147 279006 718860 279036
rect -1260 265288 43454 278060
rect -1260 264747 42152 265288
rect -1260 259575 43062 264747
rect -1260 242194 40853 259575
rect 676747 256411 718860 279006
rect 674545 254112 718860 256411
rect -1260 242164 43453 242194
rect -1260 239999 43454 242164
rect 674146 242129 718860 254112
rect -1260 237330 43626 239999
rect 674061 239339 718860 242129
rect 674143 239018 718860 239339
rect -1260 234860 43457 237330
rect 674099 236228 718860 239018
rect -1260 222088 43454 234860
rect 674146 234036 718860 236228
rect 674147 234006 718860 234036
rect -1260 221747 42152 222088
rect -1260 216575 43062 221747
rect -1260 198994 40853 216575
rect 676747 211411 718860 234006
rect 674545 208912 718860 211411
rect -1260 198964 43453 198994
rect -1260 196760 43454 198964
rect -1260 194091 43587 196760
rect 674146 196140 718860 208912
rect -1260 191660 43457 194091
rect 674143 193677 718860 196140
rect -1260 178888 43454 191660
rect 674042 191015 718860 193677
rect 674146 188836 718860 191015
rect 674147 188806 718860 188836
rect -1260 178747 42152 178888
rect -1260 173575 43062 178747
rect -1260 126460 40853 173575
rect 676747 166411 718860 188806
rect 674545 163912 718860 166411
rect 674146 151140 718860 163912
rect 674143 148603 718860 151140
rect 674146 143836 718860 148603
rect 674147 143806 718860 143836
rect -1260 108940 41260 126460
rect 676747 121411 718860 143806
rect 674545 118712 718860 121411
rect -1260 86499 40853 108940
rect 674146 105940 718860 118712
rect 674143 103403 718860 105940
rect 674146 98636 718860 103403
rect 674147 98606 718860 98636
rect -1260 66740 42960 86499
rect -1260 42060 40853 66740
rect 187150 43453 189873 43585
rect 295800 43453 298523 43624
rect 350583 43453 353306 43657
rect 405391 43453 408114 43630
rect 460222 43453 462945 43642
rect 514982 43453 517705 43597
rect 185006 43036 203803 43453
rect 293606 43036 312403 43453
rect 348406 43036 367203 43453
rect 403206 43036 422003 43453
rect 458006 43036 476803 43453
rect 512806 43036 531603 43453
rect -1260 40853 41260 42060
rect 147050 41260 152222 43036
rect 77540 40853 95060 41260
rect 131216 40853 152222 41260
rect 185006 42342 207022 43036
rect 185006 42204 208065 42342
rect 185006 40853 208478 42204
rect 237701 40853 257460 42960
rect 293606 42342 316622 43036
rect 348406 42342 371422 43036
rect 403206 42342 426222 43036
rect 458006 42342 481022 43036
rect 512806 42342 535822 43036
rect 293606 42204 316665 42342
rect 348406 42204 371465 42342
rect 403206 42204 426265 42342
rect 458006 42204 481065 42342
rect 512806 42204 535865 42342
rect 293606 40853 317078 42204
rect 348406 40853 371878 42204
rect 403206 40853 426678 42204
rect 458006 40853 481478 42204
rect 512806 40853 536278 42204
rect 676747 41260 718860 98606
rect 567740 40853 585260 41260
rect 621540 40853 639060 41260
rect 675540 40853 718860 41260
rect -1260 -1260 718860 40853
rect -1260 -1267 1261 -1260
<< error_s >>
rect 149223 18082 150855 18116
<< metal1 >>
rect 41866 995682 675734 995734
rect 41866 95347 41918 995682
rect 41525 95291 41536 95347
rect 41835 95291 41918 95347
rect 41866 41918 41918 95291
rect 675682 41918 675734 995682
rect 41866 41866 145063 41918
rect 145115 41866 145127 41918
rect 145179 41866 675734 41918
rect 140988 40073 140996 40125
rect 141048 40073 141992 40125
rect 142044 40073 143068 40125
rect 143120 40073 143437 40125
rect 143489 40073 144603 40125
rect 144655 40073 144661 40125
rect 142573 40000 142619 40073
rect 644271 20040 644277 20057
rect 644262 20012 644277 20040
rect 644271 20005 644277 20012
rect 644329 20040 644335 20057
rect 653205 20040 653211 20052
rect 644329 20012 653211 20040
rect 644329 20005 644335 20012
rect 653205 20000 653211 20012
rect 653375 20040 653381 20052
rect 653375 20012 653397 20040
rect 653375 20000 653381 20012
rect 646996 19928 647002 19940
rect 646984 19900 647002 19928
rect 646996 19888 647002 19900
rect 647054 19928 647060 19940
rect 652981 19928 652987 19940
rect 647054 19900 652987 19928
rect 647054 19888 647060 19900
rect 652981 19888 652987 19900
rect 653151 19928 653157 19940
rect 653151 19900 653173 19928
rect 653151 19888 653157 19900
rect 643999 19816 644005 19831
rect 643994 19788 644005 19816
rect 643999 19779 644005 19788
rect 644057 19816 644063 19831
rect 652757 19816 652763 19828
rect 644057 19788 652763 19816
rect 644057 19779 644063 19788
rect 652757 19776 652763 19788
rect 652927 19816 652933 19828
rect 652927 19788 652948 19816
rect 652927 19776 652933 19788
rect 643902 19480 643908 19503
rect 643896 19452 643908 19480
rect 643902 19451 643908 19452
rect 643960 19480 643966 19503
rect 652085 19480 652091 19492
rect 643960 19452 652091 19480
rect 643960 19451 643966 19452
rect 652085 19440 652091 19452
rect 652255 19440 652261 19492
rect 646111 19144 646117 19152
rect 646099 19116 646117 19144
rect 646111 19100 646117 19116
rect 646169 19144 646175 19152
rect 651413 19144 651419 19156
rect 646169 19116 651419 19144
rect 646169 19100 646175 19116
rect 651413 19104 651419 19116
rect 651583 19144 651589 19156
rect 651583 19116 651611 19144
rect 651583 19104 651589 19116
rect 643343 19032 643349 19048
rect 643335 19004 643349 19032
rect 643343 18996 643349 19004
rect 643401 19032 643407 19048
rect 651189 19032 651195 19044
rect 643401 19004 651195 19032
rect 643401 18996 643407 19004
rect 651189 18992 651195 19004
rect 651359 19032 651365 19044
rect 651359 19004 651383 19032
rect 651359 18992 651365 19004
rect 644826 18920 644832 18935
rect 644814 18892 644832 18920
rect 644826 18883 644832 18892
rect 644884 18920 644890 18935
rect 650965 18920 650971 18932
rect 644884 18892 650971 18920
rect 644884 18883 644890 18892
rect 650965 18880 650971 18892
rect 651135 18920 651141 18932
rect 651135 18892 651150 18920
rect 651135 18880 651141 18892
rect 643801 18360 643807 18373
rect 643794 18332 643807 18360
rect 643801 18321 643807 18332
rect 643859 18360 643865 18373
rect 649845 18360 649851 18372
rect 643859 18332 649851 18360
rect 643859 18321 643865 18332
rect 649845 18320 649851 18332
rect 650015 18360 650021 18372
rect 650015 18332 650037 18360
rect 650015 18320 650021 18332
rect 644104 18248 644110 18272
rect 644094 18220 644110 18248
rect 644162 18248 644168 18272
rect 649621 18248 649627 18260
rect 644162 18220 649627 18248
rect 649621 18208 649627 18220
rect 649791 18248 649797 18260
rect 649791 18220 649809 18248
rect 649791 18208 649797 18220
rect 649397 18136 649403 18148
rect 649390 18108 649403 18136
rect 649397 18096 649403 18108
rect 649567 18136 649573 18148
rect 652347 18136 652353 18145
rect 649567 18108 652353 18136
rect 649567 18096 649573 18108
rect 652347 18093 652353 18108
rect 652405 18136 652411 18145
rect 652405 18108 652422 18136
rect 652405 18093 652411 18108
rect 645376 18024 645382 18037
rect 645369 17996 645382 18024
rect 645376 17985 645382 17996
rect 645434 18024 645440 18037
rect 649173 18024 649179 18036
rect 645434 17996 649179 18024
rect 645434 17985 645440 17996
rect 649173 17984 649179 17996
rect 649343 18024 649349 18036
rect 649343 17996 649360 18024
rect 649343 17984 649349 17996
rect 648949 17912 648955 17924
rect 648943 17884 648955 17912
rect 648949 17872 648955 17884
rect 649119 17912 649125 17924
rect 652228 17912 652234 17929
rect 649119 17884 652234 17912
rect 649119 17872 649125 17884
rect 652228 17877 652234 17884
rect 652286 17912 652292 17929
rect 652286 17884 652310 17912
rect 652286 17877 652292 17884
rect 646665 17800 646671 17816
rect 646658 17772 646671 17800
rect 646665 17764 646671 17772
rect 646723 17800 646729 17816
rect 648725 17800 648731 17812
rect 646723 17772 648731 17800
rect 646723 17764 646729 17772
rect 648725 17760 648731 17772
rect 648895 17800 648901 17812
rect 648895 17772 648909 17800
rect 648895 17760 648901 17772
rect 643679 17688 643685 17698
rect 643674 17660 643685 17688
rect 643679 17646 643685 17660
rect 643737 17688 643743 17698
rect 648501 17688 648507 17700
rect 643737 17660 648507 17688
rect 643737 17646 643743 17660
rect 648501 17648 648507 17660
rect 648671 17688 648677 17700
rect 648671 17660 648683 17688
rect 648671 17648 648677 17660
rect 648277 17576 648283 17588
rect 648268 17548 648283 17576
rect 648277 17536 648283 17548
rect 648447 17576 648453 17588
rect 649859 17576 649865 17587
rect 648447 17548 649865 17576
rect 648447 17536 648453 17548
rect 649859 17535 649865 17548
rect 649917 17576 649923 17587
rect 649917 17548 649928 17576
rect 649917 17535 649923 17548
rect 648053 17464 648059 17476
rect 648043 17436 648059 17464
rect 648053 17424 648059 17436
rect 648223 17464 648229 17476
rect 649747 17464 649753 17477
rect 648223 17436 649753 17464
rect 648223 17424 648229 17436
rect 649747 17425 649753 17436
rect 649805 17464 649811 17477
rect 649805 17436 649817 17464
rect 649805 17425 649811 17436
rect 647829 17352 647835 17364
rect 647816 17324 647835 17352
rect 647829 17312 647835 17324
rect 647999 17352 648005 17364
rect 652090 17352 652096 17363
rect 647999 17324 652096 17352
rect 647999 17312 648005 17324
rect 652090 17311 652096 17324
rect 652148 17352 652154 17363
rect 652148 17324 652168 17352
rect 652148 17311 652154 17324
rect 643453 17240 643459 17254
rect 643450 17212 643459 17240
rect 643453 17202 643459 17212
rect 643511 17240 643517 17254
rect 647605 17240 647611 17252
rect 643511 17212 647611 17240
rect 643511 17202 643517 17212
rect 647605 17200 647611 17212
rect 647775 17240 647781 17252
rect 647775 17212 647794 17240
rect 647775 17200 647781 17212
rect 643565 17128 643571 17140
rect 643559 17100 643571 17128
rect 643565 17088 643571 17100
rect 643623 17128 643629 17140
rect 647381 17128 647387 17140
rect 643623 17100 647387 17128
rect 643623 17088 643629 17100
rect 647381 17088 647387 17100
rect 647551 17128 647557 17140
rect 647551 17100 647570 17128
rect 647551 17088 647557 17100
rect 646996 16891 647002 16943
rect 647054 16931 647060 16943
rect 647952 16931 647958 16943
rect 647054 16903 647958 16931
rect 647054 16891 647060 16903
rect 647952 16891 647958 16903
rect 648010 16891 648016 16943
rect 649056 16892 649062 16944
rect 649114 16932 649120 16944
rect 652632 16932 652638 16944
rect 649114 16904 652638 16932
rect 649114 16892 649120 16904
rect 652632 16892 652638 16904
rect 652690 16892 652696 16944
rect 649608 16769 649614 16821
rect 649666 16809 649672 16821
rect 653488 16809 653494 16821
rect 649666 16781 653494 16809
rect 649666 16769 649672 16781
rect 653488 16769 653494 16781
rect 653546 16769 653552 16821
rect 650123 16592 650129 16644
rect 650181 16632 650187 16644
rect 653932 16632 653938 16639
rect 650181 16604 653938 16632
rect 650181 16592 650187 16604
rect 653932 16587 653938 16604
rect 653990 16632 653996 16639
rect 653990 16604 653997 16632
rect 653990 16587 653996 16604
rect 648501 9927 648507 9979
rect 648559 9967 648565 9979
rect 652718 9967 652724 9979
rect 648559 9939 652724 9967
rect 648559 9927 648565 9939
rect 652718 9927 652724 9939
rect 652776 9927 652782 9979
rect 647209 9841 647215 9893
rect 647267 9881 647273 9893
rect 652347 9881 652353 9893
rect 647267 9853 652353 9881
rect 647267 9841 647273 9853
rect 652347 9841 652353 9853
rect 652405 9881 652411 9893
rect 652405 9853 652420 9881
rect 652405 9841 652411 9853
rect 647952 9782 647958 9794
rect 647948 9754 647958 9782
rect 647952 9742 647958 9754
rect 648010 9782 648016 9794
rect 652228 9782 652234 9794
rect 648010 9754 652234 9782
rect 648010 9742 648016 9754
rect 652228 9742 652234 9754
rect 652286 9782 652292 9794
rect 652286 9754 652296 9782
rect 652286 9742 652292 9754
rect 646664 9694 646670 9706
rect 646660 9666 646670 9694
rect 646664 9654 646670 9666
rect 646722 9694 646728 9706
rect 652090 9694 652096 9706
rect 646722 9666 652096 9694
rect 646722 9654 646728 9666
rect 652090 9654 652096 9666
rect 652148 9694 652154 9706
rect 652148 9666 652157 9694
rect 652148 9654 652154 9666
rect 645370 9551 645376 9603
rect 645428 9591 645434 9603
rect 650795 9591 650801 9603
rect 645428 9563 650801 9591
rect 645428 9551 645434 9563
rect 650795 9551 650801 9563
rect 650853 9551 650859 9603
rect 644821 9448 644827 9500
rect 644879 9488 644885 9500
rect 652508 9488 652514 9500
rect 644879 9460 652514 9488
rect 644879 9448 644885 9460
rect 652508 9448 652514 9460
rect 652566 9448 652572 9500
rect 646111 9350 646117 9402
rect 646169 9390 646175 9402
rect 652878 9390 652884 9402
rect 646169 9362 652884 9390
rect 646169 9350 646175 9362
rect 652878 9350 652884 9362
rect 652936 9350 652942 9402
<< via1 >>
rect 41536 95291 41835 95347
rect 145063 41866 145115 41918
rect 145127 41866 145179 41918
rect 140996 40073 141048 40125
rect 141992 40073 142044 40125
rect 143068 40073 143120 40125
rect 143437 40073 143489 40125
rect 144603 40073 144655 40125
rect 644277 20005 644329 20057
rect 653211 20000 653375 20052
rect 647002 19888 647054 19940
rect 652987 19888 653151 19940
rect 644005 19779 644057 19831
rect 652763 19776 652927 19828
rect 643908 19451 643960 19503
rect 652091 19440 652255 19492
rect 646117 19100 646169 19152
rect 651419 19104 651583 19156
rect 643349 18996 643401 19048
rect 651195 18992 651359 19044
rect 644832 18883 644884 18935
rect 650971 18880 651135 18932
rect 643807 18321 643859 18373
rect 649851 18320 650015 18372
rect 644110 18220 644162 18272
rect 649627 18208 649791 18260
rect 649403 18096 649567 18148
rect 652353 18093 652405 18145
rect 645382 17985 645434 18037
rect 649179 17984 649343 18036
rect 648955 17872 649119 17924
rect 652234 17877 652286 17929
rect 646671 17764 646723 17816
rect 648731 17760 648895 17812
rect 643685 17646 643737 17698
rect 648507 17648 648671 17700
rect 648283 17536 648447 17588
rect 649865 17535 649917 17587
rect 648059 17424 648223 17476
rect 649753 17425 649805 17477
rect 647835 17312 647999 17364
rect 652096 17311 652148 17363
rect 643459 17202 643511 17254
rect 647611 17200 647775 17252
rect 643571 17088 643623 17140
rect 647387 17088 647551 17140
rect 647002 16891 647054 16943
rect 647958 16891 648010 16943
rect 649062 16892 649114 16944
rect 652638 16892 652690 16944
rect 649614 16769 649666 16821
rect 653494 16769 653546 16821
rect 650129 16592 650181 16644
rect 653938 16587 653990 16639
rect 648507 9927 648559 9979
rect 652724 9927 652776 9979
rect 647215 9841 647267 9893
rect 652353 9841 652405 9893
rect 647958 9742 648010 9794
rect 652234 9742 652286 9794
rect 646670 9654 646722 9706
rect 652096 9654 652148 9706
rect 645376 9551 645428 9603
rect 650801 9551 650853 9603
rect 644827 9448 644879 9500
rect 652514 9448 652566 9500
rect 646117 9350 646169 9402
rect 652884 9350 652936 9402
<< metal2 >>
rect 69634 996754 69695 996786
rect 69634 995407 69695 996693
rect 71635 996754 71696 996786
rect 71635 995407 71696 996693
rect 120834 996754 120895 996786
rect 76497 995407 76553 995887
rect 77049 995407 77105 995887
rect 77693 995407 77749 995887
rect 78337 995407 78393 995887
rect 80177 995407 80233 995887
rect 80729 995407 80785 995887
rect 81373 995407 81429 995887
rect 82017 995407 82073 995887
rect 84501 995407 84557 995887
rect 85053 995407 85109 995887
rect 85697 995407 85753 995887
rect 86341 995407 86397 995887
rect 86893 995407 86949 995887
rect 87537 995407 87593 995887
rect 88733 995407 88789 995887
rect 89377 995407 89433 995887
rect 91217 995407 91273 995887
rect 120834 995407 120895 996693
rect 122835 996748 122896 996786
rect 122835 995407 122896 996687
rect 172034 996754 172095 996786
rect 127897 995407 127953 995887
rect 128449 995407 128505 995887
rect 129093 995407 129149 995887
rect 129737 995407 129793 995887
rect 131577 995407 131633 995887
rect 132129 995407 132185 995887
rect 132773 995407 132829 995887
rect 133417 995407 133473 995887
rect 135901 995407 135957 995887
rect 136453 995407 136509 995887
rect 137097 995407 137153 995887
rect 137741 995407 137797 995887
rect 138293 995407 138349 995887
rect 138937 995407 138993 995887
rect 140133 995407 140189 995887
rect 140777 995407 140833 995887
rect 142617 995407 142673 995887
rect 172034 995407 172095 996693
rect 174035 996757 174096 996786
rect 174035 995407 174096 996696
rect 223234 996760 223295 996786
rect 179297 995407 179353 995887
rect 179849 995407 179905 995887
rect 180493 995407 180549 995887
rect 181137 995407 181193 995887
rect 182977 995407 183033 995887
rect 183529 995407 183585 995887
rect 184173 995407 184229 995887
rect 184817 995407 184873 995887
rect 187301 995407 187357 995887
rect 187853 995407 187909 995887
rect 188497 995407 188553 995887
rect 189141 995407 189197 995887
rect 189693 995407 189749 995887
rect 190337 995407 190393 995887
rect 191533 995407 191589 995887
rect 192177 995407 192233 995887
rect 194017 995407 194073 995887
rect 223234 995407 223295 996699
rect 225235 996746 225296 996786
rect 225235 995407 225296 996685
rect 274434 996757 274495 996786
rect 230697 995407 230753 995887
rect 231249 995407 231305 995887
rect 231893 995407 231949 995887
rect 232537 995407 232593 995887
rect 234377 995407 234433 995887
rect 234929 995407 234985 995887
rect 235573 995407 235629 995887
rect 236217 995407 236273 995887
rect 238701 995407 238757 995887
rect 239253 995407 239309 995887
rect 239897 995407 239953 995887
rect 240541 995407 240597 995887
rect 241093 995407 241149 995887
rect 241737 995407 241793 995887
rect 242933 995407 242989 995887
rect 243577 995407 243633 995887
rect 245417 995407 245473 995887
rect 274434 995407 274495 996696
rect 276435 996757 276496 996786
rect 276435 995407 276496 996696
rect 378834 996763 378895 996786
rect 282297 995407 282353 995887
rect 282849 995407 282905 995887
rect 283493 995407 283549 995887
rect 284137 995407 284193 995887
rect 285977 995407 286033 995887
rect 286529 995407 286585 995887
rect 287173 995407 287229 995887
rect 287817 995407 287873 995887
rect 290301 995407 290357 995887
rect 290853 995407 290909 995887
rect 291497 995407 291553 995887
rect 292141 995407 292197 995887
rect 292693 995407 292749 995887
rect 293337 995407 293393 995887
rect 294533 995407 294589 995887
rect 295177 995407 295233 995887
rect 297017 995407 297073 995887
rect 378834 995407 378895 996702
rect 380835 996760 380896 996786
rect 380835 995407 380896 996699
rect 467834 996748 467895 996786
rect 384097 995407 384153 995887
rect 384649 995407 384705 995887
rect 385293 995407 385349 995887
rect 385937 995407 385993 995887
rect 387777 995407 387833 995887
rect 388329 995407 388385 995887
rect 388973 995407 389029 995887
rect 389617 995407 389673 995887
rect 392101 995407 392157 995887
rect 392653 995407 392709 995887
rect 393297 995407 393353 995887
rect 393941 995407 393997 995887
rect 394493 995407 394549 995887
rect 395137 995407 395193 995887
rect 396333 995407 396389 995887
rect 396977 995407 397033 995887
rect 398817 995407 398873 995887
rect 467834 995407 467895 996687
rect 469835 996751 469896 996786
rect 469835 995407 469896 996690
rect 519034 996751 519095 996786
rect 473097 995407 473153 995887
rect 473649 995407 473705 995887
rect 474293 995407 474349 995887
rect 474937 995407 474993 995887
rect 476777 995407 476833 995887
rect 477329 995407 477385 995887
rect 477973 995407 478029 995887
rect 478617 995407 478673 995887
rect 481101 995407 481157 995887
rect 481653 995407 481709 995887
rect 482297 995407 482353 995887
rect 482941 995407 482997 995887
rect 483493 995407 483549 995887
rect 484137 995407 484193 995887
rect 485333 995407 485389 995887
rect 485977 995407 486033 995887
rect 487817 995407 487873 995887
rect 519034 995407 519095 996690
rect 521035 996754 521096 996786
rect 521035 995407 521096 996693
rect 618434 996751 618495 996786
rect 524497 995407 524553 995887
rect 525049 995407 525105 995887
rect 525693 995407 525749 995887
rect 526337 995407 526393 995887
rect 528177 995407 528233 995887
rect 528729 995407 528785 995887
rect 529373 995407 529429 995887
rect 530017 995407 530073 995887
rect 532501 995407 532557 995887
rect 533053 995407 533109 995887
rect 533697 995407 533753 995887
rect 534341 995407 534397 995887
rect 534893 995407 534949 995887
rect 535537 995407 535593 995887
rect 536733 995407 536789 995887
rect 537377 995407 537433 995887
rect 539217 995407 539273 995887
rect 618434 995407 618495 996690
rect 620435 996754 620496 996786
rect 620435 995407 620496 996693
rect 626297 995407 626353 995887
rect 626849 995407 626905 995887
rect 627493 995407 627549 995887
rect 628137 995407 628193 995887
rect 629977 995407 630033 995887
rect 630529 995407 630585 995887
rect 631173 995407 631229 995887
rect 631817 995407 631873 995887
rect 634301 995407 634357 995887
rect 634853 995407 634909 995887
rect 635497 995407 635553 995887
rect 636141 995407 636197 995887
rect 636693 995407 636749 995887
rect 637337 995407 637393 995887
rect 638533 995407 638589 995887
rect 639177 995407 639233 995887
rect 641017 995407 641073 995887
rect 41863 969273 42193 969280
rect 41713 969217 42193 969273
rect 41863 969210 42193 969217
rect 41863 967433 42193 967440
rect 41713 967377 42193 967433
rect 41863 967370 42193 967377
rect 675407 967247 675887 967303
rect 41863 966789 42193 966796
rect 41713 966733 42193 966789
rect 41863 966726 42193 966733
rect 675407 966751 675737 966758
rect 675407 966695 675887 966751
rect 675407 966688 675737 966695
rect 675407 966107 675737 966114
rect 675407 966051 675887 966107
rect 675407 966044 675737 966051
rect 41863 965593 42193 965600
rect 41713 965537 42193 965593
rect 41863 965530 42193 965537
rect 675407 965463 675737 965470
rect 675407 965407 675887 965463
rect 675407 965400 675737 965407
rect 41713 964893 42193 964949
rect 41863 964397 42193 964404
rect 41713 964341 42193 964397
rect 41863 964334 42193 964341
rect 41863 963753 42193 963760
rect 41713 963697 42193 963753
rect 41863 963690 42193 963697
rect 675407 963623 675737 963630
rect 675407 963567 675887 963623
rect 675407 963560 675737 963567
rect 41863 963109 42193 963116
rect 41713 963053 42193 963109
rect 41863 963046 42193 963053
rect 675407 963071 675737 963078
rect 675407 963015 675887 963071
rect 675407 963008 675737 963015
rect 41863 962557 42193 962564
rect 41713 962501 42193 962557
rect 41863 962494 42193 962501
rect 675407 962427 675737 962434
rect 675407 962371 675887 962427
rect 675407 962364 675737 962371
rect 675407 961783 675737 961790
rect 675407 961727 675887 961783
rect 675407 961720 675737 961727
rect 41863 960073 42193 960080
rect 41713 960017 42193 960073
rect 41863 960010 42193 960017
rect 41863 959429 42193 959436
rect 41713 959373 42193 959429
rect 41863 959366 42193 959373
rect 675407 959299 675737 959306
rect 675407 959243 675887 959299
rect 675407 959236 675737 959243
rect 41863 958785 42193 958792
rect 41713 958729 42193 958785
rect 41863 958722 42193 958729
rect 675407 958747 675737 958754
rect 675407 958691 675887 958747
rect 675407 958684 675737 958691
rect 41863 958233 42193 958240
rect 41713 958177 42193 958233
rect 41863 958170 42193 958177
rect 675407 958103 675737 958110
rect 675407 958047 675887 958103
rect 675407 958040 675737 958047
rect 675407 957459 675737 957466
rect 675407 957403 675887 957459
rect 675407 957396 675737 957403
rect 675407 956851 675887 956907
rect 41863 956393 42193 956400
rect 41713 956337 42193 956393
rect 41863 956330 42193 956337
rect 675407 956263 675737 956270
rect 675407 956207 675887 956263
rect 675407 956200 675737 956207
rect 41863 955749 42193 955756
rect 41713 955693 42193 955749
rect 41863 955686 42193 955693
rect 41863 955105 42193 955112
rect 41713 955049 42193 955105
rect 41863 955042 42193 955049
rect 675407 955067 675737 955074
rect 675407 955011 675887 955067
rect 675407 955004 675737 955011
rect 41713 954497 42193 954553
rect 675407 954423 675737 954430
rect 675407 954367 675887 954423
rect 675407 954360 675737 954367
rect 675407 952583 675737 952590
rect 675407 952527 675887 952583
rect 675407 952520 675737 952527
rect 675407 878047 675887 878103
rect 675407 877551 675737 877558
rect 675407 877495 675887 877551
rect 675407 877488 675737 877495
rect 675407 876907 675737 876914
rect 675407 876851 675887 876907
rect 675407 876844 675737 876851
rect 675407 876263 675737 876270
rect 675407 876207 675887 876263
rect 675407 876200 675737 876207
rect 675407 874423 675737 874430
rect 675407 874367 675887 874423
rect 675407 874360 675737 874367
rect 675407 873871 675737 873878
rect 675407 873815 675887 873871
rect 675407 873808 675737 873815
rect 675407 873227 675737 873234
rect 675407 873171 675887 873227
rect 675407 873164 675737 873171
rect 675407 872583 675737 872590
rect 675407 872527 675887 872583
rect 675407 872520 675737 872527
rect 675407 870099 675737 870106
rect 675407 870043 675887 870099
rect 675407 870036 675737 870043
rect 675407 869547 675737 869554
rect 675407 869491 675887 869547
rect 675407 869484 675737 869491
rect 675407 868903 675737 868910
rect 675407 868847 675887 868903
rect 675407 868840 675737 868847
rect 675407 868259 675737 868266
rect 675407 868203 675887 868259
rect 675407 868196 675737 868203
rect 675407 867651 675887 867707
rect 675407 867063 675737 867070
rect 675407 867007 675887 867063
rect 675407 867000 675737 867007
rect 675407 865867 675737 865874
rect 675407 865811 675887 865867
rect 675407 865804 675737 865811
rect 675407 865223 675737 865230
rect 675407 865167 675887 865223
rect 675407 865160 675737 865167
rect 675407 863383 675737 863390
rect 675407 863327 675887 863383
rect 675407 863320 675737 863327
rect 41863 799473 42193 799480
rect 41713 799417 42193 799473
rect 41863 799410 42193 799417
rect 41863 797633 42193 797640
rect 41713 797577 42193 797633
rect 41863 797570 42193 797577
rect 41863 796989 42193 796996
rect 41713 796933 42193 796989
rect 41863 796926 42193 796933
rect 41863 795793 42193 795800
rect 41713 795737 42193 795793
rect 41863 795730 42193 795737
rect 41713 795093 42193 795149
rect 41863 794597 42193 794604
rect 41713 794541 42193 794597
rect 41863 794534 42193 794541
rect 41863 793953 42193 793960
rect 41713 793897 42193 793953
rect 41863 793890 42193 793897
rect 41863 793309 42193 793316
rect 41713 793253 42193 793309
rect 41863 793246 42193 793253
rect 41863 792757 42193 792764
rect 41713 792701 42193 792757
rect 41863 792694 42193 792701
rect 41863 790273 42193 790280
rect 41713 790217 42193 790273
rect 41863 790210 42193 790217
rect 41863 789629 42193 789636
rect 41713 789573 42193 789629
rect 41863 789566 42193 789573
rect 41863 788985 42193 788992
rect 41713 788929 42193 788985
rect 41863 788922 42193 788929
rect 675407 788847 675887 788903
rect 41863 788433 42193 788440
rect 41713 788377 42193 788433
rect 41863 788370 42193 788377
rect 675407 788351 675737 788358
rect 675407 788295 675887 788351
rect 675407 788288 675737 788295
rect 675407 787707 675737 787714
rect 675407 787651 675887 787707
rect 675407 787644 675737 787651
rect 675407 787063 675737 787070
rect 675407 787007 675887 787063
rect 675407 787000 675737 787007
rect 41863 786593 42193 786600
rect 41713 786537 42193 786593
rect 41863 786530 42193 786537
rect 41863 785949 42193 785956
rect 41713 785893 42193 785949
rect 41863 785886 42193 785893
rect 41863 785305 42193 785312
rect 41713 785249 42193 785305
rect 41863 785242 42193 785249
rect 675407 785223 675737 785230
rect 675407 785167 675887 785223
rect 675407 785160 675737 785167
rect 41713 784697 42193 784753
rect 675407 784671 675737 784678
rect 675407 784615 675887 784671
rect 675407 784608 675737 784615
rect 675407 784027 675737 784034
rect 675407 783971 675887 784027
rect 675407 783964 675737 783971
rect 675407 783383 675737 783390
rect 675407 783327 675887 783383
rect 675407 783320 675737 783327
rect 675407 780899 675737 780906
rect 675407 780843 675887 780899
rect 675407 780836 675737 780843
rect 675407 780347 675737 780354
rect 675407 780291 675887 780347
rect 675407 780284 675737 780291
rect 675407 779703 675737 779710
rect 675407 779647 675887 779703
rect 675407 779640 675737 779647
rect 675407 779059 675737 779066
rect 675407 779003 675887 779059
rect 675407 778996 675737 779003
rect 675407 778451 675887 778507
rect 675407 777863 675737 777870
rect 675407 777807 675887 777863
rect 675407 777800 675737 777807
rect 675407 776667 675737 776674
rect 675407 776611 675887 776667
rect 675407 776604 675737 776611
rect 675407 776023 675737 776030
rect 675407 775967 675887 776023
rect 675407 775960 675737 775967
rect 675407 774183 675737 774190
rect 675407 774127 675887 774183
rect 675407 774120 675737 774127
rect 41863 756273 42193 756280
rect 41713 756217 42193 756273
rect 41863 756210 42193 756217
rect 41863 754433 42193 754440
rect 41713 754377 42193 754433
rect 41863 754370 42193 754377
rect 41863 753789 42193 753796
rect 41713 753733 42193 753789
rect 41863 753726 42193 753733
rect 41863 752593 42193 752600
rect 41713 752537 42193 752593
rect 41863 752530 42193 752537
rect 41713 751893 42193 751949
rect 41863 751397 42193 751404
rect 41713 751341 42193 751397
rect 41863 751334 42193 751341
rect 41863 750753 42193 750760
rect 41713 750697 42193 750753
rect 41863 750690 42193 750697
rect 41863 750109 42193 750116
rect 41713 750053 42193 750109
rect 41863 750046 42193 750053
rect 41863 749557 42193 749564
rect 41713 749501 42193 749557
rect 41863 749494 42193 749501
rect 41863 747073 42193 747080
rect 41713 747017 42193 747073
rect 41863 747010 42193 747017
rect 41863 746429 42193 746436
rect 41713 746373 42193 746429
rect 41863 746366 42193 746373
rect 41863 745785 42193 745792
rect 41713 745729 42193 745785
rect 41863 745722 42193 745729
rect 41863 745233 42193 745240
rect 41713 745177 42193 745233
rect 41863 745170 42193 745177
rect 675407 743847 675887 743903
rect 41863 743393 42193 743400
rect 41713 743337 42193 743393
rect 41863 743330 42193 743337
rect 675407 743351 675737 743358
rect 675407 743295 675887 743351
rect 675407 743288 675737 743295
rect 41863 742749 42193 742756
rect 41713 742693 42193 742749
rect 41863 742686 42193 742693
rect 675407 742707 675737 742714
rect 675407 742651 675887 742707
rect 675407 742644 675737 742651
rect 41863 742105 42193 742112
rect 41713 742049 42193 742105
rect 41863 742042 42193 742049
rect 675407 742063 675737 742070
rect 675407 742007 675887 742063
rect 675407 742000 675737 742007
rect 41713 741497 42193 741553
rect 675407 740223 675737 740230
rect 675407 740167 675887 740223
rect 675407 740160 675737 740167
rect 675407 739671 675737 739678
rect 675407 739615 675887 739671
rect 675407 739608 675737 739615
rect 675407 739027 675737 739034
rect 675407 738971 675887 739027
rect 675407 738964 675737 738971
rect 675407 738383 675737 738390
rect 675407 738327 675887 738383
rect 675407 738320 675737 738327
rect 675407 735899 675737 735906
rect 675407 735843 675887 735899
rect 675407 735836 675737 735843
rect 675407 735347 675737 735354
rect 675407 735291 675887 735347
rect 675407 735284 675737 735291
rect 675407 734703 675737 734710
rect 675407 734647 675887 734703
rect 675407 734640 675737 734647
rect 675407 734059 675737 734066
rect 675407 734003 675887 734059
rect 675407 733996 675737 734003
rect 675407 733451 675887 733507
rect 675407 732863 675737 732870
rect 675407 732807 675887 732863
rect 675407 732800 675737 732807
rect 675407 731667 675737 731674
rect 675407 731611 675887 731667
rect 675407 731604 675737 731611
rect 675407 731023 675737 731030
rect 675407 730967 675887 731023
rect 675407 730960 675737 730967
rect 675407 729183 675737 729190
rect 675407 729127 675887 729183
rect 675407 729120 675737 729127
rect 41863 713073 42193 713080
rect 41713 713017 42193 713073
rect 41863 713010 42193 713017
rect 41863 711233 42193 711240
rect 41713 711177 42193 711233
rect 41863 711170 42193 711177
rect 41863 710589 42193 710596
rect 41713 710533 42193 710589
rect 41863 710526 42193 710533
rect 41863 709393 42193 709400
rect 41713 709337 42193 709393
rect 41863 709330 42193 709337
rect 41713 708693 42193 708749
rect 41863 708197 42193 708204
rect 41713 708141 42193 708197
rect 41863 708134 42193 708141
rect 41863 707553 42193 707560
rect 41713 707497 42193 707553
rect 41863 707490 42193 707497
rect 41863 706909 42193 706916
rect 41713 706853 42193 706909
rect 41863 706846 42193 706853
rect 41863 706357 42193 706364
rect 41713 706301 42193 706357
rect 41863 706294 42193 706301
rect 41863 703873 42193 703880
rect 41713 703817 42193 703873
rect 41863 703810 42193 703817
rect 41863 703229 42193 703236
rect 41713 703173 42193 703229
rect 41863 703166 42193 703173
rect 41863 702585 42193 702592
rect 41713 702529 42193 702585
rect 41863 702522 42193 702529
rect 41863 702033 42193 702040
rect 41713 701977 42193 702033
rect 41863 701970 42193 701977
rect 41863 700193 42193 700200
rect 41713 700137 42193 700193
rect 41863 700130 42193 700137
rect 41863 699549 42193 699556
rect 41713 699493 42193 699549
rect 41863 699486 42193 699493
rect 41863 698905 42193 698912
rect 41713 698849 42193 698905
rect 41863 698842 42193 698849
rect 675407 698847 675887 698903
rect 41713 698297 42193 698353
rect 675407 698351 675737 698358
rect 675407 698295 675887 698351
rect 675407 698288 675737 698295
rect 675407 697707 675737 697714
rect 675407 697651 675887 697707
rect 675407 697644 675737 697651
rect 675407 697063 675737 697070
rect 675407 697007 675887 697063
rect 675407 697000 675737 697007
rect 675407 695223 675737 695230
rect 675407 695167 675887 695223
rect 675407 695160 675737 695167
rect 675407 694671 675737 694678
rect 675407 694615 675887 694671
rect 675407 694608 675737 694615
rect 675407 694027 675737 694034
rect 675407 693971 675887 694027
rect 675407 693964 675737 693971
rect 675407 693383 675737 693390
rect 675407 693327 675887 693383
rect 675407 693320 675737 693327
rect 675407 690899 675737 690906
rect 675407 690843 675887 690899
rect 675407 690836 675737 690843
rect 675407 690347 675737 690354
rect 675407 690291 675887 690347
rect 675407 690284 675737 690291
rect 675407 689703 675737 689710
rect 675407 689647 675887 689703
rect 675407 689640 675737 689647
rect 675407 689059 675737 689066
rect 675407 689003 675887 689059
rect 675407 688996 675737 689003
rect 675407 688451 675887 688507
rect 675407 687863 675737 687870
rect 675407 687807 675887 687863
rect 675407 687800 675737 687807
rect 675407 686667 675737 686674
rect 675407 686611 675887 686667
rect 675407 686604 675737 686611
rect 675407 686023 675737 686030
rect 675407 685967 675887 686023
rect 675407 685960 675737 685967
rect 675407 684183 675737 684190
rect 675407 684127 675887 684183
rect 675407 684120 675737 684127
rect 41863 669873 42193 669880
rect 41713 669817 42193 669873
rect 41863 669810 42193 669817
rect 41863 668033 42193 668040
rect 41713 667977 42193 668033
rect 41863 667970 42193 667977
rect 41863 667389 42193 667396
rect 41713 667333 42193 667389
rect 41863 667326 42193 667333
rect 41863 666193 42193 666200
rect 41713 666137 42193 666193
rect 41863 666130 42193 666137
rect 41713 665493 42193 665549
rect 41863 664997 42193 665004
rect 41713 664941 42193 664997
rect 41863 664934 42193 664941
rect 41863 664353 42193 664360
rect 41713 664297 42193 664353
rect 41863 664290 42193 664297
rect 41863 663709 42193 663716
rect 41713 663653 42193 663709
rect 41863 663646 42193 663653
rect 41863 663157 42193 663164
rect 41713 663101 42193 663157
rect 41863 663094 42193 663101
rect 41863 660673 42193 660680
rect 41713 660617 42193 660673
rect 41863 660610 42193 660617
rect 41863 660029 42193 660036
rect 41713 659973 42193 660029
rect 41863 659966 42193 659973
rect 41863 659385 42193 659392
rect 41713 659329 42193 659385
rect 41863 659322 42193 659329
rect 41863 658833 42193 658840
rect 41713 658777 42193 658833
rect 41863 658770 42193 658777
rect 41863 656993 42193 657000
rect 41713 656937 42193 656993
rect 41863 656930 42193 656937
rect 41863 656349 42193 656356
rect 41713 656293 42193 656349
rect 41863 656286 42193 656293
rect 41863 655705 42193 655712
rect 41713 655649 42193 655705
rect 41863 655642 42193 655649
rect 41713 655097 42193 655153
rect 675407 653647 675887 653703
rect 675407 653151 675737 653158
rect 675407 653095 675887 653151
rect 675407 653088 675737 653095
rect 675407 652507 675737 652514
rect 675407 652451 675887 652507
rect 675407 652444 675737 652451
rect 675407 651863 675737 651870
rect 675407 651807 675887 651863
rect 675407 651800 675737 651807
rect 675407 650023 675737 650030
rect 675407 649967 675887 650023
rect 675407 649960 675737 649967
rect 675407 649471 675737 649478
rect 675407 649415 675887 649471
rect 675407 649408 675737 649415
rect 675407 648827 675737 648834
rect 675407 648771 675887 648827
rect 675407 648764 675737 648771
rect 675407 648183 675737 648190
rect 675407 648127 675887 648183
rect 675407 648120 675737 648127
rect 675407 645699 675737 645706
rect 675407 645643 675887 645699
rect 675407 645636 675737 645643
rect 675407 645147 675737 645154
rect 675407 645091 675887 645147
rect 675407 645084 675737 645091
rect 675407 644503 675737 644510
rect 675407 644447 675887 644503
rect 675407 644440 675737 644447
rect 675407 643859 675737 643866
rect 675407 643803 675887 643859
rect 675407 643796 675737 643803
rect 675407 643251 675887 643307
rect 675407 642663 675737 642670
rect 675407 642607 675887 642663
rect 675407 642600 675737 642607
rect 675407 641467 675737 641474
rect 675407 641411 675887 641467
rect 675407 641404 675737 641411
rect 675407 640823 675737 640830
rect 675407 640767 675887 640823
rect 675407 640760 675737 640767
rect 675407 638983 675737 638990
rect 675407 638927 675887 638983
rect 675407 638920 675737 638927
rect 41863 626673 42193 626680
rect 41713 626617 42193 626673
rect 41863 626610 42193 626617
rect 41863 624833 42193 624840
rect 41713 624777 42193 624833
rect 41863 624770 42193 624777
rect 41863 624189 42193 624196
rect 41713 624133 42193 624189
rect 41863 624126 42193 624133
rect 41863 622993 42193 623000
rect 41713 622937 42193 622993
rect 41863 622930 42193 622937
rect 41713 622293 42193 622349
rect 41863 621797 42193 621804
rect 41713 621741 42193 621797
rect 41863 621734 42193 621741
rect 41863 621153 42193 621160
rect 41713 621097 42193 621153
rect 41863 621090 42193 621097
rect 41863 620509 42193 620516
rect 41713 620453 42193 620509
rect 41863 620446 42193 620453
rect 41863 619957 42193 619964
rect 41713 619901 42193 619957
rect 41863 619894 42193 619901
rect 41863 617473 42193 617480
rect 41713 617417 42193 617473
rect 41863 617410 42193 617417
rect 41863 616829 42193 616836
rect 41713 616773 42193 616829
rect 41863 616766 42193 616773
rect 41863 616185 42193 616192
rect 41713 616129 42193 616185
rect 41863 616122 42193 616129
rect 41863 615633 42193 615640
rect 41713 615577 42193 615633
rect 41863 615570 42193 615577
rect 41863 613793 42193 613800
rect 41713 613737 42193 613793
rect 41863 613730 42193 613737
rect 41863 613149 42193 613156
rect 41713 613093 42193 613149
rect 41863 613086 42193 613093
rect 41863 612505 42193 612512
rect 41713 612449 42193 612505
rect 41863 612442 42193 612449
rect 41713 611897 42193 611953
rect 675407 608647 675887 608703
rect 675407 608151 675737 608158
rect 675407 608095 675887 608151
rect 675407 608088 675737 608095
rect 675407 607507 675737 607514
rect 675407 607451 675887 607507
rect 675407 607444 675737 607451
rect 675407 606863 675737 606870
rect 675407 606807 675887 606863
rect 675407 606800 675737 606807
rect 675407 605023 675737 605030
rect 675407 604967 675887 605023
rect 675407 604960 675737 604967
rect 675407 604471 675737 604478
rect 675407 604415 675887 604471
rect 675407 604408 675737 604415
rect 675407 603827 675737 603834
rect 675407 603771 675887 603827
rect 675407 603764 675737 603771
rect 675407 603183 675737 603190
rect 675407 603127 675887 603183
rect 675407 603120 675737 603127
rect 675407 600699 675737 600706
rect 675407 600643 675887 600699
rect 675407 600636 675737 600643
rect 675407 600147 675737 600154
rect 675407 600091 675887 600147
rect 675407 600084 675737 600091
rect 675407 599503 675737 599510
rect 675407 599447 675887 599503
rect 675407 599440 675737 599447
rect 675407 598859 675737 598866
rect 675407 598803 675887 598859
rect 675407 598796 675737 598803
rect 675407 597663 675737 597670
rect 675407 597607 675887 597663
rect 675407 597600 675737 597607
rect 675407 596467 675737 596474
rect 675407 596411 675887 596467
rect 675407 596404 675737 596411
rect 675407 595823 675737 595830
rect 675407 595767 675887 595823
rect 675407 595760 675737 595767
rect 675407 593983 675737 593990
rect 675407 593927 675887 593983
rect 675407 593920 675737 593927
rect 41863 583473 42193 583480
rect 41713 583417 42193 583473
rect 41863 583410 42193 583417
rect 41863 581633 42193 581640
rect 41713 581577 42193 581633
rect 41863 581570 42193 581577
rect 41863 580989 42193 580996
rect 41713 580933 42193 580989
rect 41863 580926 42193 580933
rect 41863 579793 42193 579800
rect 41713 579737 42193 579793
rect 41863 579730 42193 579737
rect 41713 579093 42193 579149
rect 41863 578597 42193 578604
rect 41713 578541 42193 578597
rect 41863 578534 42193 578541
rect 41863 577953 42193 577960
rect 41713 577897 42193 577953
rect 41863 577890 42193 577897
rect 41863 577309 42193 577316
rect 41713 577253 42193 577309
rect 41863 577246 42193 577253
rect 41863 576757 42193 576764
rect 41713 576701 42193 576757
rect 41863 576694 42193 576701
rect 41863 574273 42193 574280
rect 41713 574217 42193 574273
rect 41863 574210 42193 574217
rect 41863 573629 42193 573636
rect 41713 573573 42193 573629
rect 41863 573566 42193 573573
rect 41863 572985 42193 572992
rect 41713 572929 42193 572985
rect 41863 572922 42193 572929
rect 41863 572433 42193 572440
rect 41713 572377 42193 572433
rect 41863 572370 42193 572377
rect 41863 570593 42193 570600
rect 41713 570537 42193 570593
rect 41863 570530 42193 570537
rect 41863 569949 42193 569956
rect 41713 569893 42193 569949
rect 41863 569886 42193 569893
rect 41863 569305 42193 569312
rect 41713 569249 42193 569305
rect 41863 569242 42193 569249
rect 41713 568697 42193 568753
rect 675407 563447 675887 563503
rect 675407 562951 675737 562958
rect 675407 562895 675887 562951
rect 675407 562888 675737 562895
rect 675407 562307 675737 562314
rect 675407 562251 675887 562307
rect 675407 562244 675737 562251
rect 675407 561663 675737 561670
rect 675407 561607 675887 561663
rect 675407 561600 675737 561607
rect 675407 559823 675737 559830
rect 675407 559767 675887 559823
rect 675407 559760 675737 559767
rect 675407 559271 675737 559278
rect 675407 559215 675887 559271
rect 675407 559208 675737 559215
rect 675407 558627 675737 558634
rect 675407 558571 675887 558627
rect 675407 558564 675737 558571
rect 675407 557983 675737 557990
rect 675407 557927 675887 557983
rect 675407 557920 675737 557927
rect 675407 555499 675737 555506
rect 675407 555443 675887 555499
rect 675407 555436 675737 555443
rect 675407 554947 675737 554954
rect 675407 554891 675887 554947
rect 675407 554884 675737 554891
rect 675407 554303 675737 554310
rect 675407 554247 675887 554303
rect 675407 554240 675737 554247
rect 675407 553659 675737 553666
rect 675407 553603 675887 553659
rect 675407 553596 675737 553603
rect 675407 553051 675887 553107
rect 675407 552463 675737 552470
rect 675407 552407 675887 552463
rect 675407 552400 675737 552407
rect 675407 551267 675737 551274
rect 675407 551211 675887 551267
rect 675407 551204 675737 551211
rect 675407 550623 675737 550630
rect 675407 550567 675887 550623
rect 675407 550560 675737 550567
rect 675407 548783 675737 548790
rect 675407 548727 675887 548783
rect 675407 548720 675737 548727
rect 41863 540273 42193 540280
rect 41713 540217 42193 540273
rect 41863 540210 42193 540217
rect 41863 538433 42193 538440
rect 41713 538377 42193 538433
rect 41863 538370 42193 538377
rect 41863 537789 42193 537796
rect 41713 537733 42193 537789
rect 41863 537726 42193 537733
rect 41863 536593 42193 536600
rect 41713 536537 42193 536593
rect 41863 536530 42193 536537
rect 41713 535893 42193 535949
rect 41863 535397 42193 535404
rect 41713 535341 42193 535397
rect 41863 535334 42193 535341
rect 41863 534753 42193 534760
rect 41713 534697 42193 534753
rect 41863 534690 42193 534697
rect 41863 534109 42193 534116
rect 41713 534053 42193 534109
rect 41863 534046 42193 534053
rect 41863 533557 42193 533564
rect 41713 533501 42193 533557
rect 41863 533494 42193 533501
rect 41863 531073 42193 531080
rect 41713 531017 42193 531073
rect 41863 531010 42193 531017
rect 41863 530429 42193 530436
rect 41713 530373 42193 530429
rect 41863 530366 42193 530373
rect 41863 529785 42193 529792
rect 41713 529729 42193 529785
rect 41863 529722 42193 529729
rect 41863 529233 42193 529240
rect 41713 529177 42193 529233
rect 41863 529170 42193 529177
rect 41863 527393 42193 527400
rect 41713 527337 42193 527393
rect 41863 527330 42193 527337
rect 41863 526749 42193 526756
rect 41713 526693 42193 526749
rect 41863 526686 42193 526693
rect 41863 526105 42193 526112
rect 41713 526049 42193 526105
rect 41863 526042 42193 526049
rect 41713 525497 42193 525553
rect 41863 412673 42193 412680
rect 41713 412617 42193 412673
rect 41863 412610 42193 412617
rect 41863 410833 42193 410840
rect 41713 410777 42193 410833
rect 41863 410770 42193 410777
rect 41863 410189 42193 410196
rect 41713 410133 42193 410189
rect 41863 410126 42193 410133
rect 41863 408993 42193 409000
rect 41713 408937 42193 408993
rect 41863 408930 42193 408937
rect 41713 408293 42193 408349
rect 41863 407797 42193 407804
rect 41713 407741 42193 407797
rect 41863 407734 42193 407741
rect 41863 407153 42193 407160
rect 41713 407097 42193 407153
rect 41863 407090 42193 407097
rect 41863 406509 42193 406516
rect 41713 406453 42193 406509
rect 41863 406446 42193 406453
rect 41863 405957 42193 405964
rect 41713 405901 42193 405957
rect 41863 405894 42193 405901
rect 41863 403473 42193 403480
rect 41713 403417 42193 403473
rect 41863 403410 42193 403417
rect 41863 402829 42193 402836
rect 41713 402773 42193 402829
rect 41863 402766 42193 402773
rect 41863 402185 42193 402192
rect 41713 402129 42193 402185
rect 41863 402122 42193 402129
rect 41863 401633 42193 401640
rect 41713 401577 42193 401633
rect 41863 401570 42193 401577
rect 41863 399793 42193 399800
rect 41713 399737 42193 399793
rect 41863 399730 42193 399737
rect 41863 399149 42193 399156
rect 41713 399093 42193 399149
rect 41863 399086 42193 399093
rect 41863 398505 42193 398512
rect 41713 398449 42193 398505
rect 41863 398442 42193 398449
rect 41713 397897 42193 397953
rect 675407 386247 675887 386303
rect 675407 385751 675737 385758
rect 675407 385695 675887 385751
rect 675407 385688 675737 385695
rect 675407 385107 675737 385114
rect 675407 385051 675887 385107
rect 675407 385044 675737 385051
rect 675407 384463 675737 384470
rect 675407 384407 675887 384463
rect 675407 384400 675737 384407
rect 675407 382623 675737 382630
rect 675407 382567 675887 382623
rect 675407 382560 675737 382567
rect 675407 382071 675737 382078
rect 675407 382015 675887 382071
rect 675407 382008 675737 382015
rect 675407 381427 675737 381434
rect 675407 381371 675887 381427
rect 675407 381364 675737 381371
rect 675407 380783 675737 380790
rect 675407 380727 675887 380783
rect 675407 380720 675737 380727
rect 675407 378299 675737 378306
rect 675407 378243 675887 378299
rect 675407 378236 675737 378243
rect 675407 377747 675737 377754
rect 675407 377691 675887 377747
rect 675407 377684 675737 377691
rect 675407 377103 675737 377110
rect 675407 377047 675887 377103
rect 675407 377040 675737 377047
rect 675407 376459 675737 376466
rect 675407 376403 675887 376459
rect 675407 376396 675737 376403
rect 675407 375851 675887 375907
rect 675407 375263 675737 375270
rect 675407 375207 675887 375263
rect 675407 375200 675737 375207
rect 675407 374011 675887 374067
rect 675407 373423 675737 373430
rect 675407 373367 675887 373423
rect 675407 373360 675737 373367
rect 675407 371583 675737 371590
rect 675407 371527 675887 371583
rect 675407 371520 675737 371527
rect 41863 369473 42193 369480
rect 41713 369417 42193 369473
rect 41863 369410 42193 369417
rect 41863 367633 42193 367640
rect 41713 367577 42193 367633
rect 41863 367570 42193 367577
rect 41863 366989 42193 366996
rect 41713 366933 42193 366989
rect 41863 366926 42193 366933
rect 41863 365793 42193 365800
rect 41713 365737 42193 365793
rect 41863 365730 42193 365737
rect 41713 365093 42193 365149
rect 41863 364597 42193 364604
rect 41713 364541 42193 364597
rect 41863 364534 42193 364541
rect 41863 363953 42193 363960
rect 41713 363897 42193 363953
rect 41863 363890 42193 363897
rect 41863 363309 42193 363316
rect 41713 363253 42193 363309
rect 41863 363246 42193 363253
rect 41863 362757 42193 362764
rect 41713 362701 42193 362757
rect 41863 362694 42193 362701
rect 41863 360273 42193 360280
rect 41713 360217 42193 360273
rect 41863 360210 42193 360217
rect 41863 359629 42193 359636
rect 41713 359573 42193 359629
rect 41863 359566 42193 359573
rect 41863 358985 42193 358992
rect 41713 358929 42193 358985
rect 41863 358922 42193 358929
rect 41863 358433 42193 358440
rect 41713 358377 42193 358433
rect 41863 358370 42193 358377
rect 41863 356593 42193 356600
rect 41713 356537 42193 356593
rect 41863 356530 42193 356537
rect 41863 355949 42193 355956
rect 41713 355893 42193 355949
rect 41863 355886 42193 355893
rect 41863 355305 42193 355312
rect 41713 355249 42193 355305
rect 41863 355242 42193 355249
rect 41713 354697 42193 354753
rect 675407 341047 675887 341103
rect 675407 340551 675737 340558
rect 675407 340495 675887 340551
rect 675407 340488 675737 340495
rect 675407 339907 675737 339914
rect 675407 339851 675887 339907
rect 675407 339844 675737 339851
rect 675407 339263 675737 339270
rect 675407 339207 675887 339263
rect 675407 339200 675737 339207
rect 675407 337423 675737 337430
rect 675407 337367 675887 337423
rect 675407 337360 675737 337367
rect 675407 336871 675737 336878
rect 675407 336815 675887 336871
rect 675407 336808 675737 336815
rect 675407 336227 675737 336234
rect 675407 336171 675887 336227
rect 675407 336164 675737 336171
rect 675407 335583 675737 335590
rect 675407 335527 675887 335583
rect 675407 335520 675737 335527
rect 675407 333099 675737 333106
rect 675407 333043 675887 333099
rect 675407 333036 675737 333043
rect 675407 332547 675737 332554
rect 675407 332491 675887 332547
rect 675407 332484 675737 332491
rect 675407 331903 675737 331910
rect 675407 331847 675887 331903
rect 675407 331840 675737 331847
rect 675407 331259 675737 331266
rect 675407 331203 675887 331259
rect 675407 331196 675737 331203
rect 675407 330651 675887 330707
rect 675407 330063 675737 330070
rect 675407 330007 675887 330063
rect 675407 330000 675737 330007
rect 675407 328811 675887 328867
rect 675407 328223 675737 328230
rect 675407 328167 675887 328223
rect 675407 328160 675737 328167
rect 675407 326383 675737 326390
rect 675407 326327 675887 326383
rect 675407 326320 675737 326327
rect 41863 326273 42193 326280
rect 41713 326217 42193 326273
rect 41863 326210 42193 326217
rect 41863 324433 42193 324440
rect 41713 324377 42193 324433
rect 41863 324370 42193 324377
rect 41863 323789 42193 323796
rect 41713 323733 42193 323789
rect 41863 323726 42193 323733
rect 41863 322593 42193 322600
rect 41713 322537 42193 322593
rect 41863 322530 42193 322537
rect 41713 321893 42193 321949
rect 41863 321397 42193 321404
rect 41713 321341 42193 321397
rect 41863 321334 42193 321341
rect 41863 320753 42193 320760
rect 41713 320697 42193 320753
rect 41863 320690 42193 320697
rect 41863 320109 42193 320116
rect 41713 320053 42193 320109
rect 41863 320046 42193 320053
rect 41863 319557 42193 319564
rect 41713 319501 42193 319557
rect 41863 319494 42193 319501
rect 41863 317073 42193 317080
rect 41713 317017 42193 317073
rect 41863 317010 42193 317017
rect 41863 316429 42193 316436
rect 41713 316373 42193 316429
rect 41863 316366 42193 316373
rect 41863 315785 42193 315792
rect 41713 315729 42193 315785
rect 41863 315722 42193 315729
rect 41863 315233 42193 315240
rect 41713 315177 42193 315233
rect 41863 315170 42193 315177
rect 41863 313393 42193 313400
rect 41713 313337 42193 313393
rect 41863 313330 42193 313337
rect 41863 312749 42193 312756
rect 41713 312693 42193 312749
rect 41863 312686 42193 312693
rect 41863 312105 42193 312112
rect 41713 312049 42193 312105
rect 41863 312042 42193 312049
rect 41713 311497 42193 311553
rect 675407 296047 675887 296103
rect 675407 295551 675737 295558
rect 675407 295495 675887 295551
rect 675407 295488 675737 295495
rect 675407 294907 675737 294914
rect 675407 294851 675887 294907
rect 675407 294844 675737 294851
rect 675407 294263 675737 294270
rect 675407 294207 675887 294263
rect 675407 294200 675737 294207
rect 675407 292423 675737 292430
rect 675407 292367 675887 292423
rect 675407 292360 675737 292367
rect 675407 291871 675737 291878
rect 675407 291815 675887 291871
rect 675407 291808 675737 291815
rect 675407 291227 675737 291234
rect 675407 291171 675887 291227
rect 675407 291164 675737 291171
rect 675407 290583 675737 290590
rect 675407 290527 675887 290583
rect 675407 290520 675737 290527
rect 675407 288099 675737 288106
rect 675407 288043 675887 288099
rect 675407 288036 675737 288043
rect 675407 287547 675737 287554
rect 675407 287491 675887 287547
rect 675407 287484 675737 287491
rect 675407 286903 675737 286910
rect 675407 286847 675887 286903
rect 675407 286840 675737 286847
rect 675407 286259 675737 286266
rect 675407 286203 675887 286259
rect 675407 286196 675737 286203
rect 675407 285651 675887 285707
rect 675407 285063 675737 285070
rect 675407 285007 675887 285063
rect 675407 285000 675737 285007
rect 675407 283811 675887 283867
rect 675407 283223 675737 283230
rect 675407 283167 675887 283223
rect 675407 283160 675737 283167
rect 41863 283073 42193 283080
rect 41713 283017 42193 283073
rect 41863 283010 42193 283017
rect 675407 281383 675737 281390
rect 675407 281327 675887 281383
rect 675407 281320 675737 281327
rect 41863 281233 42193 281240
rect 41713 281177 42193 281233
rect 41863 281170 42193 281177
rect 41863 280589 42193 280596
rect 41713 280533 42193 280589
rect 41863 280526 42193 280533
rect 41863 279393 42193 279400
rect 41713 279337 42193 279393
rect 41863 279330 42193 279337
rect 41713 278693 42193 278749
rect 41863 278197 42193 278204
rect 41713 278141 42193 278197
rect 41863 278134 42193 278141
rect 41863 277553 42193 277560
rect 41713 277497 42193 277553
rect 41863 277490 42193 277497
rect 41863 276909 42193 276916
rect 41713 276853 42193 276909
rect 41863 276846 42193 276853
rect 41863 276357 42193 276364
rect 41713 276301 42193 276357
rect 41863 276294 42193 276301
rect 41863 273873 42193 273880
rect 41713 273817 42193 273873
rect 41863 273810 42193 273817
rect 41863 273229 42193 273236
rect 41713 273173 42193 273229
rect 41863 273166 42193 273173
rect 41863 272585 42193 272592
rect 41713 272529 42193 272585
rect 41863 272522 42193 272529
rect 41863 272033 42193 272040
rect 41713 271977 42193 272033
rect 41863 271970 42193 271977
rect 41863 270193 42193 270200
rect 41713 270137 42193 270193
rect 41863 270130 42193 270137
rect 41863 269549 42193 269556
rect 41713 269493 42193 269549
rect 41863 269486 42193 269493
rect 41863 268905 42193 268912
rect 41713 268849 42193 268905
rect 41863 268842 42193 268849
rect 41713 268297 42193 268353
rect 675407 251047 675887 251103
rect 675407 250551 675737 250558
rect 675407 250495 675887 250551
rect 675407 250488 675737 250495
rect 675407 249907 675737 249914
rect 675407 249851 675887 249907
rect 675407 249844 675737 249851
rect 675407 249263 675737 249270
rect 675407 249207 675887 249263
rect 675407 249200 675737 249207
rect 675407 247423 675737 247430
rect 675407 247367 675887 247423
rect 675407 247360 675737 247367
rect 675407 246871 675737 246878
rect 675407 246815 675887 246871
rect 675407 246808 675737 246815
rect 675407 246227 675737 246234
rect 675407 246171 675887 246227
rect 675407 246164 675737 246171
rect 675407 245583 675737 245590
rect 675407 245527 675887 245583
rect 675407 245520 675737 245527
rect 675407 243099 675737 243106
rect 675407 243043 675887 243099
rect 675407 243036 675737 243043
rect 675407 242547 675737 242554
rect 675407 242491 675887 242547
rect 675407 242484 675737 242491
rect 675407 241903 675737 241910
rect 675407 241847 675887 241903
rect 675407 241840 675737 241847
rect 675407 241259 675737 241266
rect 675407 241203 675887 241259
rect 675407 241196 675737 241203
rect 675407 240651 675887 240707
rect 675407 240063 675737 240070
rect 675407 240007 675887 240063
rect 675407 240000 675737 240007
rect 41863 239873 42193 239880
rect 41713 239817 42193 239873
rect 41863 239810 42193 239817
rect 675407 238811 675887 238867
rect 675407 238223 675737 238230
rect 675407 238167 675887 238223
rect 675407 238160 675737 238167
rect 41863 238033 42193 238040
rect 41713 237977 42193 238033
rect 41863 237970 42193 237977
rect 41713 237333 42193 237389
rect 675407 236383 675737 236390
rect 675407 236327 675887 236383
rect 675407 236320 675737 236327
rect 41863 236193 42193 236200
rect 41713 236137 42193 236193
rect 41863 236130 42193 236137
rect 41713 235493 42193 235549
rect 41863 234997 42193 235004
rect 41713 234941 42193 234997
rect 41863 234934 42193 234941
rect 41863 234353 42193 234360
rect 41713 234297 42193 234353
rect 41863 234290 42193 234297
rect 41863 233709 42193 233716
rect 41713 233653 42193 233709
rect 41863 233646 42193 233653
rect 41863 233157 42193 233164
rect 41713 233101 42193 233157
rect 41863 233094 42193 233101
rect 41863 230673 42193 230680
rect 41713 230617 42193 230673
rect 41863 230610 42193 230617
rect 41863 230029 42193 230036
rect 41713 229973 42193 230029
rect 41863 229966 42193 229973
rect 41863 229385 42193 229392
rect 41713 229329 42193 229385
rect 41863 229322 42193 229329
rect 41863 228833 42193 228840
rect 41713 228777 42193 228833
rect 41863 228770 42193 228777
rect 41863 226993 42193 227000
rect 41713 226937 42193 226993
rect 41863 226930 42193 226937
rect 41863 226349 42193 226356
rect 41713 226293 42193 226349
rect 41863 226286 42193 226293
rect 41863 225705 42193 225712
rect 41713 225649 42193 225705
rect 41863 225642 42193 225649
rect 41713 225097 42193 225153
rect 675407 205847 675887 205903
rect 675407 205351 675737 205358
rect 675407 205295 675887 205351
rect 675407 205288 675737 205295
rect 675407 204707 675737 204714
rect 675407 204651 675887 204707
rect 675407 204644 675737 204651
rect 675407 204063 675737 204070
rect 675407 204007 675887 204063
rect 675407 204000 675737 204007
rect 675407 202223 675737 202230
rect 675407 202167 675887 202223
rect 675407 202160 675737 202167
rect 675407 201671 675737 201678
rect 675407 201615 675887 201671
rect 675407 201608 675737 201615
rect 675407 201027 675737 201034
rect 675407 200971 675887 201027
rect 675407 200964 675737 200971
rect 675407 200383 675737 200390
rect 675407 200327 675887 200383
rect 675407 200320 675737 200327
rect 675407 197899 675737 197906
rect 675407 197843 675887 197899
rect 675407 197836 675737 197843
rect 675407 197347 675737 197354
rect 675407 197291 675887 197347
rect 675407 197284 675737 197291
rect 675407 196703 675737 196710
rect 41863 196673 42193 196680
rect 41713 196617 42193 196673
rect 675407 196647 675887 196703
rect 675407 196640 675737 196647
rect 41863 196610 42193 196617
rect 675407 196059 675737 196066
rect 675407 196003 675887 196059
rect 675407 195996 675737 196003
rect 675407 195451 675887 195507
rect 675407 194863 675737 194870
rect 41863 194833 42193 194840
rect 41713 194777 42193 194833
rect 675407 194807 675887 194863
rect 675407 194800 675737 194807
rect 41863 194770 42193 194777
rect 41713 194133 42193 194189
rect 675407 193611 675887 193667
rect 675407 193023 675737 193030
rect 41863 192993 42193 193000
rect 41713 192937 42193 192993
rect 675407 192967 675887 193023
rect 675407 192960 675737 192967
rect 41863 192930 42193 192937
rect 41713 192293 42193 192349
rect 41863 191797 42193 191804
rect 41713 191741 42193 191797
rect 41863 191734 42193 191741
rect 675407 191183 675737 191190
rect 41863 191153 42193 191160
rect 41713 191097 42193 191153
rect 675407 191127 675887 191183
rect 675407 191120 675737 191127
rect 41863 191090 42193 191097
rect 41863 190509 42193 190516
rect 41713 190453 42193 190509
rect 41863 190446 42193 190453
rect 41863 189957 42193 189964
rect 41713 189901 42193 189957
rect 41863 189894 42193 189901
rect 41863 187473 42193 187480
rect 41713 187417 42193 187473
rect 41863 187410 42193 187417
rect 41863 186829 42193 186836
rect 41713 186773 42193 186829
rect 41863 186766 42193 186773
rect 41863 186185 42193 186192
rect 41713 186129 42193 186185
rect 41863 186122 42193 186129
rect 41863 185633 42193 185640
rect 41713 185577 42193 185633
rect 41863 185570 42193 185577
rect 41863 183793 42193 183800
rect 41713 183737 42193 183793
rect 41863 183730 42193 183737
rect 41863 183149 42193 183156
rect 41713 183093 42193 183149
rect 41863 183086 42193 183093
rect 41863 182505 42193 182512
rect 41713 182449 42193 182505
rect 41863 182442 42193 182449
rect 41713 181897 42193 181953
rect 675407 160847 675887 160903
rect 675407 160351 675737 160358
rect 675407 160295 675887 160351
rect 675407 160288 675737 160295
rect 675407 159707 675737 159714
rect 675407 159651 675887 159707
rect 675407 159644 675737 159651
rect 675407 159063 675737 159070
rect 675407 159007 675887 159063
rect 675407 159000 675737 159007
rect 675407 157223 675737 157230
rect 675407 157167 675887 157223
rect 675407 157160 675737 157167
rect 675407 156671 675737 156678
rect 675407 156615 675887 156671
rect 675407 156608 675737 156615
rect 675407 156027 675737 156034
rect 675407 155971 675887 156027
rect 675407 155964 675737 155971
rect 675407 155383 675737 155390
rect 675407 155327 675887 155383
rect 675407 155320 675737 155327
rect 675407 152899 675737 152906
rect 675407 152843 675887 152899
rect 675407 152836 675737 152843
rect 675407 152347 675737 152354
rect 675407 152291 675887 152347
rect 675407 152284 675737 152291
rect 675407 151703 675737 151710
rect 675407 151647 675887 151703
rect 675407 151640 675737 151647
rect 675407 151059 675737 151066
rect 675407 151003 675887 151059
rect 675407 150996 675737 151003
rect 675407 150451 675887 150507
rect 675407 149863 675737 149870
rect 675407 149807 675887 149863
rect 675407 149800 675737 149807
rect 675407 148611 675887 148667
rect 675407 148023 675737 148030
rect 675407 147967 675887 148023
rect 675407 147960 675737 147967
rect 675407 147379 675737 147386
rect 675407 147323 675887 147379
rect 675407 147316 675737 147323
rect 675407 146183 675737 146190
rect 675407 146127 675887 146183
rect 675407 146120 675737 146127
rect 675407 115647 675887 115703
rect 675407 115151 675737 115158
rect 675407 115095 675887 115151
rect 675407 115088 675737 115095
rect 675407 114507 675737 114514
rect 675407 114451 675887 114507
rect 675407 114444 675737 114451
rect 675407 113863 675737 113870
rect 675407 113807 675887 113863
rect 675407 113800 675737 113807
rect 675407 112023 675737 112030
rect 675407 111967 675887 112023
rect 675407 111960 675737 111967
rect 675407 111471 675737 111478
rect 675407 111415 675887 111471
rect 675407 111408 675737 111415
rect 675407 110827 675737 110834
rect 675407 110771 675887 110827
rect 675407 110764 675737 110771
rect 675407 110183 675737 110190
rect 675407 110127 675887 110183
rect 675407 110120 675737 110127
rect 675407 107699 675737 107706
rect 675407 107643 675887 107699
rect 675407 107636 675737 107643
rect 675407 107147 675737 107154
rect 675407 107091 675887 107147
rect 675407 107084 675737 107091
rect 675407 106503 675737 106510
rect 675407 106447 675887 106503
rect 675407 106440 675737 106447
rect 675407 105859 675737 105866
rect 675407 105803 675887 105859
rect 675407 105796 675737 105803
rect 675407 105251 675887 105307
rect 675407 104663 675737 104670
rect 675407 104607 675887 104663
rect 675407 104600 675737 104607
rect 675407 103411 675887 103467
rect 675407 102823 675737 102830
rect 675407 102767 675887 102823
rect 675407 102760 675737 102767
rect 675407 100983 675737 100990
rect 675407 100927 675887 100983
rect 675407 100920 675737 100927
rect 18917 95739 18934 95795
rect 19194 95739 41478 95795
rect 41829 95739 41845 95795
rect 18555 95515 18569 95571
rect 18829 95515 41470 95571
rect 41821 95515 41845 95571
rect 17829 95291 17843 95347
rect 18112 95291 41467 95347
rect 41835 95291 41845 95347
rect 141708 42047 141774 42193
rect 141710 40350 141771 42047
rect 145035 41918 145207 41924
rect 145035 41866 145063 41918
rect 145115 41866 145127 41918
rect 145179 41866 145207 41918
rect 145035 41860 145207 41866
rect 140996 40125 141048 40131
rect 140996 40067 141048 40073
rect 141004 39990 141042 40067
rect 141710 40000 141771 40289
rect 141992 40125 142044 40131
rect 141986 40073 141992 40120
rect 143068 40125 143120 40131
rect 142044 40073 142050 40120
rect 141986 39998 142050 40073
rect 143407 40125 143519 40131
rect 143407 40090 143437 40125
rect 143489 40090 143519 40125
rect 144603 40125 144655 40131
rect 143068 40067 143120 40073
rect 143078 39996 143110 40067
rect 143398 40034 143435 40090
rect 143491 40034 143528 40090
rect 144603 40067 144655 40073
rect 144610 39990 144652 40067
rect 145106 39990 145136 41860
rect 145830 40874 145888 40881
rect 145828 40872 145888 40874
rect 145828 40816 145830 40872
rect 145886 40816 145888 40872
rect 145828 40803 145888 40816
rect 145852 40134 145888 40803
rect 148107 40347 148167 40356
rect 148107 40278 148167 40287
rect 145828 40132 145906 40134
rect 145828 40076 145839 40132
rect 145895 40076 145906 40132
rect 145828 40074 145906 40076
rect 148109 20494 148165 40278
rect 148109 20438 149299 20494
rect 149243 20108 149299 20438
rect 152301 17140 152357 42193
rect 187327 41713 187383 42193
rect 189167 41713 189223 42193
rect 189811 41713 189867 42193
rect 191007 41713 191063 42193
rect 191651 41713 191707 42193
rect 192203 41713 192259 42193
rect 192847 41713 192903 42193
rect 193491 41713 193547 42193
rect 194043 41713 194099 42193
rect 196527 41713 196583 42193
rect 197171 41713 197227 42193
rect 197815 41713 197871 42193
rect 198367 41713 198423 42193
rect 200207 41713 200263 42193
rect 200851 41713 200907 42193
rect 201495 41713 201551 42193
rect 202047 41713 202103 42193
rect 202717 40882 202769 42193
rect 202713 40871 202773 40882
rect 205928 40881 205980 42193
rect 295927 41713 295983 42193
rect 297767 41713 297823 42193
rect 298411 41713 298467 42193
rect 299607 41713 299663 42193
rect 300251 41713 300307 42193
rect 300803 41713 300859 42193
rect 301447 41713 301503 42193
rect 302091 41713 302147 42193
rect 302643 41713 302699 42193
rect 305127 41713 305183 42193
rect 305771 41713 305827 42193
rect 306415 41713 306471 42193
rect 306967 41713 307023 42193
rect 308807 41713 308863 42193
rect 309451 41713 309507 42193
rect 310095 41713 310151 42193
rect 310647 41713 310703 42193
rect 311317 40882 311369 42193
rect 202713 40815 202715 40871
rect 202771 40815 202773 40871
rect 202713 40804 202773 40815
rect 205924 40870 205984 40881
rect 205924 40814 205926 40870
rect 205982 40814 205984 40870
rect 205924 40803 205984 40814
rect 311313 40871 311373 40882
rect 315497 40876 315549 42193
rect 350727 41713 350783 42193
rect 352567 41713 352623 42193
rect 353211 41713 353267 42193
rect 354407 41713 354463 42193
rect 355051 41713 355107 42193
rect 355603 41713 355659 42193
rect 356247 41713 356303 42193
rect 356891 41713 356947 42193
rect 357443 41713 357499 42193
rect 359927 41713 359983 42193
rect 360571 41713 360627 42193
rect 361215 41713 361271 42193
rect 361767 41713 361823 42193
rect 363607 41713 363663 42193
rect 364251 41713 364307 42193
rect 364895 41713 364951 42193
rect 365447 41713 365503 42193
rect 366117 40882 366169 42193
rect 311313 40815 311315 40871
rect 311371 40815 311373 40871
rect 315484 40874 315562 40876
rect 315484 40818 315495 40874
rect 315551 40818 315562 40874
rect 315484 40816 315562 40818
rect 366113 40871 366173 40882
rect 370302 40881 370354 42171
rect 405527 41713 405583 42193
rect 407367 41713 407423 42193
rect 408011 41713 408067 42193
rect 409207 41713 409263 42193
rect 409851 41713 409907 42193
rect 410403 41713 410459 42193
rect 411047 41713 411103 42193
rect 411691 41713 411747 42193
rect 412243 41713 412299 42193
rect 414727 41713 414783 42193
rect 415371 41713 415427 42193
rect 416015 41713 416071 42193
rect 416567 41713 416623 42193
rect 418407 41713 418463 42193
rect 419051 41713 419107 42193
rect 419695 41713 419751 42193
rect 420247 41713 420303 42193
rect 420917 40882 420969 42193
rect 311313 40804 311373 40815
rect 366113 40815 366115 40871
rect 366171 40815 366173 40871
rect 366113 40804 366173 40815
rect 370298 40870 370358 40881
rect 370298 40814 370300 40870
rect 370356 40814 370358 40870
rect 370298 40803 370358 40814
rect 420913 40871 420973 40882
rect 420913 40815 420915 40871
rect 420971 40815 420973 40871
rect 425115 40869 425167 42193
rect 460327 41713 460383 42193
rect 462167 41713 462223 42193
rect 462811 41713 462867 42193
rect 464007 41713 464063 42193
rect 464651 41713 464707 42193
rect 465203 41713 465259 42193
rect 465847 41713 465903 42193
rect 466491 41713 466547 42193
rect 467043 41713 467099 42193
rect 469527 41713 469583 42193
rect 470171 41713 470227 42193
rect 470815 41713 470871 42193
rect 471367 41713 471423 42193
rect 473207 41713 473263 42193
rect 473851 41713 473907 42193
rect 474495 41713 474551 42193
rect 475047 41713 475103 42193
rect 475717 40882 475769 42193
rect 479915 40883 479967 42193
rect 515127 41713 515183 42193
rect 516967 41713 517023 42193
rect 517611 41713 517667 42193
rect 518807 41713 518863 42193
rect 519451 41713 519507 42193
rect 520003 41713 520059 42193
rect 520647 41713 520703 42193
rect 521291 41713 521347 42193
rect 521843 41713 521899 42193
rect 524327 41713 524383 42193
rect 524971 41713 525027 42193
rect 525615 41713 525671 42193
rect 526167 41713 526223 42193
rect 528007 41713 528063 42193
rect 528651 41713 528707 42193
rect 529295 41713 529351 42193
rect 529847 41713 529903 42193
rect 475713 40871 475773 40882
rect 420913 40804 420973 40815
rect 425111 40858 425171 40869
rect 425111 40802 425113 40858
rect 425169 40802 425171 40858
rect 475713 40815 475715 40871
rect 475771 40815 475773 40871
rect 475713 40804 475773 40815
rect 479911 40872 479971 40883
rect 530517 40882 530569 42193
rect 479911 40816 479913 40872
rect 479969 40816 479971 40872
rect 479911 40805 479971 40816
rect 530513 40871 530573 40882
rect 534772 40871 534824 42193
rect 647219 41877 647271 42193
rect 647443 41877 647495 42193
rect 647667 41877 647719 42193
rect 647891 41877 647943 42193
rect 648115 41877 648167 42193
rect 648339 41877 648391 42193
rect 648563 41877 648615 42193
rect 648787 41877 648839 42193
rect 649011 41877 649063 42193
rect 649235 41877 649287 42193
rect 649459 41877 649511 42193
rect 649683 41877 649735 42193
rect 649907 41877 649959 42193
rect 650131 41877 650183 42193
rect 650355 41877 650407 42193
rect 650579 41877 650631 42193
rect 650803 41877 650855 42193
rect 651027 41877 651079 42193
rect 651251 41877 651303 42193
rect 651475 41877 651527 42193
rect 651699 41877 651751 42193
rect 651923 41877 651975 42193
rect 652147 41877 652199 42193
rect 652371 41877 652423 42193
rect 652595 41877 652647 42193
rect 652819 41877 652871 42193
rect 653043 41877 653095 42193
rect 653267 41877 653319 42193
rect 653491 41877 653543 42193
rect 653715 41877 653767 42193
rect 653939 41877 653991 42193
rect 654163 41877 654215 42193
rect 530513 40815 530515 40871
rect 530571 40815 530573 40871
rect 530513 40804 530573 40815
rect 534768 40860 534828 40871
rect 534768 40804 534770 40860
rect 534826 40804 534828 40860
rect 425111 40791 425171 40802
rect 534768 40793 534828 40804
rect 644277 20057 644329 20063
rect 644277 19999 644329 20005
rect 644005 19831 644057 19837
rect 644005 19773 644057 19779
rect 643908 19503 643960 19509
rect 643908 19445 643960 19451
rect 643361 19054 643389 19062
rect 643349 19048 643401 19054
rect 643349 18990 643401 18996
rect 151931 17084 152357 17140
rect 643361 14515 643389 18990
rect 643807 18373 643859 18379
rect 643807 18315 643859 18321
rect 643685 17698 643737 17704
rect 643685 17640 643737 17646
rect 643459 17254 643511 17260
rect 643459 17196 643511 17202
rect 643345 14506 643405 14515
rect 643345 14437 643405 14446
rect 643471 11803 643499 17196
rect 643571 17140 643623 17146
rect 643571 17082 643623 17088
rect 643583 12616 643611 17082
rect 643697 13693 643725 17640
rect 643681 13684 643741 13693
rect 643681 13615 643741 13624
rect 643819 13326 643847 18315
rect 643920 15335 643948 19445
rect 643904 15326 643964 15335
rect 643904 15257 643964 15266
rect 643738 13298 643847 13326
rect 643567 12607 643627 12616
rect 643567 12538 643627 12547
rect 643583 12530 643611 12538
rect 643738 12383 643766 13298
rect 643455 11794 643515 11803
rect 643455 11725 643515 11734
rect 644017 11570 644045 19773
rect 644110 18272 644162 18278
rect 644110 18214 644162 18220
rect 643900 11542 644045 11570
rect 643900 10984 643928 11542
rect 643884 10975 643944 10984
rect 643884 10906 643944 10915
rect 644122 9977 644150 18214
rect 644289 16269 644317 19999
rect 647002 19940 647054 19946
rect 647002 19882 647054 19888
rect 646117 19152 646169 19158
rect 646117 19094 646169 19100
rect 644832 18935 644884 18941
rect 644832 18877 644884 18883
rect 644844 16237 644872 18877
rect 645382 18037 645434 18043
rect 645382 17979 645434 17985
rect 645394 16212 645422 17979
rect 646129 16263 646157 19094
rect 646671 17816 646723 17822
rect 646671 17758 646723 17764
rect 646683 16277 646711 17758
rect 647014 16949 647042 19882
rect 647002 16943 647054 16949
rect 647002 16885 647054 16891
rect 647230 16235 647258 41877
rect 647454 17146 647482 41877
rect 647678 17258 647706 41877
rect 647902 17370 647930 41877
rect 648126 17482 648154 41877
rect 648350 17594 648378 41877
rect 648574 17706 648602 41877
rect 648798 17818 648826 41877
rect 649022 17930 649050 41877
rect 649246 18042 649274 41877
rect 649470 18154 649498 41877
rect 649694 18266 649722 41877
rect 649918 18378 649946 41877
rect 649851 18372 650016 18378
rect 650015 18320 650016 18372
rect 649851 18314 650016 18320
rect 649918 18312 649946 18314
rect 649627 18260 649792 18266
rect 649791 18208 649792 18260
rect 649627 18202 649792 18208
rect 649694 18198 649722 18202
rect 649403 18148 649568 18154
rect 649567 18096 649568 18148
rect 649403 18090 649568 18096
rect 649470 18084 649498 18090
rect 649179 18036 649344 18042
rect 649343 17984 649344 18036
rect 649179 17978 649344 17984
rect 649246 17967 649274 17978
rect 650142 17961 650170 41877
rect 649507 17933 650170 17961
rect 648955 17924 649120 17930
rect 649119 17872 649120 17924
rect 648955 17866 649120 17872
rect 649022 17856 649050 17866
rect 648731 17812 648896 17818
rect 648895 17760 648896 17812
rect 648731 17754 648896 17760
rect 648798 17743 648826 17754
rect 648507 17700 648672 17706
rect 648671 17648 648672 17700
rect 648507 17642 648672 17648
rect 648574 17639 648602 17642
rect 648283 17588 648448 17594
rect 648447 17536 648448 17588
rect 648283 17530 648448 17536
rect 648350 17525 648378 17530
rect 648059 17476 648224 17482
rect 648223 17424 648224 17476
rect 648059 17418 648224 17424
rect 648126 17411 648154 17418
rect 649507 17399 649535 17933
rect 650366 17779 650394 41877
rect 648522 17371 649535 17399
rect 649621 17751 650394 17779
rect 647835 17364 648000 17370
rect 647999 17312 648000 17364
rect 647835 17306 648000 17312
rect 647902 17299 647930 17306
rect 647611 17252 647776 17258
rect 647775 17200 647776 17252
rect 647611 17194 647776 17200
rect 647678 17183 647706 17194
rect 647387 17140 647552 17146
rect 647551 17088 647552 17140
rect 647387 17082 647552 17088
rect 647454 17077 647482 17082
rect 647958 16943 648010 16949
rect 647958 16885 648010 16891
rect 647970 15409 647998 16885
rect 648522 15436 648550 17371
rect 649621 17291 649649 17751
rect 650590 17688 650618 41877
rect 650814 18614 650842 41877
rect 651038 18938 651066 41877
rect 651262 19050 651290 41877
rect 651486 19162 651514 41877
rect 651419 19156 651584 19162
rect 651583 19104 651584 19156
rect 651419 19098 651584 19104
rect 651486 19075 651514 19098
rect 651195 19044 651360 19050
rect 651359 18992 651360 19044
rect 651195 18986 651360 18992
rect 651262 18970 651290 18986
rect 650971 18932 651136 18938
rect 651135 18880 651136 18932
rect 650971 18874 651136 18880
rect 651038 18866 651066 18874
rect 650012 17660 650618 17688
rect 650812 18536 650842 18614
rect 649865 17587 649917 17593
rect 649865 17529 649917 17535
rect 649753 17477 649805 17483
rect 649753 17419 649805 17425
rect 649238 17263 649649 17291
rect 649062 16944 649114 16950
rect 649062 16886 649114 16892
rect 649074 15446 649102 16886
rect 649238 10031 649266 17263
rect 649614 16821 649666 16827
rect 649614 16763 649666 16769
rect 649626 15424 649654 16763
rect 649765 12892 649793 17419
rect 649877 13698 649905 17529
rect 649861 13689 649921 13698
rect 649861 13620 649921 13629
rect 649749 12883 649809 12892
rect 649749 12814 649809 12823
rect 649765 12813 649793 12814
rect 650012 10990 650040 17660
rect 650129 16644 650181 16650
rect 650129 16586 650181 16592
rect 650141 14507 650169 16586
rect 650125 14498 650185 14507
rect 650125 14429 650185 14438
rect 649996 10981 650056 10990
rect 649996 10912 650056 10921
rect 649074 10003 649266 10031
rect 648507 9979 648559 9985
rect 644122 9949 644318 9977
rect 648507 9921 648559 9927
rect 647215 9893 647267 9899
rect 647215 9835 647267 9841
rect 647958 9794 648010 9800
rect 647958 9736 648010 9742
rect 646670 9706 646722 9712
rect 646670 9648 646722 9654
rect 650812 9609 650840 18536
rect 651710 11799 651738 41877
rect 651697 11790 651758 11799
rect 651753 11734 651758 11790
rect 651697 11725 651758 11734
rect 651934 10171 651962 41877
rect 652158 19498 652186 41877
rect 652091 19492 652256 19498
rect 652255 19440 652256 19492
rect 652091 19434 652256 19440
rect 652158 19423 652186 19434
rect 652382 18451 652410 41877
rect 652606 19301 652634 41877
rect 652830 19834 652858 41877
rect 653054 19946 653082 41877
rect 653278 20058 653306 41877
rect 653211 20052 653376 20058
rect 653375 20000 653376 20052
rect 653211 19994 653376 20000
rect 653278 19991 653306 19994
rect 652987 19940 653152 19946
rect 653151 19888 653152 19940
rect 652987 19882 653152 19888
rect 652763 19828 652928 19834
rect 652927 19776 652928 19828
rect 652763 19770 652928 19776
rect 652606 19273 652678 19301
rect 652382 18423 652548 18451
rect 652353 18145 652405 18151
rect 652353 18087 652405 18093
rect 652234 17929 652286 17935
rect 652234 17871 652286 17877
rect 652096 17363 652148 17369
rect 652096 17305 652148 17311
rect 651918 10162 651978 10171
rect 651918 10093 651978 10102
rect 652108 9712 652136 17305
rect 652246 9800 652274 17871
rect 652365 9899 652393 18087
rect 652353 9893 652405 9899
rect 652353 9835 652405 9841
rect 652234 9794 652286 9800
rect 652234 9736 652286 9742
rect 652096 9706 652148 9712
rect 652096 9648 652148 9654
rect 645376 9603 645428 9609
rect 645376 9545 645428 9551
rect 650801 9603 650853 9609
rect 650801 9545 650853 9551
rect 652520 9506 652548 18423
rect 652650 16950 652678 19273
rect 652638 16944 652690 16950
rect 652638 16886 652690 16892
rect 653502 16827 653530 41877
rect 653494 16821 653546 16827
rect 653494 16763 653546 16769
rect 653726 16532 653754 41877
rect 653950 16645 653978 41877
rect 653938 16639 653990 16645
rect 653938 16581 653990 16587
rect 652735 16504 653754 16532
rect 652735 9985 652763 16504
rect 654174 16433 654202 41877
rect 652896 16405 654202 16433
rect 652724 9979 652776 9985
rect 652724 9921 652776 9927
rect 644827 9500 644879 9506
rect 644827 9442 644879 9448
rect 652514 9500 652566 9506
rect 652514 9442 652566 9448
rect 652896 9408 652924 16405
rect 646117 9402 646169 9408
rect 646117 9344 646169 9350
rect 652884 9402 652936 9408
rect 652884 9344 652936 9350
<< via2 >>
rect 69634 996693 69695 996754
rect 71635 996693 71696 996754
rect 120834 996693 120895 996754
rect 122835 996687 122896 996748
rect 172034 996693 172095 996754
rect 174035 996696 174096 996757
rect 223234 996699 223295 996760
rect 225235 996685 225296 996746
rect 274434 996696 274495 996757
rect 276435 996696 276496 996757
rect 378834 996702 378895 996763
rect 380835 996699 380896 996760
rect 467834 996687 467895 996748
rect 469835 996690 469896 996751
rect 519034 996690 519095 996751
rect 521035 996693 521096 996754
rect 618434 996690 618495 996751
rect 620435 996693 620496 996754
rect 18934 95739 19194 95795
rect 41478 95739 41829 95795
rect 18569 95515 18829 95571
rect 41470 95515 41821 95571
rect 17843 95291 18112 95347
rect 41467 95291 41536 95347
rect 41536 95291 41818 95347
rect 141710 40289 141771 40350
rect 143435 40073 143437 40090
rect 143437 40073 143489 40090
rect 143489 40073 143491 40090
rect 143435 40034 143491 40073
rect 145830 40816 145886 40872
rect 148107 40287 148167 40347
rect 145839 40076 145895 40132
rect 202715 40815 202771 40871
rect 205926 40814 205982 40870
rect 311315 40815 311371 40871
rect 315495 40818 315551 40874
rect 366115 40815 366171 40871
rect 370300 40814 370356 40870
rect 420915 40815 420971 40871
rect 425113 40802 425169 40858
rect 475715 40815 475771 40871
rect 479913 40816 479969 40872
rect 530515 40815 530571 40871
rect 534770 40804 534826 40860
rect 643345 14446 643405 14506
rect 643681 13624 643741 13684
rect 643904 15266 643964 15326
rect 643567 12547 643627 12607
rect 643455 11734 643515 11794
rect 643884 10915 643944 10975
rect 649861 13629 649921 13689
rect 649749 12823 649809 12883
rect 650125 14438 650185 14498
rect 649996 10921 650056 10981
rect 651697 11734 651753 11790
rect 651918 10102 651978 10162
<< metal3 >>
rect 71300 1006801 71750 1006864
rect 71300 1006097 71377 1006801
rect 71681 1006097 71750 1006801
rect 70733 1000260 71114 1000330
rect 70733 999556 70772 1000260
rect 71076 999556 71114 1000260
rect 70733 997902 71114 999556
rect 70733 997758 70776 997902
rect 71080 997758 71114 997902
rect 70733 997615 71114 997758
rect 71300 997901 71750 1006097
rect 122500 1006801 122950 1006864
rect 122500 1006097 122577 1006801
rect 122881 1006097 122950 1006801
rect 71300 997757 71358 997901
rect 71662 997757 71750 997901
rect 71300 997615 71750 997757
rect 121933 1000260 122314 1000330
rect 121933 999556 121972 1000260
rect 122276 999556 122314 1000260
rect 121933 997902 122314 999556
rect 121933 997758 121976 997902
rect 122280 997758 122314 997902
rect 121933 997615 122314 997758
rect 122500 997901 122950 1006097
rect 173700 1006801 174150 1006864
rect 173700 1006097 173777 1006801
rect 174081 1006097 174150 1006801
rect 122500 997757 122558 997901
rect 122862 997757 122950 997901
rect 122500 997615 122950 997757
rect 173133 1000260 173514 1000330
rect 173133 999556 173172 1000260
rect 173476 999556 173514 1000260
rect 173133 997902 173514 999556
rect 173133 997758 173176 997902
rect 173480 997758 173514 997902
rect 173133 997615 173514 997758
rect 173700 997901 174150 1006097
rect 224900 1006801 225350 1006864
rect 224900 1006097 224977 1006801
rect 225281 1006097 225350 1006801
rect 173700 997757 173758 997901
rect 174062 997757 174150 997901
rect 173700 997615 174150 997757
rect 224333 1000260 224714 1000330
rect 224333 999556 224372 1000260
rect 224676 999556 224714 1000260
rect 224333 997902 224714 999556
rect 224333 997758 224376 997902
rect 224680 997758 224714 997902
rect 224333 997615 224714 997758
rect 224900 997901 225350 1006097
rect 276100 1006801 276550 1006864
rect 276100 1006097 276177 1006801
rect 276481 1006097 276550 1006801
rect 224900 997757 224958 997901
rect 225257 997757 225350 997901
rect 224900 997615 225350 997757
rect 275533 1000260 275914 1000330
rect 275533 999556 275572 1000260
rect 275876 999556 275914 1000260
rect 275533 997902 275914 999556
rect 275533 997758 275576 997902
rect 275880 997758 275914 997902
rect 275533 997615 275914 997758
rect 276100 997901 276550 1006097
rect 380500 1006801 380950 1006864
rect 380500 1006097 380577 1006801
rect 380881 1006097 380950 1006801
rect 276100 997757 276158 997901
rect 276462 997757 276550 997901
rect 276100 997615 276550 997757
rect 379933 1000260 380314 1000330
rect 379933 999556 379972 1000260
rect 380276 999556 380314 1000260
rect 379933 997902 380314 999556
rect 379933 997758 379976 997902
rect 380280 997758 380314 997902
rect 69629 996754 69700 996759
rect 69629 996693 69634 996754
rect 69695 996693 69700 996754
rect 69629 996688 69700 996693
rect 71630 996754 71701 996759
rect 71630 996693 71635 996754
rect 71696 996693 71701 996754
rect 72383 996696 74649 996756
rect 120829 996754 120900 996759
rect 71630 996688 71701 996693
rect 120829 996693 120834 996754
rect 120895 996693 120900 996754
rect 120829 996688 120900 996693
rect 122830 996748 122901 996753
rect 122830 996687 122835 996748
rect 122896 996687 122901 996748
rect 123602 996696 126002 996756
rect 172029 996754 172100 996759
rect 172029 996693 172034 996754
rect 172095 996693 172100 996754
rect 172029 996688 172100 996693
rect 174030 996757 174101 996762
rect 174030 996696 174035 996757
rect 174096 996696 174101 996757
rect 223229 996760 223300 996765
rect 174817 996696 177414 996756
rect 223229 996699 223234 996760
rect 223295 996699 223300 996760
rect 274429 996757 274500 996762
rect 174030 996691 174101 996696
rect 223229 996694 223300 996699
rect 225230 996746 225301 996751
rect 122830 996682 122901 996687
rect 225230 996685 225235 996746
rect 225296 996685 225301 996746
rect 225983 996696 228817 996756
rect 274429 996696 274434 996757
rect 274495 996696 274500 996757
rect 274429 996691 274500 996696
rect 276430 996757 276501 996762
rect 276430 996696 276435 996757
rect 276496 996696 276501 996757
rect 277181 996696 280424 996756
rect 276430 996691 276501 996696
rect 225230 996680 225301 996685
rect 333499 995407 338279 997742
rect 343478 995407 348258 997742
rect 379933 997615 380314 997758
rect 380500 997901 380950 1006097
rect 469500 1006801 469950 1006864
rect 469500 1006097 469577 1006801
rect 469881 1006097 469950 1006801
rect 380500 997757 380558 997901
rect 380862 997757 380950 997901
rect 380500 997615 380950 997757
rect 468933 1000260 469314 1000330
rect 468933 999556 468972 1000260
rect 469276 999556 469314 1000260
rect 468933 997902 469314 999556
rect 468933 997758 468976 997902
rect 469280 997758 469314 997902
rect 468933 997615 469314 997758
rect 469500 997901 469950 1006097
rect 520700 1006801 521150 1006864
rect 520700 1006097 520777 1006801
rect 521081 1006097 521150 1006801
rect 469500 997757 469558 997901
rect 469862 997757 469950 997901
rect 469500 997615 469950 997757
rect 520133 1000260 520514 1000330
rect 520133 999556 520172 1000260
rect 520476 999556 520514 1000260
rect 520133 997902 520514 999556
rect 520133 997758 520176 997902
rect 520480 997758 520514 997902
rect 520133 997615 520514 997758
rect 520700 997901 521150 1006097
rect 620100 1006801 620550 1006864
rect 620100 1006097 620177 1006801
rect 620481 1006097 620550 1006801
rect 520700 997757 520758 997901
rect 521062 997757 521150 997901
rect 520700 997615 521150 997757
rect 619533 1000260 619914 1000330
rect 619533 999556 619572 1000260
rect 619876 999556 619914 1000260
rect 619533 997902 619914 999556
rect 619533 997758 619576 997902
rect 619880 997758 619914 997902
rect 378829 996763 378900 996768
rect 378829 996702 378834 996763
rect 378895 996702 378900 996763
rect 378829 996697 378900 996702
rect 380830 996760 380901 996765
rect 380830 996699 380835 996760
rect 380896 996699 380901 996760
rect 380830 996694 380901 996699
rect 381595 996696 382235 996756
rect 467829 996748 467900 996753
rect 467829 996687 467834 996748
rect 467895 996687 467900 996748
rect 467829 996682 467900 996687
rect 469830 996751 469901 996756
rect 469830 996690 469835 996751
rect 469896 996690 469901 996751
rect 470601 996696 471209 996756
rect 519029 996751 519100 996756
rect 469830 996685 469901 996690
rect 519029 996690 519034 996751
rect 519095 996690 519100 996751
rect 519029 996685 519100 996690
rect 521030 996754 521101 996759
rect 521030 996693 521035 996754
rect 521096 996693 521101 996754
rect 521803 996696 522603 996756
rect 521030 996688 521101 996693
rect 575699 995407 580479 997640
rect 585678 995407 590458 997664
rect 619533 997615 619914 997758
rect 620100 997901 620550 1006097
rect 620100 997757 620158 997901
rect 620462 997757 620550 997901
rect 620100 997615 620550 997757
rect 618429 996751 618500 996756
rect 618429 996690 618434 996751
rect 618495 996690 618500 996751
rect 618429 996685 618500 996690
rect 620430 996754 620501 996759
rect 620430 996693 620435 996754
rect 620496 996693 620501 996754
rect 621201 996696 624463 996756
rect 620430 996688 620501 996693
rect 675407 971144 676767 971206
rect 677626 970068 680341 970107
rect 677626 970064 679567 970068
rect 677626 969760 677649 970064
rect 677793 969764 679567 970064
rect 680271 969764 680341 970068
rect 677793 969760 680341 969764
rect 677626 969726 680341 969760
rect 677626 969463 686875 969540
rect 677626 969462 686108 969463
rect 41713 969210 42193 969280
rect 675407 969142 676797 969204
rect 677626 969158 677648 969462
rect 677792 969159 686108 969462
rect 686812 969159 686875 969463
rect 677792 969158 686875 969159
rect 677626 969090 686875 969158
rect 41713 967370 42193 967440
rect 675407 967240 675887 967310
rect 41713 966726 42193 966796
rect 675407 966688 675887 966758
rect 675407 966044 675887 966114
rect 41713 965530 42193 965600
rect 675407 965400 675887 965470
rect 41713 964886 42193 964956
rect 41713 964334 42193 964404
rect 41713 963690 42193 963760
rect 675407 963560 675887 963630
rect 41713 963046 42193 963116
rect 675407 963008 675887 963078
rect 41713 962494 42193 962564
rect 675407 962364 675887 962434
rect 675407 961720 675887 961790
rect 41713 960010 42193 960080
rect 41713 959366 42193 959436
rect 675407 959236 675887 959306
rect 41713 958722 42193 958792
rect 675407 958684 675887 958754
rect 41713 958170 42193 958240
rect 675407 958040 675887 958110
rect 675407 957396 675887 957466
rect 675407 956844 675887 956914
rect 41713 956330 42193 956400
rect 675407 956200 675887 956270
rect 41713 955686 42193 955756
rect 41713 955042 42193 955112
rect 675407 955004 675887 955074
rect 41713 954490 42193 954560
rect 675407 954360 675887 954430
rect 40832 949550 40892 952819
rect 675407 952520 675887 952590
rect 30782 948827 39885 948896
rect 30782 948523 30845 948827
rect 31549 948808 39885 948827
rect 31549 948523 39705 948808
rect 30782 948504 39705 948523
rect 39849 948504 39885 948808
rect 40810 948781 42193 948841
rect 30782 948446 39885 948504
rect 37316 948222 39885 948260
rect 37316 947918 37386 948222
rect 38090 948216 39885 948222
rect 38090 947918 39704 948216
rect 37316 947912 39704 947918
rect 39848 947912 39885 948216
rect 37316 947879 39885 947912
rect 40810 946781 42193 946841
rect 39880 926939 42193 926940
rect 39880 922151 41039 926939
rect 41837 922151 42193 926939
rect 675407 922499 677778 922500
rect 39880 921851 42193 921852
rect 39880 917191 39919 921851
rect 40717 917191 42193 921851
rect 675407 917701 675787 922499
rect 676585 917701 677778 922499
rect 675407 917700 677778 917701
rect 39880 917190 42193 917191
rect 675407 917409 677778 917410
rect 39880 916899 42193 916900
rect 39880 912101 41039 916899
rect 41837 912101 42193 916899
rect 675407 912749 676907 917409
rect 677705 912749 677778 917409
rect 675407 912748 677778 912749
rect 39880 912100 42193 912101
rect 675407 907661 675787 912449
rect 676585 907661 677778 912449
rect 675407 907660 677778 907661
rect 39913 879878 42193 884658
rect 675407 881144 676767 881206
rect 677626 880068 680341 880107
rect 677626 880064 679567 880068
rect 677626 879760 677649 880064
rect 677793 879764 679567 880064
rect 680271 879764 680341 880068
rect 677793 879760 680341 879764
rect 677626 879726 680341 879760
rect 677626 879463 686875 879540
rect 677626 879462 686108 879463
rect 675407 879142 676797 879204
rect 677626 879158 677648 879462
rect 677792 879159 686108 879462
rect 686812 879159 686875 879463
rect 677792 879158 686875 879159
rect 677626 879090 686875 879158
rect 675407 878040 675887 878110
rect 675407 877488 675887 877558
rect 675407 876844 675887 876914
rect 675407 876200 675887 876270
rect 39913 869899 42193 874679
rect 675407 874360 675887 874430
rect 675407 873808 675887 873878
rect 675407 873164 675887 873234
rect 675407 872520 675887 872590
rect 675407 870036 675887 870106
rect 675407 869484 675887 869554
rect 675407 868840 675887 868910
rect 675407 868196 675887 868266
rect 675407 867644 675887 867714
rect 675407 867000 675887 867070
rect 675407 865804 675887 865874
rect 675407 865160 675887 865230
rect 675407 863320 675887 863390
rect 39920 837678 42193 842458
rect 39920 827699 42193 832479
rect 675407 828521 677782 833301
rect 675407 818542 677782 823322
rect 41713 799410 42193 799480
rect 41713 797570 42193 797640
rect 41713 796926 42193 796996
rect 41713 795730 42193 795800
rect 41713 795086 42193 795156
rect 41713 794534 42193 794604
rect 41713 793890 42193 793960
rect 41713 793246 42193 793316
rect 41713 792694 42193 792764
rect 675407 792144 676767 792206
rect 677626 791068 680341 791107
rect 677626 791064 679567 791068
rect 677626 790760 677649 791064
rect 677793 790764 679567 791064
rect 680271 790764 680341 791068
rect 677793 790760 680341 790764
rect 677626 790726 680341 790760
rect 677626 790463 686875 790540
rect 677626 790462 686108 790463
rect 41713 790210 42193 790280
rect 675407 790142 676797 790204
rect 677626 790158 677648 790462
rect 677792 790159 686108 790462
rect 686812 790159 686875 790463
rect 677792 790158 686875 790159
rect 677626 790090 686875 790158
rect 41713 789566 42193 789636
rect 41713 788922 42193 788992
rect 675407 788840 675887 788910
rect 41713 788370 42193 788440
rect 675407 788288 675887 788358
rect 675407 787644 675887 787714
rect 675407 787000 675887 787070
rect 41713 786530 42193 786600
rect 41713 785886 42193 785956
rect 41713 785242 42193 785312
rect 675407 785160 675887 785230
rect 41713 784690 42193 784760
rect 675407 784608 675887 784678
rect 675407 783964 675887 784034
rect 675407 783320 675887 783390
rect 40832 779539 40892 783008
rect 675407 780836 675887 780906
rect 675407 780284 675887 780354
rect 675407 779640 675887 779710
rect 675407 778996 675887 779066
rect 30782 778827 39885 778896
rect 30782 778523 30845 778827
rect 31549 778808 39885 778827
rect 31549 778523 39705 778808
rect 30782 778504 39705 778523
rect 39849 778504 39885 778808
rect 40810 778781 42193 778841
rect 30782 778446 39885 778504
rect 675407 778444 675887 778514
rect 37316 778222 39885 778260
rect 37316 777918 37386 778222
rect 38090 778216 39885 778222
rect 38090 777918 39704 778216
rect 37316 777912 39704 777918
rect 39848 777912 39885 778216
rect 37316 777879 39885 777912
rect 675407 777800 675887 777870
rect 40810 776781 42193 776841
rect 675407 776604 675887 776674
rect 675407 775960 675887 776030
rect 675407 774120 675887 774190
rect 41713 756210 42193 756280
rect 41713 754370 42193 754440
rect 41713 753726 42193 753796
rect 41713 752530 42193 752600
rect 41713 751886 42193 751956
rect 41713 751334 42193 751404
rect 41713 750690 42193 750760
rect 41713 750046 42193 750116
rect 41713 749494 42193 749564
rect 675407 747144 676767 747206
rect 41713 747010 42193 747080
rect 41713 746366 42193 746436
rect 677626 746068 680341 746107
rect 677626 746064 679567 746068
rect 41713 745722 42193 745792
rect 677626 745760 677649 746064
rect 677793 745764 679567 746064
rect 680271 745764 680341 746068
rect 677793 745760 680341 745764
rect 677626 745726 680341 745760
rect 677626 745463 686875 745540
rect 677626 745462 686108 745463
rect 41713 745170 42193 745240
rect 675407 745142 676797 745204
rect 677626 745158 677648 745462
rect 677792 745159 686108 745462
rect 686812 745159 686875 745463
rect 677792 745158 686875 745159
rect 677626 745090 686875 745158
rect 675407 743840 675887 743910
rect 41713 743330 42193 743400
rect 675407 743288 675887 743358
rect 41713 742686 42193 742756
rect 675407 742644 675887 742714
rect 41713 742042 42193 742112
rect 675407 742000 675887 742070
rect 41713 741490 42193 741560
rect 675407 740160 675887 740230
rect 40832 736546 40892 739828
rect 675407 739608 675887 739678
rect 675407 738964 675887 739034
rect 675407 738320 675887 738390
rect 30782 735827 39885 735896
rect 30782 735523 30845 735827
rect 31549 735808 39885 735827
rect 31549 735523 39705 735808
rect 30782 735504 39705 735523
rect 39849 735504 39885 735808
rect 40810 735781 42193 735841
rect 675407 735836 675887 735906
rect 30782 735446 39885 735504
rect 675407 735284 675887 735354
rect 37316 735222 39885 735260
rect 37316 734918 37386 735222
rect 38090 735216 39885 735222
rect 38090 734918 39704 735216
rect 37316 734912 39704 734918
rect 39848 734912 39885 735216
rect 37316 734879 39885 734912
rect 675407 734640 675887 734710
rect 675407 733996 675887 734066
rect 40810 733781 42193 733841
rect 675407 733444 675887 733514
rect 675407 732800 675887 732870
rect 675407 731604 675887 731674
rect 675407 730960 675887 731030
rect 675407 729120 675887 729190
rect 41713 713010 42193 713080
rect 41713 711170 42193 711240
rect 41713 710526 42193 710596
rect 41713 709330 42193 709400
rect 41713 708686 42193 708756
rect 41713 708134 42193 708204
rect 41713 707490 42193 707560
rect 41713 706846 42193 706916
rect 41713 706294 42193 706364
rect 41713 703810 42193 703880
rect 41713 703166 42193 703236
rect 41713 702522 42193 702592
rect 675407 702144 676767 702206
rect 41713 701970 42193 702040
rect 677626 701068 680341 701107
rect 677626 701064 679567 701068
rect 677626 700760 677649 701064
rect 677793 700764 679567 701064
rect 680271 700764 680341 701068
rect 677793 700760 680341 700764
rect 677626 700726 680341 700760
rect 677626 700463 686875 700540
rect 677626 700462 686108 700463
rect 41713 700130 42193 700200
rect 675407 700142 676797 700204
rect 677626 700158 677648 700462
rect 677792 700159 686108 700462
rect 686812 700159 686875 700463
rect 677792 700158 686875 700159
rect 677626 700090 686875 700158
rect 41713 699486 42193 699556
rect 41713 698842 42193 698912
rect 675407 698840 675887 698910
rect 41713 698290 42193 698360
rect 675407 698288 675887 698358
rect 675407 697644 675887 697714
rect 675407 697000 675887 697070
rect 40832 693552 40892 696608
rect 675407 695160 675887 695230
rect 675407 694608 675887 694678
rect 675407 693964 675887 694034
rect 675407 693320 675887 693390
rect 30782 692827 39885 692896
rect 30782 692523 30845 692827
rect 31549 692808 39885 692827
rect 31549 692523 39705 692808
rect 30782 692504 39705 692523
rect 39849 692504 39885 692808
rect 40810 692781 42193 692841
rect 30782 692446 39885 692504
rect 37316 692222 39885 692260
rect 37316 691918 37386 692222
rect 38090 692216 39885 692222
rect 38090 691918 39704 692216
rect 37316 691912 39704 691918
rect 39848 691912 39885 692216
rect 37316 691879 39885 691912
rect 40810 690781 42193 690841
rect 675407 690836 675887 690906
rect 675407 690284 675887 690354
rect 675407 689640 675887 689710
rect 675407 688996 675887 689066
rect 675407 688444 675887 688514
rect 675407 687800 675887 687870
rect 675407 686604 675887 686674
rect 675407 685960 675887 686030
rect 675407 684120 675887 684190
rect 41713 669810 42193 669880
rect 41713 667970 42193 668040
rect 41713 667326 42193 667396
rect 41713 666130 42193 666200
rect 41713 665486 42193 665556
rect 41713 664934 42193 665004
rect 41713 664290 42193 664360
rect 41713 663646 42193 663716
rect 41713 663094 42193 663164
rect 41713 660610 42193 660680
rect 41713 659966 42193 660036
rect 41713 659322 42193 659392
rect 41713 658770 42193 658840
rect 675407 657144 676767 657206
rect 41713 656930 42193 657000
rect 41713 656286 42193 656356
rect 677626 656068 680341 656107
rect 677626 656064 679567 656068
rect 677626 655760 677649 656064
rect 677793 655764 679567 656064
rect 680271 655764 680341 656068
rect 677793 655760 680341 655764
rect 677626 655726 680341 655760
rect 41713 655642 42193 655712
rect 677626 655463 686875 655540
rect 677626 655462 686108 655463
rect 41713 655090 42193 655160
rect 675407 655142 676797 655204
rect 677626 655158 677648 655462
rect 677792 655159 686108 655462
rect 686812 655159 686875 655463
rect 677792 655158 686875 655159
rect 677626 655090 686875 655158
rect 675407 653640 675887 653710
rect 40832 650533 40892 653443
rect 675407 653088 675887 653158
rect 675407 652444 675887 652514
rect 675407 651800 675887 651870
rect 675407 649960 675887 650030
rect 30782 649827 39885 649896
rect 30782 649523 30845 649827
rect 31549 649808 39885 649827
rect 31549 649523 39705 649808
rect 30782 649504 39705 649523
rect 39849 649504 39885 649808
rect 40810 649781 42193 649841
rect 30782 649446 39885 649504
rect 675407 649408 675887 649478
rect 37316 649222 39885 649260
rect 37316 648918 37386 649222
rect 38090 649216 39885 649222
rect 38090 648918 39704 649216
rect 37316 648912 39704 648918
rect 39848 648912 39885 649216
rect 37316 648879 39885 648912
rect 675407 648764 675887 648834
rect 675407 648120 675887 648190
rect 40810 647781 42193 647841
rect 675407 645636 675887 645706
rect 675407 645084 675887 645154
rect 675407 644440 675887 644510
rect 675407 643796 675887 643866
rect 675407 643244 675887 643314
rect 675407 642600 675887 642670
rect 675407 641404 675887 641474
rect 675407 640760 675887 640830
rect 675407 638920 675887 638990
rect 41713 626610 42193 626680
rect 41713 624770 42193 624840
rect 41713 624126 42193 624196
rect 41713 622930 42193 623000
rect 41713 622286 42193 622356
rect 41713 621734 42193 621804
rect 41713 621090 42193 621160
rect 41713 620446 42193 620516
rect 41713 619894 42193 619964
rect 41713 617410 42193 617480
rect 41713 616766 42193 616836
rect 41713 616122 42193 616192
rect 41713 615570 42193 615640
rect 41713 613730 42193 613800
rect 41713 613086 42193 613156
rect 41713 612442 42193 612512
rect 675407 612144 676767 612206
rect 41713 611890 42193 611960
rect 677626 611068 680341 611107
rect 677626 611064 679567 611068
rect 677626 610760 677649 611064
rect 677793 610764 679567 611064
rect 680271 610764 680341 611068
rect 677793 610760 680341 610764
rect 677626 610726 680341 610760
rect 677626 610463 686875 610540
rect 677626 610462 686108 610463
rect 40832 607531 40892 610227
rect 675407 610142 676797 610204
rect 677626 610158 677648 610462
rect 677792 610159 686108 610462
rect 686812 610159 686875 610463
rect 677792 610158 686875 610159
rect 677626 610090 686875 610158
rect 675407 608640 675887 608710
rect 675407 608088 675887 608158
rect 675407 607444 675887 607514
rect 30782 606827 39885 606896
rect 30782 606523 30845 606827
rect 31549 606808 39885 606827
rect 31549 606523 39705 606808
rect 30782 606504 39705 606523
rect 39849 606504 39885 606808
rect 40810 606781 42193 606841
rect 675407 606800 675887 606870
rect 30782 606446 39885 606504
rect 37316 606222 39885 606260
rect 37316 605918 37386 606222
rect 38090 606216 39885 606222
rect 38090 605918 39704 606216
rect 37316 605912 39704 605918
rect 39848 605912 39885 606216
rect 37316 605879 39885 605912
rect 675407 604960 675887 605030
rect 40810 604781 42193 604841
rect 675407 604408 675887 604478
rect 675407 603764 675887 603834
rect 675407 603120 675887 603190
rect 675407 600636 675887 600706
rect 675407 600084 675887 600154
rect 675407 599440 675887 599510
rect 675407 598796 675887 598866
rect 675407 598244 675887 598314
rect 675407 597600 675887 597670
rect 675407 596404 675887 596474
rect 675407 595760 675887 595830
rect 675407 593920 675887 593990
rect 41713 583410 42193 583480
rect 41713 581570 42193 581640
rect 41713 580926 42193 580996
rect 41713 579730 42193 579800
rect 41713 579086 42193 579156
rect 41713 578534 42193 578604
rect 41713 577890 42193 577960
rect 41713 577246 42193 577316
rect 41713 576694 42193 576764
rect 41713 574210 42193 574280
rect 41713 573566 42193 573636
rect 41713 572922 42193 572992
rect 41713 572370 42193 572440
rect 41713 570530 42193 570600
rect 41713 569886 42193 569956
rect 41713 569242 42193 569312
rect 41713 568690 42193 568760
rect 675407 567144 676767 567206
rect 40832 564525 40892 567008
rect 677626 566068 680341 566107
rect 677626 566064 679567 566068
rect 677626 565760 677649 566064
rect 677793 565764 679567 566064
rect 680271 565764 680341 566068
rect 677793 565760 680341 565764
rect 677626 565726 680341 565760
rect 677626 565463 686875 565540
rect 677626 565462 686108 565463
rect 675407 565142 676797 565204
rect 677626 565158 677648 565462
rect 677792 565159 686108 565462
rect 686812 565159 686875 565463
rect 677792 565158 686875 565159
rect 677626 565090 686875 565158
rect 30782 563827 39885 563896
rect 30782 563523 30845 563827
rect 31549 563808 39885 563827
rect 31549 563523 39705 563808
rect 30782 563504 39705 563523
rect 39849 563504 39885 563808
rect 40810 563781 42193 563841
rect 30782 563446 39885 563504
rect 675407 563440 675887 563510
rect 37316 563222 39885 563260
rect 37316 562918 37386 563222
rect 38090 563216 39885 563222
rect 38090 562918 39704 563216
rect 37316 562912 39704 562918
rect 39848 562912 39885 563216
rect 37316 562879 39885 562912
rect 675407 562888 675887 562958
rect 675407 562244 675887 562314
rect 40810 561781 42193 561841
rect 675407 561600 675887 561670
rect 675407 559760 675887 559830
rect 675407 559208 675887 559278
rect 675407 558564 675887 558634
rect 675407 557920 675887 557990
rect 675407 555436 675887 555506
rect 675407 554884 675887 554954
rect 675407 554240 675887 554310
rect 675407 553596 675887 553666
rect 675407 553044 675887 553114
rect 675407 552400 675887 552470
rect 675407 551204 675887 551274
rect 675407 550560 675887 550630
rect 675407 548720 675887 548790
rect 41713 540210 42193 540280
rect 41713 538370 42193 538440
rect 41713 537726 42193 537796
rect 41713 536530 42193 536600
rect 41713 535886 42193 535956
rect 41713 535334 42193 535404
rect 41713 534690 42193 534760
rect 41713 534046 42193 534116
rect 41713 533494 42193 533564
rect 41713 531010 42193 531080
rect 41713 530366 42193 530436
rect 41713 529722 42193 529792
rect 41713 529170 42193 529240
rect 41713 527330 42193 527400
rect 41713 526686 42193 526756
rect 41713 526042 42193 526112
rect 41713 525490 42193 525560
rect 40832 521519 40892 523808
rect 30782 520827 39885 520896
rect 30782 520523 30845 520827
rect 31549 520808 39885 520827
rect 31549 520523 39705 520808
rect 30782 520504 39705 520523
rect 39849 520504 39885 520808
rect 40810 520781 42193 520841
rect 30782 520446 39885 520504
rect 37316 520222 39885 520260
rect 37316 519918 37386 520222
rect 38090 520216 39885 520222
rect 38090 519918 39704 520216
rect 37316 519912 39704 519918
rect 39848 519912 39885 520216
rect 37316 519879 39885 519912
rect 40810 518781 42193 518841
rect 675407 513921 677812 518701
rect 675407 503942 677812 508722
rect 39874 493078 42193 497858
rect 39874 483099 42193 487879
rect 675407 474699 677752 474700
rect 675407 469901 676907 474699
rect 677705 469901 677752 474699
rect 675407 469900 677752 469901
rect 675407 469599 677549 469600
rect 675407 464949 675787 469599
rect 676585 464949 677549 469599
rect 675407 459861 676907 464649
rect 677705 459861 677752 464649
rect 675407 459860 677752 459861
rect 39870 455739 42193 455740
rect 39870 450953 39919 455739
rect 40717 450953 42193 455739
rect 39870 450951 42193 450953
rect 40051 446001 41039 450651
rect 41837 446001 42193 450651
rect 40051 446000 42193 446001
rect 39870 445699 42193 445700
rect 39870 440901 39919 445699
rect 40717 440901 42193 445699
rect 39870 440900 42193 440901
rect 675407 425721 677812 430501
rect 675407 415742 677812 420522
rect 41713 412610 42193 412680
rect 41713 410770 42193 410840
rect 41713 410126 42193 410196
rect 41713 408930 42193 409000
rect 41713 408286 42193 408356
rect 41713 407734 42193 407804
rect 41713 407090 42193 407160
rect 41713 406446 42193 406516
rect 41713 405894 42193 405964
rect 41713 403410 42193 403480
rect 41713 402766 42193 402836
rect 41713 402122 42193 402192
rect 41713 401570 42193 401640
rect 41713 399730 42193 399800
rect 41713 399086 42193 399156
rect 41713 398442 42193 398512
rect 41713 397890 42193 397960
rect 40832 392553 40892 396208
rect 30782 391827 39885 391896
rect 30782 391523 30845 391827
rect 31549 391808 39885 391827
rect 31549 391523 39705 391808
rect 30782 391504 39705 391523
rect 39849 391504 39885 391808
rect 40810 391781 42193 391841
rect 30782 391446 39885 391504
rect 37316 391222 39885 391260
rect 37316 390918 37386 391222
rect 38090 391216 39885 391222
rect 38090 390918 39704 391216
rect 37316 390912 39704 390918
rect 39848 390912 39885 391216
rect 37316 390879 39885 390912
rect 675407 390144 676767 390206
rect 40810 389781 42193 389841
rect 677626 389068 680341 389107
rect 677626 389064 679567 389068
rect 677626 388760 677649 389064
rect 677793 388764 679567 389064
rect 680271 388764 680341 389068
rect 677793 388760 680341 388764
rect 677626 388726 680341 388760
rect 677626 388463 686875 388540
rect 677626 388462 686108 388463
rect 675407 388142 676797 388204
rect 677626 388158 677648 388462
rect 677792 388159 686108 388462
rect 686812 388159 686875 388463
rect 677792 388158 686875 388159
rect 677626 388090 686875 388158
rect 675407 386240 675887 386310
rect 675407 385688 675887 385758
rect 675407 385044 675887 385114
rect 675407 384400 675887 384470
rect 675407 382560 675887 382630
rect 675407 382008 675887 382078
rect 675407 381364 675887 381434
rect 675407 380720 675887 380790
rect 675407 378236 675887 378306
rect 675407 377684 675887 377754
rect 675407 377040 675887 377110
rect 675407 376396 675887 376466
rect 675407 375844 675887 375914
rect 675407 375200 675887 375270
rect 675407 374004 675887 374074
rect 675407 373360 675887 373430
rect 675407 371520 675887 371590
rect 41713 369410 42193 369480
rect 41713 367570 42193 367640
rect 41713 366926 42193 366996
rect 41713 365730 42193 365800
rect 41713 365086 42193 365156
rect 41713 364534 42193 364604
rect 41713 363890 42193 363960
rect 41713 363246 42193 363316
rect 41713 362694 42193 362764
rect 41713 360210 42193 360280
rect 41713 359566 42193 359636
rect 41713 358922 42193 358992
rect 41713 358370 42193 358440
rect 41713 356530 42193 356600
rect 41713 355886 42193 355956
rect 41713 355242 42193 355312
rect 41713 354690 42193 354760
rect 40832 349533 40892 353008
rect 30782 348827 39885 348896
rect 30782 348523 30845 348827
rect 31549 348808 39885 348827
rect 31549 348523 39705 348808
rect 30782 348504 39705 348523
rect 39849 348504 39885 348808
rect 40810 348781 42193 348841
rect 30782 348446 39885 348504
rect 37316 348222 39885 348260
rect 37316 347918 37386 348222
rect 38090 348216 39885 348222
rect 38090 347918 39704 348216
rect 37316 347912 39704 347918
rect 39848 347912 39885 348216
rect 37316 347879 39885 347912
rect 40810 346781 42193 346841
rect 675407 345144 676767 345206
rect 677626 344068 680341 344107
rect 677626 344064 679567 344068
rect 677626 343760 677649 344064
rect 677793 343764 679567 344064
rect 680271 343764 680341 344068
rect 677793 343760 680341 343764
rect 677626 343726 680341 343760
rect 677626 343463 686875 343540
rect 677626 343462 686108 343463
rect 675407 343142 676797 343204
rect 677626 343158 677648 343462
rect 677792 343159 686108 343462
rect 686812 343159 686875 343463
rect 677792 343158 686875 343159
rect 677626 343090 686875 343158
rect 675407 341040 675887 341110
rect 675407 340488 675887 340558
rect 675407 339844 675887 339914
rect 675407 339200 675887 339270
rect 675407 337360 675887 337430
rect 675407 336808 675887 336878
rect 675407 336164 675887 336234
rect 675407 335520 675887 335590
rect 675407 333036 675887 333106
rect 675407 332484 675887 332554
rect 675407 331840 675887 331910
rect 675407 331196 675887 331266
rect 675407 330644 675887 330714
rect 675407 330000 675887 330070
rect 675407 328804 675887 328874
rect 675407 328160 675887 328230
rect 675407 326320 675887 326390
rect 41713 326210 42193 326280
rect 41713 324370 42193 324440
rect 41713 323726 42193 323796
rect 41713 322530 42193 322600
rect 41713 321886 42193 321956
rect 41713 321334 42193 321404
rect 41713 320690 42193 320760
rect 41713 320046 42193 320116
rect 41713 319494 42193 319564
rect 41713 317010 42193 317080
rect 41713 316366 42193 316436
rect 41713 315722 42193 315792
rect 41713 315170 42193 315240
rect 41713 313330 42193 313400
rect 41713 312686 42193 312756
rect 41713 312042 42193 312112
rect 41713 311490 42193 311560
rect 40832 306514 40892 309808
rect 30782 305827 39885 305896
rect 30782 305523 30845 305827
rect 31549 305808 39885 305827
rect 31549 305523 39705 305808
rect 30782 305504 39705 305523
rect 39849 305504 39885 305808
rect 40810 305781 42193 305841
rect 30782 305446 39885 305504
rect 37316 305222 39885 305260
rect 37316 304918 37386 305222
rect 38090 305216 39885 305222
rect 38090 304918 39704 305216
rect 37316 304912 39704 304918
rect 39848 304912 39885 305216
rect 37316 304879 39885 304912
rect 40810 303781 42193 303841
rect 675407 300144 676767 300206
rect 677626 299068 680341 299107
rect 677626 299064 679567 299068
rect 677626 298760 677649 299064
rect 677793 298764 679567 299064
rect 680271 298764 680341 299068
rect 677793 298760 680341 298764
rect 677626 298726 680341 298760
rect 677626 298463 686875 298540
rect 677626 298462 686108 298463
rect 675407 298142 676797 298204
rect 677626 298158 677648 298462
rect 677792 298159 686108 298462
rect 686812 298159 686875 298463
rect 677792 298158 686875 298159
rect 677626 298090 686875 298158
rect 675407 296040 675887 296110
rect 675407 295488 675887 295558
rect 675407 294844 675887 294914
rect 675407 294200 675887 294270
rect 675407 292360 675887 292430
rect 675407 291808 675887 291878
rect 675407 291164 675887 291234
rect 675407 290520 675887 290590
rect 675407 288036 675887 288106
rect 675407 287484 675887 287554
rect 675407 286840 675887 286910
rect 675407 286196 675887 286266
rect 675407 285644 675887 285714
rect 675407 285000 675887 285070
rect 675407 283804 675887 283874
rect 675407 283160 675887 283230
rect 41713 283010 42193 283080
rect 675407 281320 675887 281390
rect 41713 281170 42193 281240
rect 41713 280526 42193 280596
rect 41713 279330 42193 279400
rect 41713 278686 42193 278756
rect 41713 278134 42193 278204
rect 41713 277490 42193 277560
rect 41713 276846 42193 276916
rect 41713 276294 42193 276364
rect 41713 273810 42193 273880
rect 41713 273166 42193 273236
rect 41713 272522 42193 272592
rect 41713 271970 42193 272040
rect 41713 270130 42193 270200
rect 41713 269486 42193 269556
rect 41713 268842 42193 268912
rect 41713 268290 42193 268360
rect 40832 263525 40892 266624
rect 30782 262827 39885 262896
rect 30782 262523 30845 262827
rect 31549 262808 39885 262827
rect 31549 262523 39705 262808
rect 30782 262504 39705 262523
rect 39849 262504 39885 262808
rect 40810 262781 42193 262841
rect 30782 262446 39885 262504
rect 37316 262222 39885 262260
rect 37316 261918 37386 262222
rect 38090 262216 39885 262222
rect 38090 261918 39704 262216
rect 37316 261912 39704 261918
rect 39848 261912 39885 262216
rect 37316 261879 39885 261912
rect 40810 260781 42193 260841
rect 675407 255144 676767 255206
rect 677626 254068 680341 254107
rect 677626 254064 679567 254068
rect 677626 253760 677649 254064
rect 677793 253764 679567 254064
rect 680271 253764 680341 254068
rect 677793 253760 680341 253764
rect 677626 253726 680341 253760
rect 677626 253463 686875 253540
rect 677626 253462 686108 253463
rect 675407 253142 676797 253204
rect 677626 253158 677648 253462
rect 677792 253159 686108 253462
rect 686812 253159 686875 253463
rect 677792 253158 686875 253159
rect 677626 253090 686875 253158
rect 675407 251040 675887 251110
rect 675407 250488 675887 250558
rect 675407 249844 675887 249914
rect 675407 249200 675887 249270
rect 675407 247360 675887 247430
rect 675407 246808 675887 246878
rect 675407 246164 675887 246234
rect 675407 245520 675887 245590
rect 675407 243036 675887 243106
rect 675407 242484 675887 242554
rect 675407 241840 675887 241910
rect 675407 241196 675887 241266
rect 675407 240644 675887 240714
rect 675407 240000 675887 240070
rect 41713 239810 42193 239880
rect 675407 238804 675887 238874
rect 675407 238160 675887 238230
rect 41713 237970 42193 238040
rect 41713 237326 42193 237396
rect 675407 236320 675887 236390
rect 41713 236130 42193 236200
rect 41713 235486 42193 235556
rect 41713 234934 42193 235004
rect 41713 234290 42193 234360
rect 41713 233646 42193 233716
rect 41713 233094 42193 233164
rect 41713 230610 42193 230680
rect 41713 229966 42193 230036
rect 41713 229322 42193 229392
rect 41713 228770 42193 228840
rect 41713 226930 42193 227000
rect 41713 226286 42193 226356
rect 41713 225642 42193 225712
rect 41713 225090 42193 225160
rect 40832 220519 40892 223429
rect 30782 219827 39885 219896
rect 30782 219523 30845 219827
rect 31549 219808 39885 219827
rect 31549 219523 39705 219808
rect 30782 219504 39705 219523
rect 39849 219504 39885 219808
rect 40810 219781 42193 219841
rect 30782 219446 39885 219504
rect 37316 219222 39885 219260
rect 37316 218918 37386 219222
rect 38090 219216 39885 219222
rect 38090 218918 39704 219216
rect 37316 218912 39704 218918
rect 39848 218912 39885 219216
rect 37316 218879 39885 218912
rect 40810 217781 42193 217841
rect 675407 210144 676767 210206
rect 677626 209068 680341 209107
rect 677626 209064 679567 209068
rect 677626 208760 677649 209064
rect 677793 208764 679567 209064
rect 680271 208764 680341 209068
rect 677793 208760 680341 208764
rect 677626 208726 680341 208760
rect 677626 208463 686875 208540
rect 677626 208462 686108 208463
rect 675407 208142 676797 208204
rect 677626 208158 677648 208462
rect 677792 208159 686108 208462
rect 686812 208159 686875 208463
rect 677792 208158 686875 208159
rect 677626 208090 686875 208158
rect 675407 205840 675887 205910
rect 675407 205288 675887 205358
rect 675407 204644 675887 204714
rect 675407 204000 675887 204070
rect 675407 202160 675887 202230
rect 675407 201608 675887 201678
rect 675407 200964 675887 201034
rect 675407 200320 675887 200390
rect 675407 197836 675887 197906
rect 675407 197284 675887 197354
rect 41713 196610 42193 196680
rect 675407 196640 675887 196710
rect 675407 195996 675887 196066
rect 675407 195444 675887 195514
rect 41713 194770 42193 194840
rect 675407 194800 675887 194870
rect 41713 194126 42193 194196
rect 675407 193604 675887 193674
rect 41713 192930 42193 193000
rect 675407 192960 675887 193030
rect 41713 192286 42193 192356
rect 41713 191734 42193 191804
rect 41713 191090 42193 191160
rect 675407 191120 675887 191190
rect 41713 190446 42193 190516
rect 41713 189894 42193 189964
rect 41713 187410 42193 187480
rect 41713 186766 42193 186836
rect 41713 186122 42193 186192
rect 41713 185570 42193 185640
rect 41713 183730 42193 183800
rect 41713 183086 42193 183156
rect 41713 182442 42193 182512
rect 41713 181890 42193 181960
rect 40832 177543 40892 180230
rect 30782 176827 39885 176896
rect 30782 176523 30845 176827
rect 31549 176808 39885 176827
rect 31549 176523 39705 176808
rect 30782 176504 39705 176523
rect 39849 176504 39885 176808
rect 40810 176781 42193 176841
rect 30782 176446 39885 176504
rect 37316 176222 39885 176260
rect 37316 175918 37386 176222
rect 38090 176216 39885 176222
rect 38090 175918 39704 176216
rect 37316 175912 39704 175918
rect 39848 175912 39885 176216
rect 37316 175879 39885 175912
rect 40810 174781 42193 174841
rect 675407 165144 676767 165206
rect 677626 164068 680341 164107
rect 677626 164064 679567 164068
rect 677626 163760 677649 164064
rect 677793 163764 679567 164064
rect 680271 163764 680341 164068
rect 677793 163760 680341 163764
rect 677626 163726 680341 163760
rect 677626 163463 686875 163540
rect 677626 163462 686108 163463
rect 675407 163142 676797 163204
rect 677626 163158 677648 163462
rect 677792 163159 686108 163462
rect 686812 163159 686875 163463
rect 677792 163158 686875 163159
rect 677626 163090 686875 163158
rect 675407 160840 675887 160910
rect 675407 160288 675887 160358
rect 675407 159644 675887 159714
rect 675407 159000 675887 159070
rect 675407 157160 675887 157230
rect 675407 156608 675887 156678
rect 675407 155964 675887 156034
rect 675407 155320 675887 155390
rect 675407 152836 675887 152906
rect 675407 152284 675887 152354
rect 675407 151640 675887 151710
rect 675407 150996 675887 151066
rect 675407 150444 675887 150514
rect 675407 149800 675887 149870
rect 675407 148604 675887 148674
rect 675407 147960 675887 148030
rect 675407 146120 675887 146190
rect 39790 120278 42193 125058
rect 675407 120144 676744 120206
rect 677626 119068 680341 119107
rect 677626 119064 679567 119068
rect 677626 118760 677649 119064
rect 677793 118764 679567 119064
rect 680271 118764 680341 119068
rect 677793 118760 680341 118764
rect 677626 118726 680341 118760
rect 677626 118463 686875 118540
rect 677626 118462 686108 118463
rect 675407 118142 676716 118204
rect 677626 118158 677648 118462
rect 677792 118159 686108 118462
rect 686812 118159 686875 118463
rect 677792 118158 686875 118159
rect 677626 118090 686875 118158
rect 675407 115640 675887 115710
rect 675407 115088 675887 115158
rect 39790 110299 42193 115079
rect 675407 114444 675887 114514
rect 675407 113800 675887 113870
rect 675407 111960 675887 112030
rect 675407 111408 675887 111478
rect 675407 110764 675887 110834
rect 675407 110120 675887 110190
rect 675407 107636 675887 107706
rect 675407 107084 675887 107154
rect 675407 106440 675887 106510
rect 675407 105796 675887 105866
rect 675407 105244 675887 105314
rect 675407 104600 675887 104670
rect 675407 103404 675887 103474
rect 675407 102760 675887 102830
rect 19586 101323 31666 101352
rect 19586 99489 30809 101323
rect 31637 99489 31666 101323
rect 675407 100920 675887 100990
rect 19586 99457 31666 99489
rect 17843 95353 17912 95915
rect 18569 95576 18629 95915
rect 18934 95800 18994 95915
rect 18929 95795 19201 95800
rect 18929 95739 18934 95795
rect 19194 95739 19201 95795
rect 18929 95729 19201 95739
rect 41447 95795 42193 95802
rect 41447 95739 41478 95795
rect 41829 95739 42193 95795
rect 41447 95732 42193 95739
rect 18563 95571 18835 95576
rect 18563 95515 18569 95571
rect 18829 95515 18835 95571
rect 18563 95505 18835 95515
rect 41447 95571 42193 95579
rect 41447 95515 41470 95571
rect 41821 95515 42193 95571
rect 41447 95509 42193 95515
rect 17837 95347 18118 95353
rect 17837 95291 17843 95347
rect 18112 95291 18118 95347
rect 17837 95283 18118 95291
rect 41447 95347 42193 95354
rect 41447 95291 41467 95347
rect 41818 95291 42193 95347
rect 41447 95284 42193 95291
rect 19024 94481 38186 94499
rect 19024 92770 19050 94481
rect 19352 94456 38186 94481
rect 19352 92802 37362 94456
rect 38160 92802 38186 94456
rect 19352 92770 38186 92802
rect 19024 92753 38186 92770
rect 39566 78151 42193 82940
rect 39566 68100 42193 72900
rect 78942 39820 83722 42193
rect 88921 39820 93701 42194
rect 145825 40874 145891 40877
rect 145825 40872 148252 40874
rect 145825 40816 145830 40872
rect 145886 40816 148252 40872
rect 145825 40814 148252 40816
rect 202708 40873 202778 40878
rect 202708 40871 203064 40873
rect 202708 40815 202715 40871
rect 202771 40815 203064 40871
rect 205919 40870 205989 40877
rect 145825 40811 145891 40814
rect 202708 40813 203064 40815
rect 205764 40814 205926 40870
rect 205982 40814 205989 40870
rect 202708 40808 202778 40813
rect 205764 40810 205989 40814
rect 205919 40807 205989 40810
rect 141705 40352 141776 40355
rect 141705 40350 148181 40352
rect 141705 40289 141710 40350
rect 141771 40347 148181 40350
rect 141771 40292 148107 40347
rect 141771 40289 141776 40292
rect 141705 40284 141776 40289
rect 148102 40287 148107 40292
rect 148167 40292 148181 40347
rect 148167 40287 148172 40292
rect 148102 40282 148172 40287
rect 133094 40158 144010 40218
rect 133094 39984 133154 40158
rect 143407 40095 143519 40097
rect 143402 40090 143524 40095
rect 143402 40034 143435 40090
rect 143491 40034 143524 40090
rect 143402 39992 143524 40034
rect 143950 39984 144010 40158
rect 145832 40132 145902 40148
rect 145832 40076 145839 40132
rect 145895 40076 145902 40132
rect 145832 39982 145902 40076
rect 148901 39873 149351 39914
rect 148901 39729 148969 39873
rect 149273 39729 149351 39873
rect 148901 31573 149351 39729
rect 149537 39872 149918 39914
rect 149537 39728 149571 39872
rect 149875 39728 149918 39872
rect 149537 38114 149918 39728
rect 203701 39873 204151 39895
rect 203701 39729 203769 39873
rect 204073 39729 204151 39873
rect 149537 37410 149575 38114
rect 149879 37410 149918 38114
rect 149537 37340 149918 37410
rect 153624 38176 154090 38249
rect 153624 37340 153655 38176
rect 154064 37340 154090 38176
rect 153024 34784 153490 34873
rect 153024 33947 153046 34784
rect 153462 33947 153490 34784
rect 148901 30869 148970 31573
rect 149274 30869 149351 31573
rect 148901 30806 149351 30869
rect 152424 31631 152890 31723
rect 152424 30800 152457 31631
rect 152858 30800 152890 31631
rect 152424 20597 152890 30800
rect 152424 20133 152445 20597
rect 152866 20133 152890 20597
rect 152424 20111 152890 20133
rect 153024 20597 153490 33947
rect 153024 20133 153045 20597
rect 153466 20133 153490 20597
rect 153024 20111 153490 20133
rect 153624 20597 154090 37340
rect 153624 20133 153642 20597
rect 154063 20133 154090 20597
rect 153624 20111 154090 20133
rect 154224 35989 154690 36081
rect 154224 35178 154268 35989
rect 154659 35178 154690 35989
rect 154224 20600 154690 35178
rect 203701 31573 204151 39729
rect 204337 39872 204718 39895
rect 204337 39728 204371 39872
rect 204675 39728 204718 39872
rect 204337 38114 204718 39728
rect 241420 39564 246049 42193
rect 251300 39564 256100 42193
rect 311308 40873 311378 40878
rect 315488 40874 315558 40881
rect 315488 40873 315495 40874
rect 311308 40871 312684 40873
rect 311308 40815 311315 40871
rect 311371 40815 312684 40871
rect 311308 40813 312684 40815
rect 315360 40818 315495 40873
rect 315551 40818 315558 40874
rect 315360 40813 315558 40818
rect 311308 40808 311378 40813
rect 315488 40811 315558 40813
rect 366108 40873 366178 40878
rect 366108 40871 367484 40873
rect 366108 40815 366115 40871
rect 366171 40815 367484 40871
rect 370293 40870 370363 40877
rect 370293 40869 370300 40870
rect 366108 40813 367484 40815
rect 370159 40814 370300 40869
rect 370356 40814 370363 40870
rect 366108 40808 366178 40813
rect 370159 40809 370363 40814
rect 370293 40807 370363 40809
rect 420908 40873 420978 40878
rect 475708 40873 475778 40878
rect 420908 40871 422262 40873
rect 420908 40815 420915 40871
rect 420971 40815 422262 40871
rect 475708 40871 477055 40873
rect 425106 40864 425176 40865
rect 420908 40813 422262 40815
rect 424960 40858 425176 40864
rect 420908 40808 420978 40813
rect 424960 40804 425113 40858
rect 425106 40802 425113 40804
rect 425169 40802 425176 40858
rect 475708 40815 475715 40871
rect 475771 40815 477055 40871
rect 479906 40872 479976 40879
rect 479906 40869 479913 40872
rect 475708 40813 477055 40815
rect 479767 40816 479913 40869
rect 479969 40816 479976 40872
rect 475708 40808 475778 40813
rect 479767 40809 479976 40816
rect 530508 40873 530578 40878
rect 530508 40871 531856 40873
rect 530508 40815 530515 40871
rect 530571 40815 531856 40871
rect 534763 40863 534833 40867
rect 530508 40813 531856 40815
rect 534569 40860 534833 40863
rect 530508 40808 530578 40813
rect 534569 40804 534770 40860
rect 534826 40804 534833 40860
rect 534569 40803 534833 40804
rect 425106 40795 425176 40802
rect 534763 40797 534833 40803
rect 313301 39873 313751 39895
rect 313301 39729 313369 39873
rect 313673 39729 313751 39873
rect 204337 37410 204375 38114
rect 204679 37410 204718 38114
rect 204337 37340 204718 37410
rect 203701 30869 203770 31573
rect 204074 30869 204151 31573
rect 203701 30806 204151 30869
rect 313301 31573 313751 39729
rect 313937 39872 314318 39895
rect 313937 39728 313971 39872
rect 314275 39728 314318 39872
rect 313937 38114 314318 39728
rect 313937 37410 313975 38114
rect 314279 37410 314318 38114
rect 313937 37340 314318 37410
rect 368101 39873 368551 39895
rect 368101 39729 368169 39873
rect 368473 39729 368551 39873
rect 313301 30869 313370 31573
rect 313674 30869 313751 31573
rect 313301 30806 313751 30869
rect 368101 31573 368551 39729
rect 368737 39872 369118 39895
rect 368737 39728 368771 39872
rect 369075 39728 369118 39872
rect 368737 38114 369118 39728
rect 368737 37410 368775 38114
rect 369079 37410 369118 38114
rect 368737 37340 369118 37410
rect 422901 39873 423351 39895
rect 422901 39729 422969 39873
rect 423273 39729 423351 39873
rect 368101 30869 368170 31573
rect 368474 30869 368551 31573
rect 368101 30806 368551 30869
rect 422901 31573 423351 39729
rect 423537 39872 423918 39895
rect 423537 39728 423571 39872
rect 423875 39728 423918 39872
rect 423537 38114 423918 39728
rect 423537 37410 423575 38114
rect 423879 37410 423918 38114
rect 423537 37340 423918 37410
rect 477701 39873 478151 39895
rect 477701 39729 477769 39873
rect 478073 39729 478151 39873
rect 422901 30869 422970 31573
rect 423274 30869 423351 31573
rect 422901 30806 423351 30869
rect 477701 31573 478151 39729
rect 478337 39872 478718 39895
rect 478337 39728 478371 39872
rect 478675 39728 478718 39872
rect 478337 38114 478718 39728
rect 478337 37410 478375 38114
rect 478679 37410 478718 38114
rect 478337 37340 478718 37410
rect 532501 39873 532951 39895
rect 532501 39729 532569 39873
rect 532873 39729 532951 39873
rect 477701 30869 477770 31573
rect 478074 30869 478151 31573
rect 477701 30806 478151 30869
rect 532501 31573 532951 39729
rect 533137 39872 533518 39895
rect 533137 39728 533171 39872
rect 533475 39728 533518 39872
rect 569142 39844 573922 42193
rect 579121 39844 583901 42193
rect 622942 39906 627722 42193
rect 632921 39906 637701 42193
rect 533137 38114 533518 39728
rect 533137 37410 533175 38114
rect 533479 37410 533518 38114
rect 533137 37340 533518 37410
rect 640496 38118 641506 38169
rect 640496 37380 640578 38118
rect 641436 37380 641506 38118
rect 532501 30869 532570 31573
rect 532874 30869 532951 31573
rect 532501 30806 532951 30869
rect 154224 20136 154248 20600
rect 154669 20136 154690 20600
rect 154224 20111 154690 20136
rect 640496 16570 641506 37380
rect 640496 15710 640542 16570
rect 641444 15710 641506 16570
rect 640496 15658 641506 15710
rect 642098 32580 643108 32640
rect 642098 32020 642152 32580
rect 643060 32020 643108 32580
rect 642098 16566 643108 32020
rect 642098 15706 642146 16566
rect 643048 15706 643108 16566
rect 642098 15658 643108 15706
rect 643899 15326 643969 15331
rect 643899 15266 643904 15326
rect 643964 15266 643969 15326
rect 643899 15261 643969 15266
rect 643340 14506 643410 14511
rect 643340 14446 643345 14506
rect 643405 14446 643410 14506
rect 643340 14441 643410 14446
rect 650120 14498 650190 14503
rect 650120 14438 650125 14498
rect 650185 14438 650190 14498
rect 650120 14433 650190 14438
rect 649856 13689 649926 13694
rect 643676 13684 643746 13689
rect 643676 13624 643681 13684
rect 643741 13624 643746 13684
rect 649856 13629 649861 13689
rect 649921 13629 649926 13689
rect 649856 13624 649926 13629
rect 643676 13619 643746 13624
rect 649744 12883 649814 12888
rect 649744 12823 649749 12883
rect 649809 12823 649814 12883
rect 649744 12818 649814 12823
rect 643562 12607 643632 12612
rect 643562 12547 643567 12607
rect 643627 12547 643632 12607
rect 643562 12542 643632 12547
rect 643450 11794 643520 11799
rect 643450 11734 643455 11794
rect 643515 11734 643520 11794
rect 651692 11792 651758 11795
rect 643450 11729 643520 11734
rect 650182 11790 651758 11792
rect 650182 11734 651697 11790
rect 651753 11734 651758 11790
rect 650182 11732 651758 11734
rect 651692 11729 651758 11732
rect 649991 10981 650061 10986
rect 643879 10975 643949 10980
rect 643879 10915 643884 10975
rect 643944 10915 643949 10975
rect 649991 10921 649996 10981
rect 650056 10921 650061 10981
rect 649991 10916 650061 10921
rect 643879 10910 643949 10915
rect 651913 10162 651983 10167
rect 651913 10161 651918 10162
rect 650163 10102 651918 10161
rect 651978 10102 651983 10162
rect 650163 10101 651983 10102
rect 651913 10097 651983 10101
<< via3 >>
rect 71377 1006097 71681 1006801
rect 70772 999556 71076 1000260
rect 70776 997758 71080 997902
rect 122577 1006097 122881 1006801
rect 71358 997757 71662 997901
rect 121972 999556 122276 1000260
rect 121976 997758 122280 997902
rect 173777 1006097 174081 1006801
rect 122558 997757 122862 997901
rect 173172 999556 173476 1000260
rect 173176 997758 173480 997902
rect 224977 1006097 225281 1006801
rect 173758 997757 174062 997901
rect 224372 999556 224676 1000260
rect 224376 997758 224680 997902
rect 276177 1006097 276481 1006801
rect 224958 997757 225257 997901
rect 275572 999556 275876 1000260
rect 275576 997758 275880 997902
rect 380577 1006097 380881 1006801
rect 276158 997757 276462 997901
rect 379972 999556 380276 1000260
rect 379976 997758 380280 997902
rect 469577 1006097 469881 1006801
rect 380558 997757 380862 997901
rect 468972 999556 469276 1000260
rect 468976 997758 469280 997902
rect 520777 1006097 521081 1006801
rect 469558 997757 469862 997901
rect 520172 999556 520476 1000260
rect 520176 997758 520480 997902
rect 620177 1006097 620481 1006801
rect 520758 997757 521062 997901
rect 619572 999556 619876 1000260
rect 619576 997758 619880 997902
rect 620158 997757 620462 997901
rect 677649 969760 677793 970064
rect 679567 969764 680271 970068
rect 677648 969158 677792 969462
rect 686108 969159 686812 969463
rect 30845 948523 31549 948827
rect 39705 948504 39849 948808
rect 37386 947918 38090 948222
rect 39704 947912 39848 948216
rect 41039 922151 41837 926939
rect 39919 917191 40717 921851
rect 675787 917701 676585 922499
rect 41039 912101 41837 916899
rect 676907 912749 677705 917409
rect 675787 907661 676585 912449
rect 677649 879760 677793 880064
rect 679567 879764 680271 880068
rect 677648 879158 677792 879462
rect 686108 879159 686812 879463
rect 677649 790760 677793 791064
rect 679567 790764 680271 791068
rect 677648 790158 677792 790462
rect 686108 790159 686812 790463
rect 30845 778523 31549 778827
rect 39705 778504 39849 778808
rect 37386 777918 38090 778222
rect 39704 777912 39848 778216
rect 677649 745760 677793 746064
rect 679567 745764 680271 746068
rect 677648 745158 677792 745462
rect 686108 745159 686812 745463
rect 30845 735523 31549 735827
rect 39705 735504 39849 735808
rect 37386 734918 38090 735222
rect 39704 734912 39848 735216
rect 677649 700760 677793 701064
rect 679567 700764 680271 701068
rect 677648 700158 677792 700462
rect 686108 700159 686812 700463
rect 30845 692523 31549 692827
rect 39705 692504 39849 692808
rect 37386 691918 38090 692222
rect 39704 691912 39848 692216
rect 677649 655760 677793 656064
rect 679567 655764 680271 656068
rect 677648 655158 677792 655462
rect 686108 655159 686812 655463
rect 30845 649523 31549 649827
rect 39705 649504 39849 649808
rect 37386 648918 38090 649222
rect 39704 648912 39848 649216
rect 677649 610760 677793 611064
rect 679567 610764 680271 611068
rect 677648 610158 677792 610462
rect 686108 610159 686812 610463
rect 30845 606523 31549 606827
rect 39705 606504 39849 606808
rect 37386 605918 38090 606222
rect 39704 605912 39848 606216
rect 677649 565760 677793 566064
rect 679567 565764 680271 566068
rect 677648 565158 677792 565462
rect 686108 565159 686812 565463
rect 30845 563523 31549 563827
rect 39705 563504 39849 563808
rect 37386 562918 38090 563222
rect 39704 562912 39848 563216
rect 30845 520523 31549 520827
rect 39705 520504 39849 520808
rect 37386 519918 38090 520222
rect 39704 519912 39848 520216
rect 676907 469901 677705 474699
rect 675787 464949 676585 469599
rect 676907 459861 677705 464649
rect 39919 450953 40717 455739
rect 41039 446001 41837 450651
rect 39919 440901 40717 445699
rect 30845 391523 31549 391827
rect 39705 391504 39849 391808
rect 37386 390918 38090 391222
rect 39704 390912 39848 391216
rect 677649 388760 677793 389064
rect 679567 388764 680271 389068
rect 677648 388158 677792 388462
rect 686108 388159 686812 388463
rect 30845 348523 31549 348827
rect 39705 348504 39849 348808
rect 37386 347918 38090 348222
rect 39704 347912 39848 348216
rect 677649 343760 677793 344064
rect 679567 343764 680271 344068
rect 677648 343158 677792 343462
rect 686108 343159 686812 343463
rect 30845 305523 31549 305827
rect 39705 305504 39849 305808
rect 37386 304918 38090 305222
rect 39704 304912 39848 305216
rect 677649 298760 677793 299064
rect 679567 298764 680271 299068
rect 677648 298158 677792 298462
rect 686108 298159 686812 298463
rect 30845 262523 31549 262827
rect 39705 262504 39849 262808
rect 37386 261918 38090 262222
rect 39704 261912 39848 262216
rect 677649 253760 677793 254064
rect 679567 253764 680271 254068
rect 677648 253158 677792 253462
rect 686108 253159 686812 253463
rect 30845 219523 31549 219827
rect 39705 219504 39849 219808
rect 37386 218918 38090 219222
rect 39704 218912 39848 219216
rect 677649 208760 677793 209064
rect 679567 208764 680271 209068
rect 677648 208158 677792 208462
rect 686108 208159 686812 208463
rect 30845 176523 31549 176827
rect 39705 176504 39849 176808
rect 37386 175918 38090 176222
rect 39704 175912 39848 176216
rect 677649 163760 677793 164064
rect 679567 163764 680271 164068
rect 677648 163158 677792 163462
rect 686108 163159 686812 163463
rect 677649 118760 677793 119064
rect 679567 118764 680271 119068
rect 677648 118158 677792 118462
rect 686108 118159 686812 118463
rect 30809 99489 31637 101323
rect 19050 92770 19352 94481
rect 37362 92802 38160 94456
rect 148969 39729 149273 39873
rect 149571 39728 149875 39872
rect 203769 39729 204073 39873
rect 149575 37410 149879 38114
rect 153655 37340 154064 38176
rect 153046 33947 153462 34784
rect 148970 30869 149274 31573
rect 152457 30800 152858 31631
rect 152445 20133 152866 20597
rect 153045 20133 153466 20597
rect 153642 20133 154063 20597
rect 154268 35178 154659 35989
rect 204371 39728 204675 39872
rect 313369 39729 313673 39873
rect 204375 37410 204679 38114
rect 203770 30869 204074 31573
rect 313971 39728 314275 39872
rect 313975 37410 314279 38114
rect 368169 39729 368473 39873
rect 313370 30869 313674 31573
rect 368771 39728 369075 39872
rect 368775 37410 369079 38114
rect 422969 39729 423273 39873
rect 368170 30869 368474 31573
rect 423571 39728 423875 39872
rect 423575 37410 423879 38114
rect 477769 39729 478073 39873
rect 422970 30869 423274 31573
rect 478371 39728 478675 39872
rect 478375 37410 478679 38114
rect 532569 39729 532873 39873
rect 477770 30869 478074 31573
rect 533171 39728 533475 39872
rect 533175 37410 533479 38114
rect 640578 37380 641436 38118
rect 532570 30869 532874 31573
rect 154248 20136 154669 20600
rect 640542 15710 641444 16570
rect 642152 32020 643060 32580
rect 642146 15706 643048 16566
<< metal4 >>
rect 71346 1006801 71711 1006827
rect 71346 1006097 71377 1006801
rect 71681 1006097 71711 1006801
rect 71346 1006070 71711 1006097
rect 122546 1006801 122911 1006827
rect 122546 1006097 122577 1006801
rect 122881 1006097 122911 1006801
rect 122546 1006070 122911 1006097
rect 173746 1006801 174111 1006827
rect 173746 1006097 173777 1006801
rect 174081 1006097 174111 1006801
rect 173746 1006070 174111 1006097
rect 224946 1006801 225311 1006827
rect 224946 1006097 224977 1006801
rect 225281 1006097 225311 1006801
rect 224946 1006070 225311 1006097
rect 276146 1006801 276511 1006827
rect 276146 1006097 276177 1006801
rect 276481 1006097 276511 1006801
rect 276146 1006070 276511 1006097
rect 380546 1006801 380911 1006827
rect 380546 1006097 380577 1006801
rect 380881 1006097 380911 1006801
rect 380546 1006070 380911 1006097
rect 469546 1006801 469911 1006827
rect 469546 1006097 469577 1006801
rect 469881 1006097 469911 1006801
rect 469546 1006070 469911 1006097
rect 520746 1006801 521111 1006827
rect 520746 1006097 520777 1006801
rect 521081 1006097 521111 1006801
rect 520746 1006070 521111 1006097
rect 620146 1006801 620511 1006827
rect 620146 1006097 620177 1006801
rect 620481 1006097 620511 1006801
rect 620146 1006070 620511 1006097
rect 70760 1000260 71088 1000298
rect 70760 999556 70772 1000260
rect 71076 999556 71088 1000260
rect 70760 999517 71088 999556
rect 121960 1000260 122288 1000298
rect 121960 999556 121972 1000260
rect 122276 999556 122288 1000260
rect 121960 999517 122288 999556
rect 173160 1000260 173488 1000298
rect 173160 999556 173172 1000260
rect 173476 999556 173488 1000260
rect 173160 999517 173488 999556
rect 224360 1000260 224688 1000298
rect 224360 999556 224372 1000260
rect 224676 999556 224688 1000260
rect 224360 999517 224688 999556
rect 275560 1000260 275888 1000298
rect 275560 999556 275572 1000260
rect 275876 999556 275888 1000260
rect 275560 999517 275888 999556
rect 379960 1000260 380288 1000298
rect 379960 999556 379972 1000260
rect 380276 999556 380288 1000260
rect 379960 999517 380288 999556
rect 468960 1000260 469288 1000298
rect 468960 999556 468972 1000260
rect 469276 999556 469288 1000260
rect 468960 999517 469288 999556
rect 520160 1000260 520488 1000298
rect 520160 999556 520172 1000260
rect 520476 999556 520488 1000260
rect 520160 999517 520488 999556
rect 619560 1000260 619888 1000298
rect 619560 999556 619572 1000260
rect 619876 999556 619888 1000260
rect 619560 999517 619888 999556
rect 70766 997902 71085 997909
rect 70766 997758 70776 997902
rect 71080 997758 71085 997902
rect 71353 997901 71672 997909
rect 70766 997752 71085 997758
rect 71337 997757 71358 997901
rect 71662 997757 71672 997901
rect 71337 997752 71672 997757
rect 121969 997902 122286 997907
rect 121969 997758 121976 997902
rect 122280 997758 122286 997902
rect 122553 997901 122870 997906
rect 121969 997754 122286 997758
rect 122537 997757 122558 997901
rect 122862 997757 122870 997901
rect 70837 997522 71017 997752
rect 71337 997522 71517 997752
rect 122037 997522 122217 997754
rect 122537 997753 122870 997757
rect 173169 997902 173485 997907
rect 173169 997758 173176 997902
rect 173480 997758 173485 997902
rect 173753 997901 174069 997909
rect 122537 997522 122717 997753
rect 173169 997751 173485 997758
rect 173737 997757 173758 997901
rect 174062 997757 174069 997901
rect 173737 997753 174069 997757
rect 224373 997902 224683 997905
rect 224373 997758 224376 997902
rect 224680 997758 224683 997902
rect 224952 997901 225262 997903
rect 224373 997755 224683 997758
rect 224937 997757 224958 997901
rect 225257 997757 225262 997901
rect 173237 997522 173417 997751
rect 173737 997522 173917 997753
rect 224437 997522 224617 997755
rect 224937 997753 225262 997757
rect 275572 997902 275883 997905
rect 275572 997758 275576 997902
rect 275880 997758 275883 997902
rect 276155 997901 276466 997905
rect 275572 997754 275883 997758
rect 276137 997757 276158 997901
rect 276462 997757 276466 997901
rect 276137 997754 276466 997757
rect 379971 997902 380285 997905
rect 379971 997758 379976 997902
rect 380280 997758 380285 997902
rect 380555 997901 380869 997905
rect 224937 997522 225117 997753
rect 275637 997522 275817 997754
rect 276137 997522 276317 997754
rect 379971 997753 380285 997758
rect 380537 997757 380558 997901
rect 380862 997757 380869 997901
rect 380537 997753 380869 997757
rect 468973 997902 469283 997904
rect 468973 997758 468976 997902
rect 469280 997758 469283 997902
rect 469555 997901 469864 997904
rect 468973 997754 469283 997758
rect 469537 997757 469558 997901
rect 469862 997757 469864 997901
rect 469537 997754 469864 997757
rect 520172 997902 520482 997906
rect 520172 997758 520176 997902
rect 520480 997758 520482 997902
rect 520754 997901 521064 997906
rect 380037 997522 380217 997753
rect 380537 997522 380717 997753
rect 469037 997522 469217 997754
rect 469537 997522 469717 997754
rect 520172 997753 520482 997758
rect 520737 997757 520758 997901
rect 521062 997757 521064 997901
rect 520737 997753 521064 997757
rect 619572 997902 619883 997905
rect 619572 997758 619576 997902
rect 619880 997758 619883 997902
rect 620154 997901 620465 997904
rect 619572 997754 619883 997758
rect 620137 997757 620158 997901
rect 620462 997757 620465 997901
rect 520237 997522 520417 997753
rect 520737 997522 520917 997753
rect 619637 997522 619817 997754
rect 620137 997753 620465 997757
rect 620137 997522 620317 997753
rect 677642 970064 677801 970072
rect 677642 970003 677649 970064
rect 677533 969823 677649 970003
rect 677642 969760 677649 969823
rect 677793 969760 677801 970064
rect 677642 969754 677801 969760
rect 679528 970068 680309 970080
rect 679528 969764 679567 970068
rect 680271 969764 680309 970068
rect 679528 969752 680309 969764
rect 677533 969469 677792 969503
rect 677533 969462 677803 969469
rect 677533 969323 677648 969462
rect 677644 969158 677648 969323
rect 677792 969158 677803 969462
rect 677644 969151 677803 969158
rect 686081 969463 686838 969494
rect 686081 969159 686108 969463
rect 686812 969159 686838 969463
rect 686081 969129 686838 969159
rect 30819 948827 31576 948857
rect 30819 948523 30845 948827
rect 31549 948523 31576 948827
rect 30819 948492 31576 948523
rect 39698 948808 39857 948813
rect 39698 948504 39705 948808
rect 39849 948663 39857 948808
rect 39849 948504 40124 948663
rect 39698 948494 40124 948504
rect 39705 948483 40124 948494
rect 37348 948222 38129 948234
rect 37348 947918 37386 948222
rect 38090 947918 38129 948222
rect 37348 947906 38129 947918
rect 39697 948216 39856 948224
rect 39697 947912 39704 948216
rect 39848 948163 39856 948216
rect 39848 947983 40124 948163
rect 39848 947912 39856 947983
rect 39697 947905 39856 947912
rect 41038 926939 41838 926940
rect 41038 922151 41039 926939
rect 41837 922151 41838 926939
rect 41038 922150 41838 922151
rect 675786 922499 676586 922500
rect 39918 921851 40718 921852
rect 39918 917191 39919 921851
rect 40717 917191 40718 921851
rect 675786 917701 675787 922499
rect 676585 917701 676586 922499
rect 675786 917700 676586 917701
rect 39918 917190 40718 917191
rect 676906 917409 677706 917410
rect 41038 916899 41838 916900
rect 41038 912101 41039 916899
rect 41837 912101 41838 916899
rect 676906 912749 676907 917409
rect 677705 912749 677706 917409
rect 676906 912748 677706 912749
rect 41038 912100 41838 912101
rect 675786 912449 676586 912450
rect 675786 907661 675787 912449
rect 676585 907661 676586 912449
rect 675786 907660 676586 907661
rect 677643 880064 677800 880074
rect 677643 880003 677649 880064
rect 677533 879823 677649 880003
rect 677643 879760 677649 879823
rect 677793 879760 677800 880064
rect 677643 879754 677800 879760
rect 679528 880068 680309 880080
rect 679528 879764 679567 880068
rect 680271 879764 680309 880068
rect 679528 879752 680309 879764
rect 677533 879470 677792 879503
rect 677533 879462 677799 879470
rect 677533 879323 677648 879462
rect 677642 879158 677648 879323
rect 677792 879158 677799 879462
rect 677642 879150 677799 879158
rect 686081 879463 686838 879494
rect 686081 879159 686108 879463
rect 686812 879159 686838 879463
rect 686081 879129 686838 879159
rect 677642 791064 677798 791075
rect 677642 791003 677649 791064
rect 677533 790823 677649 791003
rect 677642 790760 677649 790823
rect 677793 790760 677798 791064
rect 677642 790755 677798 790760
rect 679528 791068 680309 791080
rect 679528 790764 679567 791068
rect 680271 790764 680309 791068
rect 679528 790752 680309 790764
rect 677533 790472 677792 790503
rect 677533 790462 677798 790472
rect 677533 790323 677648 790462
rect 677642 790158 677648 790323
rect 677792 790158 677798 790462
rect 677642 790152 677798 790158
rect 686081 790463 686838 790494
rect 686081 790159 686108 790463
rect 686812 790159 686838 790463
rect 686081 790129 686838 790159
rect 30819 778827 31576 778857
rect 30819 778523 30845 778827
rect 31549 778523 31576 778827
rect 30819 778492 31576 778523
rect 39695 778808 39861 778822
rect 39695 778504 39705 778808
rect 39849 778663 39861 778808
rect 39849 778504 40124 778663
rect 39695 778494 40124 778504
rect 39705 778483 40124 778494
rect 37348 778222 38129 778234
rect 37348 777918 37386 778222
rect 38090 777918 38129 778222
rect 37348 777906 38129 777918
rect 39688 778216 39854 778230
rect 39688 777912 39704 778216
rect 39848 778163 39854 778216
rect 39848 777983 40124 778163
rect 39848 777912 39854 777983
rect 39688 777902 39854 777912
rect 677642 746064 677799 746073
rect 677642 746003 677649 746064
rect 677533 745823 677649 746003
rect 677642 745760 677649 745823
rect 677793 745760 677799 746064
rect 677642 745752 677799 745760
rect 679528 746068 680309 746080
rect 679528 745764 679567 746068
rect 680271 745764 680309 746068
rect 679528 745752 680309 745764
rect 677533 745471 677792 745503
rect 677533 745462 677799 745471
rect 677533 745323 677648 745462
rect 677642 745158 677648 745323
rect 677792 745158 677799 745462
rect 677642 745150 677799 745158
rect 686081 745463 686838 745494
rect 686081 745159 686108 745463
rect 686812 745159 686838 745463
rect 686081 745129 686838 745159
rect 30819 735827 31576 735857
rect 30819 735523 30845 735827
rect 31549 735523 31576 735827
rect 30819 735492 31576 735523
rect 39699 735808 39862 735816
rect 39699 735504 39705 735808
rect 39849 735663 39862 735808
rect 39849 735504 40124 735663
rect 39699 735495 40124 735504
rect 39705 735483 40124 735495
rect 37348 735222 38129 735234
rect 37348 734918 37386 735222
rect 38090 734918 38129 735222
rect 37348 734906 38129 734918
rect 39695 735216 39858 735227
rect 39695 734912 39704 735216
rect 39848 735163 39858 735216
rect 39848 734983 40124 735163
rect 39848 734912 39858 734983
rect 39695 734906 39858 734912
rect 677643 701064 677803 701071
rect 677643 701003 677649 701064
rect 677533 700823 677649 701003
rect 677643 700760 677649 700823
rect 677793 700760 677803 701064
rect 677643 700754 677803 700760
rect 679528 701068 680309 701080
rect 679528 700764 679567 701068
rect 680271 700764 680309 701068
rect 679528 700752 680309 700764
rect 677533 700469 677792 700503
rect 677533 700462 677801 700469
rect 677533 700323 677648 700462
rect 677641 700158 677648 700323
rect 677792 700158 677801 700462
rect 677641 700152 677801 700158
rect 686081 700463 686838 700494
rect 686081 700159 686108 700463
rect 686812 700159 686838 700463
rect 686081 700129 686838 700159
rect 30819 692827 31576 692857
rect 30819 692523 30845 692827
rect 31549 692523 31576 692827
rect 30819 692492 31576 692523
rect 39699 692808 39859 692829
rect 39699 692504 39705 692808
rect 39849 692663 39859 692808
rect 39849 692504 40124 692663
rect 39699 692496 40124 692504
rect 39705 692483 40124 692496
rect 37348 692222 38129 692234
rect 37348 691918 37386 692222
rect 38090 691918 38129 692222
rect 37348 691906 38129 691918
rect 39695 692216 39855 692234
rect 39695 691912 39704 692216
rect 39848 692163 39855 692216
rect 39848 691983 40124 692163
rect 39848 691912 39855 691983
rect 39695 691901 39855 691912
rect 677644 656064 677802 656073
rect 677644 656003 677649 656064
rect 677533 655823 677649 656003
rect 677644 655760 677649 655823
rect 677793 655760 677802 656064
rect 677644 655753 677802 655760
rect 679528 656068 680309 656080
rect 679528 655764 679567 656068
rect 680271 655764 680309 656068
rect 679528 655752 680309 655764
rect 677533 655469 677792 655503
rect 677533 655462 677799 655469
rect 677533 655323 677648 655462
rect 677641 655158 677648 655323
rect 677792 655158 677799 655462
rect 677641 655149 677799 655158
rect 686081 655463 686838 655494
rect 686081 655159 686108 655463
rect 686812 655159 686838 655463
rect 686081 655129 686838 655159
rect 30819 649827 31576 649857
rect 30819 649523 30845 649827
rect 31549 649523 31576 649827
rect 30819 649492 31576 649523
rect 39697 649808 39859 649817
rect 39697 649504 39705 649808
rect 39849 649663 39859 649808
rect 39849 649504 40124 649663
rect 39697 649493 40124 649504
rect 39705 649483 40124 649493
rect 37348 649222 38129 649234
rect 37348 648918 37386 649222
rect 38090 648918 38129 649222
rect 37348 648906 38129 648918
rect 39694 649216 39856 649225
rect 39694 648912 39704 649216
rect 39848 649163 39856 649216
rect 39848 648983 40124 649163
rect 39848 648912 39856 648983
rect 39694 648901 39856 648912
rect 677643 611064 677805 611072
rect 677643 611003 677649 611064
rect 677533 610823 677649 611003
rect 677643 610760 677649 610823
rect 677793 610760 677805 611064
rect 677643 610752 677805 610760
rect 679528 611068 680309 611080
rect 679528 610764 679567 611068
rect 680271 610764 680309 611068
rect 679528 610752 680309 610764
rect 677533 610470 677792 610503
rect 677533 610462 677801 610470
rect 677533 610323 677648 610462
rect 677639 610158 677648 610323
rect 677792 610158 677801 610462
rect 677639 610150 677801 610158
rect 686081 610463 686838 610494
rect 686081 610159 686108 610463
rect 686812 610159 686838 610463
rect 686081 610129 686838 610159
rect 30819 606827 31576 606857
rect 30819 606523 30845 606827
rect 31549 606523 31576 606827
rect 30819 606492 31576 606523
rect 39697 606808 39858 606818
rect 39697 606504 39705 606808
rect 39849 606663 39858 606808
rect 39849 606504 40124 606663
rect 39697 606496 40124 606504
rect 39705 606483 40124 606496
rect 37348 606222 38129 606234
rect 37348 605918 37386 606222
rect 38090 605918 38129 606222
rect 37348 605906 38129 605918
rect 39695 606216 39856 606226
rect 39695 605912 39704 606216
rect 39848 606163 39856 606216
rect 39848 605983 40124 606163
rect 39848 605912 39856 605983
rect 39695 605904 39856 605912
rect 677645 566064 677799 566076
rect 677645 566003 677649 566064
rect 677533 565823 677649 566003
rect 677645 565760 677649 565823
rect 677793 565760 677799 566064
rect 677645 565756 677799 565760
rect 679528 566068 680309 566080
rect 679528 565764 679567 566068
rect 680271 565764 680309 566068
rect 679528 565752 680309 565764
rect 677533 565467 677792 565503
rect 677533 565462 677797 565467
rect 677533 565323 677648 565462
rect 677643 565158 677648 565323
rect 677792 565158 677797 565462
rect 677643 565147 677797 565158
rect 686081 565463 686838 565494
rect 686081 565159 686108 565463
rect 686812 565159 686838 565463
rect 686081 565129 686838 565159
rect 30819 563827 31576 563857
rect 30819 563523 30845 563827
rect 31549 563523 31576 563827
rect 30819 563492 31576 563523
rect 39696 563808 39856 563824
rect 39696 563504 39705 563808
rect 39849 563663 39856 563808
rect 39849 563504 40124 563663
rect 39696 563495 40124 563504
rect 39705 563483 40124 563495
rect 37348 563222 38129 563234
rect 37348 562918 37386 563222
rect 38090 562918 38129 563222
rect 37348 562906 38129 562918
rect 39692 563216 39852 563228
rect 39692 562912 39704 563216
rect 39848 563163 39852 563216
rect 39848 562983 40124 563163
rect 39848 562912 39852 562983
rect 39692 562899 39852 562912
rect 30819 520827 31576 520857
rect 30819 520523 30845 520827
rect 31549 520523 31576 520827
rect 30819 520492 31576 520523
rect 39697 520808 39860 520818
rect 39697 520504 39705 520808
rect 39849 520663 39860 520808
rect 39849 520504 40124 520663
rect 39697 520497 40124 520504
rect 39705 520483 40124 520497
rect 37348 520222 38129 520234
rect 37348 519918 37386 520222
rect 38090 519918 38129 520222
rect 37348 519906 38129 519918
rect 39695 520216 39858 520224
rect 39695 519912 39704 520216
rect 39848 520163 39858 520216
rect 39848 519983 40124 520163
rect 39848 519912 39858 519983
rect 39695 519903 39858 519912
rect 676906 474699 677706 474700
rect 676906 469901 676907 474699
rect 677705 469901 677706 474699
rect 676906 469900 677706 469901
rect 675786 469599 676586 469600
rect 675786 464949 675787 469599
rect 676585 464949 676586 469599
rect 675786 464948 676586 464949
rect 676906 464649 677706 464650
rect 676906 459861 676907 464649
rect 677705 459861 677706 464649
rect 676906 459860 677706 459861
rect 680587 459800 681277 459993
rect 688881 459800 688947 474800
rect 0 455645 4843 456094
rect 28653 440800 28719 455800
rect 32933 455546 33623 455800
rect 36323 455607 37013 455799
rect 38503 455546 39593 455800
rect 39918 455739 40718 455740
rect 39918 450953 39919 455739
rect 40717 450953 40718 455739
rect 39918 450952 40718 450953
rect 41038 450651 41838 450652
rect 41038 446001 41039 450651
rect 41837 446001 41838 450651
rect 41038 446000 41838 446001
rect 39918 445699 40718 445700
rect 39918 440901 39919 445699
rect 40717 440901 40718 445699
rect 39918 440900 40718 440901
rect 30819 391827 31576 391857
rect 30819 391523 30845 391827
rect 31549 391523 31576 391827
rect 30819 391492 31576 391523
rect 39697 391808 39858 391823
rect 39697 391504 39705 391808
rect 39849 391663 39858 391808
rect 39849 391504 40124 391663
rect 39697 391497 40124 391504
rect 39705 391483 40124 391497
rect 37348 391222 38129 391234
rect 37348 390918 37386 391222
rect 38090 390918 38129 391222
rect 37348 390906 38129 390918
rect 39694 391216 39855 391226
rect 39694 390912 39704 391216
rect 39848 391163 39855 391216
rect 39848 390983 40124 391163
rect 39848 390912 39855 390983
rect 39694 390900 39855 390912
rect 677643 389064 677798 389078
rect 677643 389003 677649 389064
rect 677533 388823 677649 389003
rect 677643 388760 677649 388823
rect 677793 388760 677798 389064
rect 677643 388755 677798 388760
rect 679528 389068 680309 389080
rect 679528 388764 679567 389068
rect 680271 388764 680309 389068
rect 679528 388752 680309 388764
rect 677533 388470 677792 388503
rect 677533 388462 677796 388470
rect 677533 388323 677648 388462
rect 677641 388158 677648 388323
rect 677792 388158 677796 388462
rect 677641 388147 677796 388158
rect 686081 388463 686838 388494
rect 686081 388159 686108 388463
rect 686812 388159 686838 388463
rect 686081 388129 686838 388159
rect 30819 348827 31576 348857
rect 30819 348523 30845 348827
rect 31549 348523 31576 348827
rect 30819 348492 31576 348523
rect 39692 348808 39854 348820
rect 39692 348504 39705 348808
rect 39849 348663 39854 348808
rect 39849 348504 40124 348663
rect 39692 348495 40124 348504
rect 39705 348483 40124 348495
rect 37348 348222 38129 348234
rect 37348 347918 37386 348222
rect 38090 347918 38129 348222
rect 37348 347906 38129 347918
rect 39695 348216 39857 348228
rect 39695 347912 39704 348216
rect 39848 348163 39857 348216
rect 39848 347983 40124 348163
rect 39848 347912 39857 347983
rect 39695 347903 39857 347912
rect 677643 344064 677802 344076
rect 677643 344003 677649 344064
rect 677533 343823 677649 344003
rect 677643 343760 677649 343823
rect 677793 343760 677802 344064
rect 677643 343754 677802 343760
rect 679528 344068 680309 344080
rect 679528 343764 679567 344068
rect 680271 343764 680309 344068
rect 679528 343752 680309 343764
rect 677533 343471 677792 343503
rect 677533 343462 677800 343471
rect 677533 343323 677648 343462
rect 677641 343158 677648 343323
rect 677792 343158 677800 343462
rect 677641 343149 677800 343158
rect 686081 343463 686838 343494
rect 686081 343159 686108 343463
rect 686812 343159 686838 343463
rect 686081 343129 686838 343159
rect 30819 305827 31576 305857
rect 30819 305523 30845 305827
rect 31549 305523 31576 305827
rect 30819 305492 31576 305523
rect 39695 305808 39860 305822
rect 39695 305504 39705 305808
rect 39849 305663 39860 305808
rect 39849 305504 40124 305663
rect 39695 305496 40124 305504
rect 39705 305483 40124 305496
rect 37348 305222 38129 305234
rect 37348 304918 37386 305222
rect 38090 304918 38129 305222
rect 37348 304906 38129 304918
rect 39691 305216 39856 305229
rect 39691 304912 39704 305216
rect 39848 305163 39856 305216
rect 39848 304983 40124 305163
rect 39848 304912 39856 304983
rect 39691 304903 39856 304912
rect 677641 299064 677803 299072
rect 677641 299003 677649 299064
rect 677533 298823 677649 299003
rect 677641 298760 677649 298823
rect 677793 298760 677803 299064
rect 677641 298752 677803 298760
rect 679528 299068 680309 299080
rect 679528 298764 679567 299068
rect 680271 298764 680309 299068
rect 679528 298752 680309 298764
rect 677533 298472 677792 298503
rect 677533 298462 677801 298472
rect 677533 298323 677648 298462
rect 677639 298158 677648 298323
rect 677792 298158 677801 298462
rect 677639 298152 677801 298158
rect 686081 298463 686838 298494
rect 686081 298159 686108 298463
rect 686812 298159 686838 298463
rect 686081 298129 686838 298159
rect 30819 262827 31576 262857
rect 30819 262523 30845 262827
rect 31549 262523 31576 262827
rect 30819 262492 31576 262523
rect 39695 262808 39854 262816
rect 39695 262504 39705 262808
rect 39849 262663 39854 262808
rect 39849 262504 40124 262663
rect 39695 262498 40124 262504
rect 39705 262483 40124 262498
rect 37348 262222 38129 262234
rect 37348 261918 37386 262222
rect 38090 261918 38129 262222
rect 37348 261906 38129 261918
rect 39697 262216 39856 262225
rect 39697 261912 39704 262216
rect 39848 262163 39856 262216
rect 39848 261983 40124 262163
rect 39848 261912 39856 261983
rect 39697 261907 39856 261912
rect 677643 254064 677800 254075
rect 677643 254003 677649 254064
rect 677533 253823 677649 254003
rect 677643 253760 677649 253823
rect 677793 253760 677800 254064
rect 677643 253755 677800 253760
rect 679528 254068 680309 254080
rect 679528 253764 679567 254068
rect 680271 253764 680309 254068
rect 679528 253752 680309 253764
rect 677533 253468 677792 253503
rect 677533 253462 677799 253468
rect 677533 253323 677648 253462
rect 677642 253158 677648 253323
rect 677792 253158 677799 253462
rect 677642 253148 677799 253158
rect 686081 253463 686838 253494
rect 686081 253159 686108 253463
rect 686812 253159 686838 253463
rect 686081 253129 686838 253159
rect 30819 219827 31576 219857
rect 30819 219523 30845 219827
rect 31549 219523 31576 219827
rect 30819 219492 31576 219523
rect 39698 219808 39854 219820
rect 39698 219504 39705 219808
rect 39849 219663 39854 219808
rect 39849 219504 40124 219663
rect 39698 219498 40124 219504
rect 39705 219483 40124 219498
rect 37348 219222 38129 219234
rect 37348 218918 37386 219222
rect 38090 218918 38129 219222
rect 37348 218906 38129 218918
rect 39697 219216 39853 219226
rect 39697 218912 39704 219216
rect 39848 219163 39853 219216
rect 39848 218983 40124 219163
rect 39848 218912 39853 218983
rect 39697 218904 39853 218912
rect 677641 209064 677796 209073
rect 677641 209003 677649 209064
rect 677533 208823 677649 209003
rect 677641 208760 677649 208823
rect 677793 208760 677796 209064
rect 677641 208755 677796 208760
rect 679528 209068 680309 209080
rect 679528 208764 679567 209068
rect 680271 208764 680309 209068
rect 679528 208752 680309 208764
rect 677533 208470 677792 208503
rect 677533 208462 677796 208470
rect 677533 208323 677648 208462
rect 677641 208158 677648 208323
rect 677792 208158 677796 208462
rect 677641 208152 677796 208158
rect 686081 208463 686838 208494
rect 686081 208159 686108 208463
rect 686812 208159 686838 208463
rect 686081 208129 686838 208159
rect 30819 176827 31576 176857
rect 30819 176523 30845 176827
rect 31549 176523 31576 176827
rect 30819 176492 31576 176523
rect 39697 176808 39853 176817
rect 39697 176504 39705 176808
rect 39849 176663 39853 176808
rect 39849 176504 40124 176663
rect 39697 176483 40124 176504
rect 39697 176480 39853 176483
rect 37348 176222 38129 176234
rect 37348 175918 37386 176222
rect 38090 175918 38129 176222
rect 37348 175906 38129 175918
rect 39698 176216 39853 176224
rect 39698 175912 39704 176216
rect 39848 176163 39853 176216
rect 39848 175983 40124 176163
rect 39848 175912 39853 175983
rect 39698 175901 39853 175912
rect 677643 164064 677799 164072
rect 677643 164003 677649 164064
rect 677533 163823 677649 164003
rect 677643 163760 677649 163823
rect 677793 163760 677799 164064
rect 677643 163752 677799 163760
rect 679528 164068 680309 164080
rect 679528 163764 679567 164068
rect 680271 163764 680309 164068
rect 679528 163752 680309 163764
rect 677533 163470 677792 163503
rect 677533 163462 677798 163470
rect 677533 163323 677648 163462
rect 677642 163158 677648 163323
rect 677792 163158 677798 163462
rect 677642 163150 677798 163158
rect 686081 163463 686838 163494
rect 686081 163159 686108 163463
rect 686812 163159 686838 163463
rect 686081 163129 686838 163159
rect 677644 119064 677803 119073
rect 677644 119003 677649 119064
rect 677533 118823 677649 119003
rect 677644 118760 677649 118823
rect 677793 118760 677803 119064
rect 677644 118753 677803 118760
rect 679528 119068 680309 119080
rect 679528 118764 679567 119068
rect 680271 118764 680309 119068
rect 679528 118752 680309 118764
rect 677533 118474 677792 118503
rect 677533 118462 677801 118474
rect 677533 118323 677648 118462
rect 677642 118158 677648 118323
rect 677792 118158 677801 118462
rect 677642 118154 677801 118158
rect 686081 118463 686838 118494
rect 686081 118159 686108 118463
rect 686812 118159 686838 118463
rect 686081 118129 686838 118159
rect 4570 107636 18733 108632
rect 18333 107186 18733 107636
rect 19043 107655 21342 108633
rect 19043 107186 19361 107655
rect 30773 101323 31662 101349
rect 30773 99489 30809 101323
rect 31637 99489 31662 101323
rect 30773 99457 31662 99489
rect 19040 94481 19369 96114
rect 19040 92770 19050 94481
rect 19352 92770 19369 94481
rect 19040 92731 19369 92770
rect 37315 94456 38198 94497
rect 37315 92802 37362 94456
rect 38160 92802 38198 94456
rect 37315 92755 38198 92802
rect 149134 39886 149314 40149
rect 149634 39886 149814 40149
rect 148962 39873 149314 39886
rect 148962 39729 148969 39873
rect 149273 39729 149314 39873
rect 149564 39872 149883 39886
rect 203934 39881 204114 40148
rect 204434 39885 204614 40148
rect 148962 39718 149281 39729
rect 149564 39728 149571 39872
rect 149875 39728 149883 39872
rect 149564 39718 149883 39728
rect 203765 39873 204114 39881
rect 203765 39729 203769 39873
rect 204073 39729 204114 39873
rect 204363 39872 204676 39885
rect 313534 39883 313714 40148
rect 203765 39717 204078 39729
rect 204363 39728 204371 39872
rect 204675 39728 204676 39872
rect 204363 39721 204676 39728
rect 313358 39873 313714 39883
rect 314034 39879 314214 40148
rect 368334 39879 368514 40148
rect 313358 39729 313369 39873
rect 313673 39729 313714 39873
rect 313961 39872 314283 39879
rect 313358 39723 313680 39729
rect 313961 39728 313971 39872
rect 314275 39728 314283 39872
rect 313961 39719 314283 39728
rect 368161 39873 368514 39879
rect 368834 39878 369014 40148
rect 423134 39880 423314 40148
rect 368161 39729 368169 39873
rect 368473 39729 368514 39873
rect 368763 39872 369084 39878
rect 368161 39721 368482 39729
rect 368763 39728 368771 39872
rect 369075 39728 369084 39872
rect 368763 39720 369084 39728
rect 422962 39873 423314 39880
rect 423634 39878 423814 40148
rect 477934 39884 478114 40148
rect 478434 39884 478614 40148
rect 422962 39729 422969 39873
rect 423273 39729 423314 39873
rect 423566 39872 423885 39878
rect 422962 39723 423281 39729
rect 423566 39728 423571 39872
rect 423875 39728 423885 39872
rect 423566 39721 423885 39728
rect 477762 39873 478114 39884
rect 477762 39729 477769 39873
rect 478073 39729 478114 39873
rect 478364 39872 478682 39884
rect 532734 39881 532914 40148
rect 533234 39882 533414 40148
rect 477762 39721 478080 39729
rect 478364 39728 478371 39872
rect 478675 39728 478682 39872
rect 478364 39721 478682 39728
rect 532563 39873 532914 39881
rect 532563 39729 532569 39873
rect 532873 39729 532914 39873
rect 533164 39872 533482 39882
rect 532563 39722 532881 39729
rect 533164 39728 533171 39872
rect 533475 39728 533482 39872
rect 533164 39723 533482 39728
rect 153640 38176 154074 38190
rect 149563 38114 149891 38153
rect 149563 37410 149575 38114
rect 149879 37410 149891 38114
rect 149563 37372 149891 37410
rect 153640 37340 153655 38176
rect 154064 37340 154074 38176
rect 204363 38114 204691 38153
rect 204363 37410 204375 38114
rect 204679 37410 204691 38114
rect 204363 37372 204691 37410
rect 313963 38114 314291 38153
rect 313963 37410 313975 38114
rect 314279 37410 314291 38114
rect 313963 37372 314291 37410
rect 368763 38114 369091 38153
rect 368763 37410 368775 38114
rect 369079 37410 369091 38114
rect 368763 37372 369091 37410
rect 423563 38114 423891 38153
rect 423563 37410 423575 38114
rect 423879 37410 423891 38114
rect 423563 37372 423891 37410
rect 478363 38114 478691 38153
rect 478363 37410 478375 38114
rect 478679 37410 478691 38114
rect 478363 37372 478691 37410
rect 533163 38114 533491 38153
rect 533163 37410 533175 38114
rect 533479 37410 533491 38114
rect 533163 37372 533491 37410
rect 640508 38118 641494 38170
rect 640508 37380 640578 38118
rect 641436 37380 641494 38118
rect 153640 37327 154074 37340
rect 640508 37328 641494 37380
rect 154241 35989 154677 36003
rect 154241 35178 154268 35989
rect 154659 35178 154677 35989
rect 154241 35148 154677 35178
rect 153032 34784 153474 34802
rect 153032 33947 153046 34784
rect 153462 33947 153474 34784
rect 153032 33933 153474 33947
rect 642100 32580 643096 32626
rect 642100 32020 642152 32580
rect 643060 32020 643096 32580
rect 642100 31988 643096 32020
rect 152438 31631 152880 31651
rect 148940 31573 149305 31600
rect 148940 30869 148970 31573
rect 149274 30869 149305 31573
rect 148940 30843 149305 30869
rect 152438 30800 152457 31631
rect 152858 30800 152880 31631
rect 203740 31573 204105 31600
rect 203740 30869 203770 31573
rect 204074 30869 204105 31573
rect 203740 30843 204105 30869
rect 313340 31573 313705 31600
rect 313340 30869 313370 31573
rect 313674 30869 313705 31573
rect 313340 30843 313705 30869
rect 368140 31573 368505 31600
rect 368140 30869 368170 31573
rect 368474 30869 368505 31573
rect 368140 30843 368505 30869
rect 422940 31573 423305 31600
rect 422940 30869 422970 31573
rect 423274 30869 423305 31573
rect 422940 30843 423305 30869
rect 477740 31573 478105 31600
rect 477740 30869 477770 31573
rect 478074 30869 478105 31573
rect 477740 30843 478105 30869
rect 532540 31573 532905 31600
rect 532540 30869 532570 31573
rect 532874 30869 532905 31573
rect 532540 30843 532905 30869
rect 152438 30782 152880 30800
rect 152424 20597 152890 20619
rect 152424 20133 152445 20597
rect 152866 20133 152890 20597
rect 152424 19693 152890 20133
rect 152424 19414 152450 19693
rect 152862 19414 152890 19693
rect 152424 19368 152890 19414
rect 153024 20597 153490 20619
rect 153024 20133 153045 20597
rect 153466 20133 153490 20597
rect 153024 18987 153490 20133
rect 153024 18710 153051 18987
rect 153463 18710 153490 18987
rect 153024 18659 153490 18710
rect 153624 20597 154090 20619
rect 153624 20133 153642 20597
rect 154063 20133 154090 20597
rect 153624 18294 154090 20133
rect 153624 18015 153652 18294
rect 154064 18015 154090 18294
rect 153624 17958 154090 18015
rect 154224 20600 154690 20619
rect 154224 20136 154248 20600
rect 154669 20136 154690 20600
rect 154224 17594 154690 20136
rect 154224 17316 154253 17594
rect 154665 17316 154690 17594
rect 154224 17251 154690 17316
rect 640486 16570 641502 16616
rect 640486 15710 640542 16570
rect 641444 15710 641502 16570
rect 640486 14496 641502 15710
rect 640486 14230 640518 14496
rect 641476 14230 641502 14496
rect 640486 12868 641502 14230
rect 640486 12608 640508 12868
rect 641466 12608 641502 12868
rect 640486 11238 641502 12608
rect 640486 10966 640520 11238
rect 641478 10966 641502 11238
rect 640486 10844 641502 10966
rect 642090 16566 643106 16622
rect 642090 15706 642146 16566
rect 643048 15706 643106 16566
rect 642090 13676 643106 15706
rect 642090 13414 642124 13676
rect 643082 13414 643106 13676
rect 642090 12050 643106 13414
rect 642090 11782 642110 12050
rect 643068 11782 643106 12050
rect 642090 10844 643106 11782
<< via4 >>
rect 41063 922151 41813 926939
rect 39943 917191 40693 921851
rect 675811 917701 676561 922499
rect 41063 912101 41813 916899
rect 676931 912749 677681 917409
rect 675811 907661 676561 912449
rect 676931 469901 677681 474699
rect 675811 464949 676561 469599
rect 676931 459861 677681 464649
rect 39943 450953 40693 455739
rect 41063 446001 41813 450651
rect 39943 440901 40693 445699
rect 149433 19411 149685 19693
rect 152450 19414 152862 19693
rect 150241 18712 150493 18994
rect 153051 18710 153463 18987
rect 150733 18010 150985 18292
rect 153652 18015 154064 18294
rect 151541 17311 151793 17593
rect 154253 17316 154665 17594
rect 640518 14230 641476 14496
rect 640508 12608 641466 12868
rect 640520 10966 641478 11238
rect 642124 13414 643082 13676
rect 642110 11782 643068 12050
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181241 1018512 193760 1031002
rect 232641 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030788
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030788
rect 628240 1018512 640760 1031002
rect 348400 1007147 348466 1008947
rect 348400 1004968 348466 1005617
rect 348400 1000607 348527 1001257
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19619 924934
rect 39918 921851 40718 927310
rect 39918 917191 39943 921851
rect 40693 917191 40718 921851
rect 6811 871210 18975 883378
rect 6811 829010 18975 841178
rect 6598 786640 19088 799160
rect 6598 743440 19088 755960
rect 6598 700240 19088 712760
rect 6598 657040 19088 669560
rect 6598 613840 19088 626360
rect 6598 570641 19088 583160
rect 6598 527441 19088 539960
rect 6811 484410 18975 496578
rect 39918 455739 40718 917191
rect 6167 442854 19619 453734
rect 39918 450953 39943 455739
rect 40693 450953 40718 455739
rect 39918 445699 40718 450953
rect 39918 440901 39943 445699
rect 40693 440901 40718 445699
rect 39918 440658 40718 440901
rect 41038 926939 41838 927310
rect 41038 922151 41063 926939
rect 41813 922151 41838 926939
rect 41038 916899 41838 922151
rect 41038 912101 41063 916899
rect 41813 912101 41838 916899
rect 41038 450651 41838 912101
rect 675786 922499 676586 922776
rect 675786 917701 675811 922499
rect 676561 917701 676586 922499
rect 675786 912449 676586 917701
rect 675786 907661 675811 912449
rect 676561 907661 676586 912449
rect 675786 469599 676586 907661
rect 675786 464949 675811 469599
rect 676561 464949 676586 469599
rect 675786 459306 676586 464949
rect 676906 917409 677706 922776
rect 676906 912749 676931 917409
rect 677681 912749 677706 917409
rect 676906 474699 677706 912749
rect 697980 909666 711432 920546
rect 698512 863640 711002 876160
rect 698624 819822 710788 831990
rect 698512 774440 711002 786960
rect 698512 729440 711002 741960
rect 698512 684440 711002 696960
rect 698512 639240 711002 651760
rect 698512 594240 711002 606760
rect 698512 549040 711002 561560
rect 698624 505222 710788 517390
rect 676906 469901 676931 474699
rect 677681 469901 677706 474699
rect 676906 464649 677706 469901
rect 676906 459861 676931 464649
rect 677681 459861 677706 464649
rect 697980 461866 711432 472746
rect 676906 459306 677706 459861
rect 41038 446001 41063 450651
rect 41813 446001 41838 450651
rect 41038 440658 41838 446001
rect 698624 417022 710788 429190
rect 6598 399841 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203959
rect 698512 146440 711002 158959
rect 6811 111610 18975 123778
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 149388 19693 152916 19718
rect 149388 19411 149433 19693
rect 149685 19414 152450 19693
rect 152862 19414 152916 19693
rect 149685 19411 152916 19414
rect 149388 19386 152916 19411
rect 150180 18994 153515 19018
rect 80222 6811 92390 18975
rect 150180 18712 150241 18994
rect 150493 18987 153515 18994
rect 150493 18712 153051 18987
rect 150180 18710 153051 18712
rect 153463 18710 153515 18987
rect 150180 18686 153515 18710
rect 136713 7143 144149 18309
rect 150671 18294 154113 18318
rect 150671 18292 153652 18294
rect 150671 18010 150733 18292
rect 150985 18015 153652 18292
rect 154064 18015 154113 18294
rect 150985 18010 154113 18015
rect 150671 17986 154113 18010
rect 151506 17594 154712 17618
rect 151506 17593 154253 17594
rect 151506 17311 151541 17593
rect 151793 17316 154253 17593
rect 154665 17316 154712 17594
rect 151793 17311 154712 17316
rect 151506 17286 154712 17311
rect 187640 6598 200159 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
rect 640396 14496 644288 14526
rect 640396 14230 640518 14496
rect 641476 14230 644288 14496
rect 640396 14206 644288 14230
rect 640396 13676 644288 13710
rect 640396 13414 642124 13676
rect 643082 13414 644288 13676
rect 640396 13390 644288 13414
rect 640396 12868 644288 12894
rect 640396 12608 640508 12868
rect 641466 12608 644288 12868
rect 640396 12574 644288 12608
rect 640396 12050 644288 12078
rect 640396 11782 642110 12050
rect 643068 11782 644288 12050
rect 640396 11758 644288 11782
rect 640396 11238 644288 11262
rect 640396 10966 640520 11238
rect 641478 10966 644288 11238
rect 640396 10942 644288 10966
<< comment >>
rect 42097 995463 675503 995503
rect 42097 42137 42137 995463
rect 675463 42137 675503 995463
rect 42097 42097 675503 42137
use sky130_ef_io__gpiov2_pad_wrapped  area0_gpio_pad[0] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform -1 0 202400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area0_gpio_pad[1]
timestamp 1683647856
transform -1 0 311000 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area0_gpio_pad[2]
timestamp 1683647856
transform -1 0 365800 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area0_gpio_pad[3]
timestamp 1683647856
transform -1 0 420600 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area0_gpio_pad[4]
timestamp 1683647856
transform -1 0 475400 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area0_gpio_pad[5]
timestamp 1683647856
transform -1 0 530200 0 -1 42193
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[0]
timestamp 1683647856
transform 1 0 282000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[1]
timestamp 1683647856
transform 1 0 230400 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[2]
timestamp 1683647856
transform 1 0 179000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[3]
timestamp 1683647856
transform 1 0 127600 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[4]
timestamp 1683647856
transform 1 0 76200 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[5]
timestamp 1683647856
transform 0 -1 42193 1 0 954200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[6]
timestamp 1683647856
transform 0 -1 42193 1 0 784400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[7]
timestamp 1683647856
transform 0 -1 42193 1 0 741200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[8]
timestamp 1683647856
transform 0 -1 42193 1 0 698000
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[9]
timestamp 1683647856
transform 0 1 675407 -1 0 654000
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[10]
timestamp 1683647856
transform 0 1 675407 -1 0 699200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[11]
timestamp 1683647856
transform 0 1 675407 -1 0 744200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[12]
timestamp 1683647856
transform 0 1 675407 -1 0 789200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[13]
timestamp 1683647856
transform 0 1 675407 -1 0 878400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[14]
timestamp 1683647856
transform 0 1 675407 -1 0 967600
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[15]
timestamp 1683647856
transform 1 0 626000 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[16]
timestamp 1683647856
transform 1 0 524200 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[17]
timestamp 1683647856
transform 1 0 472800 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  area1_gpio_pad[18]
timestamp 1683647856
transform 1 0 383800 0 1 995407
box -143 0 16134 42193
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_1 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform -1 0 51400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_2
timestamp 1683647856
transform -1 0 55400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_3
timestamp 1683647856
transform -1 0 59400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_4
timestamp 1683647856
transform -1 0 63400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_5
timestamp 1683647856
transform -1 0 67400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_6
timestamp 1683647856
transform -1 0 71400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_7
timestamp 1683647856
transform -1 0 105200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_8
timestamp 1683647856
transform -1 0 109200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_9
timestamp 1683647856
transform -1 0 113200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_10
timestamp 1683647856
transform -1 0 117200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_11
timestamp 1683647856
transform -1 0 121200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_12
timestamp 1683647856
transform -1 0 125200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_13
timestamp 1683647856
transform -1 0 159000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_14
timestamp 1683647856
transform -1 0 163000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_15
timestamp 1683647856
transform -1 0 167000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_16
timestamp 1683647856
transform -1 0 171000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_17
timestamp 1683647856
transform -1 0 175000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_18
timestamp 1683647856
transform -1 0 179000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_19
timestamp 1683647856
transform -1 0 213800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_20
timestamp 1683647856
transform -1 0 217800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_21
timestamp 1683647856
transform -1 0 221800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_22
timestamp 1683647856
transform -1 0 225800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_23
timestamp 1683647856
transform -1 0 229800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_24
timestamp 1683647856
transform -1 0 233800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_25
timestamp 1683647856
transform -1 0 267600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_26
timestamp 1683647856
transform -1 0 271600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_27
timestamp 1683647856
transform -1 0 275600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_28
timestamp 1683647856
transform -1 0 279600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_29
timestamp 1683647856
transform -1 0 283600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_30
timestamp 1683647856
transform -1 0 287600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_31
timestamp 1683647856
transform -1 0 322400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_32
timestamp 1683647856
transform -1 0 326400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_33
timestamp 1683647856
transform -1 0 330400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_34
timestamp 1683647856
transform -1 0 334400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_35
timestamp 1683647856
transform -1 0 338400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_36
timestamp 1683647856
transform -1 0 342400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_37
timestamp 1683647856
transform -1 0 377200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_38
timestamp 1683647856
transform -1 0 381200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_39
timestamp 1683647856
transform -1 0 385200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_40
timestamp 1683647856
transform -1 0 389200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_41
timestamp 1683647856
transform -1 0 393200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_42
timestamp 1683647856
transform -1 0 397200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_43
timestamp 1683647856
transform -1 0 432000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_44
timestamp 1683647856
transform -1 0 436000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_45
timestamp 1683647856
transform -1 0 440000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_46
timestamp 1683647856
transform -1 0 444000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_47
timestamp 1683647856
transform -1 0 448000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_48
timestamp 1683647856
transform -1 0 452000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_49
timestamp 1683647856
transform -1 0 486800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_50
timestamp 1683647856
transform -1 0 490800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_51
timestamp 1683647856
transform -1 0 494800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_52
timestamp 1683647856
transform -1 0 498800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_53
timestamp 1683647856
transform -1 0 502800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_54
timestamp 1683647856
transform -1 0 506800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_55
timestamp 1683647856
transform -1 0 541600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_56
timestamp 1683647856
transform -1 0 545600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_57
timestamp 1683647856
transform -1 0 549600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_58
timestamp 1683647856
transform -1 0 553600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_59
timestamp 1683647856
transform -1 0 557600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_60
timestamp 1683647856
transform -1 0 561600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_61
timestamp 1683647856
transform -1 0 595400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_62
timestamp 1683647856
transform -1 0 599400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_63
timestamp 1683647856
transform -1 0 603400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_64
timestamp 1683647856
transform -1 0 607400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_65
timestamp 1683647856
transform -1 0 611400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_66
timestamp 1683647856
transform -1 0 615400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_67
timestamp 1683647856
transform -1 0 649200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_68
timestamp 1683647856
transform -1 0 653200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_69
timestamp 1683647856
transform -1 0 657200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_70
timestamp 1683647856
transform -1 0 661200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_71
timestamp 1683647856
transform -1 0 665200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um  bus_tie_72
timestamp 1683647856
transform -1 0 669200 0 -1 39593
box 0 0 4000 39593
use caravel_logo  caravel_logo_0
timestamp 1638586901
transform 1 0 215294 0 1 5119
box -2520 0 15000 15560
use caravel_motto  caravel_motto_0
timestamp 1637698310
transform 1 0 -108943 0 1 -4710
box 373080 14838 395618 19242
use chip_io_gpio_connects  chip_io_gpio_connects_0
timestamp 1686151263
transform 0 -1 742000 1 0 320000
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_1
timestamp 1686151263
transform 0 -1 640200 1 0 320000
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_2
timestamp 1686151263
transform 0 -1 588800 1 0 320000
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_3
timestamp 1686151263
transform 0 -1 499800 1 0 320000
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_4
timestamp 1686151263
transform 0 -1 398000 1 0 320000
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_5
timestamp 1686151263
transform 0 -1 346400 1 0 320000
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_6
timestamp 1686151263
transform 0 -1 295000 1 0 320000
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_7
timestamp 1686151263
transform 0 -1 243600 1 0 320000
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_8
timestamp 1686151263
transform 0 -1 192200 1 0 320000
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_35
timestamp 1686151263
transform 0 1 86400 -1 0 717600
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_39
timestamp 1686151263
transform 0 1 195000 -1 0 717600
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_40
timestamp 1686151263
transform 0 1 249800 -1 0 717600
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_41
timestamp 1686151263
transform 0 1 304600 -1 0 717600
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_42
timestamp 1686151263
transform 0 1 359400 -1 0 717600
box 675407 99896 676763 117658
use chip_io_gpio_connects  chip_io_gpio_connects_43
timestamp 1686151263
transform 0 1 414200 -1 0 717600
box 675407 99896 676763 117658
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_0
timestamp 1686151263
transform 1 0 0 0 1 0
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_1
timestamp 1686151263
transform 1 0 0 0 1 45200
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_2
timestamp 1686151263
transform 1 0 0 0 1 90200
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_3
timestamp 1686151263
transform 1 0 0 0 1 135400
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_4
timestamp 1686151263
transform 1 0 0 0 1 180400
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_5
timestamp 1686151263
transform 1 0 0 0 1 225400
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_6
timestamp 1686151263
transform 1 0 0 0 1 270600
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_7
timestamp 1686151263
transform 1 0 0 0 1 447800
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_8
timestamp 1686151263
transform 1 0 0 0 1 493000
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_9
timestamp 1686151263
transform 1 0 0 0 1 538000
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_10
timestamp 1686151263
transform 1 0 0 0 1 583200
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_11
timestamp 1686151263
transform 1 0 0 0 1 628200
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_12
timestamp 1686151263
transform 1 0 0 0 1 673200
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_13
timestamp 1686151263
transform 1 0 0 0 1 762400
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_14
timestamp 1686151263
transform 1 0 0 0 1 851600
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_15
timestamp 1686151263
transform -1 0 717600 0 -1 1070200
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_16
timestamp 1686151263
transform -1 0 717600 0 -1 900400
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_17
timestamp 1686151263
transform -1 0 717600 0 -1 857200
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_18
timestamp 1686151263
transform -1 0 717600 0 -1 814000
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_19
timestamp 1686151263
transform -1 0 717600 0 -1 770800
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_20
timestamp 1686151263
transform -1 0 717600 0 -1 727600
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_21
timestamp 1686151263
transform -1 0 717600 0 -1 684400
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_22
timestamp 1686151263
transform -1 0 717600 0 -1 641200
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_23
timestamp 1686151263
transform -1 0 717600 0 -1 513600
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_24
timestamp 1686151263
transform -1 0 717600 0 -1 470400
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_25
timestamp 1686151263
transform -1 0 717600 0 -1 427200
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_26
timestamp 1686151263
transform -1 0 717600 0 -1 384000
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_27
timestamp 1686151263
transform -1 0 717600 0 -1 340800
box 675406 99896 676777 117452
use chip_io_gpio_connects_horiz  chip_io_gpio_connects_horiz_28
timestamp 1686151263
transform -1 0 717600 0 -1 297600
box 675406 99896 676777 117452
use constant_block  constant_value_inst[0]
timestamp 1665254080
transform 0 -1 678029 -1 0 120205
box 0 496 2800 2224
use constant_block  constant_value_inst[1]
timestamp 1665254080
transform 0 -1 678029 -1 0 165205
box 0 496 2800 2224
use constant_block  constant_value_inst[2]
timestamp 1665254080
transform 0 -1 678029 -1 0 210205
box 0 496 2800 2224
use constant_block  constant_value_inst[3]
timestamp 1665254080
transform 0 -1 678029 -1 0 255205
box 0 496 2800 2224
use constant_block  constant_value_inst[4]
timestamp 1665254080
transform 0 -1 678029 -1 0 300205
box 0 496 2800 2224
use constant_block  constant_value_inst[5]
timestamp 1665254080
transform 0 -1 678029 -1 0 345205
box 0 496 2800 2224
use constant_block  constant_value_inst[6]
timestamp 1665254080
transform 0 -1 678029 -1 0 390205
box 0 496 2800 2224
use constant_block  constant_value_inst[7]
timestamp 1665254080
transform 0 -1 678029 -1 0 567205
box 0 496 2800 2224
use constant_block  constant_value_inst[8]
timestamp 1665254080
transform 0 -1 678029 -1 0 612205
box 0 496 2800 2224
use constant_block  constant_value_inst[9]
timestamp 1665254080
transform 0 -1 678029 -1 0 657205
box 0 496 2800 2224
use constant_block  constant_value_inst[10]
timestamp 1665254080
transform 0 -1 678029 -1 0 702205
box 0 496 2800 2224
use constant_block  constant_value_inst[11]
timestamp 1665254080
transform 0 -1 678029 -1 0 747205
box 0 496 2800 2224
use constant_block  constant_value_inst[12]
timestamp 1665254080
transform 0 -1 678029 -1 0 792205
box 0 496 2800 2224
use constant_block  constant_value_inst[13]
timestamp 1665254080
transform 0 -1 678029 -1 0 881205
box 0 496 2800 2224
use constant_block  constant_value_inst[14]
timestamp 1665254080
transform 0 -1 678029 -1 0 971205
box 0 496 2800 2224
use constant_block  constant_value_inst[15]
timestamp 1665254080
transform 1 0 618435 0 -1 998018
box 0 496 2800 2224
use constant_block  constant_value_inst[16]
timestamp 1665254080
transform 1 0 519035 0 -1 998018
box 0 496 2800 2224
use constant_block  constant_value_inst[17]
timestamp 1665254080
transform 1 0 467835 0 -1 998018
box 0 496 2800 2224
use constant_block  constant_value_inst[18]
timestamp 1665254080
transform 1 0 378835 0 -1 998018
box 0 496 2800 2224
use constant_block  constant_value_inst[19]
timestamp 1665254080
transform 1 0 274435 0 -1 998018
box 0 496 2800 2224
use constant_block  constant_value_inst[20]
timestamp 1665254080
transform 1 0 223235 0 -1 998018
box 0 496 2800 2224
use constant_block  constant_value_inst[21]
timestamp 1665254080
transform 1 0 172035 0 -1 998018
box 0 496 2800 2224
use constant_block  constant_value_inst[22]
timestamp 1665254080
transform 1 0 120835 0 -1 998018
box 0 496 2800 2224
use constant_block  constant_value_inst[23]
timestamp 1665254080
transform 1 0 69635 0 -1 998018
box 0 496 2800 2224
use constant_block  constant_value_inst[24]
timestamp 1665254080
transform 0 1 39578 1 0 946781
box 0 496 2800 2224
use constant_block  constant_value_inst[25]
timestamp 1665254080
transform 0 1 39578 1 0 776781
box 0 496 2800 2224
use constant_block  constant_value_inst[26]
timestamp 1665254080
transform 0 1 39578 1 0 733781
box 0 496 2800 2224
use constant_block  constant_value_inst[27]
timestamp 1665254080
transform 0 1 39578 1 0 690781
box 0 496 2800 2224
use constant_block  constant_value_inst[28]
timestamp 1665254080
transform 0 1 39578 1 0 647781
box 0 496 2800 2224
use constant_block  constant_value_inst[29]
timestamp 1665254080
transform 0 1 39578 1 0 604781
box 0 496 2800 2224
use constant_block  constant_value_inst[30]
timestamp 1665254080
transform 0 1 39578 1 0 561781
box 0 496 2800 2224
use constant_block  constant_value_inst[31]
timestamp 1665254080
transform 0 1 39578 1 0 518781
box 0 496 2800 2224
use constant_block  constant_value_inst[32]
timestamp 1665254080
transform 0 1 39578 1 0 389781
box 0 496 2800 2224
use constant_block  constant_value_inst[33]
timestamp 1665254080
transform 0 1 39578 1 0 346781
box 0 496 2800 2224
use constant_block  constant_value_inst[34]
timestamp 1665254080
transform 0 1 39578 1 0 303781
box 0 496 2800 2224
use constant_block  constant_value_inst[35]
timestamp 1665254080
transform 0 1 39578 1 0 260781
box 0 496 2800 2224
use constant_block  constant_value_inst[36]
timestamp 1665254080
transform 0 1 39578 1 0 217781
box 0 496 2800 2224
use constant_block  constant_value_inst[37]
timestamp 1665254080
transform 0 1 39578 1 0 174781
box 0 496 2800 2224
use constant_block  constant_value_inst[38]
timestamp 1665254080
transform -1 0 205816 0 1 39552
box 0 496 2800 2224
use constant_block  constant_value_inst[39]
timestamp 1665254080
transform -1 0 315416 0 1 39552
box 0 496 2800 2224
use constant_block  constant_value_inst[40]
timestamp 1665254080
transform -1 0 370216 0 1 39552
box 0 496 2800 2224
use constant_block  constant_value_inst[41]
timestamp 1665254080
transform -1 0 425016 0 1 39552
box 0 496 2800 2224
use constant_block  constant_value_inst[42]
timestamp 1665254080
transform -1 0 479816 0 1 39552
box 0 496 2800 2224
use constant_block  constant_value_inst[43]
timestamp 1665254080
transform -1 0 534616 0 1 39552
box 0 496 2800 2224
use constant_block  constant_value_xres_inst
timestamp 1665254080
transform -1 0 151016 0 1 39552
box 0 496 2800 2224
use copyright_block_of  copyright_block_of_0
timestamp 1680028979
transform 1 0 95817 0 1 16746
box -262 -10348 35048 2764
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform 1 0 348400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_1
timestamp 1683647856
transform 0 1 678007 -1 0 70000
box 0 0 1000 39593
use sky130_ef_io__disconnect_vdda_slice_5um  disconnect_vdda_2
timestamp 1683647856
transform 0 -1 39593 1 0 152400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_5 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform 1 0 40800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_6
timestamp 1683647856
transform 1 0 44800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_7
timestamp 1683647856
transform 1 0 48800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_8
timestamp 1683647856
transform 1 0 52800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_9
timestamp 1683647856
transform 1 0 56800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_10
timestamp 1683647856
transform 1 0 60800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_11
timestamp 1683647856
transform 1 0 64800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_12
timestamp 1683647856
transform 1 0 68800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_13 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform 1 0 72800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_14 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform 1 0 74800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_15 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform 1 0 75800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_16
timestamp 1683647856
transform 1 0 76000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_18
timestamp 1683647856
transform 1 0 92200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_19
timestamp 1683647856
transform 1 0 96200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_20
timestamp 1683647856
transform 1 0 100200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_21
timestamp 1683647856
transform 1 0 104200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_22
timestamp 1683647856
transform 1 0 108200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_23
timestamp 1683647856
transform 1 0 112200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_24
timestamp 1683647856
transform 1 0 116200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_25
timestamp 1683647856
transform 1 0 120200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_26
timestamp 1683647856
transform 1 0 124200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_27
timestamp 1683647856
transform 1 0 126200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_28
timestamp 1683647856
transform 1 0 127200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_29
timestamp 1683647856
transform 1 0 127400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_31
timestamp 1683647856
transform 1 0 143600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_32
timestamp 1683647856
transform 1 0 147600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_33
timestamp 1683647856
transform 1 0 151600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_34
timestamp 1683647856
transform 1 0 155600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_35
timestamp 1683647856
transform 1 0 159600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_36
timestamp 1683647856
transform 1 0 163600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_37
timestamp 1683647856
transform 1 0 167600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_38
timestamp 1683647856
transform 1 0 171600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_39
timestamp 1683647856
transform 1 0 175600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_40
timestamp 1683647856
transform 1 0 177600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_41
timestamp 1683647856
transform 1 0 178600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_42
timestamp 1683647856
transform 1 0 178800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_44
timestamp 1683647856
transform 1 0 195000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_45
timestamp 1683647856
transform 1 0 199000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_46
timestamp 1683647856
transform 1 0 203000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_47
timestamp 1683647856
transform 1 0 207000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_48
timestamp 1683647856
transform 1 0 211000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_49
timestamp 1683647856
transform 1 0 215000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_50
timestamp 1683647856
transform 1 0 219000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_51
timestamp 1683647856
transform 1 0 223000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_52
timestamp 1683647856
transform 1 0 227000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_53
timestamp 1683647856
transform 1 0 229000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_54
timestamp 1683647856
transform 1 0 230000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_55
timestamp 1683647856
transform 1 0 230200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_57
timestamp 1683647856
transform 1 0 246400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_58
timestamp 1683647856
transform 1 0 250400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_59
timestamp 1683647856
transform 1 0 254400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_60
timestamp 1683647856
transform 1 0 258400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_61
timestamp 1683647856
transform 1 0 262400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_62
timestamp 1683647856
transform 1 0 266400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_63
timestamp 1683647856
transform 1 0 270400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_64
timestamp 1683647856
transform 1 0 274400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_65
timestamp 1683647856
transform 1 0 278400 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_66
timestamp 1683647856
transform 1 0 280400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_67
timestamp 1683647856
transform 1 0 281400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_68
timestamp 1683647856
transform 1 0 281600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_69
timestamp 1683647856
transform 1 0 281800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_71
timestamp 1683647856
transform 1 0 298000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_72
timestamp 1683647856
transform 1 0 302000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_73
timestamp 1683647856
transform 1 0 306000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_74
timestamp 1683647856
transform 1 0 310000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_75
timestamp 1683647856
transform 1 0 314000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_76
timestamp 1683647856
transform 1 0 318000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_77
timestamp 1683647856
transform 1 0 322000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_78
timestamp 1683647856
transform 1 0 326000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_79
timestamp 1683647856
transform 1 0 330000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_80
timestamp 1683647856
transform 1 0 332000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_81
timestamp 1683647856
transform 1 0 333000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_82
timestamp 1683647856
transform 1 0 333200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_86
timestamp 1683647856
transform 1 0 350400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_87
timestamp 1683647856
transform 1 0 354400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_88
timestamp 1683647856
transform 1 0 358400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_89
timestamp 1683647856
transform 1 0 362400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_90
timestamp 1683647856
transform 1 0 366400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_91
timestamp 1683647856
transform 1 0 370400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_92
timestamp 1683647856
transform 1 0 374400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_93
timestamp 1683647856
transform 1 0 378400 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_94
timestamp 1683647856
transform 1 0 382400 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_95
timestamp 1683647856
transform 1 0 383400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_96
timestamp 1683647856
transform 1 0 383600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_98
timestamp 1683647856
transform 1 0 399800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_99
timestamp 1683647856
transform 1 0 403800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_100
timestamp 1683647856
transform 1 0 407800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_101
timestamp 1683647856
transform 1 0 411800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_102
timestamp 1683647856
transform 1 0 415800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_103
timestamp 1683647856
transform 1 0 419800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_104
timestamp 1683647856
transform 1 0 423800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_105
timestamp 1683647856
transform 1 0 427800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_106
timestamp 1683647856
transform 1 0 431800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_107
timestamp 1683647856
transform 1 0 435800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_108
timestamp 1683647856
transform 1 0 439800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_109
timestamp 1683647856
transform 1 0 443800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_110
timestamp 1683647856
transform 1 0 447800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_111
timestamp 1683647856
transform 1 0 451800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_112
timestamp 1683647856
transform 1 0 455800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_113
timestamp 1683647856
transform 1 0 459800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_114
timestamp 1683647856
transform 1 0 463800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_115
timestamp 1683647856
transform 1 0 467800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_116
timestamp 1683647856
transform 1 0 471800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_118
timestamp 1683647856
transform 1 0 488800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_119
timestamp 1683647856
transform 1 0 492800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_120
timestamp 1683647856
transform 1 0 496800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_121
timestamp 1683647856
transform 1 0 500800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_122
timestamp 1683647856
transform 1 0 504800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_123
timestamp 1683647856
transform 1 0 508800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_124
timestamp 1683647856
transform 1 0 512800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_125
timestamp 1683647856
transform 1 0 516800 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_126
timestamp 1683647856
transform 1 0 520800 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_127
timestamp 1683647856
transform 1 0 522800 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_128
timestamp 1683647856
transform 1 0 523800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_129
timestamp 1683647856
transform 1 0 524000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_131
timestamp 1683647856
transform 1 0 540200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_132
timestamp 1683647856
transform 1 0 544200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_133
timestamp 1683647856
transform 1 0 548200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_134
timestamp 1683647856
transform 1 0 552200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_135
timestamp 1683647856
transform 1 0 556200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_136
timestamp 1683647856
transform 1 0 560200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_137
timestamp 1683647856
transform 1 0 564200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_138
timestamp 1683647856
transform 1 0 568200 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_139
timestamp 1683647856
transform 1 0 572200 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_140
timestamp 1683647856
transform 1 0 574200 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_141
timestamp 1683647856
transform 1 0 575200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_142
timestamp 1683647856
transform 1 0 575400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_144
timestamp 1683647856
transform 1 0 590600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_145
timestamp 1683647856
transform 1 0 594600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_146
timestamp 1683647856
transform 1 0 598600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_147
timestamp 1683647856
transform 1 0 602600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_148
timestamp 1683647856
transform 1 0 606600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_149
timestamp 1683647856
transform 1 0 610600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_150
timestamp 1683647856
transform 1 0 614600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_151
timestamp 1683647856
transform 1 0 618600 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_152
timestamp 1683647856
transform 1 0 622600 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_153
timestamp 1683647856
transform 1 0 624600 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_154
timestamp 1683647856
transform 1 0 625600 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_155
timestamp 1683647856
transform 1 0 625800 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_157
timestamp 1683647856
transform 1 0 642000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_158
timestamp 1683647856
transform 1 0 646000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_159
timestamp 1683647856
transform 1 0 650000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_160
timestamp 1683647856
transform 1 0 654000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_161
timestamp 1683647856
transform 1 0 658000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_162
timestamp 1683647856
transform 1 0 662000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_163
timestamp 1683647856
transform 1 0 666000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_164
timestamp 1683647856
transform 1 0 670000 0 1 998007
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_165
timestamp 1683647856
transform 1 0 674000 0 1 998007
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_166
timestamp 1683647856
transform 1 0 676000 0 1 998007
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_167
timestamp 1683647856
transform 1 0 677000 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_168
timestamp 1683647856
transform 1 0 677200 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_169
timestamp 1683647856
transform 1 0 677400 0 1 998007
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_170
timestamp 1683647856
transform -1 0 44000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_171
timestamp 1683647856
transform -1 0 46000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_172
timestamp 1683647856
transform -1 0 47000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_173
timestamp 1683647856
transform -1 0 47200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_174
timestamp 1683647856
transform -1 0 47400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_181
timestamp 1683647856
transform -1 0 75400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_182
timestamp 1683647856
transform -1 0 77400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_183
timestamp 1683647856
transform -1 0 78400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_184
timestamp 1683647856
transform -1 0 78600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_185
timestamp 1683647856
transform -1 0 78800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_187
timestamp 1683647856
transform -1 0 97800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_188
timestamp 1683647856
transform -1 0 99800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_189
timestamp 1683647856
transform -1 0 100800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_190
timestamp 1683647856
transform -1 0 101000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_191
timestamp 1683647856
transform -1 0 101200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_198
timestamp 1683647856
transform -1 0 129200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_199
timestamp 1683647856
transform -1 0 131200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_200
timestamp 1683647856
transform -1 0 132200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_201
timestamp 1683647856
transform -1 0 132400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_202
timestamp 1683647856
transform -1 0 132600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_204
timestamp 1683647856
transform -1 0 151600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_205
timestamp 1683647856
transform -1 0 153600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_206
timestamp 1683647856
transform -1 0 154600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_207
timestamp 1683647856
transform -1 0 154800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_208
timestamp 1683647856
transform -1 0 155000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_215
timestamp 1683647856
transform -1 0 183000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_216
timestamp 1683647856
transform -1 0 185000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_217
timestamp 1683647856
transform -1 0 186000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_218
timestamp 1683647856
transform -1 0 186200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_219
timestamp 1683647856
transform -1 0 186400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_221
timestamp 1683647856
transform -1 0 206400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_222
timestamp 1683647856
transform -1 0 208400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_223
timestamp 1683647856
transform -1 0 209400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_224
timestamp 1683647856
transform -1 0 209600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_225
timestamp 1683647856
transform -1 0 209800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_232
timestamp 1683647856
transform -1 0 237800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_233
timestamp 1683647856
transform -1 0 239800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_234
timestamp 1683647856
transform -1 0 240800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_235
timestamp 1683647856
transform -1 0 241000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_236
timestamp 1683647856
transform -1 0 241200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_238
timestamp 1683647856
transform -1 0 260200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_239
timestamp 1683647856
transform -1 0 262200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_240
timestamp 1683647856
transform -1 0 263200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_241
timestamp 1683647856
transform -1 0 263400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_242
timestamp 1683647856
transform -1 0 263600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_249
timestamp 1683647856
transform -1 0 291600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_250
timestamp 1683647856
transform -1 0 293600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_251
timestamp 1683647856
transform -1 0 294600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_252
timestamp 1683647856
transform -1 0 294800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_253
timestamp 1683647856
transform -1 0 295000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_255
timestamp 1683647856
transform -1 0 315000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_256
timestamp 1683647856
transform -1 0 317000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_257
timestamp 1683647856
transform -1 0 318000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_258
timestamp 1683647856
transform -1 0 318200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_259
timestamp 1683647856
transform -1 0 318400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_266
timestamp 1683647856
transform -1 0 346400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_267
timestamp 1683647856
transform -1 0 348400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_268
timestamp 1683647856
transform -1 0 349400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_269
timestamp 1683647856
transform -1 0 349600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_270
timestamp 1683647856
transform -1 0 349800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_272
timestamp 1683647856
transform -1 0 369800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_273
timestamp 1683647856
transform -1 0 371800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_274
timestamp 1683647856
transform -1 0 372800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_275
timestamp 1683647856
transform -1 0 373000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_276
timestamp 1683647856
transform -1 0 373200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_283
timestamp 1683647856
transform -1 0 401200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_284
timestamp 1683647856
transform -1 0 403200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_285
timestamp 1683647856
transform -1 0 404200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_286
timestamp 1683647856
transform -1 0 404400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_287
timestamp 1683647856
transform -1 0 404600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_289
timestamp 1683647856
transform -1 0 424600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_290
timestamp 1683647856
transform -1 0 426600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_291
timestamp 1683647856
transform -1 0 427600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_292
timestamp 1683647856
transform -1 0 427800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_293
timestamp 1683647856
transform -1 0 428000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_300
timestamp 1683647856
transform -1 0 456000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_301
timestamp 1683647856
transform -1 0 458000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_302
timestamp 1683647856
transform -1 0 459000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_303
timestamp 1683647856
transform -1 0 459200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_304
timestamp 1683647856
transform -1 0 459400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_306
timestamp 1683647856
transform -1 0 479400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_307
timestamp 1683647856
transform -1 0 481400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_308
timestamp 1683647856
transform -1 0 482400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_309
timestamp 1683647856
transform -1 0 482600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_310
timestamp 1683647856
transform -1 0 482800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_317
timestamp 1683647856
transform -1 0 510800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_318
timestamp 1683647856
transform -1 0 512800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_319
timestamp 1683647856
transform -1 0 513800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_320
timestamp 1683647856
transform -1 0 514000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_321
timestamp 1683647856
transform -1 0 514200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_323
timestamp 1683647856
transform -1 0 534200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_324
timestamp 1683647856
transform -1 0 536200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_325
timestamp 1683647856
transform -1 0 537200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_326
timestamp 1683647856
transform -1 0 537400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_327
timestamp 1683647856
transform -1 0 537600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_334
timestamp 1683647856
transform -1 0 565600 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_335
timestamp 1683647856
transform -1 0 567600 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_336
timestamp 1683647856
transform -1 0 568600 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_337
timestamp 1683647856
transform -1 0 568800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_338
timestamp 1683647856
transform -1 0 569000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_340
timestamp 1683647856
transform -1 0 588000 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_341
timestamp 1683647856
transform -1 0 590000 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_342
timestamp 1683647856
transform -1 0 591000 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_343
timestamp 1683647856
transform -1 0 591200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_344
timestamp 1683647856
transform -1 0 591400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_351
timestamp 1683647856
transform -1 0 619400 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_352
timestamp 1683647856
transform -1 0 621400 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_353
timestamp 1683647856
transform -1 0 622400 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_354
timestamp 1683647856
transform -1 0 622600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_355
timestamp 1683647856
transform -1 0 622800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_357
timestamp 1683647856
transform -1 0 641800 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_358
timestamp 1683647856
transform -1 0 643800 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_359
timestamp 1683647856
transform -1 0 644800 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_360
timestamp 1683647856
transform -1 0 645000 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_361
timestamp 1683647856
transform -1 0 645200 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_368
timestamp 1683647856
transform -1 0 673200 0 -1 39593
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_369
timestamp 1683647856
transform -1 0 675200 0 -1 39593
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_370
timestamp 1683647856
transform -1 0 676200 0 -1 39593
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_371
timestamp 1683647856
transform -1 0 676400 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_372
timestamp 1683647856
transform -1 0 676600 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_373
timestamp 1683647856
transform -1 0 676800 0 -1 39593
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_374
timestamp 1683647856
transform 0 -1 39593 1 0 40800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_375
timestamp 1683647856
transform 0 -1 39593 1 0 44800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_376
timestamp 1683647856
transform 0 -1 39593 1 0 48800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_377
timestamp 1683647856
transform 0 -1 39593 1 0 52800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_378
timestamp 1683647856
transform 0 -1 39593 1 0 56800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_379
timestamp 1683647856
transform 0 -1 39593 1 0 60800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_380
timestamp 1683647856
transform 0 -1 39593 1 0 64800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_381
timestamp 1683647856
transform 0 -1 39593 1 0 66800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_382
timestamp 1683647856
transform 0 -1 39593 1 0 67800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_384
timestamp 1683647856
transform 0 -1 39593 1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_385
timestamp 1683647856
transform 0 -1 39593 1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_386
timestamp 1683647856
transform 0 -1 39593 1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_387
timestamp 1683647856
transform 0 -1 39593 1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_388
timestamp 1683647856
transform 0 -1 39593 1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_389
timestamp 1683647856
transform 0 -1 39593 1 0 103000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_390
timestamp 1683647856
transform 0 -1 39593 1 0 107000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_391
timestamp 1683647856
transform 0 -1 39593 1 0 109000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_392
timestamp 1683647856
transform 0 -1 39593 1 0 110000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_394
timestamp 1683647856
transform 0 -1 39593 1 0 125200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_395
timestamp 1683647856
transform 0 -1 39593 1 0 129200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_396
timestamp 1683647856
transform 0 -1 39593 1 0 133200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_397
timestamp 1683647856
transform 0 -1 39593 1 0 137200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_398
timestamp 1683647856
transform 0 -1 39593 1 0 141200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_399
timestamp 1683647856
transform 0 -1 39593 1 0 145200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_400
timestamp 1683647856
transform 0 -1 39593 1 0 149200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_401
timestamp 1683647856
transform 0 -1 39593 1 0 151200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_402
timestamp 1683647856
transform 0 -1 39593 1 0 152200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_405
timestamp 1683647856
transform 0 -1 39593 1 0 154400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_406
timestamp 1683647856
transform 0 -1 39593 1 0 158400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_407
timestamp 1683647856
transform 0 -1 39593 1 0 162400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_408
timestamp 1683647856
transform 0 -1 39593 1 0 166400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_409
timestamp 1683647856
transform 0 -1 39593 1 0 170400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_410
timestamp 1683647856
transform 0 -1 39593 1 0 174400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_411
timestamp 1683647856
transform 0 -1 39593 1 0 178400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_412
timestamp 1683647856
transform 0 -1 39593 1 0 180400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_413
timestamp 1683647856
transform 0 -1 39593 1 0 181400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_415
timestamp 1683647856
transform 0 -1 39593 1 0 197600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_416
timestamp 1683647856
transform 0 -1 39593 1 0 201600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_417
timestamp 1683647856
transform 0 -1 39593 1 0 205600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_418
timestamp 1683647856
transform 0 -1 39593 1 0 209600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_419
timestamp 1683647856
transform 0 -1 39593 1 0 213600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_420
timestamp 1683647856
transform 0 -1 39593 1 0 217600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_421
timestamp 1683647856
transform 0 -1 39593 1 0 221600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_422
timestamp 1683647856
transform 0 -1 39593 1 0 223600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_423
timestamp 1683647856
transform 0 -1 39593 1 0 224600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_425
timestamp 1683647856
transform 0 -1 39593 1 0 240800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_426
timestamp 1683647856
transform 0 -1 39593 1 0 244800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_427
timestamp 1683647856
transform 0 -1 39593 1 0 248800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_428
timestamp 1683647856
transform 0 -1 39593 1 0 252800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_429
timestamp 1683647856
transform 0 -1 39593 1 0 256800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_430
timestamp 1683647856
transform 0 -1 39593 1 0 260800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_431
timestamp 1683647856
transform 0 -1 39593 1 0 264800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_432
timestamp 1683647856
transform 0 -1 39593 1 0 266800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_433
timestamp 1683647856
transform 0 -1 39593 1 0 267800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_435
timestamp 1683647856
transform 0 -1 39593 1 0 284000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_436
timestamp 1683647856
transform 0 -1 39593 1 0 288000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_437
timestamp 1683647856
transform 0 -1 39593 1 0 292000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_438
timestamp 1683647856
transform 0 -1 39593 1 0 296000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_439
timestamp 1683647856
transform 0 -1 39593 1 0 300000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_440
timestamp 1683647856
transform 0 -1 39593 1 0 304000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_441
timestamp 1683647856
transform 0 -1 39593 1 0 308000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_442
timestamp 1683647856
transform 0 -1 39593 1 0 310000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_443
timestamp 1683647856
transform 0 -1 39593 1 0 311000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_445
timestamp 1683647856
transform 0 -1 39593 1 0 327200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_446
timestamp 1683647856
transform 0 -1 39593 1 0 331200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_447
timestamp 1683647856
transform 0 -1 39593 1 0 335200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_448
timestamp 1683647856
transform 0 -1 39593 1 0 339200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_449
timestamp 1683647856
transform 0 -1 39593 1 0 343200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_450
timestamp 1683647856
transform 0 -1 39593 1 0 347200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_451
timestamp 1683647856
transform 0 -1 39593 1 0 351200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_452
timestamp 1683647856
transform 0 -1 39593 1 0 353200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_453
timestamp 1683647856
transform 0 -1 39593 1 0 354200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_455
timestamp 1683647856
transform 0 -1 39593 1 0 370400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_456
timestamp 1683647856
transform 0 -1 39593 1 0 374400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_457
timestamp 1683647856
transform 0 -1 39593 1 0 378400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_458
timestamp 1683647856
transform 0 -1 39593 1 0 382400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_459
timestamp 1683647856
transform 0 -1 39593 1 0 386400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_460
timestamp 1683647856
transform 0 -1 39593 1 0 390400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_461
timestamp 1683647856
transform 0 -1 39593 1 0 394400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_462
timestamp 1683647856
transform 0 -1 39593 1 0 396400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_463
timestamp 1683647856
transform 0 -1 39593 1 0 397400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_465
timestamp 1683647856
transform 0 -1 39593 1 0 413600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_466
timestamp 1683647856
transform 0 -1 39593 1 0 417600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_467
timestamp 1683647856
transform 0 -1 39593 1 0 421600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_468
timestamp 1683647856
transform 0 -1 39593 1 0 425600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_469
timestamp 1683647856
transform 0 -1 39593 1 0 429600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_470
timestamp 1683647856
transform 0 -1 39593 1 0 433600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_471
timestamp 1683647856
transform 0 -1 39593 1 0 437600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_472
timestamp 1683647856
transform 0 -1 39593 1 0 439600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_473
timestamp 1683647856
transform 0 -1 39593 1 0 440600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_475
timestamp 1683647856
transform 0 -1 39593 1 0 455800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_476
timestamp 1683647856
transform 0 -1 39593 1 0 459800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_477
timestamp 1683647856
transform 0 -1 39593 1 0 463800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_478
timestamp 1683647856
transform 0 -1 39593 1 0 467800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_479
timestamp 1683647856
transform 0 -1 39593 1 0 471800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_480
timestamp 1683647856
transform 0 -1 39593 1 0 475800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_481
timestamp 1683647856
transform 0 -1 39593 1 0 479800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_482
timestamp 1683647856
transform 0 -1 39593 1 0 481800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_483
timestamp 1683647856
transform 0 -1 39593 1 0 482800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_485
timestamp 1683647856
transform 0 -1 39593 1 0 498000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_486
timestamp 1683647856
transform 0 -1 39593 1 0 502000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_487
timestamp 1683647856
transform 0 -1 39593 1 0 506000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_488
timestamp 1683647856
transform 0 -1 39593 1 0 510000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_489
timestamp 1683647856
transform 0 -1 39593 1 0 514000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_490
timestamp 1683647856
transform 0 -1 39593 1 0 518000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_491
timestamp 1683647856
transform 0 -1 39593 1 0 522000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_492
timestamp 1683647856
transform 0 -1 39593 1 0 524000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_493
timestamp 1683647856
transform 0 -1 39593 1 0 525000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_495
timestamp 1683647856
transform 0 -1 39593 1 0 541200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_496
timestamp 1683647856
transform 0 -1 39593 1 0 545200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_497
timestamp 1683647856
transform 0 -1 39593 1 0 549200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_498
timestamp 1683647856
transform 0 -1 39593 1 0 553200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_499
timestamp 1683647856
transform 0 -1 39593 1 0 557200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_500
timestamp 1683647856
transform 0 -1 39593 1 0 561200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_501
timestamp 1683647856
transform 0 -1 39593 1 0 565200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_502
timestamp 1683647856
transform 0 -1 39593 1 0 567200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_503
timestamp 1683647856
transform 0 -1 39593 1 0 568200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_505
timestamp 1683647856
transform 0 -1 39593 1 0 584400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_506
timestamp 1683647856
transform 0 -1 39593 1 0 588400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_507
timestamp 1683647856
transform 0 -1 39593 1 0 592400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_508
timestamp 1683647856
transform 0 -1 39593 1 0 596400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_509
timestamp 1683647856
transform 0 -1 39593 1 0 600400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_510
timestamp 1683647856
transform 0 -1 39593 1 0 604400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_511
timestamp 1683647856
transform 0 -1 39593 1 0 608400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_512
timestamp 1683647856
transform 0 -1 39593 1 0 610400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_513
timestamp 1683647856
transform 0 -1 39593 1 0 611400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_515
timestamp 1683647856
transform 0 -1 39593 1 0 627600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_516
timestamp 1683647856
transform 0 -1 39593 1 0 631600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_517
timestamp 1683647856
transform 0 -1 39593 1 0 635600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_518
timestamp 1683647856
transform 0 -1 39593 1 0 639600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_519
timestamp 1683647856
transform 0 -1 39593 1 0 643600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_520
timestamp 1683647856
transform 0 -1 39593 1 0 647600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_521
timestamp 1683647856
transform 0 -1 39593 1 0 651600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_522
timestamp 1683647856
transform 0 -1 39593 1 0 653600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_523
timestamp 1683647856
transform 0 -1 39593 1 0 654600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_525
timestamp 1683647856
transform 0 -1 39593 1 0 670800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_526
timestamp 1683647856
transform 0 -1 39593 1 0 674800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_527
timestamp 1683647856
transform 0 -1 39593 1 0 678800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_528
timestamp 1683647856
transform 0 -1 39593 1 0 682800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_529
timestamp 1683647856
transform 0 -1 39593 1 0 686800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_530
timestamp 1683647856
transform 0 -1 39593 1 0 690800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_531
timestamp 1683647856
transform 0 -1 39593 1 0 694800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_532
timestamp 1683647856
transform 0 -1 39593 1 0 696800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_533
timestamp 1683647856
transform 0 -1 39593 1 0 697800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_535
timestamp 1683647856
transform 0 -1 39593 1 0 714000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_536
timestamp 1683647856
transform 0 -1 39593 1 0 718000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_537
timestamp 1683647856
transform 0 -1 39593 1 0 722000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_538
timestamp 1683647856
transform 0 -1 39593 1 0 726000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_539
timestamp 1683647856
transform 0 -1 39593 1 0 730000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_540
timestamp 1683647856
transform 0 -1 39593 1 0 734000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_541
timestamp 1683647856
transform 0 -1 39593 1 0 738000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_542
timestamp 1683647856
transform 0 -1 39593 1 0 740000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_543
timestamp 1683647856
transform 0 -1 39593 1 0 741000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_545
timestamp 1683647856
transform 0 -1 39593 1 0 757200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_546
timestamp 1683647856
transform 0 -1 39593 1 0 761200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_547
timestamp 1683647856
transform 0 -1 39593 1 0 765200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_548
timestamp 1683647856
transform 0 -1 39593 1 0 769200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_549
timestamp 1683647856
transform 0 -1 39593 1 0 773200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_550
timestamp 1683647856
transform 0 -1 39593 1 0 777200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_551
timestamp 1683647856
transform 0 -1 39593 1 0 781200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_552
timestamp 1683647856
transform 0 -1 39593 1 0 783200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_553
timestamp 1683647856
transform 0 -1 39593 1 0 784200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_555
timestamp 1683647856
transform 0 -1 39593 1 0 800400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_556
timestamp 1683647856
transform 0 -1 39593 1 0 804400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_557
timestamp 1683647856
transform 0 -1 39593 1 0 808400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_558
timestamp 1683647856
transform 0 -1 39593 1 0 812400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_559
timestamp 1683647856
transform 0 -1 39593 1 0 816400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_560
timestamp 1683647856
transform 0 -1 39593 1 0 820400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_561
timestamp 1683647856
transform 0 -1 39593 1 0 824400
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_562
timestamp 1683647856
transform 0 -1 39593 1 0 826400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_563
timestamp 1683647856
transform 0 -1 39593 1 0 827400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_565
timestamp 1683647856
transform 0 -1 39593 1 0 842600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_566
timestamp 1683647856
transform 0 -1 39593 1 0 846600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_567
timestamp 1683647856
transform 0 -1 39593 1 0 850600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_568
timestamp 1683647856
transform 0 -1 39593 1 0 854600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_569
timestamp 1683647856
transform 0 -1 39593 1 0 858600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_570
timestamp 1683647856
transform 0 -1 39593 1 0 862600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_571
timestamp 1683647856
transform 0 -1 39593 1 0 866600
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_572
timestamp 1683647856
transform 0 -1 39593 1 0 868600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_573
timestamp 1683647856
transform 0 -1 39593 1 0 869600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_575
timestamp 1683647856
transform 0 -1 39593 1 0 884800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_576
timestamp 1683647856
transform 0 -1 39593 1 0 888800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_577
timestamp 1683647856
transform 0 -1 39593 1 0 892800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_578
timestamp 1683647856
transform 0 -1 39593 1 0 896800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_579
timestamp 1683647856
transform 0 -1 39593 1 0 900800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_580
timestamp 1683647856
transform 0 -1 39593 1 0 904800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_581
timestamp 1683647856
transform 0 -1 39593 1 0 908800
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_582
timestamp 1683647856
transform 0 -1 39593 1 0 910800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_583
timestamp 1683647856
transform 0 -1 39593 1 0 911800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_585
timestamp 1683647856
transform 0 -1 39593 1 0 927000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_586
timestamp 1683647856
transform 0 -1 39593 1 0 931000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_587
timestamp 1683647856
transform 0 -1 39593 1 0 935000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_588
timestamp 1683647856
transform 0 -1 39593 1 0 939000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_589
timestamp 1683647856
transform 0 -1 39593 1 0 943000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_590
timestamp 1683647856
transform 0 -1 39593 1 0 947000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_591
timestamp 1683647856
transform 0 -1 39593 1 0 951000
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_592
timestamp 1683647856
transform 0 -1 39593 1 0 953000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_593
timestamp 1683647856
transform 0 -1 39593 1 0 954000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_595
timestamp 1683647856
transform 0 -1 39593 1 0 970200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_596
timestamp 1683647856
transform 0 -1 39593 1 0 974200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_597
timestamp 1683647856
transform 0 -1 39593 1 0 978200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_598
timestamp 1683647856
transform 0 -1 39593 1 0 982200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_599
timestamp 1683647856
transform 0 -1 39593 1 0 986200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_600
timestamp 1683647856
transform 0 -1 39593 1 0 990200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_10um  FILLER_601
timestamp 1683647856
transform 0 -1 39593 1 0 994200
box 0 0 2000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_602
timestamp 1683647856
transform 0 -1 39593 1 0 996200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_603
timestamp 1683647856
transform 0 -1 39593 1 0 997200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_604
timestamp 1683647856
transform 0 -1 39593 1 0 997400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_605
timestamp 1683647856
transform 0 1 678007 -1 0 44000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_606
timestamp 1683647856
transform 0 1 678007 -1 0 48000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_607
timestamp 1683647856
transform 0 1 678007 -1 0 52000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_608
timestamp 1683647856
transform 0 1 678007 -1 0 56000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_609
timestamp 1683647856
transform 0 1 678007 -1 0 60000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_610
timestamp 1683647856
transform 0 1 678007 -1 0 64000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_611
timestamp 1683647856
transform 0 1 678007 -1 0 68000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_612
timestamp 1683647856
transform 0 1 678007 -1 0 69000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_615
timestamp 1683647856
transform 0 1 678007 -1 0 75000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_616
timestamp 1683647856
transform 0 1 678007 -1 0 79000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_617
timestamp 1683647856
transform 0 1 678007 -1 0 83000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_618
timestamp 1683647856
transform 0 1 678007 -1 0 87000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_619
timestamp 1683647856
transform 0 1 678007 -1 0 91000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_620
timestamp 1683647856
transform 0 1 678007 -1 0 95000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_621
timestamp 1683647856
transform 0 1 678007 -1 0 99000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_622
timestamp 1683647856
transform 0 1 678007 -1 0 100000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_624
timestamp 1683647856
transform 0 1 678007 -1 0 120000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_625
timestamp 1683647856
transform 0 1 678007 -1 0 124000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_626
timestamp 1683647856
transform 0 1 678007 -1 0 128000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_627
timestamp 1683647856
transform 0 1 678007 -1 0 132000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_628
timestamp 1683647856
transform 0 1 678007 -1 0 136000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_629
timestamp 1683647856
transform 0 1 678007 -1 0 140000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_630
timestamp 1683647856
transform 0 1 678007 -1 0 144000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_631
timestamp 1683647856
transform 0 1 678007 -1 0 145000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_632
timestamp 1683647856
transform 0 1 678007 -1 0 145200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_634
timestamp 1683647856
transform 0 1 678007 -1 0 165200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_635
timestamp 1683647856
transform 0 1 678007 -1 0 169200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_636
timestamp 1683647856
transform 0 1 678007 -1 0 173200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_637
timestamp 1683647856
transform 0 1 678007 -1 0 177200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_638
timestamp 1683647856
transform 0 1 678007 -1 0 181200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_639
timestamp 1683647856
transform 0 1 678007 -1 0 185200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_640
timestamp 1683647856
transform 0 1 678007 -1 0 189200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_641
timestamp 1683647856
transform 0 1 678007 -1 0 190200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_643
timestamp 1683647856
transform 0 1 678007 -1 0 210200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_644
timestamp 1683647856
transform 0 1 678007 -1 0 214200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_645
timestamp 1683647856
transform 0 1 678007 -1 0 218200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_646
timestamp 1683647856
transform 0 1 678007 -1 0 222200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_647
timestamp 1683647856
transform 0 1 678007 -1 0 226200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_648
timestamp 1683647856
transform 0 1 678007 -1 0 230200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_649
timestamp 1683647856
transform 0 1 678007 -1 0 234200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_650
timestamp 1683647856
transform 0 1 678007 -1 0 235200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_651
timestamp 1683647856
transform 0 1 678007 -1 0 235400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_653
timestamp 1683647856
transform 0 1 678007 -1 0 255400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_654
timestamp 1683647856
transform 0 1 678007 -1 0 259400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_655
timestamp 1683647856
transform 0 1 678007 -1 0 263400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_656
timestamp 1683647856
transform 0 1 678007 -1 0 267400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_657
timestamp 1683647856
transform 0 1 678007 -1 0 271400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_658
timestamp 1683647856
transform 0 1 678007 -1 0 275400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_659
timestamp 1683647856
transform 0 1 678007 -1 0 279400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_660
timestamp 1683647856
transform 0 1 678007 -1 0 280400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_662
timestamp 1683647856
transform 0 1 678007 -1 0 300400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_663
timestamp 1683647856
transform 0 1 678007 -1 0 304400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_664
timestamp 1683647856
transform 0 1 678007 -1 0 308400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_665
timestamp 1683647856
transform 0 1 678007 -1 0 312400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_666
timestamp 1683647856
transform 0 1 678007 -1 0 316400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_667
timestamp 1683647856
transform 0 1 678007 -1 0 320400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_668
timestamp 1683647856
transform 0 1 678007 -1 0 324400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_669
timestamp 1683647856
transform 0 1 678007 -1 0 325400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_671
timestamp 1683647856
transform 0 1 678007 -1 0 345400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_672
timestamp 1683647856
transform 0 1 678007 -1 0 349400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_673
timestamp 1683647856
transform 0 1 678007 -1 0 353400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_674
timestamp 1683647856
transform 0 1 678007 -1 0 357400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_675
timestamp 1683647856
transform 0 1 678007 -1 0 361400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_676
timestamp 1683647856
transform 0 1 678007 -1 0 365400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_677
timestamp 1683647856
transform 0 1 678007 -1 0 369400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_678
timestamp 1683647856
transform 0 1 678007 -1 0 370400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_679
timestamp 1683647856
transform 0 1 678007 -1 0 370600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_681
timestamp 1683647856
transform 0 1 678007 -1 0 390600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_682
timestamp 1683647856
transform 0 1 678007 -1 0 394600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_683
timestamp 1683647856
transform 0 1 678007 -1 0 398600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_684
timestamp 1683647856
transform 0 1 678007 -1 0 402600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_685
timestamp 1683647856
transform 0 1 678007 -1 0 406600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_686
timestamp 1683647856
transform 0 1 678007 -1 0 410600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_687
timestamp 1683647856
transform 0 1 678007 -1 0 414600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_688
timestamp 1683647856
transform 0 1 678007 -1 0 415600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_690
timestamp 1683647856
transform 0 1 678007 -1 0 434600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_691
timestamp 1683647856
transform 0 1 678007 -1 0 438600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_692
timestamp 1683647856
transform 0 1 678007 -1 0 442600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_693
timestamp 1683647856
transform 0 1 678007 -1 0 446600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_694
timestamp 1683647856
transform 0 1 678007 -1 0 450600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_695
timestamp 1683647856
transform 0 1 678007 -1 0 454600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_696
timestamp 1683647856
transform 0 1 678007 -1 0 458600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_697
timestamp 1683647856
transform 0 1 678007 -1 0 459600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_698
timestamp 1683647856
transform 0 1 678007 -1 0 459800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_700
timestamp 1683647856
transform 0 1 678007 -1 0 478800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_701
timestamp 1683647856
transform 0 1 678007 -1 0 482800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_702
timestamp 1683647856
transform 0 1 678007 -1 0 486800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_703
timestamp 1683647856
transform 0 1 678007 -1 0 490800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_704
timestamp 1683647856
transform 0 1 678007 -1 0 494800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_705
timestamp 1683647856
transform 0 1 678007 -1 0 498800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_706
timestamp 1683647856
transform 0 1 678007 -1 0 502800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_707
timestamp 1683647856
transform 0 1 678007 -1 0 503800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_709
timestamp 1683647856
transform 0 1 678007 -1 0 522800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_710
timestamp 1683647856
transform 0 1 678007 -1 0 526800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_711
timestamp 1683647856
transform 0 1 678007 -1 0 530800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_712
timestamp 1683647856
transform 0 1 678007 -1 0 534800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_713
timestamp 1683647856
transform 0 1 678007 -1 0 538800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_714
timestamp 1683647856
transform 0 1 678007 -1 0 542800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_715
timestamp 1683647856
transform 0 1 678007 -1 0 546800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_716
timestamp 1683647856
transform 0 1 678007 -1 0 547800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_718
timestamp 1683647856
transform 0 1 678007 -1 0 567800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_719
timestamp 1683647856
transform 0 1 678007 -1 0 571800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_720
timestamp 1683647856
transform 0 1 678007 -1 0 575800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_721
timestamp 1683647856
transform 0 1 678007 -1 0 579800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_722
timestamp 1683647856
transform 0 1 678007 -1 0 583800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_723
timestamp 1683647856
transform 0 1 678007 -1 0 587800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_724
timestamp 1683647856
transform 0 1 678007 -1 0 591800
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_725
timestamp 1683647856
transform 0 1 678007 -1 0 592800
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_726
timestamp 1683647856
transform 0 1 678007 -1 0 593000
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_728
timestamp 1683647856
transform 0 1 678007 -1 0 613000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_729
timestamp 1683647856
transform 0 1 678007 -1 0 617000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_730
timestamp 1683647856
transform 0 1 678007 -1 0 621000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_731
timestamp 1683647856
transform 0 1 678007 -1 0 625000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_732
timestamp 1683647856
transform 0 1 678007 -1 0 629000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_733
timestamp 1683647856
transform 0 1 678007 -1 0 633000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_734
timestamp 1683647856
transform 0 1 678007 -1 0 637000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_735
timestamp 1683647856
transform 0 1 678007 -1 0 638000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_737
timestamp 1683647856
transform 0 1 678007 -1 0 658000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_738
timestamp 1683647856
transform 0 1 678007 -1 0 662000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_739
timestamp 1683647856
transform 0 1 678007 -1 0 666000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_740
timestamp 1683647856
transform 0 1 678007 -1 0 670000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_741
timestamp 1683647856
transform 0 1 678007 -1 0 674000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_742
timestamp 1683647856
transform 0 1 678007 -1 0 678000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_743
timestamp 1683647856
transform 0 1 678007 -1 0 682000
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_744
timestamp 1683647856
transform 0 1 678007 -1 0 683000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_745
timestamp 1683647856
transform 0 1 678007 -1 0 683200
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_747
timestamp 1683647856
transform 0 1 678007 -1 0 703200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_748
timestamp 1683647856
transform 0 1 678007 -1 0 707200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_749
timestamp 1683647856
transform 0 1 678007 -1 0 711200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_750
timestamp 1683647856
transform 0 1 678007 -1 0 715200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_751
timestamp 1683647856
transform 0 1 678007 -1 0 719200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_752
timestamp 1683647856
transform 0 1 678007 -1 0 723200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_753
timestamp 1683647856
transform 0 1 678007 -1 0 727200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_754
timestamp 1683647856
transform 0 1 678007 -1 0 728200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_756
timestamp 1683647856
transform 0 1 678007 -1 0 748200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_757
timestamp 1683647856
transform 0 1 678007 -1 0 752200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_758
timestamp 1683647856
transform 0 1 678007 -1 0 756200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_759
timestamp 1683647856
transform 0 1 678007 -1 0 760200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_760
timestamp 1683647856
transform 0 1 678007 -1 0 764200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_761
timestamp 1683647856
transform 0 1 678007 -1 0 768200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_762
timestamp 1683647856
transform 0 1 678007 -1 0 772200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_763
timestamp 1683647856
transform 0 1 678007 -1 0 773200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_765
timestamp 1683647856
transform 0 1 678007 -1 0 793200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_766
timestamp 1683647856
transform 0 1 678007 -1 0 797200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_767
timestamp 1683647856
transform 0 1 678007 -1 0 801200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_768
timestamp 1683647856
transform 0 1 678007 -1 0 805200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_769
timestamp 1683647856
transform 0 1 678007 -1 0 809200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_770
timestamp 1683647856
transform 0 1 678007 -1 0 813200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_771
timestamp 1683647856
transform 0 1 678007 -1 0 817200
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_772
timestamp 1683647856
transform 0 1 678007 -1 0 818200
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_773
timestamp 1683647856
transform 0 1 678007 -1 0 818400
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_775
timestamp 1683647856
transform 0 1 678007 -1 0 837400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_776
timestamp 1683647856
transform 0 1 678007 -1 0 841400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_777
timestamp 1683647856
transform 0 1 678007 -1 0 845400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_778
timestamp 1683647856
transform 0 1 678007 -1 0 849400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_779
timestamp 1683647856
transform 0 1 678007 -1 0 853400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_780
timestamp 1683647856
transform 0 1 678007 -1 0 857400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_781
timestamp 1683647856
transform 0 1 678007 -1 0 861400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_782
timestamp 1683647856
transform 0 1 678007 -1 0 862400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_784
timestamp 1683647856
transform 0 1 678007 -1 0 882400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_785
timestamp 1683647856
transform 0 1 678007 -1 0 886400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_786
timestamp 1683647856
transform 0 1 678007 -1 0 890400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_787
timestamp 1683647856
transform 0 1 678007 -1 0 894400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_788
timestamp 1683647856
transform 0 1 678007 -1 0 898400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_789
timestamp 1683647856
transform 0 1 678007 -1 0 902400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_790
timestamp 1683647856
transform 0 1 678007 -1 0 906400
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_791
timestamp 1683647856
transform 0 1 678007 -1 0 907400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_792
timestamp 1683647856
transform 0 1 678007 -1 0 907600
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_794
timestamp 1683647856
transform 0 1 678007 -1 0 926600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_795
timestamp 1683647856
transform 0 1 678007 -1 0 930600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_796
timestamp 1683647856
transform 0 1 678007 -1 0 934600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_797
timestamp 1683647856
transform 0 1 678007 -1 0 938600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_798
timestamp 1683647856
transform 0 1 678007 -1 0 942600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_799
timestamp 1683647856
transform 0 1 678007 -1 0 946600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_800
timestamp 1683647856
transform 0 1 678007 -1 0 950600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_801
timestamp 1683647856
transform 0 1 678007 -1 0 951600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_803
timestamp 1683647856
transform 0 1 678007 -1 0 971600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_804
timestamp 1683647856
transform 0 1 678007 -1 0 975600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_805
timestamp 1683647856
transform 0 1 678007 -1 0 979600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_806
timestamp 1683647856
transform 0 1 678007 -1 0 983600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_807
timestamp 1683647856
transform 0 1 678007 -1 0 987600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_808
timestamp 1683647856
transform 0 1 678007 -1 0 991600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_20um  FILLER_809
timestamp 1683647856
transform 0 1 678007 -1 0 995600
box 0 0 4000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_810
timestamp 1683647856
transform 0 1 678007 -1 0 996600
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_1um  FILLER_811
timestamp 1683647856
transform 0 1 678007 -1 0 996800
box 0 0 200 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB1
timestamp 1683647856
transform 0 1 678007 -1 0 71000
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB2
timestamp 1683647856
transform 0 -1 39593 1 0 153400
box 0 0 1000 39593
use sky130_ef_io__com_bus_slice_5um  FILLER_SB3
timestamp 1683647856
transform 1 0 349400 0 1 998007
box 0 0 1000 39593
use sky130_fd_io__top_xres4v2  master_resetb_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform -1 0 147600 0 -1 40000
box -103 0 15124 40000
use sky130_ef_io__vccd_lvc_clamped_pad  mgmt_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform 0 -1 39593 1 0 68000
box 0 -2107 17239 39593
use sky130_ef_io__vdda_hvc_clamped_pad  mgmt_vdda_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform -1 0 637800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform 0 -1 39593 1 0 110200
box 0 -407 15000 39593
use sky130_ef_io__vddio_hvc_clamped_pad  mgmt_vddio_hvclamp_pad\[1\]
timestamp 1683647856
transform 0 -1 39593 1 0 869800
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  mgmt_vssa_hvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform -1 0 93800 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped_pad  mgmt_vssd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform -1 0 256200 0 -1 39593
box 0 -2107 17239 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[0\] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform -1 0 584000 0 -1 39593
box 0 -407 15000 39593
use sky130_ef_io__vssio_hvc_clamped_pad  mgmt_vssio_hvclamp_pad\[1\]
timestamp 1683647856
transform 1 0 333400 0 1 998007
box 0 -407 15000 39593
use open_source  open_source_0
timestamp 1666123577
transform 1 0 155011 0 1 2193
box 752 5164 29030 16242
use simple_por  por
timestamp 1680223961
transform 0 1 11078 -1 0 107236
box -52 -62 11344 8684
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_0
timestamp 1683647856
transform 0 -1 42193 1 0 181600
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_1
timestamp 1683647856
transform 0 -1 42193 1 0 224800
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_2
timestamp 1683647856
transform 0 -1 42193 1 0 268000
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_3
timestamp 1683647856
transform 0 -1 42193 1 0 311200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_4
timestamp 1683647856
transform 0 -1 42193 1 0 354400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_5
timestamp 1683647856
transform 0 -1 42193 1 0 397600
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_6
timestamp 1683647856
transform 0 -1 42193 1 0 525200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_7
timestamp 1683647856
transform 0 -1 42193 1 0 568400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_8
timestamp 1683647856
transform 0 -1 42193 1 0 611600
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_9
timestamp 1683647856
transform 0 -1 42193 1 0 654800
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_10
timestamp 1683647856
transform 0 1 675407 -1 0 609000
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_11
timestamp 1683647856
transform 0 1 675407 -1 0 563800
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_12
timestamp 1683647856
transform 0 1 675407 -1 0 386600
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_13
timestamp 1683647856
transform 0 1 675407 -1 0 341400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_14
timestamp 1683647856
transform 0 1 675407 -1 0 296400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_15
timestamp 1683647856
transform 0 1 675407 -1 0 251400
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_16
timestamp 1683647856
transform 0 1 675407 -1 0 206200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_17
timestamp 1683647856
transform 0 1 675407 -1 0 161200
box -143 0 16134 42193
use sky130_ef_io__gpiov2_pad_wrapped  sky130_ef_io__gpiov2_pad_wrapped_18
timestamp 1683647856
transform 0 1 675407 -1 0 116000
box -143 0 16134 42193
use sky130_ef_io__corner_pad  user0_corner[0] $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform -1 0 40000 0 -1 40800
box 0 0 40000 40800
use sky130_ef_io__corner_pad  user0_corner[1]
timestamp 1683647856
transform 0 1 676800 -1 0 40000
box 0 0 40000 40800
use sky130_ef_io__corner_pad  user1_corner
timestamp 1683647856
transform 1 0 677600 0 1 996800
box 0 0 40000 40800
use sky130_ef_io__vccd_lvc_clamped3_pad  user1_vccd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform 0 1 678007 -1 0 922600
box 0 -2177 17187 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[0\]
timestamp 1683647856
transform 0 1 678007 -1 0 833400
box 0 -407 15000 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user1_vdda_hvclamp_pad\[1\]
timestamp 1683647856
transform 0 1 678007 -1 0 518800
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[0\]
timestamp 1683647856
transform 1 0 575600 0 1 998007
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user1_vssa_hvclamp_pad\[1\]
timestamp 1683647856
transform 0 1 678007 -1 0 430600
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  user1_vssd_lvclamp_pad $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1683647856
transform 0 1 678007 -1 0 474800
box 0 -2177 17187 39593
use sky130_ef_io__corner_pad  user2_corner
timestamp 1683647856
transform 0 -1 40800 1 0 997600
box 0 0 40000 40800
use sky130_ef_io__vccd_lvc_clamped3_pad  user2_vccd_lvclamp_pad
timestamp 1683647856
transform 0 -1 39593 1 0 912000
box 0 -2177 17187 39593
use sky130_ef_io__vdda_hvc_clamped_pad  user2_vdda_hvclamp_pad
timestamp 1683647856
transform 0 -1 39593 1 0 483000
box 0 -407 15000 39593
use sky130_ef_io__vssa_hvc_clamped_pad  user2_vssa_hvclamp_pad
timestamp 1683647856
transform 0 -1 39593 1 0 827600
box 0 -407 15000 39593
use sky130_ef_io__vssd_lvc_clamped3_pad  user2_vssd_lvclamp_pad
timestamp 1683647856
transform 0 -1 39593 1 0 440800
box 0 -2177 17187 39593
use user_id_textblock  user_id_textblock_0
timestamp 1608324878
transform 1 0 42717 0 1 6915
box -656 1508 33720 10344
use user_id_programming  user_id_value
timestamp 1650371074
transform 1 0 643154 0 1 9246
box 0 0 7109 7077
use xres_buf  xres_buf_0
timestamp 1678062433
transform -1 0 152583 0 1 16471
box 0 -400 4000 3800
<< labels >>
flabel metal3 s 675407 778996 675887 779066 0 FreeSans 400 0 0 0 gpio_analog_en[12]
port 453 nsew
flabel metal3 s 675407 780284 675887 780354 0 FreeSans 400 0 0 0 gpio_analog_pol[12]
port 541 nsew
flabel metal3 s 675407 783320 675887 783390 0 FreeSans 400 0 0 0 gpio_analog_sel[12]
port 497 nsew
flabel metal3 s 675407 779640 675887 779710 0 FreeSans 400 0 0 0 gpio_dm0[12]
port 585 nsew
flabel metal3 s 675407 777800 675887 777870 0 FreeSans 400 0 0 0 gpio_dm1[12]
port 629 nsew
flabel metal3 s 675407 783964 675887 784034 0 FreeSans 400 0 0 0 gpio_dm2[12]
port 673 nsew
flabel metal3 s 675407 784608 675887 784678 0 FreeSans 400 0 0 0 gpio_holdover[12]
port 409 nsew
flabel metal3 s 675407 787644 675887 787714 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[12]
port 277 nsew
flabel metal3 s 675407 780836 675887 780906 0 FreeSans 400 0 0 0 gpio_inp_dis[12]
port 233 nsew
flabel metal3 s 675407 788288 675887 788358 0 FreeSans 400 0 0 0 gpio_oeb[12]
port 189 nsew
flabel metal3 s 675407 785160 675887 785230 0 FreeSans 400 0 0 0 gpio_out[12]
port 145 nsew
flabel metal3 s 675407 775960 675887 776030 0 FreeSans 400 0 0 0 gpio_slow_sel[12]
port 365 nsew
flabel metal3 s 675407 787000 675887 787070 0 FreeSans 400 0 0 0 gpio_vtrip_sel[12]
port 321 nsew
flabel metal3 s 675407 774120 675887 774190 0 FreeSans 400 0 0 0 gpio_in[12]
port 717 nsew
flabel metal3 s 675407 868196 675887 868266 0 FreeSans 400 0 0 0 gpio_analog_en[13]
port 452 nsew
flabel metal3 s 675407 869484 675887 869554 0 FreeSans 400 0 0 0 gpio_analog_pol[13]
port 540 nsew
flabel metal3 s 675407 872520 675887 872590 0 FreeSans 400 0 0 0 gpio_analog_sel[13]
port 496 nsew
flabel metal3 s 675407 868840 675887 868910 0 FreeSans 400 0 0 0 gpio_dm0[13]
port 584 nsew
flabel metal3 s 675407 867000 675887 867070 0 FreeSans 400 0 0 0 gpio_dm1[13]
port 628 nsew
flabel metal3 s 675407 873164 675887 873234 0 FreeSans 400 0 0 0 gpio_dm2[13]
port 672 nsew
flabel metal3 s 675407 873808 675887 873878 0 FreeSans 400 0 0 0 gpio_holdover[13]
port 408 nsew
flabel metal3 s 675407 876844 675887 876914 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[13]
port 276 nsew
flabel metal3 s 675407 870036 675887 870106 0 FreeSans 400 0 0 0 gpio_inp_dis[13]
port 232 nsew
flabel metal3 s 675407 877488 675887 877558 0 FreeSans 400 0 0 0 gpio_oeb[13]
port 188 nsew
flabel metal3 s 675407 874360 675887 874430 0 FreeSans 400 0 0 0 gpio_out[13]
port 144 nsew
flabel metal3 s 675407 865160 675887 865230 0 FreeSans 400 0 0 0 gpio_slow_sel[13]
port 364 nsew
flabel metal3 s 675407 876200 675887 876270 0 FreeSans 400 0 0 0 gpio_vtrip_sel[13]
port 320 nsew
flabel metal3 s 675407 863320 675887 863390 0 FreeSans 400 0 0 0 gpio_in[13]
port 716 nsew
flabel metal3 s 675407 957396 675887 957466 0 FreeSans 400 0 0 0 gpio_analog_en[14]
port 451 nsew
flabel metal3 s 675407 958684 675887 958754 0 FreeSans 400 0 0 0 gpio_analog_pol[14]
port 539 nsew
flabel metal3 s 675407 961720 675887 961790 0 FreeSans 400 0 0 0 gpio_analog_sel[14]
port 495 nsew
flabel metal3 s 675407 958040 675887 958110 0 FreeSans 400 0 0 0 gpio_dm0[14]
port 583 nsew
flabel metal3 s 675407 956200 675887 956270 0 FreeSans 400 0 0 0 gpio_dm1[14]
port 627 nsew
flabel metal3 s 675407 962364 675887 962434 0 FreeSans 400 0 0 0 gpio_dm2[14]
port 671 nsew
flabel metal3 s 675407 963008 675887 963078 0 FreeSans 400 0 0 0 gpio_holdover[14]
port 407 nsew
flabel metal3 s 675407 966044 675887 966114 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[14]
port 275 nsew
flabel metal3 s 675407 959236 675887 959306 0 FreeSans 400 0 0 0 gpio_inp_dis[14]
port 231 nsew
flabel metal3 s 675407 966688 675887 966758 0 FreeSans 400 0 0 0 gpio_oeb[14]
port 187 nsew
flabel metal3 s 675407 963560 675887 963630 0 FreeSans 400 0 0 0 gpio_out[14]
port 143 nsew
flabel metal3 s 675407 954360 675887 954430 0 FreeSans 400 0 0 0 gpio_slow_sel[14]
port 363 nsew
flabel metal3 s 675407 965400 675887 965470 0 FreeSans 400 0 0 0 gpio_vtrip_sel[14]
port 319 nsew
flabel metal3 s 675407 952520 675887 952590 0 FreeSans 400 0 0 0 gpio_in[14]
port 715 nsew
flabel metal2 s 636141 995407 636197 995887 0 FreeSans 400 90 0 0 gpio_analog_en[15]
port 450 nsew
flabel metal2 s 634853 995407 634909 995887 0 FreeSans 400 90 0 0 gpio_analog_pol[15]
port 538 nsew
flabel metal2 s 631817 995407 631873 995887 0 FreeSans 400 90 0 0 gpio_analog_sel[15]
port 494 nsew
flabel metal2 s 635497 995407 635553 995887 0 FreeSans 400 90 0 0 gpio_dm0[15]
port 582 nsew
flabel metal2 s 637337 995407 637393 995887 0 FreeSans 400 90 0 0 gpio_dm1[15]
port 626 nsew
flabel metal2 s 631173 995407 631229 995887 0 FreeSans 400 90 0 0 gpio_dm2[15]
port 670 nsew
flabel metal2 s 630529 995407 630585 995887 0 FreeSans 400 90 0 0 gpio_holdover[15]
port 406 nsew
flabel metal2 s 627493 995407 627549 995887 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[15]
port 274 nsew
flabel metal2 s 634301 995407 634357 995887 0 FreeSans 400 90 0 0 gpio_inp_dis[15]
port 230 nsew
flabel metal2 s 626849 995407 626905 995887 0 FreeSans 400 90 0 0 gpio_oeb[15]
port 186 nsew
flabel metal2 s 629977 995407 630033 995887 0 FreeSans 400 90 0 0 gpio_out[15]
port 142 nsew
flabel metal2 s 639177 995407 639233 995887 0 FreeSans 400 90 0 0 gpio_slow_sel[15]
port 362 nsew
flabel metal2 s 628137 995407 628193 995887 0 FreeSans 400 90 0 0 gpio_vtrip_sel[15]
port 318 nsew
flabel metal2 s 641017 995407 641073 995887 0 FreeSans 400 90 0 0 gpio_in[15]
port 714 nsew
flabel metal2 s 534341 995407 534397 995887 0 FreeSans 400 90 0 0 gpio_analog_en[16]
port 449 nsew
flabel metal2 s 533053 995407 533109 995887 0 FreeSans 400 90 0 0 gpio_analog_pol[16]
port 537 nsew
flabel metal2 s 530017 995407 530073 995887 0 FreeSans 400 90 0 0 gpio_analog_sel[16]
port 493 nsew
flabel metal2 s 533697 995407 533753 995887 0 FreeSans 400 90 0 0 gpio_dm0[16]
port 581 nsew
flabel metal2 s 535537 995407 535593 995887 0 FreeSans 400 90 0 0 gpio_dm1[16]
port 625 nsew
flabel metal2 s 529373 995407 529429 995887 0 FreeSans 400 90 0 0 gpio_dm2[16]
port 669 nsew
flabel metal2 s 528729 995407 528785 995887 0 FreeSans 400 90 0 0 gpio_holdover[16]
port 405 nsew
flabel metal2 s 525693 995407 525749 995887 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[16]
port 273 nsew
flabel metal2 s 532501 995407 532557 995887 0 FreeSans 400 90 0 0 gpio_inp_dis[16]
port 229 nsew
flabel metal2 s 525049 995407 525105 995887 0 FreeSans 400 90 0 0 gpio_oeb[16]
port 185 nsew
flabel metal2 s 528177 995407 528233 995887 0 FreeSans 400 90 0 0 gpio_out[16]
port 141 nsew
flabel metal2 s 537377 995407 537433 995887 0 FreeSans 400 90 0 0 gpio_slow_sel[16]
port 361 nsew
flabel metal2 s 526337 995407 526393 995887 0 FreeSans 400 90 0 0 gpio_vtrip_sel[16]
port 317 nsew
flabel metal2 s 539217 995407 539273 995887 0 FreeSans 400 90 0 0 gpio_in[16]
port 713 nsew
flabel metal2 s 484137 995407 484193 995887 0 FreeSans 400 90 0 0 gpio_dm1[17]
port 624 nsew
flabel metal2 s 477973 995407 478029 995887 0 FreeSans 400 90 0 0 gpio_dm2[17]
port 668 nsew
flabel metal2 s 477329 995407 477385 995887 0 FreeSans 400 90 0 0 gpio_holdover[17]
port 404 nsew
flabel metal2 s 474293 995407 474349 995887 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[17]
port 272 nsew
flabel metal2 s 481101 995407 481157 995887 0 FreeSans 400 90 0 0 gpio_inp_dis[17]
port 228 nsew
flabel metal2 s 473649 995407 473705 995887 0 FreeSans 400 90 0 0 gpio_oeb[17]
port 184 nsew
flabel metal2 s 476777 995407 476833 995887 0 FreeSans 400 90 0 0 gpio_out[17]
port 140 nsew
flabel metal2 s 485977 995407 486033 995887 0 FreeSans 400 90 0 0 gpio_slow_sel[17]
port 360 nsew
flabel metal2 s 474937 995407 474993 995887 0 FreeSans 400 90 0 0 gpio_vtrip_sel[17]
port 316 nsew
flabel metal2 s 487817 995407 487873 995887 0 FreeSans 400 90 0 0 gpio_in[17]
port 712 nsew
flabel metal2 s 393941 995407 393997 995887 0 FreeSans 400 90 0 0 gpio_analog_en[18]
port 447 nsew
flabel metal2 s 392653 995407 392709 995887 0 FreeSans 400 90 0 0 gpio_analog_pol[18]
port 535 nsew
flabel metal2 s 389617 995407 389673 995887 0 FreeSans 400 90 0 0 gpio_analog_sel[18]
port 491 nsew
flabel metal2 s 393297 995407 393353 995887 0 FreeSans 400 90 0 0 gpio_dm0[18]
port 579 nsew
flabel metal2 s 395137 995407 395193 995887 0 FreeSans 400 90 0 0 gpio_dm1[18]
port 623 nsew
flabel metal2 s 388973 995407 389029 995887 0 FreeSans 400 90 0 0 gpio_dm2[18]
port 667 nsew
flabel metal2 s 388329 995407 388385 995887 0 FreeSans 400 90 0 0 gpio_holdover[18]
port 403 nsew
flabel metal2 s 385293 995407 385349 995887 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[18]
port 271 nsew
flabel metal2 s 392101 995407 392157 995887 0 FreeSans 400 90 0 0 gpio_inp_dis[18]
port 227 nsew
flabel metal2 s 384649 995407 384705 995887 0 FreeSans 400 90 0 0 gpio_oeb[18]
port 183 nsew
flabel metal2 s 387777 995407 387833 995887 0 FreeSans 400 90 0 0 gpio_out[18]
port 139 nsew
flabel metal2 s 396977 995407 397033 995887 0 FreeSans 400 90 0 0 gpio_slow_sel[18]
port 359 nsew
flabel metal2 s 385937 995407 385993 995887 0 FreeSans 400 90 0 0 gpio_vtrip_sel[18]
port 315 nsew
flabel metal2 s 398817 995407 398873 995887 0 FreeSans 400 90 0 0 gpio_in[18]
port 711 nsew
flabel metal2 s 482941 995407 482997 995887 0 FreeSans 400 90 0 0 gpio_analog_en[17]
port 448 nsew
flabel metal2 s 481653 995407 481709 995887 0 FreeSans 400 90 0 0 gpio_analog_pol[17]
port 536 nsew
flabel metal2 s 478617 995407 478673 995887 0 FreeSans 400 90 0 0 gpio_analog_sel[17]
port 492 nsew
flabel metal2 s 482297 995407 482353 995887 0 FreeSans 400 90 0 0 gpio_dm0[17]
port 580 nsew
flabel metal3 s 675407 739608 675887 739678 0 FreeSans 400 0 0 0 gpio_holdover[11]
port 410 nsew
flabel metal3 s 675407 742644 675887 742714 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[11]
port 278 nsew
flabel metal3 s 675407 735836 675887 735906 0 FreeSans 400 0 0 0 gpio_inp_dis[11]
port 234 nsew
flabel metal3 s 675407 743288 675887 743358 0 FreeSans 400 0 0 0 gpio_oeb[11]
port 190 nsew
flabel metal3 s 675407 740160 675887 740230 0 FreeSans 400 0 0 0 gpio_out[11]
port 146 nsew
flabel metal3 s 675407 730960 675887 731030 0 FreeSans 400 0 0 0 gpio_slow_sel[11]
port 366 nsew
flabel metal3 s 675407 742000 675887 742070 0 FreeSans 400 0 0 0 gpio_vtrip_sel[11]
port 322 nsew
flabel metal3 s 675407 729120 675887 729190 0 FreeSans 400 0 0 0 gpio_in[11]
port 718 nsew
flabel metal3 s 675407 688996 675887 689066 0 FreeSans 400 0 0 0 gpio_analog_en[10]
port 455 nsew
flabel metal3 s 675407 690284 675887 690354 0 FreeSans 400 0 0 0 gpio_analog_pol[10]
port 543 nsew
flabel metal3 s 675407 693320 675887 693390 0 FreeSans 400 0 0 0 gpio_analog_sel[10]
port 499 nsew
flabel metal3 s 675407 689640 675887 689710 0 FreeSans 400 0 0 0 gpio_dm0[10]
port 587 nsew
flabel metal3 s 675407 687800 675887 687870 0 FreeSans 400 0 0 0 gpio_dm1[10]
port 631 nsew
flabel metal3 s 675407 693964 675887 694034 0 FreeSans 400 0 0 0 gpio_dm2[10]
port 675 nsew
flabel metal3 s 675407 694608 675887 694678 0 FreeSans 400 0 0 0 gpio_holdover[10]
port 411 nsew
flabel metal3 s 675407 697644 675887 697714 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[10]
port 279 nsew
flabel metal3 s 675407 690836 675887 690906 0 FreeSans 400 0 0 0 gpio_inp_dis[10]
port 235 nsew
flabel metal3 s 675407 698288 675887 698358 0 FreeSans 400 0 0 0 gpio_oeb[10]
port 191 nsew
flabel metal3 s 675407 695160 675887 695230 0 FreeSans 400 0 0 0 gpio_out[10]
port 147 nsew
flabel metal3 s 675407 685960 675887 686030 0 FreeSans 400 0 0 0 gpio_slow_sel[10]
port 367 nsew
flabel metal3 s 675407 697000 675887 697070 0 FreeSans 400 0 0 0 gpio_vtrip_sel[10]
port 323 nsew
flabel metal3 s 675407 684120 675887 684190 0 FreeSans 400 0 0 0 gpio_in[10]
port 719 nsew
flabel metal3 s 675407 553596 675887 553666 0 FreeSans 400 0 0 0 gpio_analog_en[7]
port 458 nsew
flabel metal3 s 675407 554884 675887 554954 0 FreeSans 400 0 0 0 gpio_analog_pol[7]
port 546 nsew
flabel metal3 s 675407 557920 675887 557990 0 FreeSans 400 0 0 0 gpio_analog_sel[7]
port 502 nsew
flabel metal3 s 675407 554240 675887 554310 0 FreeSans 400 0 0 0 gpio_dm0[7]
port 590 nsew
flabel metal3 s 675407 552400 675887 552470 0 FreeSans 400 0 0 0 gpio_dm1[7]
port 634 nsew
flabel metal3 s 675407 558564 675887 558634 0 FreeSans 400 0 0 0 gpio_dm2[7]
port 678 nsew
flabel metal3 s 675407 559208 675887 559278 0 FreeSans 400 0 0 0 gpio_holdover[7]
port 414 nsew
flabel metal3 s 675407 562244 675887 562314 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[7]
port 282 nsew
flabel metal3 s 675407 555436 675887 555506 0 FreeSans 400 0 0 0 gpio_inp_dis[7]
port 238 nsew
flabel metal3 s 675407 562888 675887 562958 0 FreeSans 400 0 0 0 gpio_oeb[7]
port 194 nsew
flabel metal3 s 675407 559760 675887 559830 0 FreeSans 400 0 0 0 gpio_out[7]
port 150 nsew
flabel metal3 s 675407 550560 675887 550630 0 FreeSans 400 0 0 0 gpio_slow_sel[7]
port 370 nsew
flabel metal3 s 675407 561600 675887 561670 0 FreeSans 400 0 0 0 gpio_vtrip_sel[7]
port 326 nsew
flabel metal3 s 675407 548720 675887 548790 0 FreeSans 400 0 0 0 gpio_in[7]
port 722 nsew
flabel metal3 s 675407 598796 675887 598866 0 FreeSans 400 0 0 0 gpio_analog_en[8]
port 457 nsew
flabel metal3 s 675407 600084 675887 600154 0 FreeSans 400 0 0 0 gpio_analog_pol[8]
port 545 nsew
flabel metal3 s 675407 603120 675887 603190 0 FreeSans 400 0 0 0 gpio_analog_sel[8]
port 501 nsew
flabel metal3 s 675407 599440 675887 599510 0 FreeSans 400 0 0 0 gpio_dm0[8]
port 589 nsew
flabel metal3 s 675407 597600 675887 597670 0 FreeSans 400 0 0 0 gpio_dm1[8]
port 633 nsew
flabel metal3 s 675407 603764 675887 603834 0 FreeSans 400 0 0 0 gpio_dm2[8]
port 677 nsew
flabel metal3 s 675407 604408 675887 604478 0 FreeSans 400 0 0 0 gpio_holdover[8]
port 413 nsew
flabel metal3 s 675407 607444 675887 607514 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[8]
port 281 nsew
flabel metal3 s 675407 600636 675887 600706 0 FreeSans 400 0 0 0 gpio_inp_dis[8]
port 237 nsew
flabel metal3 s 675407 608088 675887 608158 0 FreeSans 400 0 0 0 gpio_oeb[8]
port 193 nsew
flabel metal3 s 675407 604960 675887 605030 0 FreeSans 400 0 0 0 gpio_out[8]
port 149 nsew
flabel metal3 s 675407 595760 675887 595830 0 FreeSans 400 0 0 0 gpio_slow_sel[8]
port 369 nsew
flabel metal3 s 675407 606800 675887 606870 0 FreeSans 400 0 0 0 gpio_vtrip_sel[8]
port 325 nsew
flabel metal3 s 675407 593920 675887 593990 0 FreeSans 400 0 0 0 gpio_in[8]
port 721 nsew
flabel metal3 s 675407 643796 675887 643866 0 FreeSans 400 0 0 0 gpio_analog_en[9]
port 456 nsew
flabel metal3 s 675407 645084 675887 645154 0 FreeSans 400 0 0 0 gpio_analog_pol[9]
port 544 nsew
flabel metal3 s 675407 648120 675887 648190 0 FreeSans 400 0 0 0 gpio_analog_sel[9]
port 500 nsew
flabel metal3 s 675407 644440 675887 644510 0 FreeSans 400 0 0 0 gpio_dm0[9]
port 588 nsew
flabel metal3 s 675407 642600 675887 642670 0 FreeSans 400 0 0 0 gpio_dm1[9]
port 632 nsew
flabel metal3 s 675407 648764 675887 648834 0 FreeSans 400 0 0 0 gpio_dm2[9]
port 676 nsew
flabel metal3 s 675407 649408 675887 649478 0 FreeSans 400 0 0 0 gpio_holdover[9]
port 412 nsew
flabel metal3 s 675407 652444 675887 652514 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[9]
port 280 nsew
flabel metal3 s 675407 645636 675887 645706 0 FreeSans 400 0 0 0 gpio_inp_dis[9]
port 236 nsew
flabel metal3 s 675407 653088 675887 653158 0 FreeSans 400 0 0 0 gpio_oeb[9]
port 192 nsew
flabel metal3 s 675407 649960 675887 650030 0 FreeSans 400 0 0 0 gpio_out[9]
port 148 nsew
flabel metal3 s 675407 640760 675887 640830 0 FreeSans 400 0 0 0 gpio_slow_sel[9]
port 368 nsew
flabel metal3 s 675407 651800 675887 651870 0 FreeSans 400 0 0 0 gpio_vtrip_sel[9]
port 324 nsew
flabel metal3 s 675407 638920 675887 638990 0 FreeSans 400 0 0 0 gpio_in[9]
port 720 nsew
flabel metal3 s 675407 733996 675887 734066 0 FreeSans 400 0 0 0 gpio_analog_en[11]
port 454 nsew
flabel metal3 s 675407 735284 675887 735354 0 FreeSans 400 0 0 0 gpio_analog_pol[11]
port 542 nsew
flabel metal3 s 675407 738320 675887 738390 0 FreeSans 400 0 0 0 gpio_analog_sel[11]
port 498 nsew
flabel metal3 s 675407 734640 675887 734710 0 FreeSans 400 0 0 0 gpio_dm0[11]
port 586 nsew
flabel metal3 s 675407 732800 675887 732870 0 FreeSans 400 0 0 0 gpio_dm1[11]
port 630 nsew
flabel metal3 s 675407 738964 675887 739034 0 FreeSans 400 0 0 0 gpio_dm2[11]
port 674 nsew
flabel metal2 s 295177 995407 295233 995887 0 FreeSans 400 90 0 0 gpio_slow_sel[19]
port 358 nsew
flabel metal2 s 284137 995407 284193 995887 0 FreeSans 400 90 0 0 gpio_vtrip_sel[19]
port 314 nsew
flabel metal2 s 297017 995407 297073 995887 0 FreeSans 400 90 0 0 gpio_in[19]
port 710 nsew
flabel metal2 s 240541 995407 240597 995887 0 FreeSans 400 90 0 0 gpio_analog_en[20]
port 445 nsew
flabel metal2 s 239253 995407 239309 995887 0 FreeSans 400 90 0 0 gpio_analog_pol[20]
port 533 nsew
flabel metal2 s 236217 995407 236273 995887 0 FreeSans 400 90 0 0 gpio_analog_sel[20]
port 489 nsew
flabel metal2 s 239897 995407 239953 995887 0 FreeSans 400 90 0 0 gpio_dm0[20]
port 577 nsew
flabel metal2 s 241737 995407 241793 995887 0 FreeSans 400 90 0 0 gpio_dm1[20]
port 621 nsew
flabel metal2 s 235573 995407 235629 995887 0 FreeSans 400 90 0 0 gpio_dm2[20]
port 665 nsew
flabel metal2 s 234929 995407 234985 995887 0 FreeSans 400 90 0 0 gpio_holdover[20]
port 401 nsew
flabel metal2 s 231893 995407 231949 995887 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[20]
port 269 nsew
flabel metal2 s 238701 995407 238757 995887 0 FreeSans 400 90 0 0 gpio_inp_dis[20]
port 225 nsew
flabel metal2 s 231249 995407 231305 995887 0 FreeSans 400 90 0 0 gpio_oeb[20]
port 181 nsew
flabel metal2 s 234377 995407 234433 995887 0 FreeSans 400 90 0 0 gpio_out[20]
port 137 nsew
flabel metal2 s 243577 995407 243633 995887 0 FreeSans 400 90 0 0 gpio_slow_sel[20]
port 357 nsew
flabel metal2 s 232537 995407 232593 995887 0 FreeSans 400 90 0 0 gpio_vtrip_sel[20]
port 313 nsew
flabel metal2 s 245417 995407 245473 995887 0 FreeSans 400 90 0 0 gpio_in[20]
port 709 nsew
flabel metal2 s 292141 995407 292197 995887 0 FreeSans 400 90 0 0 gpio_analog_en[19]
port 446 nsew
flabel metal2 s 290853 995407 290909 995887 0 FreeSans 400 90 0 0 gpio_analog_pol[19]
port 534 nsew
flabel metal2 s 287817 995407 287873 995887 0 FreeSans 400 90 0 0 gpio_analog_sel[19]
port 490 nsew
flabel metal2 s 291497 995407 291553 995887 0 FreeSans 400 90 0 0 gpio_dm0[19]
port 578 nsew
flabel metal2 s 293337 995407 293393 995887 0 FreeSans 400 90 0 0 gpio_dm1[19]
port 622 nsew
flabel metal2 s 287173 995407 287229 995887 0 FreeSans 400 90 0 0 gpio_dm2[19]
port 666 nsew
flabel metal2 s 286529 995407 286585 995887 0 FreeSans 400 90 0 0 gpio_holdover[19]
port 402 nsew
flabel metal2 s 283493 995407 283549 995887 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[19]
port 270 nsew
flabel metal2 s 290301 995407 290357 995887 0 FreeSans 400 90 0 0 gpio_inp_dis[19]
port 226 nsew
flabel metal2 s 282849 995407 282905 995887 0 FreeSans 400 90 0 0 gpio_oeb[19]
port 182 nsew
flabel metal2 s 285977 995407 286033 995887 0 FreeSans 400 90 0 0 gpio_out[19]
port 138 nsew
flabel metal2 s 194017 995407 194073 995887 0 FreeSans 400 90 0 0 gpio_in[21]
port 708 nsew
flabel metal2 s 137741 995407 137797 995887 0 FreeSans 400 90 0 0 gpio_analog_en[22]
port 443 nsew
flabel metal2 s 136453 995407 136509 995887 0 FreeSans 400 90 0 0 gpio_analog_pol[22]
port 531 nsew
flabel metal2 s 133417 995407 133473 995887 0 FreeSans 400 90 0 0 gpio_analog_sel[22]
port 487 nsew
flabel metal2 s 137097 995407 137153 995887 0 FreeSans 400 90 0 0 gpio_dm0[22]
port 575 nsew
flabel metal2 s 138937 995407 138993 995887 0 FreeSans 400 90 0 0 gpio_dm1[22]
port 619 nsew
flabel metal2 s 132773 995407 132829 995887 0 FreeSans 400 90 0 0 gpio_dm2[22]
port 663 nsew
flabel metal2 s 132129 995407 132185 995887 0 FreeSans 400 90 0 0 gpio_holdover[22]
port 399 nsew
flabel metal2 s 129093 995407 129149 995887 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[22]
port 267 nsew
flabel metal2 s 135901 995407 135957 995887 0 FreeSans 400 90 0 0 gpio_inp_dis[22]
port 223 nsew
flabel metal2 s 128449 995407 128505 995887 0 FreeSans 400 90 0 0 gpio_oeb[22]
port 179 nsew
flabel metal2 s 131577 995407 131633 995887 0 FreeSans 400 90 0 0 gpio_out[22]
port 135 nsew
flabel metal2 s 140777 995407 140833 995887 0 FreeSans 400 90 0 0 gpio_slow_sel[22]
port 355 nsew
flabel metal2 s 129737 995407 129793 995887 0 FreeSans 400 90 0 0 gpio_vtrip_sel[22]
port 311 nsew
flabel metal2 s 142617 995407 142673 995887 0 FreeSans 400 90 0 0 gpio_in[22]
port 707 nsew
flabel metal2 s 86341 995407 86397 995887 0 FreeSans 400 90 0 0 gpio_analog_en[23]
port 442 nsew
flabel metal2 s 85053 995407 85109 995887 0 FreeSans 400 90 0 0 gpio_analog_pol[23]
port 530 nsew
flabel metal2 s 82017 995407 82073 995887 0 FreeSans 400 90 0 0 gpio_analog_sel[23]
port 486 nsew
flabel metal2 s 85697 995407 85753 995887 0 FreeSans 400 90 0 0 gpio_dm0[23]
port 574 nsew
flabel metal2 s 87537 995407 87593 995887 0 FreeSans 400 90 0 0 gpio_dm1[23]
port 618 nsew
flabel metal2 s 81373 995407 81429 995887 0 FreeSans 400 90 0 0 gpio_dm2[23]
port 662 nsew
flabel metal2 s 80729 995407 80785 995887 0 FreeSans 400 90 0 0 gpio_holdover[23]
port 398 nsew
flabel metal2 s 77693 995407 77749 995887 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[23]
port 266 nsew
flabel metal2 s 84501 995407 84557 995887 0 FreeSans 400 90 0 0 gpio_inp_dis[23]
port 222 nsew
flabel metal2 s 77049 995407 77105 995887 0 FreeSans 400 90 0 0 gpio_oeb[23]
port 178 nsew
flabel metal2 s 80177 995407 80233 995887 0 FreeSans 400 90 0 0 gpio_out[23]
port 134 nsew
flabel metal2 s 89377 995407 89433 995887 0 FreeSans 400 90 0 0 gpio_slow_sel[23]
port 354 nsew
flabel metal2 s 78337 995407 78393 995887 0 FreeSans 400 90 0 0 gpio_vtrip_sel[23]
port 310 nsew
flabel metal2 s 91217 995407 91273 995887 0 FreeSans 400 90 0 0 gpio_in[23]
port 706 nsew
flabel metal3 s 41713 964334 42193 964404 0 FreeSans 400 0 0 0 gpio_analog_en[24]
port 441 nsew
flabel metal3 s 41713 963046 42193 963116 0 FreeSans 400 0 0 0 gpio_analog_pol[24]
port 529 nsew
flabel metal3 s 41713 960010 42193 960080 0 FreeSans 400 0 0 0 gpio_analog_sel[24]
port 485 nsew
flabel metal3 s 41713 963690 42193 963760 0 FreeSans 400 0 0 0 gpio_dm0[24]
port 573 nsew
flabel metal3 s 41713 965530 42193 965600 0 FreeSans 400 0 0 0 gpio_dm1[24]
port 617 nsew
flabel metal3 s 41713 959366 42193 959436 0 FreeSans 400 0 0 0 gpio_dm2[24]
port 661 nsew
flabel metal3 s 41713 958722 42193 958792 0 FreeSans 400 0 0 0 gpio_holdover[24]
port 397 nsew
flabel metal3 s 41713 955686 42193 955756 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[24]
port 265 nsew
flabel metal3 s 41713 962494 42193 962564 0 FreeSans 400 0 0 0 gpio_inp_dis[24]
port 221 nsew
flabel metal3 s 41713 955042 42193 955112 0 FreeSans 400 0 0 0 gpio_oeb[24]
port 177 nsew
flabel metal3 s 41713 958170 42193 958240 0 FreeSans 400 0 0 0 gpio_out[24]
port 133 nsew
flabel metal3 s 41713 967370 42193 967440 0 FreeSans 400 0 0 0 gpio_slow_sel[24]
port 353 nsew
flabel metal3 s 41713 956330 42193 956400 0 FreeSans 400 0 0 0 gpio_vtrip_sel[24]
port 309 nsew
flabel metal3 s 41713 969210 42193 969280 0 FreeSans 400 0 0 0 gpio_in[24]
port 705 nsew
flabel metal3 s 41713 794534 42193 794604 0 FreeSans 400 0 0 0 gpio_analog_en[25]
port 440 nsew
flabel metal3 s 41713 793246 42193 793316 0 FreeSans 400 0 0 0 gpio_analog_pol[25]
port 528 nsew
flabel metal3 s 41713 790210 42193 790280 0 FreeSans 400 0 0 0 gpio_analog_sel[25]
port 484 nsew
flabel metal3 s 41713 793890 42193 793960 0 FreeSans 400 0 0 0 gpio_dm0[25]
port 572 nsew
flabel metal3 s 41713 795730 42193 795800 0 FreeSans 400 0 0 0 gpio_dm1[25]
port 616 nsew
flabel metal3 s 41713 789566 42193 789636 0 FreeSans 400 0 0 0 gpio_dm2[25]
port 660 nsew
flabel metal3 s 41713 788922 42193 788992 0 FreeSans 400 0 0 0 gpio_holdover[25]
port 396 nsew
flabel metal3 s 41713 785886 42193 785956 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[25]
port 264 nsew
flabel metal3 s 41713 792694 42193 792764 0 FreeSans 400 0 0 0 gpio_inp_dis[25]
port 220 nsew
flabel metal3 s 41713 785242 42193 785312 0 FreeSans 400 0 0 0 gpio_oeb[25]
port 176 nsew
flabel metal3 s 41713 788370 42193 788440 0 FreeSans 400 0 0 0 gpio_out[25]
port 132 nsew
flabel metal3 s 41713 797570 42193 797640 0 FreeSans 400 0 0 0 gpio_slow_sel[25]
port 352 nsew
flabel metal3 s 41713 786530 42193 786600 0 FreeSans 400 0 0 0 gpio_vtrip_sel[25]
port 308 nsew
flabel metal3 s 41713 799410 42193 799480 0 FreeSans 400 0 0 0 gpio_in[25]
port 704 nsew
flabel metal2 s 189141 995407 189197 995887 0 FreeSans 400 90 0 0 gpio_analog_en[21]
port 444 nsew
flabel metal2 s 187853 995407 187909 995887 0 FreeSans 400 90 0 0 gpio_analog_pol[21]
port 532 nsew
flabel metal2 s 184817 995407 184873 995887 0 FreeSans 400 90 0 0 gpio_analog_sel[21]
port 488 nsew
flabel metal2 s 188497 995407 188553 995887 0 FreeSans 400 90 0 0 gpio_dm0[21]
port 576 nsew
flabel metal2 s 190337 995407 190393 995887 0 FreeSans 400 90 0 0 gpio_dm1[21]
port 620 nsew
flabel metal2 s 184173 995407 184229 995887 0 FreeSans 400 90 0 0 gpio_dm2[21]
port 664 nsew
flabel metal2 s 183529 995407 183585 995887 0 FreeSans 400 90 0 0 gpio_holdover[21]
port 400 nsew
flabel metal2 s 180493 995407 180549 995887 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[21]
port 268 nsew
flabel metal2 s 187301 995407 187357 995887 0 FreeSans 400 90 0 0 gpio_inp_dis[21]
port 224 nsew
flabel metal2 s 179849 995407 179905 995887 0 FreeSans 400 90 0 0 gpio_oeb[21]
port 180 nsew
flabel metal2 s 182977 995407 183033 995887 0 FreeSans 400 90 0 0 gpio_out[21]
port 136 nsew
flabel metal2 s 192177 995407 192233 995887 0 FreeSans 400 90 0 0 gpio_slow_sel[21]
port 356 nsew
flabel metal2 s 181137 995407 181193 995887 0 FreeSans 400 90 0 0 gpio_vtrip_sel[21]
port 312 nsew
flabel metal3 s 41713 577890 42193 577960 0 FreeSans 400 0 0 0 gpio_dm0[30]
port 567 nsew
flabel metal3 s 41713 579730 42193 579800 0 FreeSans 400 0 0 0 gpio_dm1[30]
port 611 nsew
flabel metal3 s 41713 573566 42193 573636 0 FreeSans 400 0 0 0 gpio_dm2[30]
port 655 nsew
flabel metal3 s 41713 572922 42193 572992 0 FreeSans 400 0 0 0 gpio_holdover[30]
port 391 nsew
flabel metal3 s 41713 569886 42193 569956 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[30]
port 259 nsew
flabel metal3 s 41713 576694 42193 576764 0 FreeSans 400 0 0 0 gpio_inp_dis[30]
port 215 nsew
flabel metal3 s 41713 569242 42193 569312 0 FreeSans 400 0 0 0 gpio_oeb[30]
port 171 nsew
flabel metal3 s 41713 572370 42193 572440 0 FreeSans 400 0 0 0 gpio_out[30]
port 127 nsew
flabel metal3 s 41713 581570 42193 581640 0 FreeSans 400 0 0 0 gpio_slow_sel[30]
port 347 nsew
flabel metal3 s 41713 570530 42193 570600 0 FreeSans 400 0 0 0 gpio_vtrip_sel[30]
port 303 nsew
flabel metal3 s 41713 583410 42193 583480 0 FreeSans 400 0 0 0 gpio_in[30]
port 699 nsew
flabel metal3 s 41713 535334 42193 535404 0 FreeSans 400 0 0 0 gpio_analog_en[31]
port 434 nsew
flabel metal3 s 41713 534046 42193 534116 0 FreeSans 400 0 0 0 gpio_analog_pol[31]
port 522 nsew
flabel metal3 s 41713 531010 42193 531080 0 FreeSans 400 0 0 0 gpio_analog_sel[31]
port 478 nsew
flabel metal3 s 41713 534690 42193 534760 0 FreeSans 400 0 0 0 gpio_dm0[31]
port 566 nsew
flabel metal3 s 41713 536530 42193 536600 0 FreeSans 400 0 0 0 gpio_dm1[31]
port 610 nsew
flabel metal3 s 41713 530366 42193 530436 0 FreeSans 400 0 0 0 gpio_dm2[31]
port 654 nsew
flabel metal3 s 41713 529722 42193 529792 0 FreeSans 400 0 0 0 gpio_holdover[31]
port 390 nsew
flabel metal3 s 41713 526686 42193 526756 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[31]
port 258 nsew
flabel metal3 s 41713 533494 42193 533564 0 FreeSans 400 0 0 0 gpio_inp_dis[31]
port 214 nsew
flabel metal3 s 41713 526042 42193 526112 0 FreeSans 400 0 0 0 gpio_oeb[31]
port 170 nsew
flabel metal3 s 41713 529170 42193 529240 0 FreeSans 400 0 0 0 gpio_out[31]
port 126 nsew
flabel metal3 s 41713 538370 42193 538440 0 FreeSans 400 0 0 0 gpio_slow_sel[31]
port 346 nsew
flabel metal3 s 41713 527330 42193 527400 0 FreeSans 400 0 0 0 gpio_vtrip_sel[31]
port 302 nsew
flabel metal3 s 41713 540210 42193 540280 0 FreeSans 400 0 0 0 gpio_in[31]
port 698 nsew
flabel metal3 s 41713 751334 42193 751404 0 FreeSans 400 0 0 0 gpio_analog_en[26]
port 439 nsew
flabel metal3 s 41713 750046 42193 750116 0 FreeSans 400 0 0 0 gpio_analog_pol[26]
port 527 nsew
flabel metal3 s 41713 747010 42193 747080 0 FreeSans 400 0 0 0 gpio_analog_sel[26]
port 483 nsew
flabel metal3 s 41713 750690 42193 750760 0 FreeSans 400 0 0 0 gpio_dm0[26]
port 571 nsew
flabel metal3 s 41713 752530 42193 752600 0 FreeSans 400 0 0 0 gpio_dm1[26]
port 615 nsew
flabel metal3 s 41713 746366 42193 746436 0 FreeSans 400 0 0 0 gpio_dm2[26]
port 659 nsew
flabel metal3 s 41713 745722 42193 745792 0 FreeSans 400 0 0 0 gpio_holdover[26]
port 395 nsew
flabel metal3 s 41713 742686 42193 742756 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[26]
port 263 nsew
flabel metal3 s 41713 749494 42193 749564 0 FreeSans 400 0 0 0 gpio_inp_dis[26]
port 219 nsew
flabel metal3 s 41713 742042 42193 742112 0 FreeSans 400 0 0 0 gpio_oeb[26]
port 175 nsew
flabel metal3 s 41713 745170 42193 745240 0 FreeSans 400 0 0 0 gpio_out[26]
port 131 nsew
flabel metal3 s 41713 754370 42193 754440 0 FreeSans 400 0 0 0 gpio_slow_sel[26]
port 351 nsew
flabel metal3 s 41713 743330 42193 743400 0 FreeSans 400 0 0 0 gpio_vtrip_sel[26]
port 307 nsew
flabel metal3 s 41713 756210 42193 756280 0 FreeSans 400 0 0 0 gpio_in[26]
port 703 nsew
flabel metal3 s 41713 708134 42193 708204 0 FreeSans 400 0 0 0 gpio_analog_en[27]
port 438 nsew
flabel metal3 s 41713 706846 42193 706916 0 FreeSans 400 0 0 0 gpio_analog_pol[27]
port 526 nsew
flabel metal3 s 41713 703810 42193 703880 0 FreeSans 400 0 0 0 gpio_analog_sel[27]
port 482 nsew
flabel metal3 s 41713 707490 42193 707560 0 FreeSans 400 0 0 0 gpio_dm0[27]
port 570 nsew
flabel metal3 s 41713 709330 42193 709400 0 FreeSans 400 0 0 0 gpio_dm1[27]
port 614 nsew
flabel metal3 s 41713 703166 42193 703236 0 FreeSans 400 0 0 0 gpio_dm2[27]
port 658 nsew
flabel metal3 s 41713 702522 42193 702592 0 FreeSans 400 0 0 0 gpio_holdover[27]
port 394 nsew
flabel metal3 s 41713 699486 42193 699556 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[27]
port 262 nsew
flabel metal3 s 41713 706294 42193 706364 0 FreeSans 400 0 0 0 gpio_inp_dis[27]
port 218 nsew
flabel metal3 s 41713 698842 42193 698912 0 FreeSans 400 0 0 0 gpio_oeb[27]
port 174 nsew
flabel metal3 s 41713 701970 42193 702040 0 FreeSans 400 0 0 0 gpio_out[27]
port 130 nsew
flabel metal3 s 41713 711170 42193 711240 0 FreeSans 400 0 0 0 gpio_slow_sel[27]
port 350 nsew
flabel metal3 s 41713 700130 42193 700200 0 FreeSans 400 0 0 0 gpio_vtrip_sel[27]
port 306 nsew
flabel metal3 s 41713 713010 42193 713080 0 FreeSans 400 0 0 0 gpio_in[27]
port 702 nsew
flabel metal3 s 41713 664934 42193 665004 0 FreeSans 400 0 0 0 gpio_analog_en[28]
port 437 nsew
flabel metal3 s 41713 663646 42193 663716 0 FreeSans 400 0 0 0 gpio_analog_pol[28]
port 525 nsew
flabel metal3 s 41713 660610 42193 660680 0 FreeSans 400 0 0 0 gpio_analog_sel[28]
port 481 nsew
flabel metal3 s 41713 664290 42193 664360 0 FreeSans 400 0 0 0 gpio_dm0[28]
port 569 nsew
flabel metal3 s 41713 666130 42193 666200 0 FreeSans 400 0 0 0 gpio_dm1[28]
port 613 nsew
flabel metal3 s 41713 659966 42193 660036 0 FreeSans 400 0 0 0 gpio_dm2[28]
port 657 nsew
flabel metal3 s 41713 659322 42193 659392 0 FreeSans 400 0 0 0 gpio_holdover[28]
port 393 nsew
flabel metal3 s 41713 656286 42193 656356 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[28]
port 261 nsew
flabel metal3 s 41713 663094 42193 663164 0 FreeSans 400 0 0 0 gpio_inp_dis[28]
port 217 nsew
flabel metal3 s 41713 655642 42193 655712 0 FreeSans 400 0 0 0 gpio_oeb[28]
port 173 nsew
flabel metal3 s 41713 658770 42193 658840 0 FreeSans 400 0 0 0 gpio_out[28]
port 129 nsew
flabel metal3 s 41713 667970 42193 668040 0 FreeSans 400 0 0 0 gpio_slow_sel[28]
port 349 nsew
flabel metal3 s 41713 656930 42193 657000 0 FreeSans 400 0 0 0 gpio_vtrip_sel[28]
port 305 nsew
flabel metal3 s 41713 669810 42193 669880 0 FreeSans 400 0 0 0 gpio_in[28]
port 701 nsew
flabel metal3 s 41713 621734 42193 621804 0 FreeSans 400 0 0 0 gpio_analog_en[29]
port 436 nsew
flabel metal3 s 41713 620446 42193 620516 0 FreeSans 400 0 0 0 gpio_analog_pol[29]
port 524 nsew
flabel metal3 s 41713 617410 42193 617480 0 FreeSans 400 0 0 0 gpio_analog_sel[29]
port 480 nsew
flabel metal3 s 41713 621090 42193 621160 0 FreeSans 400 0 0 0 gpio_dm0[29]
port 568 nsew
flabel metal3 s 41713 622930 42193 623000 0 FreeSans 400 0 0 0 gpio_dm1[29]
port 612 nsew
flabel metal3 s 41713 616766 42193 616836 0 FreeSans 400 0 0 0 gpio_dm2[29]
port 656 nsew
flabel metal3 s 41713 616122 42193 616192 0 FreeSans 400 0 0 0 gpio_holdover[29]
port 392 nsew
flabel metal3 s 41713 613086 42193 613156 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[29]
port 260 nsew
flabel metal3 s 41713 619894 42193 619964 0 FreeSans 400 0 0 0 gpio_inp_dis[29]
port 216 nsew
flabel metal3 s 41713 612442 42193 612512 0 FreeSans 400 0 0 0 gpio_oeb[29]
port 172 nsew
flabel metal3 s 41713 615570 42193 615640 0 FreeSans 400 0 0 0 gpio_out[29]
port 128 nsew
flabel metal3 s 41713 624770 42193 624840 0 FreeSans 400 0 0 0 gpio_slow_sel[29]
port 348 nsew
flabel metal3 s 41713 613730 42193 613800 0 FreeSans 400 0 0 0 gpio_vtrip_sel[29]
port 304 nsew
flabel metal3 s 41713 626610 42193 626680 0 FreeSans 400 0 0 0 gpio_in[29]
port 700 nsew
flabel metal3 s 41713 578534 42193 578604 0 FreeSans 400 0 0 0 gpio_analog_en[30]
port 435 nsew
flabel metal3 s 41713 577246 42193 577316 0 FreeSans 400 0 0 0 gpio_analog_pol[30]
port 523 nsew
flabel metal3 s 41713 574210 42193 574280 0 FreeSans 400 0 0 0 gpio_analog_sel[30]
port 479 nsew
flabel metal3 s 41713 236130 42193 236200 0 FreeSans 400 0 0 0 gpio_dm1[36]
port 605 nsew
flabel metal3 s 41713 229966 42193 230036 0 FreeSans 400 0 0 0 gpio_dm2[36]
port 649 nsew
flabel metal3 s 41713 229322 42193 229392 0 FreeSans 400 0 0 0 gpio_holdover[36]
port 385 nsew
flabel metal3 s 41713 226286 42193 226356 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[36]
port 253 nsew
flabel metal3 s 41713 233094 42193 233164 0 FreeSans 400 0 0 0 gpio_inp_dis[36]
port 209 nsew
flabel metal3 s 41713 225642 42193 225712 0 FreeSans 400 0 0 0 gpio_oeb[36]
port 165 nsew
flabel metal3 s 41713 228770 42193 228840 0 FreeSans 400 0 0 0 gpio_out[36]
port 121 nsew
flabel metal3 s 41713 237970 42193 238040 0 FreeSans 400 0 0 0 gpio_slow_sel[36]
port 341 nsew
flabel metal3 s 41713 226930 42193 227000 0 FreeSans 400 0 0 0 gpio_vtrip_sel[36]
port 297 nsew
flabel metal3 s 41713 239810 42193 239880 0 FreeSans 400 0 0 0 gpio_in[36]
port 693 nsew
flabel metal3 s 41713 191734 42193 191804 0 FreeSans 400 0 0 0 gpio_analog_en[37]
port 428 nsew
flabel metal3 s 41713 190446 42193 190516 0 FreeSans 400 0 0 0 gpio_analog_pol[37]
port 516 nsew
flabel metal3 s 41713 187410 42193 187480 0 FreeSans 400 0 0 0 gpio_analog_sel[37]
port 472 nsew
flabel metal3 s 41713 191090 42193 191160 0 FreeSans 400 0 0 0 gpio_dm0[37]
port 560 nsew
flabel metal3 s 41713 192930 42193 193000 0 FreeSans 400 0 0 0 gpio_dm1[37]
port 604 nsew
flabel metal3 s 41713 186766 42193 186836 0 FreeSans 400 0 0 0 gpio_dm2[37]
port 648 nsew
flabel metal3 s 41713 186122 42193 186192 0 FreeSans 400 0 0 0 gpio_holdover[37]
port 384 nsew
flabel metal3 s 41713 183086 42193 183156 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[37]
port 252 nsew
flabel metal3 s 41713 182442 42193 182512 0 FreeSans 400 0 0 0 gpio_oeb[37]
port 164 nsew
flabel metal3 s 41713 185570 42193 185640 0 FreeSans 400 0 0 0 gpio_out[37]
port 120 nsew
flabel metal3 s 41713 194770 42193 194840 0 FreeSans 400 0 0 0 gpio_slow_sel[37]
port 340 nsew
flabel metal3 s 41713 183730 42193 183800 0 FreeSans 400 0 0 0 gpio_vtrip_sel[37]
port 296 nsew
flabel metal3 s 41713 196610 42193 196680 0 FreeSans 400 0 0 0 gpio_in[37]
port 692 nsew
flabel metal3 s 41713 407734 42193 407804 0 FreeSans 400 0 0 0 gpio_analog_en[32]
port 433 nsew
flabel metal3 s 41713 406446 42193 406516 0 FreeSans 400 0 0 0 gpio_analog_pol[32]
port 521 nsew
flabel metal3 s 41713 403410 42193 403480 0 FreeSans 400 0 0 0 gpio_analog_sel[32]
port 477 nsew
flabel metal3 s 41713 407090 42193 407160 0 FreeSans 400 0 0 0 gpio_dm0[32]
port 565 nsew
flabel metal3 s 41713 408930 42193 409000 0 FreeSans 400 0 0 0 gpio_dm1[32]
port 609 nsew
flabel metal3 s 41713 402766 42193 402836 0 FreeSans 400 0 0 0 gpio_dm2[32]
port 653 nsew
flabel metal3 s 41713 402122 42193 402192 0 FreeSans 400 0 0 0 gpio_holdover[32]
port 389 nsew
flabel metal3 s 41713 399086 42193 399156 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[32]
port 257 nsew
flabel metal3 s 41713 405894 42193 405964 0 FreeSans 400 0 0 0 gpio_inp_dis[32]
port 213 nsew
flabel metal3 s 41713 398442 42193 398512 0 FreeSans 400 0 0 0 gpio_oeb[32]
port 169 nsew
flabel metal3 s 41713 401570 42193 401640 0 FreeSans 400 0 0 0 gpio_out[32]
port 125 nsew
flabel metal3 s 41713 410770 42193 410840 0 FreeSans 400 0 0 0 gpio_slow_sel[32]
port 345 nsew
flabel metal3 s 41713 399730 42193 399800 0 FreeSans 400 0 0 0 gpio_vtrip_sel[32]
port 301 nsew
flabel metal3 s 41713 412610 42193 412680 0 FreeSans 400 0 0 0 gpio_in[32]
port 697 nsew
flabel metal3 s 41713 364534 42193 364604 0 FreeSans 400 0 0 0 gpio_analog_en[33]
port 432 nsew
flabel metal3 s 41713 363246 42193 363316 0 FreeSans 400 0 0 0 gpio_analog_pol[33]
port 520 nsew
flabel metal3 s 41713 360210 42193 360280 0 FreeSans 400 0 0 0 gpio_analog_sel[33]
port 476 nsew
flabel metal3 s 41713 365730 42193 365800 0 FreeSans 400 0 0 0 gpio_dm1[33]
port 608 nsew
flabel metal3 s 41713 359566 42193 359636 0 FreeSans 400 0 0 0 gpio_dm2[33]
port 652 nsew
flabel metal3 s 41713 363890 42193 363960 0 FreeSans 400 0 0 0 gpio_dm0[33]
port 564 nsew
flabel metal3 s 41713 358922 42193 358992 0 FreeSans 400 0 0 0 gpio_holdover[33]
port 388 nsew
flabel metal3 s 41713 355886 42193 355956 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[33]
port 256 nsew
flabel metal3 s 41713 362694 42193 362764 0 FreeSans 400 0 0 0 gpio_inp_dis[33]
port 212 nsew
flabel metal3 s 41713 355242 42193 355312 0 FreeSans 400 0 0 0 gpio_oeb[33]
port 168 nsew
flabel metal3 s 41713 358370 42193 358440 0 FreeSans 400 0 0 0 gpio_out[33]
port 124 nsew
flabel metal3 s 41713 367570 42193 367640 0 FreeSans 400 0 0 0 gpio_slow_sel[33]
port 344 nsew
flabel metal3 s 41713 356530 42193 356600 0 FreeSans 400 0 0 0 gpio_vtrip_sel[33]
port 300 nsew
flabel metal3 s 41713 369410 42193 369480 0 FreeSans 400 0 0 0 gpio_in[33]
port 696 nsew
flabel metal3 s 41713 321334 42193 321404 0 FreeSans 400 0 0 0 gpio_analog_en[34]
port 431 nsew
flabel metal3 s 41713 320046 42193 320116 0 FreeSans 400 0 0 0 gpio_analog_pol[34]
port 519 nsew
flabel metal3 s 41713 317010 42193 317080 0 FreeSans 400 0 0 0 gpio_analog_sel[34]
port 475 nsew
flabel metal3 s 41713 320690 42193 320760 0 FreeSans 400 0 0 0 gpio_dm0[34]
port 563 nsew
flabel metal3 s 41713 322530 42193 322600 0 FreeSans 400 0 0 0 gpio_dm1[34]
port 607 nsew
flabel metal3 s 41713 316366 42193 316436 0 FreeSans 400 0 0 0 gpio_dm2[34]
port 651 nsew
flabel metal3 s 41713 315722 42193 315792 0 FreeSans 400 0 0 0 gpio_holdover[34]
port 387 nsew
flabel metal3 s 41713 312686 42193 312756 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[34]
port 255 nsew
flabel metal3 s 41713 319494 42193 319564 0 FreeSans 400 0 0 0 gpio_inp_dis[34]
port 211 nsew
flabel metal3 s 41713 312042 42193 312112 0 FreeSans 400 0 0 0 gpio_oeb[34]
port 167 nsew
flabel metal3 s 41713 315170 42193 315240 0 FreeSans 400 0 0 0 gpio_out[34]
port 123 nsew
flabel metal3 s 41713 324370 42193 324440 0 FreeSans 400 0 0 0 gpio_slow_sel[34]
port 343 nsew
flabel metal3 s 41713 313330 42193 313400 0 FreeSans 400 0 0 0 gpio_vtrip_sel[34]
port 299 nsew
flabel metal3 s 41713 326210 42193 326280 0 FreeSans 400 0 0 0 gpio_in[34]
port 695 nsew
flabel metal3 s 41713 278134 42193 278204 0 FreeSans 400 0 0 0 gpio_analog_en[35]
port 430 nsew
flabel metal3 s 41713 276846 42193 276916 0 FreeSans 400 0 0 0 gpio_analog_pol[35]
port 518 nsew
flabel metal3 s 41713 273810 42193 273880 0 FreeSans 400 0 0 0 gpio_analog_sel[35]
port 474 nsew
flabel metal3 s 41713 277490 42193 277560 0 FreeSans 400 0 0 0 gpio_dm0[35]
port 562 nsew
flabel metal3 s 41713 279330 42193 279400 0 FreeSans 400 0 0 0 gpio_dm1[35]
port 606 nsew
flabel metal3 s 41713 273166 42193 273236 0 FreeSans 400 0 0 0 gpio_dm2[35]
port 650 nsew
flabel metal3 s 41713 272522 42193 272592 0 FreeSans 400 0 0 0 gpio_holdover[35]
port 386 nsew
flabel metal3 s 41713 269486 42193 269556 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[35]
port 254 nsew
flabel metal3 s 41713 276294 42193 276364 0 FreeSans 400 0 0 0 gpio_inp_dis[35]
port 210 nsew
flabel metal3 s 41713 268842 42193 268912 0 FreeSans 400 0 0 0 gpio_oeb[35]
port 166 nsew
flabel metal3 s 41713 271970 42193 272040 0 FreeSans 400 0 0 0 gpio_out[35]
port 122 nsew
flabel metal3 s 41713 281170 42193 281240 0 FreeSans 400 0 0 0 gpio_slow_sel[35]
port 342 nsew
flabel metal3 s 41713 270130 42193 270200 0 FreeSans 400 0 0 0 gpio_vtrip_sel[35]
port 298 nsew
flabel metal3 s 41713 283010 42193 283080 0 FreeSans 400 0 0 0 gpio_in[35]
port 694 nsew
flabel metal3 s 41713 234934 42193 235004 0 FreeSans 400 0 0 0 gpio_analog_en[36]
port 429 nsew
flabel metal3 s 41713 233646 42193 233716 0 FreeSans 400 0 0 0 gpio_analog_pol[36]
port 517 nsew
flabel metal3 s 41713 230610 42193 230680 0 FreeSans 400 0 0 0 gpio_analog_sel[36]
port 473 nsew
flabel metal3 s 41713 234290 42193 234360 0 FreeSans 400 0 0 0 gpio_dm0[36]
port 561 nsew
flabel metal3 s 675407 286196 675887 286266 0 FreeSans 400 0 0 0 gpio_analog_en[4]
port 461 nsew
flabel metal3 s 675407 287484 675887 287554 0 FreeSans 400 0 0 0 gpio_analog_pol[4]
port 549 nsew
flabel metal3 s 675407 290520 675887 290590 0 FreeSans 400 0 0 0 gpio_analog_sel[4]
port 505 nsew
flabel metal3 s 675407 286840 675887 286910 0 FreeSans 400 0 0 0 gpio_dm0[4]
port 593 nsew
flabel metal3 s 675407 285000 675887 285070 0 FreeSans 400 0 0 0 gpio_dm1[4]
port 637 nsew
flabel metal3 s 675407 291164 675887 291234 0 FreeSans 400 0 0 0 gpio_dm2[4]
port 681 nsew
flabel metal3 s 675407 291808 675887 291878 0 FreeSans 400 0 0 0 gpio_holdover[4]
port 417 nsew
flabel metal3 s 675407 294844 675887 294914 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[4]
port 285 nsew
flabel metal3 s 675407 288036 675887 288106 0 FreeSans 400 0 0 0 gpio_inp_dis[4]
port 241 nsew
flabel metal3 s 675407 295488 675887 295558 0 FreeSans 400 0 0 0 gpio_oeb[4]
port 197 nsew
flabel metal3 s 675407 292360 675887 292430 0 FreeSans 400 0 0 0 gpio_out[4]
port 153 nsew
flabel metal3 s 675407 283160 675887 283230 0 FreeSans 400 0 0 0 gpio_slow_sel[4]
port 373 nsew
flabel metal3 s 675407 294200 675887 294270 0 FreeSans 400 0 0 0 gpio_vtrip_sel[4]
port 329 nsew
flabel metal3 s 675407 281320 675887 281390 0 FreeSans 400 0 0 0 gpio_in[4]
port 725 nsew
flabel metal3 s 675407 331196 675887 331266 0 FreeSans 400 0 0 0 gpio_analog_en[5]
port 460 nsew
flabel metal3 s 675407 332484 675887 332554 0 FreeSans 400 0 0 0 gpio_analog_pol[5]
port 548 nsew
flabel metal3 s 675407 335520 675887 335590 0 FreeSans 400 0 0 0 gpio_analog_sel[5]
port 504 nsew
flabel metal3 s 675407 331840 675887 331910 0 FreeSans 400 0 0 0 gpio_dm0[5]
port 592 nsew
flabel metal3 s 675407 330000 675887 330070 0 FreeSans 400 0 0 0 gpio_dm1[5]
port 636 nsew
flabel metal3 s 675407 336164 675887 336234 0 FreeSans 400 0 0 0 gpio_dm2[5]
port 680 nsew
flabel metal3 s 675407 336808 675887 336878 0 FreeSans 400 0 0 0 gpio_holdover[5]
port 416 nsew
flabel metal3 s 675407 339844 675887 339914 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[5]
port 284 nsew
flabel metal3 s 675407 333036 675887 333106 0 FreeSans 400 0 0 0 gpio_inp_dis[5]
port 240 nsew
flabel metal3 s 675407 340488 675887 340558 0 FreeSans 400 0 0 0 gpio_oeb[5]
port 196 nsew
flabel metal3 s 675407 337360 675887 337430 0 FreeSans 400 0 0 0 gpio_out[5]
port 152 nsew
flabel metal3 s 675407 328160 675887 328230 0 FreeSans 400 0 0 0 gpio_slow_sel[5]
port 372 nsew
flabel metal3 s 675407 339200 675887 339270 0 FreeSans 400 0 0 0 gpio_vtrip_sel[5]
port 328 nsew
flabel metal3 s 675407 376396 675887 376466 0 FreeSans 400 0 0 0 gpio_analog_en[6]
port 459 nsew
flabel metal3 s 675407 377684 675887 377754 0 FreeSans 400 0 0 0 gpio_analog_pol[6]
port 547 nsew
flabel metal3 s 675407 380720 675887 380790 0 FreeSans 400 0 0 0 gpio_analog_sel[6]
port 503 nsew
flabel metal3 s 675407 377040 675887 377110 0 FreeSans 400 0 0 0 gpio_dm0[6]
port 591 nsew
flabel metal3 s 675407 375200 675887 375270 0 FreeSans 400 0 0 0 gpio_dm1[6]
port 635 nsew
flabel metal3 s 675407 381364 675887 381434 0 FreeSans 400 0 0 0 gpio_dm2[6]
port 679 nsew
flabel metal3 s 675407 382008 675887 382078 0 FreeSans 400 0 0 0 gpio_holdover[6]
port 415 nsew
flabel metal3 s 675407 385044 675887 385114 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[6]
port 283 nsew
flabel metal3 s 675407 378236 675887 378306 0 FreeSans 400 0 0 0 gpio_inp_dis[6]
port 239 nsew
flabel metal3 s 675407 385688 675887 385758 0 FreeSans 400 0 0 0 gpio_oeb[6]
port 195 nsew
flabel metal3 s 675407 382560 675887 382630 0 FreeSans 400 0 0 0 gpio_out[6]
port 151 nsew
flabel metal3 s 675407 373360 675887 373430 0 FreeSans 400 0 0 0 gpio_slow_sel[6]
port 371 nsew
flabel metal3 s 675407 384400 675887 384470 0 FreeSans 400 0 0 0 gpio_vtrip_sel[6]
port 327 nsew
flabel metal3 s 675407 371520 675887 371590 0 FreeSans 400 0 0 0 gpio_in[6]
port 723 nsew
flabel metal3 s 675407 150996 675887 151066 0 FreeSans 400 0 0 0 gpio_analog_en[1]
port 464 nsew
flabel metal3 s 675407 152284 675887 152354 0 FreeSans 400 0 0 0 gpio_analog_pol[1]
port 552 nsew
flabel metal3 s 675407 155320 675887 155390 0 FreeSans 400 0 0 0 gpio_analog_sel[1]
port 508 nsew
flabel metal3 s 675407 151640 675887 151710 0 FreeSans 400 0 0 0 gpio_dm0[1]
port 596 nsew
flabel metal3 s 675407 149800 675887 149870 0 FreeSans 400 0 0 0 gpio_dm1[1]
port 640 nsew
flabel metal3 s 675407 155964 675887 156034 0 FreeSans 400 0 0 0 gpio_dm2[1]
port 684 nsew
flabel metal3 s 675407 156608 675887 156678 0 FreeSans 400 0 0 0 gpio_holdover[1]
port 420 nsew
flabel metal3 s 675407 159644 675887 159714 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[1]
port 288 nsew
flabel metal3 s 675407 152836 675887 152906 0 FreeSans 400 0 0 0 gpio_inp_dis[1]
port 244 nsew
flabel metal3 s 675407 160288 675887 160358 0 FreeSans 400 0 0 0 gpio_oeb[1]
port 200 nsew
flabel metal3 s 675407 157160 675887 157230 0 FreeSans 400 0 0 0 gpio_out[1]
port 156 nsew
flabel metal3 s 675407 147960 675887 148030 0 FreeSans 400 0 0 0 gpio_slow_sel[1]
port 376 nsew
flabel metal3 s 675407 159000 675887 159070 0 FreeSans 400 0 0 0 gpio_vtrip_sel[1]
port 332 nsew
flabel metal3 s 675407 146120 675887 146190 0 FreeSans 400 0 0 0 gpio_in[1]
port 728 nsew
flabel metal3 s 675407 195996 675887 196066 0 FreeSans 400 0 0 0 gpio_analog_en[2]
port 463 nsew
flabel metal3 s 675407 197284 675887 197354 0 FreeSans 400 0 0 0 gpio_analog_pol[2]
port 551 nsew
flabel metal3 s 675407 200320 675887 200390 0 FreeSans 400 0 0 0 gpio_analog_sel[2]
port 507 nsew
flabel metal3 s 675407 196640 675887 196710 0 FreeSans 400 0 0 0 gpio_dm0[2]
port 595 nsew
flabel metal3 s 675407 194800 675887 194870 0 FreeSans 400 0 0 0 gpio_dm1[2]
port 639 nsew
flabel metal3 s 675407 200964 675887 201034 0 FreeSans 400 0 0 0 gpio_dm2[2]
port 683 nsew
flabel metal3 s 675407 201608 675887 201678 0 FreeSans 400 0 0 0 gpio_holdover[2]
port 419 nsew
flabel metal3 s 675407 204644 675887 204714 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[2]
port 287 nsew
flabel metal3 s 675407 197836 675887 197906 0 FreeSans 400 0 0 0 gpio_inp_dis[2]
port 243 nsew
flabel metal3 s 675407 205288 675887 205358 0 FreeSans 400 0 0 0 gpio_oeb[2]
port 199 nsew
flabel metal3 s 675407 202160 675887 202230 0 FreeSans 400 0 0 0 gpio_out[2]
port 155 nsew
flabel metal3 s 675407 192960 675887 193030 0 FreeSans 400 0 0 0 gpio_slow_sel[2]
port 375 nsew
flabel metal3 s 675407 204000 675887 204070 0 FreeSans 400 0 0 0 gpio_vtrip_sel[2]
port 331 nsew
flabel metal3 s 675407 191120 675887 191190 0 FreeSans 400 0 0 0 gpio_in[2]
port 727 nsew
flabel metal3 s 675407 241196 675887 241266 0 FreeSans 400 0 0 0 gpio_analog_en[3]
port 462 nsew
flabel metal3 s 675407 242484 675887 242554 0 FreeSans 400 0 0 0 gpio_analog_pol[3]
port 550 nsew
flabel metal3 s 675407 245520 675887 245590 0 FreeSans 400 0 0 0 gpio_analog_sel[3]
port 506 nsew
flabel metal3 s 675407 240000 675887 240070 0 FreeSans 400 0 0 0 gpio_dm1[3]
port 638 nsew
flabel metal3 s 675407 246164 675887 246234 0 FreeSans 400 0 0 0 gpio_dm2[3]
port 682 nsew
flabel metal3 s 675407 241840 675887 241910 0 FreeSans 400 0 0 0 gpio_dm0[3]
port 594 nsew
flabel metal3 s 675407 246808 675887 246878 0 FreeSans 400 0 0 0 gpio_holdover[3]
port 418 nsew
flabel metal3 s 675407 249844 675887 249914 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[3]
port 286 nsew
flabel metal3 s 675407 243036 675887 243106 0 FreeSans 400 0 0 0 gpio_inp_dis[3]
port 242 nsew
flabel metal3 s 675407 250488 675887 250558 0 FreeSans 400 0 0 0 gpio_oeb[3]
port 198 nsew
flabel metal3 s 675407 247360 675887 247430 0 FreeSans 400 0 0 0 gpio_out[3]
port 154 nsew
flabel metal3 s 675407 238160 675887 238230 0 FreeSans 400 0 0 0 gpio_slow_sel[3]
port 374 nsew
flabel metal3 s 675407 249200 675887 249270 0 FreeSans 400 0 0 0 gpio_vtrip_sel[3]
port 330 nsew
flabel metal3 s 675407 105796 675887 105866 0 FreeSans 400 0 0 0 gpio_analog_en[0]
port 465 nsew
flabel metal3 s 675407 107084 675887 107154 0 FreeSans 400 0 0 0 gpio_analog_pol[0]
port 553 nsew
flabel metal3 s 675407 110120 675887 110190 0 FreeSans 400 0 0 0 gpio_analog_sel[0]
port 509 nsew
flabel metal3 s 675407 106440 675887 106510 0 FreeSans 400 0 0 0 gpio_dm0[0]
port 597 nsew
flabel metal3 s 675407 104600 675887 104670 0 FreeSans 400 0 0 0 gpio_dm1[0]
port 641 nsew
flabel metal3 s 675407 110764 675887 110834 0 FreeSans 400 0 0 0 gpio_dm2[0]
port 685 nsew
flabel metal3 s 675407 111408 675887 111478 0 FreeSans 400 0 0 0 gpio_holdover[0]
port 421 nsew
flabel metal3 s 675407 107636 675887 107706 0 FreeSans 400 0 0 0 gpio_inp_dis[0]
port 245 nsew
flabel metal3 s 675407 115088 675887 115158 0 FreeSans 400 0 0 0 gpio_oeb[0]
port 201 nsew
flabel metal3 s 675407 111960 675887 112030 0 FreeSans 400 0 0 0 gpio_out[0]
port 157 nsew
flabel metal3 s 675407 102760 675887 102830 0 FreeSans 400 0 0 0 gpio_slow_sel[0]
port 377 nsew
flabel metal3 s 675407 100920 675887 100990 0 FreeSans 400 0 0 0 gpio_in[0]
port 729 nsew
flabel metal3 s 675407 236320 675887 236390 0 FreeSans 400 0 0 0 gpio_in[3]
port 726 nsew
rlabel metal1 s 142538 40100 142538 40100 4 xres_vss_loop
flabel metal4 s 36323 455607 37013 455799 6 FreeSans 400 0 0 0 vdda2
port 25 nsew
flabel metal4 s 28653 440800 28719 455800 6 FreeSans 400 0 0 0 vssa2
port 27 nsew
flabel metal4 s 38503 455546 39593 455800 0 FreeSans 400 0 0 0 vccd
port 20 nsew
flabel metal4 s 680587 459800 681277 459993 0 FreeSans 400 0 0 0 vdda1
port 24 nsew
flabel metal4 s 32933 455546 33623 455800 0 FreeSans 400 0 0 0 vddio
port 18 nsew
flabel metal4 s 688881 459800 688947 474800 0 FreeSans 400 0 0 0 vssa1
port 26 nsew
flabel metal4 s 0 455645 4843 456094 0 FreeSans 400 0 0 0 vssio
port 19 nsew
flabel metal5 s 187640 6598 200160 19088 0 FreeSans 16000 0 0 0 gpio[38]
port 75 nsew
flabel metal5 s 296240 6598 308760 19088 0 FreeSans 16000 0 0 0 gpio[39]
port 74 nsew
flabel metal5 s 351040 6598 363560 19088 0 FreeSans 16000 0 0 0 gpio[40]
port 73 nsew
flabel metal5 s 405840 6598 418360 19088 0 FreeSans 16000 0 0 0 gpio[41]
port 72 nsew
flabel metal5 s 460640 6598 473160 19088 0 FreeSans 16000 0 0 0 gpio[42]
port 71 nsew
flabel metal5 s 515440 6598 527960 19088 0 FreeSans 16000 0 0 0 gpio[43]
port 70 nsew
flabel metal5 s 6167 70054 19619 80934 0 FreeSans 16000 0 0 0 vccd_pad
port 5 nsew
flabel metal5 s 624222 6811 636390 18975 0 FreeSans 16000 0 0 0 vdda_pad
port 7 nsew
flabel metal5 s 6811 111610 18975 123778 0 FreeSans 16000 0 0 0 vddio_pad
port 1 nsew
flabel metal5 s 6811 871210 18975 883378 0 FreeSans 16000 0 0 0 vddio_pad2
port 2 nsew
flabel metal5 s 80222 6811 92390 18975 0 FreeSans 16000 0 0 0 vssa_pad
port 8 nsew
flabel metal5 s 243266 6167 254146 19619 0 FreeSans 16000 0 0 0 vssd_pad
port 6 nsew
flabel metal5 s 570422 6811 582590 18975 0 FreeSans 16000 0 0 0 vssio_pad
port 3 nsew
flabel metal5 s 334810 1018624 346978 1030788 0 FreeSans 16000 0 0 0 vssio_pad2
port 4 nsew
flabel metal5 s 698512 684440 711002 696960 0 FreeSans 16000 0 0 0 gpio[10]
port 103 nsew
flabel metal5 s 698512 729440 711002 741960 0 FreeSans 16000 0 0 0 gpio[11]
port 102 nsew
flabel metal5 s 698512 774440 711002 786960 0 FreeSans 16000 0 0 0 gpio[12]
port 101 nsew
flabel metal5 s 698512 863640 711002 876160 0 FreeSans 16000 0 0 0 gpio[13]
port 100 nsew
flabel metal5 s 628240 1018512 640760 1031002 0 FreeSans 16000 0 0 0 gpio[15]
port 98 nsew
flabel metal5 s 526440 1018512 538960 1031002 0 FreeSans 16000 0 0 0 gpio[16]
port 97 nsew
flabel metal5 s 475040 1018512 487560 1031002 0 FreeSans 16000 0 0 0 gpio[17]
port 96 nsew
flabel metal5 s 386040 1018512 398560 1031002 0 FreeSans 16000 0 0 0 gpio[18]
port 95 nsew
flabel metal5 s 698512 146440 711002 158960 0 FreeSans 16000 0 0 0 gpio[1]
port 112 nsew
flabel metal5 s 698512 191440 711002 203960 0 FreeSans 16000 0 0 0 gpio[2]
port 111 nsew
flabel metal5 s 698512 236640 711002 249160 0 FreeSans 16000 0 0 0 gpio[3]
port 110 nsew
flabel metal5 s 698512 281640 711002 294160 0 FreeSans 16000 0 0 0 gpio[4]
port 109 nsew
flabel metal5 s 698512 326640 711002 339160 0 FreeSans 16000 0 0 0 gpio[5]
port 108 nsew
flabel metal5 s 698512 371840 711002 384360 0 FreeSans 16000 0 0 0 gpio[6]
port 107 nsew
flabel metal5 s 698512 549040 711002 561560 0 FreeSans 16000 0 0 0 gpio[7]
port 106 nsew
flabel metal5 s 698512 594240 711002 606760 0 FreeSans 16000 0 0 0 gpio[8]
port 105 nsew
flabel metal5 s 698512 639240 711002 651760 0 FreeSans 16000 0 0 0 gpio[9]
port 104 nsew
flabel metal5 s 284240 1018512 296760 1031002 0 FreeSans 16000 0 0 0 gpio[19]
port 94 nsew
flabel metal5 s 6598 613840 19088 626360 0 FreeSans 16000 0 0 0 gpio[29]
port 84 nsew
flabel metal5 s 6598 570640 19088 583160 0 FreeSans 16000 0 0 0 gpio[30]
port 83 nsew
flabel metal5 s 6598 527440 19088 539960 0 FreeSans 16000 0 0 0 gpio[31]
port 82 nsew
flabel metal5 s 6598 399840 19088 412360 0 FreeSans 16000 0 0 0 gpio[32]
port 81 nsew
flabel metal5 s 6598 356640 19088 369160 0 FreeSans 16000 0 0 0 gpio[33]
port 80 nsew
flabel metal5 s 6598 313440 19088 325960 0 FreeSans 16000 0 0 0 gpio[34]
port 79 nsew
flabel metal5 s 6598 270240 19088 282760 0 FreeSans 16000 0 0 0 gpio[35]
port 78 nsew
flabel metal5 s 6598 227040 19088 239560 0 FreeSans 16000 0 0 0 gpio[36]
port 77 nsew
flabel metal5 s 232640 1018512 245160 1031002 0 FreeSans 16000 0 0 0 gpio[20]
port 93 nsew
flabel metal5 s 181240 1018512 193760 1031002 0 FreeSans 16000 0 0 0 gpio[21]
port 92 nsew
flabel metal5 s 129840 1018512 142360 1031002 0 FreeSans 16000 0 0 0 gpio[22]
port 91 nsew
flabel metal5 s 78440 1018512 90960 1031002 0 FreeSans 16000 0 0 0 gpio[23]
port 90 nsew
flabel metal5 s 6598 956440 19088 968960 0 FreeSans 16000 0 0 0 gpio[24]
port 89 nsew
flabel metal5 s 6598 786640 19088 799160 0 FreeSans 16000 0 0 0 gpio[25]
port 88 nsew
flabel metal5 s 6598 743440 19088 755960 0 FreeSans 16000 0 0 0 gpio[26]
port 87 nsew
flabel metal5 s 6598 700240 19088 712760 0 FreeSans 16000 0 0 0 gpio[27]
port 86 nsew
flabel metal5 s 6598 657040 19088 669560 0 FreeSans 16000 0 0 0 gpio[28]
port 85 nsew
flabel metal5 s 136713 7143 144149 18309 0 FreeSans 16000 0 0 0 resetb_pad
port 32 nsew
flabel metal5 s 697980 909666 711432 920546 0 FreeSans 16000 0 0 0 vccd1_pad
port 14 nsew
flabel metal5 s 698624 819822 710788 831990 0 FreeSans 16000 0 0 0 vdda1_pad
port 9 nsew
flabel metal5 s 698624 505222 710788 517390 0 FreeSans 16000 0 0 0 vdda1_pad2
port 10 nsew
flabel metal5 s 577010 1018624 589178 1030788 0 FreeSans 16000 0 0 0 vssa1_pad
port 11 nsew
flabel metal5 s 698624 417022 710788 429190 0 FreeSans 16000 0 0 0 vssa1_pad2
port 12 nsew
flabel metal5 s 697980 461866 711432 472746 0 FreeSans 16000 0 0 0 vssd1_pad
port 16 nsew
flabel metal5 s 6167 914054 19619 924934 0 FreeSans 16000 0 0 0 vccd2_pad
port 15 nsew
flabel metal5 s 6811 484410 18975 496578 0 FreeSans 16000 0 0 0 vdda2_pad
port 2569 nsew
flabel metal5 s 6811 829010 18975 841178 0 FreeSans 16000 0 0 0 vssa2_pad
port 13 nsew
flabel metal5 s 6167 442854 19619 453734 0 FreeSans 16000 0 0 0 vssd2_pad
port 17 nsew
rlabel metal3 s 140494 40183 140494 40183 4 xresloop
flabel metal5 s 6598 183840 19088 196360 0 FreeSans 16000 0 0 0 gpio[37]
port 76 nsew
flabel metal5 s 698512 101240 711002 113760 0 FreeSans 16000 0 0 0 gpio[0]
port 113 nsew
flabel metal3 s 41713 189894 42193 189964 0 FreeSans 400 0 0 0 gpio_inp_dis[37]
port 208 nsew
flabel metal2 187327 41713 187383 42193 0 FreeSans 400 270 0 0 gpio_in[38]
port 691 nsew
flabel metal2 189167 41713 189223 42193 0 FreeSans 400 270 0 0 gpio_slow_sel[38]
port 339 nsew
flabel metal2 191007 41713 191063 42193 0 FreeSans 400 270 0 0 gpio_dm0[38]
port 559 nsew
flabel metal2 192847 41713 192903 42193 0 FreeSans 400 270 0 0 gpio_dm1[38]
port 603 nsew
flabel metal2 193491 41713 193547 42193 0 FreeSans 400 270 0 0 gpio_analog_pol[38]
port 515 nsew
flabel metal2 192203 41713 192259 42193 0 FreeSans 400 270 0 0 gpio_analog_en[38]
port 427 nsew
flabel metal2 194043 41713 194099 42193 0 FreeSans 400 270 0 0 gpio_inp_dis[38]
port 207 nsew
flabel metal2 196527 41713 196583 42193 0 FreeSans 400 270 0 0 gpio_analog_sel[38]
port 471 nsew
flabel metal2 197171 41713 197227 42193 0 FreeSans 400 270 0 0 gpio_dm2[38]
port 647 nsew
flabel metal2 197815 41713 197871 42193 0 FreeSans 400 270 0 0 gpio_holdover[38]
port 383 nsew
flabel metal2 198367 41713 198423 42193 0 FreeSans 400 270 0 0 gpio_out[38]
port 119 nsew
flabel metal2 200207 41713 200263 42193 0 FreeSans 400 270 0 0 gpio_vtrip_sel[38]
port 295 nsew
flabel metal2 200851 41713 200907 42193 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[38]
port 251 nsew
flabel metal2 201495 41713 201551 42193 0 FreeSans 400 270 0 0 gpio_oeb[38]
port 163 nsew
flabel metal2 295927 41713 295983 42193 0 FreeSans 400 270 0 0 gpio_in[39]
port 690 nsew
flabel metal2 297767 41713 297823 42193 0 FreeSans 400 270 0 0 gpio_slow_sel[39]
port 338 nsew
flabel metal2 299607 41713 299663 42193 0 FreeSans 400 270 0 0 gpio_dm1[39]
port 602 nsew
flabel metal2 301447 41713 301503 42193 0 FreeSans 400 270 0 0 gpio_dm0[39]
port 558 nsew
flabel metal2 302091 41713 302147 42193 0 FreeSans 400 270 0 0 gpio_analog_pol[39]
port 514 nsew
flabel metal2 300803 41713 300859 42193 0 FreeSans 400 270 0 0 gpio_analog_en[39]
port 426 nsew
flabel metal2 302643 41713 302699 42193 0 FreeSans 400 270 0 0 gpio_inp_dis[39]
port 206 nsew
flabel metal2 305127 41713 305183 42193 0 FreeSans 400 270 0 0 gpio_analog_sel[39]
port 470 nsew
flabel metal2 305771 41713 305827 42193 0 FreeSans 400 270 0 0 gpio_dm2[39]
port 646 nsew
flabel metal2 306415 41713 306471 42193 0 FreeSans 400 270 0 0 gpio_holdover[39]
port 382 nsew
flabel metal2 306967 41713 307023 42193 0 FreeSans 400 270 0 0 gpio_out[39]
port 118 nsew
flabel metal2 308807 41713 308863 42193 0 FreeSans 400 270 0 0 gpio_vtrip_sel[39]
port 294 nsew
flabel metal2 309451 41713 309507 42193 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[39]
port 250 nsew
flabel metal2 310095 41713 310151 42193 0 FreeSans 400 270 0 0 gpio_oeb[39]
port 162 nsew
flabel metal2 350727 41713 350783 42193 0 FreeSans 400 270 0 0 gpio_in[40]
port 689 nsew
flabel metal2 352567 41713 352623 42193 0 FreeSans 400 270 0 0 gpio_slow_sel[40]
port 337 nsew
flabel metal2 354407 41713 354463 42193 0 FreeSans 400 270 0 0 gpio_dm1[40]
port 601 nsew
flabel metal2 356247 41713 356303 42193 0 FreeSans 400 270 0 0 gpio_dm0[40]
port 557 nsew
flabel metal2 356891 41713 356947 42193 0 FreeSans 400 270 0 0 gpio_analog_pol[40]
port 513 nsew
flabel metal2 355603 41713 355659 42193 0 FreeSans 400 270 0 0 gpio_analog_en[40]
port 425 nsew
flabel metal2 357443 41713 357499 42193 0 FreeSans 400 270 0 0 gpio_inp_dis[40]
port 205 nsew
flabel metal2 359927 41713 359983 42193 0 FreeSans 400 270 0 0 gpio_analog_sel[40]
port 469 nsew
flabel metal2 360571 41713 360627 42193 0 FreeSans 400 270 0 0 gpio_dm2[40]
port 645 nsew
flabel metal2 361215 41713 361271 42193 0 FreeSans 400 270 0 0 gpio_holdover[40]
port 381 nsew
flabel metal2 361767 41713 361823 42193 0 FreeSans 400 270 0 0 gpio_out[40]
port 117 nsew
flabel metal2 363607 41713 363663 42193 0 FreeSans 400 270 0 0 gpio_vtrip_sel[40]
port 293 nsew
flabel metal2 364251 41713 364307 42193 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[40]
port 249 nsew
flabel metal2 364895 41713 364951 42193 0 FreeSans 400 270 0 0 gpio_oeb[40]
port 161 nsew
flabel metal2 405527 41713 405583 42193 0 FreeSans 400 270 0 0 gpio_in[41]
port 688 nsew
flabel metal2 407367 41713 407423 42193 0 FreeSans 400 270 0 0 gpio_slow_sel[41]
port 336 nsew
flabel metal2 409207 41713 409263 42193 0 FreeSans 400 270 0 0 gpio_dm1[41]
port 600 nsew
flabel metal2 411047 41713 411103 42193 0 FreeSans 400 270 0 0 gpio_dm0[41]
port 556 nsew
flabel metal2 411691 41713 411747 42193 0 FreeSans 400 270 0 0 gpio_analog_pol[41]
port 512 nsew
flabel metal2 410403 41713 410459 42193 0 FreeSans 400 270 0 0 gpio_analog_en[41]
port 424 nsew
flabel metal2 412243 41713 412299 42193 0 FreeSans 400 270 0 0 gpio_inp_dis[41]
port 204 nsew
flabel metal2 414727 41713 414783 42193 0 FreeSans 400 270 0 0 gpio_analog_sel[41]
port 468 nsew
flabel metal2 415371 41713 415427 42193 0 FreeSans 400 270 0 0 gpio_dm2[41]
port 644 nsew
flabel metal2 416015 41713 416071 42193 0 FreeSans 400 270 0 0 gpio_holdover[41]
port 380 nsew
flabel metal2 416567 41713 416623 42193 0 FreeSans 400 270 0 0 gpio_out[41]
port 116 nsew
flabel metal2 418407 41713 418463 42193 0 FreeSans 400 270 0 0 gpio_vtrip_sel[41]
port 292 nsew
flabel metal2 419051 41713 419107 42193 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[41]
port 248 nsew
flabel metal2 419695 41713 419751 42193 0 FreeSans 400 270 0 0 gpio_oeb[41]
port 160 nsew
flabel metal2 460327 41713 460383 42193 0 FreeSans 400 270 0 0 gpio_in[42]
port 687 nsew
flabel metal2 462167 41713 462223 42193 0 FreeSans 400 270 0 0 gpio_slow_sel[42]
port 335 nsew
flabel metal2 464007 41713 464063 42193 0 FreeSans 400 270 0 0 gpio_dm1[42]
port 599 nsew
flabel metal2 465847 41713 465903 42193 0 FreeSans 400 270 0 0 gpio_dm0[42]
port 555 nsew
flabel metal2 466491 41713 466547 42193 0 FreeSans 400 270 0 0 gpio_analog_pol[42]
port 511 nsew
flabel metal2 465203 41713 465259 42193 0 FreeSans 400 270 0 0 gpio_analog_en[42]
port 423 nsew
flabel metal2 467043 41713 467099 42193 0 FreeSans 400 270 0 0 gpio_inp_dis[42]
port 203 nsew
flabel metal2 469527 41713 469583 42193 0 FreeSans 400 270 0 0 gpio_analog_sel[42]
port 467 nsew
flabel metal2 470171 41713 470227 42193 0 FreeSans 400 270 0 0 gpio_dm2[42]
port 643 nsew
flabel metal2 470815 41713 470871 42193 0 FreeSans 400 270 0 0 gpio_holdover[42]
port 379 nsew
flabel metal2 471367 41713 471423 42193 0 FreeSans 400 270 0 0 gpio_out[42]
port 115 nsew
flabel metal2 473207 41713 473263 42193 0 FreeSans 400 270 0 0 gpio_vtrip_sel[42]
port 291 nsew
flabel metal2 473851 41713 473907 42193 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[42]
port 247 nsew
flabel metal2 474495 41713 474551 42193 0 FreeSans 400 270 0 0 gpio_oeb[42]
port 159 nsew
flabel metal2 515127 41713 515183 42193 0 FreeSans 400 270 0 0 gpio_in[43]
port 686 nsew
flabel metal2 516967 41713 517023 42193 0 FreeSans 400 270 0 0 gpio_slow_sel[43]
port 334 nsew
flabel metal2 518807 41713 518863 42193 0 FreeSans 400 270 0 0 gpio_dm1[43]
port 598 nsew
flabel metal2 520647 41713 520703 42193 0 FreeSans 400 270 0 0 gpio_dm0[43]
port 554 nsew
flabel metal2 521291 41713 521347 42193 0 FreeSans 400 270 0 0 gpio_analog_pol[43]
port 510 nsew
flabel metal2 520003 41713 520059 42193 0 FreeSans 400 270 0 0 gpio_analog_en[43]
port 422 nsew
flabel metal2 521843 41713 521899 42193 0 FreeSans 400 270 0 0 gpio_inp_dis[43]
port 202 nsew
flabel metal2 524327 41713 524383 42193 0 FreeSans 400 270 0 0 gpio_analog_sel[43]
port 466 nsew
flabel metal2 524971 41713 525027 42193 0 FreeSans 400 270 0 0 gpio_dm2[43]
port 642 nsew
flabel metal2 525615 41713 525671 42193 0 FreeSans 400 270 0 0 gpio_holdover[43]
port 378 nsew
flabel metal2 526167 41713 526223 42193 0 FreeSans 400 270 0 0 gpio_out[43]
port 114 nsew
flabel metal2 528007 41713 528063 42193 0 FreeSans 400 270 0 0 gpio_vtrip_sel[43]
port 290 nsew
flabel metal2 528651 41713 528707 42193 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[43]
port 246 nsew
flabel metal2 529295 41713 529351 42193 0 FreeSans 400 270 0 0 gpio_oeb[43]
port 158 nsew
flabel metal3 675407 103404 675887 103474 0 FreeSans 400 0 0 0 analog_io[0]
port 905 nsew
flabel metal3 675407 105244 675887 105314 0 FreeSans 400 0 0 0 analog_noesd_io[0]
port 949 nsew
flabel metal3 675407 150444 675887 150514 0 FreeSans 400 0 0 0 analog_noesd_io[1]
port 948 nsew
flabel metal3 675407 148604 675887 148674 0 FreeSans 400 0 0 0 analog_io[1]
port 904 nsew
flabel metal3 675407 115640 675887 115710 0 FreeSans 400 0 0 0 gpio_in_h[0]
port 773 nsew
flabel metal3 675407 160840 675887 160910 0 FreeSans 400 0 0 0 gpio_in_h[1]
port 772 nsew
flabel metal3 675407 193604 675887 193674 0 FreeSans 400 0 0 0 analog_io[2]
port 903 nsew
flabel metal3 675407 195444 675887 195514 0 FreeSans 400 0 0 0 analog_noesd_io[2]
port 947 nsew
flabel metal3 675407 205840 675887 205910 0 FreeSans 400 0 0 0 gpio_in_h[2]
port 771 nsew
flabel metal3 675407 238804 675887 238874 0 FreeSans 400 0 0 0 analog_io[3]
port 902 nsew
flabel metal3 675407 251040 675887 251110 0 FreeSans 400 0 0 0 gpio_in_h[3]
port 770 nsew
flabel metal3 675407 283804 675887 283874 0 FreeSans 400 0 0 0 analog_io[4]
port 901 nsew
flabel metal3 675407 285644 675887 285714 0 FreeSans 400 0 0 0 analog_noesd_io[4]
port 945 nsew
flabel metal3 675407 296040 675887 296110 0 FreeSans 400 0 0 0 gpio_in_h[4]
port 769 nsew
flabel metal3 675407 328804 675887 328874 0 FreeSans 400 0 0 0 analog_io[5]
port 900 nsew
flabel metal3 675407 330644 675887 330714 0 FreeSans 400 0 0 0 analog_noesd_io[5]
port 944 nsew
flabel metal3 675407 341040 675887 341110 0 FreeSans 400 0 0 0 gpio_in_h[5]
port 768 nsew
flabel metal3 675407 374004 675887 374074 0 FreeSans 400 0 0 0 analog_io[6]
port 899 nsew
flabel metal3 675407 375844 675887 375914 0 FreeSans 400 0 0 0 analog_noesd_io[6]
port 943 nsew
flabel metal3 675407 386240 675887 386310 0 FreeSans 400 0 0 0 gpio_in_h[6]
port 767 nsew
flabel metal3 s 675407 551204 675887 551274 0 FreeSans 400 0 0 0 analog_io[7]
port 898 nsew
flabel metal3 s 675407 553044 675887 553114 0 FreeSans 400 0 0 0 analog_noesd_io[7]
port 942 nsew
flabel metal3 s 675407 563440 675887 563510 0 FreeSans 400 0 0 0 gpio_in_h[7]
port 766 nsew
flabel metal3 s 675407 596404 675887 596474 0 FreeSans 400 0 0 0 analog_io[8]
port 897 nsew
flabel metal3 s 675407 598244 675887 598314 0 FreeSans 400 0 0 0 analog_noesd_io[8]
port 941 nsew
flabel metal3 s 675407 608640 675887 608710 0 FreeSans 400 0 0 0 gpio_in_h[8]
port 765 nsew
flabel metal3 s 675407 641404 675887 641474 0 FreeSans 400 0 0 0 analog_io[9]
port 896 nsew
flabel metal3 s 675407 643244 675887 643314 0 FreeSans 400 0 0 0 analog_noesd_io[9]
port 940 nsew
flabel metal3 s 675407 653640 675887 653710 0 FreeSans 400 0 0 0 gpio_in_h[9]
port 764 nsew
flabel metal3 s 675407 686604 675887 686674 0 FreeSans 400 0 0 0 analog_io[10]
port 895 nsew
flabel metal3 s 675407 688444 675887 688514 0 FreeSans 400 0 0 0 analog_noesd_io[10]
port 939 nsew
flabel metal3 s 675407 698840 675887 698910 0 FreeSans 400 0 0 0 gpio_in_h[10]
port 763 nsew
flabel metal3 s 675407 731604 675887 731674 0 FreeSans 400 0 0 0 analog_io[11]
port 894 nsew
flabel metal3 s 675407 733444 675887 733514 0 FreeSans 400 0 0 0 analog_noesd_io[11]
port 938 nsew
flabel metal3 s 675407 743840 675887 743910 0 FreeSans 400 0 0 0 gpio_in_h[11]
port 762 nsew
flabel metal3 s 675407 788840 675887 788910 0 FreeSans 400 0 0 0 gpio_in_h[12]
port 761 nsew
flabel metal3 s 675407 878040 675887 878110 0 FreeSans 400 0 0 0 gpio_in_h[13]
port 760 nsew
flabel metal3 s 675407 967240 675887 967310 0 FreeSans 400 0 0 0 gpio_in_h[14]
port 759 nsew
flabel metal2 s 626297 995407 626353 995887 0 FreeSans 400 90 0 0 gpio_in_h[15]
port 758 nsew
flabel metal2 s 524497 995407 524553 995887 0 FreeSans 400 90 0 0 gpio_in_h[16]
port 757 nsew
flabel metal2 s 473097 995407 473153 995887 0 FreeSans 400 90 0 0 gpio_in_h[17]
port 756 nsew
flabel metal2 s 384097 995407 384153 995887 0 FreeSans 400 90 0 0 gpio_in_h[18]
port 755 nsew
flabel metal2 s 282297 995407 282353 995887 0 FreeSans 400 90 0 0 gpio_in_h[19]
port 754 nsew
flabel metal2 s 230697 995407 230753 995887 0 FreeSans 400 90 0 0 gpio_in_h[20]
port 753 nsew
flabel metal2 s 179297 995407 179353 995887 0 FreeSans 400 90 0 0 gpio_in_h[21]
port 752 nsew
flabel metal2 s 127897 995407 127953 995887 0 FreeSans 400 90 0 0 gpio_in_h[22]
port 751 nsew
flabel metal2 s 76497 995407 76553 995887 0 FreeSans 400 90 0 0 gpio_in_h[23]
port 750 nsew
flabel metal3 s 41713 954490 42193 954560 0 FreeSans 400 0 0 0 gpio_in_h[24]
port 749 nsew
flabel metal3 s 41713 784690 42193 784760 0 FreeSans 400 0 0 0 gpio_in_h[25]
port 748 nsew
flabel metal3 s 41713 741490 42193 741560 0 FreeSans 400 0 0 0 gpio_in_h[26]
port 747 nsew
flabel metal3 s 41713 698290 42193 698360 0 FreeSans 400 0 0 0 gpio_in_h[27]
port 746 nsew
flabel metal3 s 41713 655090 42193 655160 0 FreeSans 400 0 0 0 gpio_in_h[28]
port 745 nsew
flabel metal3 s 41713 611890 42193 611960 0 FreeSans 400 0 0 0 gpio_in_h[29]
port 744 nsew
flabel metal3 s 41713 568690 42193 568760 0 FreeSans 400 0 0 0 gpio_in_h[30]
port 743 nsew
flabel metal3 s 41713 525490 42193 525560 0 FreeSans 400 0 0 0 gpio_in_h[31]
port 742 nsew
flabel metal3 s 41713 397890 42193 397960 0 FreeSans 400 0 0 0 gpio_in_h[32]
port 741 nsew
flabel metal3 s 41713 354690 42193 354760 0 FreeSans 400 0 0 0 gpio_in_h[33]
port 740 nsew
flabel metal3 s 41713 311490 42193 311560 0 FreeSans 400 0 0 0 gpio_in_h[34]
port 739 nsew
flabel metal3 s 41713 268290 42193 268360 0 FreeSans 400 0 0 0 gpio_in_h[35]
port 738 nsew
flabel metal3 s 41713 225090 42193 225160 0 FreeSans 400 0 0 0 gpio_in_h[36]
port 737 nsew
flabel metal3 s 41713 181890 42193 181960 0 FreeSans 400 0 0 0 gpio_in_h[37]
port 736 nsew
flabel metal2 s 202047 41713 202103 42193 0 FreeSans 400 90 0 0 gpio_in_h[38]
port 735 nsew
flabel metal2 s 310647 41713 310703 42193 0 FreeSans 400 90 0 0 gpio_in_h[39]
port 734 nsew
flabel metal2 s 365447 41713 365503 42193 0 FreeSans 400 90 0 0 gpio_in_h[40]
port 733 nsew
flabel metal2 s 420247 41713 420303 42193 0 FreeSans 400 90 0 0 gpio_in_h[41]
port 732 nsew
flabel metal2 s 475047 41713 475103 42193 0 FreeSans 400 90 0 0 gpio_in_h[42]
port 731 nsew
flabel metal2 s 529847 41713 529903 42193 0 FreeSans 400 90 0 0 gpio_in_h[43]
port 730 nsew
flabel metal3 s 675407 776604 675887 776674 0 FreeSans 400 0 0 0 analog_io[12]
port 893 nsew
flabel metal3 s 675407 865804 675887 865874 0 FreeSans 400 0 0 0 analog_io[13]
port 892 nsew
flabel metal3 s 675407 955004 675887 955074 0 FreeSans 400 0 0 0 analog_io[14]
port 891 nsew
flabel metal2 s 638533 995407 638589 995887 0 FreeSans 400 90 0 0 analog_io[15]
port 890 nsew
flabel metal2 s 536733 995407 536789 995887 0 FreeSans 400 90 0 0 analog_io[16]
port 889 nsew
flabel metal2 s 485333 995407 485389 995887 0 FreeSans 400 90 0 0 analog_io[17]
port 888 nsew
flabel metal2 s 396333 995407 396389 995887 0 FreeSans 400 90 0 0 analog_io[18]
port 887 nsew
flabel metal2 s 294533 995407 294589 995887 0 FreeSans 400 90 0 0 analog_io[19]
port 886 nsew
flabel metal2 s 242933 995407 242989 995887 0 FreeSans 400 90 0 0 analog_io[20]
port 885 nsew
flabel metal2 s 191533 995407 191589 995887 0 FreeSans 400 90 0 0 analog_io[21]
port 884 nsew
flabel metal2 s 140133 995407 140189 995887 0 FreeSans 400 90 0 0 analog_io[22]
port 883 nsew
flabel metal2 s 88733 995407 88789 995887 0 FreeSans 400 90 0 0 analog_io[23]
port 882 nsew
flabel metal3 s 41713 966726 42193 966796 0 FreeSans 400 0 0 0 analog_io[24]
port 881 nsew
flabel metal3 s 41713 796926 42193 796996 0 FreeSans 400 0 0 0 analog_io[25]
port 880 nsew
flabel metal3 s 41713 753726 42193 753796 0 FreeSans 400 0 0 0 analog_io[26]
port 879 nsew
flabel metal3 s 41713 710526 42193 710596 0 FreeSans 400 0 0 0 analog_io[27]
port 878 nsew
flabel metal3 s 41713 667326 42193 667396 0 FreeSans 400 0 0 0 analog_io[28]
port 877 nsew
flabel metal3 s 41713 624126 42193 624196 0 FreeSans 400 0 0 0 analog_io[29]
port 876 nsew
flabel metal3 s 41713 580926 42193 580996 0 FreeSans 400 0 0 0 analog_io[30]
port 875 nsew
flabel metal3 s 41713 537726 42193 537796 0 FreeSans 400 0 0 0 analog_io[31]
port 874 nsew
flabel metal3 s 41713 410126 42193 410196 0 FreeSans 400 0 0 0 analog_io[32]
port 873 nsew
flabel metal3 s 41713 366926 42193 366996 0 FreeSans 400 0 0 0 analog_io[33]
port 872 nsew
flabel metal3 s 41713 323726 42193 323796 0 FreeSans 400 0 0 0 analog_io[34]
port 871 nsew
flabel metal3 s 41713 280526 42193 280596 0 FreeSans 400 0 0 0 analog_io[35]
port 870 nsew
flabel metal3 s 41713 237326 42193 237396 0 FreeSans 400 0 0 0 analog_io[36]
port 869 nsew
flabel metal3 s 41713 194126 42193 194196 0 FreeSans 400 0 0 0 analog_io[37]
port 868 nsew
flabel metal2 s 189811 41713 189867 42193 0 FreeSans 400 90 0 0 analog_io[38]
port 867 nsew
flabel metal2 s 298411 41713 298467 42193 0 FreeSans 400 90 0 0 analog_io[39]
port 866 nsew
flabel metal2 s 353211 41713 353267 42193 0 FreeSans 400 90 0 0 analog_io[40]
port 865 nsew
flabel metal2 s 408011 41713 408067 42193 0 FreeSans 400 90 0 0 analog_io[41]
port 864 nsew
flabel metal2 s 462811 41713 462867 42193 0 FreeSans 400 90 0 0 analog_io[42]
port 863 nsew
flabel metal2 s 517611 41713 517667 42193 0 FreeSans 400 90 0 0 analog_io[43]
port 862 nsew
flabel metal3 s 675407 778444 675887 778514 0 FreeSans 400 0 0 0 analog_noesd_io[12]
port 937 nsew
flabel metal3 s 675407 867644 675887 867714 0 FreeSans 400 0 0 0 analog_noesd_io[13]
port 936 nsew
flabel metal3 s 675407 956844 675887 956914 0 FreeSans 400 0 0 0 analog_noesd_io[14]
port 935 nsew
flabel metal2 s 636693 995407 636749 995887 0 FreeSans 400 90 0 0 analog_noesd_io[15]
port 934 nsew
flabel metal2 s 534893 995407 534949 995887 0 FreeSans 400 90 0 0 analog_noesd_io[16]
port 933 nsew
flabel metal2 s 483493 995407 483549 995887 0 FreeSans 400 90 0 0 analog_noesd_io[17]
port 932 nsew
flabel metal2 s 394493 995407 394549 995887 0 FreeSans 400 90 0 0 analog_noesd_io[18]
port 931 nsew
flabel metal2 s 292693 995407 292749 995887 0 FreeSans 400 90 0 0 analog_noesd_io[19]
port 930 nsew
flabel metal2 s 241093 995407 241149 995887 0 FreeSans 400 90 0 0 analog_noesd_io[20]
port 929 nsew
flabel metal2 s 189693 995407 189749 995887 0 FreeSans 400 90 0 0 analog_noesd_io[21]
port 928 nsew
flabel metal2 s 138293 995407 138349 995887 0 FreeSans 400 90 0 0 analog_noesd_io[22]
port 927 nsew
flabel metal2 s 86893 995407 86949 995887 0 FreeSans 400 90 0 0 analog_noesd_io[23]
port 926 nsew
flabel metal3 s 41713 964886 42193 964956 0 FreeSans 400 0 0 0 analog_noesd_io[24]
port 925 nsew
flabel metal3 s 41713 795086 42193 795156 0 FreeSans 400 0 0 0 analog_noesd_io[25]
port 924 nsew
flabel metal3 s 41713 751886 42193 751956 0 FreeSans 400 0 0 0 analog_noesd_io[26]
port 923 nsew
flabel metal3 s 41713 708686 42193 708756 0 FreeSans 400 0 0 0 analog_noesd_io[27]
port 922 nsew
flabel metal3 s 41713 665486 42193 665556 0 FreeSans 400 0 0 0 analog_noesd_io[28]
port 921 nsew
flabel metal3 s 41713 622286 42193 622356 0 FreeSans 400 0 0 0 analog_noesd_io[29]
port 920 nsew
flabel metal3 s 41713 579086 42193 579156 0 FreeSans 400 0 0 0 analog_noesd_io[30]
port 919 nsew
flabel metal3 s 41713 535886 42193 535956 0 FreeSans 400 0 0 0 analog_noesd_io[31]
port 918 nsew
flabel metal3 s 41713 408286 42193 408356 0 FreeSans 400 0 0 0 analog_noesd_io[32]
port 917 nsew
flabel metal3 s 41713 365086 42193 365156 0 FreeSans 400 0 0 0 analog_noesd_io[33]
port 916 nsew
flabel metal3 s 41713 321886 42193 321956 0 FreeSans 400 0 0 0 analog_noesd_io[34]
port 915 nsew
flabel metal3 s 41713 278686 42193 278756 0 FreeSans 400 0 0 0 analog_noesd_io[35]
port 914 nsew
flabel metal3 s 41713 235486 42193 235556 0 FreeSans 400 0 0 0 analog_noesd_io[36]
port 913 nsew
flabel metal3 s 41713 192286 42193 192356 0 FreeSans 400 0 0 0 analog_noesd_io[37]
port 912 nsew
flabel metal2 s 191651 41713 191707 42193 0 FreeSans 400 90 0 0 analog_noesd_io[38]
port 911 nsew
flabel metal2 s 300251 41713 300307 42193 0 FreeSans 400 90 0 0 analog_noesd_io[39]
port 910 nsew
flabel metal2 s 355051 41713 355107 42193 0 FreeSans 400 90 0 0 analog_noesd_io[40]
port 909 nsew
flabel metal2 s 409851 41713 409907 42193 0 FreeSans 400 90 0 0 analog_noesd_io[41]
port 908 nsew
flabel metal2 s 464651 41713 464707 42193 0 FreeSans 400 90 0 0 analog_noesd_io[42]
port 907 nsew
flabel metal2 s 519451 41713 519507 42193 0 FreeSans 400 90 0 0 analog_noesd_io[43]
port 906 nsew
flabel metal3 41873 948781 42193 948841 0 FreeSans 400 0 0 0 gpio_loopback_one[24]
port 837 nsew
flabel metal3 41873 778781 42193 778841 0 FreeSans 400 0 0 0 gpio_loopback_one[25]
port 836 nsew
flabel metal3 41873 735781 42193 735841 0 FreeSans 400 0 0 0 gpio_loopback_one[26]
port 835 nsew
flabel metal3 41873 692781 42193 692841 0 FreeSans 400 0 0 0 gpio_loopback_one[27]
port 834 nsew
flabel metal3 41873 649781 42193 649841 0 FreeSans 400 0 0 0 gpio_loopback_one[28]
port 833 nsew
flabel metal3 41873 606781 42193 606841 0 FreeSans 400 0 0 0 gpio_loopback_one[29]
port 832 nsew
flabel metal3 41873 563781 42193 563841 0 FreeSans 400 0 0 0 gpio_loopback_one[30]
port 831 nsew
flabel metal3 41873 520781 42193 520841 0 FreeSans 400 0 0 0 gpio_loopback_one[31]
port 830 nsew
flabel metal3 41873 391781 42193 391841 0 FreeSans 400 0 0 0 gpio_loopback_one[32]
port 829 nsew
flabel metal3 41873 348781 42193 348841 0 FreeSans 400 0 0 0 gpio_loopback_one[33]
port 828 nsew
flabel metal3 41873 305781 42193 305841 0 FreeSans 400 0 0 0 gpio_loopback_one[34]
port 827 nsew
flabel metal3 41873 262781 42193 262841 0 FreeSans 400 0 0 0 gpio_loopback_one[35]
port 826 nsew
flabel metal3 41873 219781 42193 219841 0 FreeSans 400 0 0 0 gpio_loopback_one[36]
port 825 nsew
flabel metal3 41873 176781 42193 176841 0 FreeSans 400 0 0 0 gpio_loopback_one[37]
port 824 nsew
flabel metal2 s 530517 41877 530569 42193 0 FreeSans 400 90 0 0 gpio_loopback_one[43]
port 818 nsew
flabel metal2 s 534772 41877 534824 42193 0 FreeSans 400 90 0 0 gpio_loopback_zero[43]
port 774 nsew
flabel metal2 s 475717 41877 475769 42193 0 FreeSans 400 90 0 0 gpio_loopback_one[42]
port 819 nsew
flabel metal2 s 479915 41877 479967 42193 0 FreeSans 400 90 0 0 gpio_loopback_zero[42]
port 775 nsew
flabel metal2 s 420917 41877 420969 42193 0 FreeSans 400 90 0 0 gpio_loopback_one[41]
port 820 nsew
flabel metal2 s 425115 41877 425167 42193 0 FreeSans 400 90 0 0 gpio_loopback_zero[41]
port 776 nsew
flabel metal2 s 366117 41877 366169 42193 0 FreeSans 400 90 0 0 gpio_loopback_one[40]
port 821 nsew
flabel metal2 s 370302 41855 370354 42171 0 FreeSans 400 90 0 0 gpio_loopback_zero[40]
port 777 nsew
flabel metal2 s 311317 41877 311369 42193 0 FreeSans 400 90 0 0 gpio_loopback_one[39]
port 822 nsew
flabel metal2 s 315497 41877 315549 42193 0 FreeSans 400 90 0 0 gpio_loopback_zero[39]
port 778 nsew
flabel metal2 s 202717 41877 202769 42193 0 FreeSans 400 90 0 0 gpio_loopback_one[38]
port 823 nsew
flabel metal2 s 205928 41878 205980 42194 0 FreeSans 400 90 0 0 gpio_loopback_zero[38]
port 779 nsew
flabel metal2 s 152301 42021 152357 42193 0 FreeSans 400 90 0 0 resetb_l
port 37 nsew
flabel metal2 s 141708 42047 141774 42193 0 FreeSans 400 90 0 0 resetb_h
port 36 nsew
flabel metal3 41854 95509 42193 95579 0 FreeSans 400 0 0 0 por_l
port 35 nsew
flabel metal3 41854 95732 42193 95802 0 FreeSans 400 0 0 0 porb_l
port 34 nsew
flabel metal2 s 647219 41877 647271 42193 0 FreeSans 400 90 0 0 mask_rev[0]
port 69 nsew
flabel metal3 41854 95284 42193 95354 0 FreeSans 400 0 0 0 porb_h
port 33 nsew
flabel metal2 620435 995407 620496 995727 0 FreeSans 400 90 0 0 gpio_loopback_one[15]
port 846 nsew
flabel metal2 521035 995407 521096 995727 0 FreeSans 400 90 0 0 gpio_loopback_one[16]
port 845 nsew
flabel metal2 469835 995407 469896 995727 0 FreeSans 400 90 0 0 gpio_loopback_one[17]
port 844 nsew
flabel metal2 380835 995407 380896 995727 0 FreeSans 400 90 0 0 gpio_loopback_one[18]
port 843 nsew
flabel metal2 276435 995407 276496 995727 0 FreeSans 400 90 0 0 gpio_loopback_one[19]
port 842 nsew
flabel metal2 225235 995407 225296 995727 0 FreeSans 400 90 0 0 gpio_loopback_one[20]
port 841 nsew
flabel metal2 174035 995407 174096 995727 0 FreeSans 400 90 0 0 gpio_loopback_one[21]
port 840 nsew
flabel metal2 122835 995407 122896 995727 0 FreeSans 400 90 0 0 gpio_loopback_one[22]
port 839 nsew
flabel metal2 71635 995407 71696 995727 0 FreeSans 400 90 0 0 gpio_loopback_one[23]
port 838 nsew
flabel metal3 675407 969142 675727 969204 0 FreeSans 400 0 0 0 gpio_loopback_one[14]
port 847 nsew
flabel metal3 675407 879142 675727 879204 0 FreeSans 400 0 0 0 gpio_loopback_one[13]
port 848 nsew
flabel metal3 675407 790142 675727 790204 0 FreeSans 400 0 0 0 gpio_loopback_one[12]
port 849 nsew
flabel metal3 675407 745142 675727 745204 0 FreeSans 400 0 0 0 gpio_loopback_one[11]
port 850 nsew
flabel metal3 675407 700142 675727 700204 0 FreeSans 400 0 0 0 gpio_loopback_one[10]
port 851 nsew
flabel metal3 675407 655142 675727 655204 0 FreeSans 400 0 0 0 gpio_loopback_one[9]
port 852 nsew
flabel metal3 675407 610142 675727 610204 0 FreeSans 400 0 0 0 gpio_loopback_one[8]
port 853 nsew
flabel metal3 675407 565142 675727 565204 0 FreeSans 400 0 0 0 gpio_loopback_one[7]
port 854 nsew
flabel metal3 675407 388142 675727 388204 0 FreeSans 400 0 0 0 gpio_loopback_one[6]
port 855 nsew
flabel metal3 675407 343142 675727 343204 0 FreeSans 400 0 0 0 gpio_loopback_one[5]
port 856 nsew
flabel metal3 675407 298142 675727 298204 0 FreeSans 400 0 0 0 gpio_loopback_one[4]
port 857 nsew
flabel metal3 675407 253142 675727 253204 0 FreeSans 400 0 0 0 gpio_loopback_one[3]
port 858 nsew
flabel metal3 675407 208142 675727 208204 0 FreeSans 400 0 0 0 gpio_loopback_one[2]
port 859 nsew
flabel metal3 675407 163142 675727 163204 0 FreeSans 400 0 0 0 gpio_loopback_one[1]
port 860 nsew
flabel metal3 675407 118142 675727 118204 0 FreeSans 400 0 0 0 gpio_loopback_one[0]
port 861 nsew
flabel metal3 632921 41693 637701 42193 0 FreeSans 3200 0 0 0 vdda
port 22 nsew
flabel metal3 622942 41693 627722 42193 0 FreeSans 3200 0 0 0 vdda
port 22 nsew
flabel metal3 569142 41693 573922 42193 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 579121 41693 583901 42193 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 241420 41693 246049 42193 0 FreeSans 3200 0 0 0 vssd
port 21 nsew
flabel metal3 251300 41693 256100 42193 0 FreeSans 3200 0 0 0 vssd
port 21 nsew
flabel metal3 78942 41693 83722 42193 0 FreeSans 3200 0 0 0 vssa
port 23 nsew
flabel metal3 88921 41694 93701 42194 0 FreeSans 3200 0 0 0 vssa
port 23 nsew
flabel metal3 41693 68100 42193 72900 0 FreeSans 3200 90 0 0 vccd
port 20 nsew
flabel metal3 41693 78151 42193 82940 0 FreeSans 3200 90 0 0 vccd
port 20 nsew
flabel metal3 41693 110299 42193 115079 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 41693 120278 42193 125058 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 41693 440900 42193 445700 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 41693 450951 42193 455740 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 41693 446000 42193 450651 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 41693 483099 42193 487879 0 FreeSans 3200 90 0 0 vdda2
port 25 nsew
flabel metal3 41693 493078 42193 497858 0 FreeSans 3200 90 0 0 vdda2
port 25 nsew
flabel metal3 41693 827699 42193 832479 0 FreeSans 3200 90 0 0 vssa2
port 27 nsew
flabel metal3 41693 837678 42193 842458 0 FreeSans 3200 90 0 0 vssa2
port 27 nsew
flabel metal3 41693 869899 42193 874679 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 41693 879878 42193 884658 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 41693 912100 42193 916900 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 41693 922151 42193 926940 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 41693 917190 42193 921852 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 333499 995407 338279 995907 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 343478 995407 348258 995907 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 s 575699 995407 580479 995907 0 FreeSans 3200 0 0 0 vssa1
port 26 nsew
flabel metal3 s 585678 995407 590458 995907 0 FreeSans 3200 0 0 0 vssa1
port 26 nsew
flabel metal3 s 675407 415742 675907 420522 0 FreeSans 3200 0 0 0 vssa1
port 26 nsew
flabel metal3 s 675407 425721 675907 430501 0 FreeSans 3200 0 0 0 vssa1
port 26 nsew
flabel metal3 s 675407 503942 675907 508722 0 FreeSans 3200 0 0 0 vdda1
port 24 nsew
flabel metal3 s 675407 513921 675907 518701 0 FreeSans 3200 0 0 0 vdda1
port 24 nsew
flabel metal3 s 675407 818542 675907 823322 0 FreeSans 3200 0 0 0 vdda1
port 24 nsew
flabel metal3 s 675407 828521 675907 833301 0 FreeSans 3200 0 0 0 vdda1
port 24 nsew
flabel metal3 s 675407 907660 675907 912449 0 FreeSans 3200 0 0 0 vccd1
port 28 nsew
flabel metal3 s 675407 917700 675907 922500 0 FreeSans 3200 0 0 0 vccd1
port 28 nsew
flabel metal3 s 675407 912748 675907 917410 0 FreeSans 3200 0 0 0 vssd1
port 30 nsew
flabel metal3 675407 459860 675907 464649 0 FreeSans 3200 90 0 0 vssd1
port 30 nsew
flabel metal3 675407 469900 675907 474700 0 FreeSans 3200 90 0 0 vssd1
port 30 nsew
flabel metal3 675407 464949 675907 469600 0 FreeSans 3200 90 0 0 vccd1
port 28 nsew
flabel metal2 s 648115 41877 648167 42193 0 FreeSans 400 90 0 0 mask_rev[4]
port 65 nsew
flabel metal2 s 648339 41877 648391 42193 0 FreeSans 400 90 0 0 mask_rev[5]
port 64 nsew
flabel metal2 s 648563 41877 648615 42193 0 FreeSans 400 90 0 0 mask_rev[6]
port 63 nsew
flabel metal2 s 648787 41877 648839 42193 0 FreeSans 400 90 0 0 mask_rev[7]
port 62 nsew
flabel metal2 s 649011 41877 649063 42193 0 FreeSans 400 90 0 0 mask_rev[8]
port 61 nsew
flabel metal2 s 649235 41877 649287 42193 0 FreeSans 400 90 0 0 mask_rev[9]
port 60 nsew
flabel metal2 s 649459 41877 649511 42193 0 FreeSans 400 90 0 0 mask_rev[10]
port 59 nsew
flabel metal2 s 649683 41877 649735 42193 0 FreeSans 400 90 0 0 mask_rev[11]
port 58 nsew
flabel metal2 s 649907 41877 649959 42193 0 FreeSans 400 90 0 0 mask_rev[12]
port 57 nsew
flabel metal2 s 650131 41877 650183 42193 0 FreeSans 400 90 0 0 mask_rev[13]
port 56 nsew
flabel metal2 s 650355 41877 650407 42193 0 FreeSans 400 90 0 0 mask_rev[14]
port 55 nsew
flabel metal2 s 650579 41877 650631 42193 0 FreeSans 400 90 0 0 mask_rev[15]
port 54 nsew
flabel metal2 s 650803 41877 650855 42193 0 FreeSans 400 90 0 0 mask_rev[16]
port 53 nsew
flabel metal2 s 651027 41877 651079 42193 0 FreeSans 400 90 0 0 mask_rev[17]
port 52 nsew
flabel metal2 s 651251 41877 651303 42193 0 FreeSans 400 90 0 0 mask_rev[18]
port 51 nsew
flabel metal2 s 651475 41877 651527 42193 0 FreeSans 400 90 0 0 mask_rev[19]
port 50 nsew
flabel metal2 s 651699 41877 651751 42193 0 FreeSans 400 90 0 0 mask_rev[20]
port 49 nsew
flabel metal2 s 651923 41877 651975 42193 0 FreeSans 400 90 0 0 mask_rev[21]
port 48 nsew
flabel metal2 s 652147 41877 652199 42193 0 FreeSans 400 90 0 0 mask_rev[22]
port 47 nsew
flabel metal2 s 652371 41877 652423 42193 0 FreeSans 400 90 0 0 mask_rev[23]
port 46 nsew
flabel metal2 s 652595 41877 652647 42193 0 FreeSans 400 90 0 0 mask_rev[24]
port 45 nsew
flabel metal2 s 652819 41877 652871 42193 0 FreeSans 400 90 0 0 mask_rev[25]
port 44 nsew
flabel metal2 s 653043 41877 653095 42193 0 FreeSans 400 90 0 0 mask_rev[26]
port 43 nsew
flabel metal2 s 653267 41877 653319 42193 0 FreeSans 400 90 0 0 mask_rev[27]
port 42 nsew
flabel metal2 s 653491 41877 653543 42193 0 FreeSans 400 90 0 0 mask_rev[28]
port 41 nsew
flabel metal2 s 653715 41877 653767 42193 0 FreeSans 400 90 0 0 mask_rev[29]
port 40 nsew
flabel metal2 s 653939 41877 653991 42193 0 FreeSans 400 90 0 0 mask_rev[30]
port 39 nsew
flabel metal2 s 654163 41877 654215 42193 0 FreeSans 400 90 0 0 mask_rev[31]
port 38 nsew
flabel metal2 s 647891 41877 647943 42193 0 FreeSans 400 90 0 0 mask_rev[3]
port 66 nsew
flabel metal2 s 647667 41877 647719 42193 0 FreeSans 400 90 0 0 mask_rev[2]
port 67 nsew
flabel metal2 s 647443 41877 647495 42193 0 FreeSans 400 90 0 0 mask_rev[1]
port 68 nsew
flabel metal5 s 698512 952840 711002 965360 0 FreeSans 16000 0 0 0 gpio[14]
port 99 nsew
flabel metal3 675407 120144 675727 120206 0 FreeSans 400 0 0 0 gpio_loopback_zero[0]
port 817 nsew
flabel metal3 675407 165144 675727 165206 0 FreeSans 400 0 0 0 gpio_loopback_zero[1]
port 816 nsew
flabel metal3 675407 210144 675727 210206 0 FreeSans 400 0 0 0 gpio_loopback_zero[2]
port 815 nsew
flabel metal3 675407 255144 675727 255206 0 FreeSans 400 0 0 0 gpio_loopback_zero[3]
port 814 nsew
flabel metal3 675407 300144 675727 300206 0 FreeSans 400 0 0 0 gpio_loopback_zero[4]
port 813 nsew
flabel metal3 675407 345144 675727 345206 0 FreeSans 400 0 0 0 gpio_loopback_zero[5]
port 812 nsew
flabel metal3 675407 390144 675727 390206 0 FreeSans 400 0 0 0 gpio_loopback_zero[6]
port 811 nsew
flabel metal3 675407 567144 675727 567206 0 FreeSans 400 0 0 0 gpio_loopback_zero[7]
port 810 nsew
flabel metal3 675407 612144 675727 612206 0 FreeSans 400 0 0 0 gpio_loopback_zero[8]
port 809 nsew
flabel metal3 675407 657144 675727 657206 0 FreeSans 400 0 0 0 gpio_loopback_zero[9]
port 808 nsew
flabel metal3 675407 702144 675727 702206 0 FreeSans 400 0 0 0 gpio_loopback_zero[10]
port 807 nsew
flabel metal3 675407 747144 675727 747206 0 FreeSans 400 0 0 0 gpio_loopback_zero[11]
port 806 nsew
flabel metal3 675407 792144 675727 792206 0 FreeSans 400 0 0 0 gpio_loopback_zero[12]
port 805 nsew
flabel metal3 675407 881144 675727 881206 0 FreeSans 400 0 0 0 gpio_loopback_zero[13]
port 804 nsew
flabel metal3 675407 971144 675727 971206 0 FreeSans 400 0 0 0 gpio_loopback_zero[14]
port 803 nsew
flabel metal3 41873 776781 42193 776841 0 FreeSans 400 0 0 0 gpio_loopback_zero[25]
port 792 nsew
flabel metal3 41873 690781 42193 690841 0 FreeSans 400 0 0 0 gpio_loopback_zero[27]
port 790 nsew
flabel metal3 41873 604781 42193 604841 0 FreeSans 400 0 0 0 gpio_loopback_zero[29]
port 788 nsew
flabel metal3 41873 518781 42193 518841 0 FreeSans 400 0 0 0 gpio_loopback_zero[31]
port 786 nsew
flabel metal3 41873 346781 42193 346841 0 FreeSans 400 0 0 0 gpio_loopback_zero[33]
port 784 nsew
flabel metal3 41873 260781 42193 260841 0 FreeSans 400 0 0 0 gpio_loopback_zero[35]
port 782 nsew
flabel metal3 41873 174781 42193 174841 0 FreeSans 400 0 0 0 gpio_loopback_zero[37]
port 780 nsew
flabel metal3 41873 946781 42193 946841 0 FreeSans 400 0 0 0 gpio_loopback_zero[24]
port 793 nsew
flabel metal3 41873 733781 42193 733841 0 FreeSans 400 0 0 0 gpio_loopback_zero[26]
port 791 nsew
flabel metal3 41873 647781 42193 647841 0 FreeSans 400 0 0 0 gpio_loopback_zero[28]
port 789 nsew
flabel metal3 41873 561781 42193 561841 0 FreeSans 400 0 0 0 gpio_loopback_zero[30]
port 787 nsew
flabel metal3 41873 389781 42193 389841 0 FreeSans 400 0 0 0 gpio_loopback_zero[32]
port 785 nsew
flabel metal3 41873 303781 42193 303841 0 FreeSans 400 0 0 0 gpio_loopback_zero[34]
port 783 nsew
flabel metal3 41873 217781 42193 217841 0 FreeSans 400 0 0 0 gpio_loopback_zero[36]
port 781 nsew
flabel metal2 69634 995407 69695 995727 0 FreeSans 400 90 0 0 gpio_loopback_zero[23]
port 794 nsew
flabel metal2 120834 995407 120895 995727 0 FreeSans 400 90 0 0 gpio_loopback_zero[22]
port 795 nsew
flabel metal2 172034 995407 172095 995727 0 FreeSans 400 90 0 0 gpio_loopback_zero[21]
port 796 nsew
flabel metal2 223234 995407 223295 995727 0 FreeSans 400 90 0 0 gpio_loopback_zero[20]
port 797 nsew
flabel metal2 274434 995407 274495 995727 0 FreeSans 400 90 0 0 gpio_loopback_zero[19]
port 798 nsew
flabel metal2 378834 995407 378895 995727 0 FreeSans 400 90 0 0 gpio_loopback_zero[18]
port 799 nsew
flabel metal2 467834 995407 467895 995727 0 FreeSans 400 90 0 0 gpio_loopback_zero[17]
port 800 nsew
flabel metal2 519034 995407 519095 995727 0 FreeSans 400 90 0 0 gpio_loopback_zero[16]
port 801 nsew
flabel metal2 618434 995407 618495 995727 0 FreeSans 400 90 0 0 gpio_loopback_zero[15]
port 802 nsew
flabel metal3 s 675407 114444 675887 114514 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[0]
port 289 nsew
flabel metal3 s 675407 113800 675887 113870 0 FreeSans 400 0 0 0 gpio_vtrip_sel[0]
port 333 nsew
flabel metal3 675407 240644 675887 240714 0 FreeSans 400 0 0 0 analog_noesd_io[3]
port 946 nsew
flabel metal3 s 675407 326320 675887 326390 0 FreeSans 400 0 0 0 gpio_in[5]
port 724 nsew
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
