*---------------------------------------------------------------------------
* SPDX-FileCopyrightText: 2020 Efabless Corporation
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0
*---------------------------------------------------------------------------
* Threshold test for POR circuit
* Determine gate voltage at which the HV NFET draws 240nA nominal
*
* Result:  0.7575V
*-------------------------------------------------------------------

.lib /home/tim/projects/efabless/tech/SW/sky130A/libs.tech/ngspice/sky130.lib.spice tt


*----------------------------
* Testbench circuit
*----------------------------
Rtest vdda mir1 1MEG
Xm1 mir1 vin vss vss sky130_fd_pr__nfet_g5v0d10v5 w=2 l=0.8

Vgate vin vss DC=0
Vpwr vdda vss DC=3.3
Rgnd vss 0 0.1

*----------------------------
* Testbench control
*----------------------------
.control
* DC sweep from 0.7 to 0.8V
dc Vgate 0.7 0.8 0.001
wrdata test.data Vpwr#branch vin

.endc

.end

