VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_clocking
  CLASS BLOCK ;
  FOREIGN caravel_clocking ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 60.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 23.270 2.480 24.870 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.770 2.480 40.370 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.270 2.480 55.870 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.770 2.480 71.370 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 85.270 2.480 86.870 54.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 21.340 94.540 22.940 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 38.240 94.540 39.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.520 2.480 17.120 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.020 2.480 32.620 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.520 2.480 48.120 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.020 2.480 63.620 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 77.520 2.480 79.120 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.020 2.480 94.620 54.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 12.890 94.620 14.490 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 29.790 94.620 31.390 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.680 46.690 94.620 48.290 ;
    END
  END VPWR
  PIN core_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 56.000 35.790 60.000 ;
    END
  END core_clk
  PIN ext_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 56.000 21.530 60.000 ;
    END
  END ext_clk
  PIN ext_clk_sel
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 3.440 100.000 4.040 ;
    END
  END ext_clk_sel
  PIN ext_reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 55.800 100.000 56.400 ;
    END
  END ext_reset
  PIN pll_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 56.000 78.570 60.000 ;
    END
  END pll_clk
  PIN pll_clk90
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 56.000 92.830 60.000 ;
    END
  END pll_clk90
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 56.000 7.270 60.000 ;
    END
  END resetb
  PIN resetb_sync
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 56.000 64.310 60.000 ;
    END
  END resetb_sync
  PIN sel2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 33.360 100.000 33.960 ;
    END
  END sel2[0]
  PIN sel2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 40.840 100.000 41.440 ;
    END
  END sel2[1]
  PIN sel2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 48.320 100.000 48.920 ;
    END
  END sel2[2]
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 10.920 100.000 11.520 ;
    END
  END sel[0]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 18.400 100.000 19.000 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 25.880 100.000 26.480 ;
    END
  END sel[2]
  PIN user_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 56.000 50.050 60.000 ;
    END
  END user_clk
  OBS
      LAYER li1 ;
        RECT 0.920 2.635 94.300 54.485 ;
      LAYER met1 ;
        RECT 0.920 0.380 96.070 57.080 ;
      LAYER met2 ;
        RECT 2.400 55.720 6.710 57.110 ;
        RECT 7.550 55.720 20.970 57.110 ;
        RECT 21.810 55.720 35.230 57.110 ;
        RECT 36.070 55.720 49.490 57.110 ;
        RECT 50.330 55.720 63.750 57.110 ;
        RECT 64.590 55.720 78.010 57.110 ;
        RECT 78.850 55.720 92.270 57.110 ;
        RECT 93.110 55.720 96.040 57.110 ;
        RECT 2.400 0.350 96.040 55.720 ;
      LAYER met3 ;
        RECT 2.825 55.400 95.600 56.250 ;
        RECT 2.825 49.320 96.000 55.400 ;
        RECT 2.825 47.920 95.600 49.320 ;
        RECT 2.825 41.840 96.000 47.920 ;
        RECT 2.825 40.440 95.600 41.840 ;
        RECT 2.825 34.360 96.000 40.440 ;
        RECT 2.825 32.960 95.600 34.360 ;
        RECT 2.825 26.880 96.000 32.960 ;
        RECT 2.825 25.480 95.600 26.880 ;
        RECT 2.825 19.400 96.000 25.480 ;
        RECT 2.825 18.000 95.600 19.400 ;
        RECT 2.825 11.920 96.000 18.000 ;
        RECT 2.825 10.520 95.600 11.920 ;
        RECT 2.825 4.440 96.000 10.520 ;
        RECT 2.825 3.040 95.600 4.440 ;
        RECT 2.825 2.555 96.000 3.040 ;
      LAYER met4 ;
        RECT 72.055 4.935 77.120 42.665 ;
        RECT 79.520 4.935 84.870 42.665 ;
        RECT 87.270 4.935 88.025 42.665 ;
  END
END caravel_clocking
END LIBRARY

