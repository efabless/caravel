magic
tech sky130A
timestamp 1725322974
use sky130_ef_sc_hd__fill_4  sky130_ef_sc_hd__fill_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1720120574
transform 1 0 0 0 1 0
box -19 -24 203 296
use sky130_ef_sc_hd__fill_8  sky130_ef_sc_hd__fill_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1720120574
transform 1 0 184 0 1 0
box -19 -24 387 296
<< labels >>
flabel metal1 s 14 -8 31 8 0 FreeSans 200 0 0 0 VGND
port 2 nsew
flabel metal1 s 14 263 31 280 0 FreeSans 200 0 0 0 VPWR
port 3 nsew
flabel nwell s 14 263 31 280 0 FreeSans 200 0 0 0 VPB
port 4 nsew
flabel pwell s 14 -8 31 8 0 FreeSans 200 0 0 0 VNB
port 5 nsew
rlabel comment s 0 0 0 0 4 EF_fill_4_8
<< properties >>
string FIXED_BBOX 0 0 552 272
<< end >>
