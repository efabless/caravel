magic
tech sky130A
magscale 1 2
timestamp 1666279203
<< metal1 >>
rect 676030 897104 676036 897116
rect 663766 897076 676036 897104
rect 652018 896996 652024 897048
rect 652076 897036 652082 897048
rect 663766 897036 663794 897076
rect 676030 897064 676036 897076
rect 676088 897064 676094 897116
rect 652076 897008 663794 897036
rect 652076 896996 652082 897008
rect 654778 895772 654784 895824
rect 654836 895812 654842 895824
rect 675846 895812 675852 895824
rect 654836 895784 675852 895812
rect 654836 895772 654842 895784
rect 675846 895772 675852 895784
rect 675904 895772 675910 895824
rect 672718 895636 672724 895688
rect 672776 895676 672782 895688
rect 676030 895676 676036 895688
rect 672776 895648 676036 895676
rect 672776 895636 672782 895648
rect 676030 895636 676036 895648
rect 676088 895636 676094 895688
rect 671062 894412 671068 894464
rect 671120 894452 671126 894464
rect 675846 894452 675852 894464
rect 671120 894424 675852 894452
rect 671120 894412 671126 894424
rect 675846 894412 675852 894424
rect 675904 894412 675910 894464
rect 671890 894276 671896 894328
rect 671948 894316 671954 894328
rect 676030 894316 676036 894328
rect 671948 894288 676036 894316
rect 671948 894276 671954 894288
rect 676030 894276 676036 894288
rect 676088 894276 676094 894328
rect 672902 892984 672908 893036
rect 672960 893024 672966 893036
rect 676030 893024 676036 893036
rect 672960 892996 676036 893024
rect 672960 892984 672966 892996
rect 676030 892984 676036 892996
rect 676088 892984 676094 893036
rect 672534 892848 672540 892900
rect 672592 892888 672598 892900
rect 675846 892888 675852 892900
rect 672592 892860 675852 892888
rect 672592 892848 672598 892860
rect 675846 892848 675852 892860
rect 675904 892848 675910 892900
rect 675018 890332 675024 890384
rect 675076 890372 675082 890384
rect 676030 890372 676036 890384
rect 675076 890344 676036 890372
rect 675076 890332 675082 890344
rect 676030 890332 676036 890344
rect 676088 890332 676094 890384
rect 676214 890128 676220 890180
rect 676272 890168 676278 890180
rect 676858 890168 676864 890180
rect 676272 890140 676864 890168
rect 676272 890128 676278 890140
rect 676858 890128 676864 890140
rect 676916 890128 676922 890180
rect 674650 888904 674656 888956
rect 674708 888944 674714 888956
rect 676030 888944 676036 888956
rect 674708 888916 676036 888944
rect 674708 888904 674714 888916
rect 676030 888904 676036 888916
rect 676088 888904 676094 888956
rect 676214 888700 676220 888752
rect 676272 888740 676278 888752
rect 677042 888740 677048 888752
rect 676272 888712 677048 888740
rect 676272 888700 676278 888712
rect 677042 888700 677048 888712
rect 677100 888700 677106 888752
rect 674374 888496 674380 888548
rect 674432 888536 674438 888548
rect 676030 888536 676036 888548
rect 674432 888508 676036 888536
rect 674432 888496 674438 888508
rect 676030 888496 676036 888508
rect 676088 888496 676094 888548
rect 674190 887272 674196 887324
rect 674248 887312 674254 887324
rect 676030 887312 676036 887324
rect 674248 887284 676036 887312
rect 674248 887272 674254 887284
rect 676030 887272 676036 887284
rect 676088 887272 676094 887324
rect 670878 886864 670884 886916
rect 670936 886904 670942 886916
rect 676030 886904 676036 886916
rect 670936 886876 676036 886904
rect 670936 886864 670942 886876
rect 676030 886864 676036 886876
rect 676088 886864 676094 886916
rect 673086 885640 673092 885692
rect 673144 885680 673150 885692
rect 676030 885680 676036 885692
rect 673144 885652 676036 885680
rect 673144 885640 673150 885652
rect 676030 885640 676036 885652
rect 676088 885640 676094 885692
rect 653398 880472 653404 880524
rect 653456 880512 653462 880524
rect 653456 880484 666554 880512
rect 653456 880472 653462 880484
rect 666526 880376 666554 880484
rect 675386 880376 675392 880388
rect 666526 880348 675392 880376
rect 675386 880336 675392 880348
rect 675444 880336 675450 880388
rect 675018 879628 675024 879640
rect 674576 879600 675024 879628
rect 674576 879084 674604 879600
rect 675018 879588 675024 879600
rect 675076 879588 675082 879640
rect 677042 879492 677048 879504
rect 674760 879464 677048 879492
rect 674760 879232 674788 879464
rect 677042 879452 677048 879464
rect 677100 879452 677106 879504
rect 675938 879316 675944 879368
rect 675996 879356 676002 879368
rect 676858 879356 676864 879368
rect 675996 879328 676864 879356
rect 675996 879316 676002 879328
rect 676858 879316 676864 879328
rect 676916 879316 676922 879368
rect 674742 879180 674748 879232
rect 674800 879180 674806 879232
rect 674576 879056 675432 879084
rect 675404 878824 675432 879056
rect 675754 879044 675760 879096
rect 675812 879084 675818 879096
rect 678238 879084 678244 879096
rect 675812 879056 678244 879084
rect 675812 879044 675818 879056
rect 678238 879044 678244 879056
rect 678296 879044 678302 879096
rect 675202 878812 675208 878824
rect 674944 878784 675208 878812
rect 674944 878212 674972 878784
rect 675202 878772 675208 878784
rect 675260 878772 675266 878824
rect 675386 878772 675392 878824
rect 675444 878772 675450 878824
rect 676398 878608 676404 878620
rect 675312 878580 676404 878608
rect 674926 878160 674932 878212
rect 674984 878160 674990 878212
rect 675312 877928 675340 878580
rect 676398 878568 676404 878580
rect 676456 878568 676462 878620
rect 675938 878432 675944 878484
rect 675996 878432 676002 878484
rect 675956 878200 675984 878432
rect 675220 877900 675340 877928
rect 675588 878172 675984 878200
rect 675220 877804 675248 877900
rect 675202 877752 675208 877804
rect 675260 877752 675266 877804
rect 675588 877384 675616 878172
rect 675496 877356 675616 877384
rect 675496 877260 675524 877356
rect 675478 877208 675484 877260
rect 675536 877208 675542 877260
rect 674834 874148 674840 874200
rect 674892 874188 674898 874200
rect 675294 874188 675300 874200
rect 674892 874160 675300 874188
rect 674892 874148 674898 874160
rect 675294 874148 675300 874160
rect 675352 874148 675358 874200
rect 674374 872108 674380 872160
rect 674432 872148 674438 872160
rect 674834 872148 674840 872160
rect 674432 872120 674840 872148
rect 674432 872108 674438 872120
rect 674834 872108 674840 872120
rect 674892 872108 674898 872160
rect 657538 869388 657544 869440
rect 657596 869428 657602 869440
rect 675018 869428 675024 869440
rect 657596 869400 675024 869428
rect 657596 869388 657602 869400
rect 675018 869388 675024 869400
rect 675076 869388 675082 869440
rect 651466 868844 651472 868896
rect 651524 868884 651530 868896
rect 654778 868884 654784 868896
rect 651524 868856 654784 868884
rect 651524 868844 651530 868856
rect 654778 868844 654784 868856
rect 654836 868844 654842 868896
rect 674190 868708 674196 868760
rect 674248 868748 674254 868760
rect 675294 868748 675300 868760
rect 674248 868720 675300 868748
rect 674248 868708 674254 868720
rect 675294 868708 675300 868720
rect 675352 868708 675358 868760
rect 654134 868028 654140 868080
rect 654192 868068 654198 868080
rect 674834 868068 674840 868080
rect 654192 868040 674840 868068
rect 654192 868028 654198 868040
rect 674834 868028 674840 868040
rect 674892 868028 674898 868080
rect 651466 866600 651472 866652
rect 651524 866640 651530 866652
rect 672718 866640 672724 866652
rect 651524 866612 672724 866640
rect 651524 866600 651530 866612
rect 672718 866600 672724 866612
rect 672776 866600 672782 866652
rect 651374 865172 651380 865224
rect 651432 865212 651438 865224
rect 653398 865212 653404 865224
rect 651432 865184 653404 865212
rect 651432 865172 651438 865184
rect 653398 865172 653404 865184
rect 653456 865172 653462 865224
rect 651466 863812 651472 863864
rect 651524 863852 651530 863864
rect 657538 863852 657544 863864
rect 651524 863824 657544 863852
rect 651524 863812 651530 863824
rect 657538 863812 657544 863824
rect 657596 863812 657602 863864
rect 651466 862452 651472 862504
rect 651524 862492 651530 862504
rect 654134 862492 654140 862504
rect 651524 862464 654140 862492
rect 651524 862452 651530 862464
rect 654134 862452 654140 862464
rect 654192 862452 654198 862504
rect 35802 817096 35808 817148
rect 35860 817136 35866 817148
rect 44818 817136 44824 817148
rect 35860 817108 44824 817136
rect 35860 817096 35866 817108
rect 44818 817096 44824 817108
rect 44876 817096 44882 817148
rect 35618 816960 35624 817012
rect 35676 817000 35682 817012
rect 61378 817000 61384 817012
rect 35676 816972 61384 817000
rect 35676 816960 35682 816972
rect 61378 816960 61384 816972
rect 61436 816960 61442 817012
rect 35802 815736 35808 815788
rect 35860 815776 35866 815788
rect 43070 815776 43076 815788
rect 35860 815748 43076 815776
rect 35860 815736 35866 815748
rect 43070 815736 43076 815748
rect 43128 815736 43134 815788
rect 35434 815600 35440 815652
rect 35492 815640 35498 815652
rect 43438 815640 43444 815652
rect 35492 815612 43444 815640
rect 35492 815600 35498 815612
rect 43438 815600 43444 815612
rect 43496 815600 43502 815652
rect 35618 814376 35624 814428
rect 35676 814416 35682 814428
rect 42886 814416 42892 814428
rect 35676 814388 42892 814416
rect 35676 814376 35682 814388
rect 42886 814376 42892 814388
rect 42944 814376 42950 814428
rect 35802 814240 35808 814292
rect 35860 814280 35866 814292
rect 44174 814280 44180 814292
rect 35860 814252 44180 814280
rect 35860 814240 35866 814252
rect 44174 814240 44180 814252
rect 44232 814240 44238 814292
rect 41322 812812 41328 812864
rect 41380 812852 41386 812864
rect 44450 812852 44456 812864
rect 41380 812824 44456 812852
rect 41380 812812 41386 812824
rect 44450 812812 44456 812824
rect 44508 812812 44514 812864
rect 40954 811384 40960 811436
rect 41012 811424 41018 811436
rect 42610 811424 42616 811436
rect 41012 811396 42616 811424
rect 41012 811384 41018 811396
rect 42610 811384 42616 811396
rect 42668 811384 42674 811436
rect 40678 808596 40684 808648
rect 40736 808636 40742 808648
rect 41782 808636 41788 808648
rect 40736 808608 41788 808636
rect 40736 808596 40742 808608
rect 41782 808596 41788 808608
rect 41840 808596 41846 808648
rect 41138 808052 41144 808104
rect 41196 808092 41202 808104
rect 41598 808092 41604 808104
rect 41196 808064 41604 808092
rect 41196 808052 41202 808064
rect 41598 808052 41604 808064
rect 41656 808052 41662 808104
rect 43438 807916 43444 807968
rect 43496 807956 43502 807968
rect 62942 807956 62948 807968
rect 43496 807928 62948 807956
rect 43496 807916 43502 807928
rect 62942 807916 62948 807928
rect 63000 807916 63006 807968
rect 41138 807304 41144 807356
rect 41196 807344 41202 807356
rect 44634 807344 44640 807356
rect 41196 807316 44640 807344
rect 41196 807304 41202 807316
rect 44634 807304 44640 807316
rect 44692 807304 44698 807356
rect 41322 806080 41328 806132
rect 41380 806120 41386 806132
rect 50338 806120 50344 806132
rect 41380 806092 50344 806120
rect 41380 806080 41386 806092
rect 50338 806080 50344 806092
rect 50396 806080 50402 806132
rect 41138 805944 41144 805996
rect 41196 805984 41202 805996
rect 62666 805984 62672 805996
rect 41196 805956 62672 805984
rect 41196 805944 41202 805956
rect 62666 805944 62672 805956
rect 62724 805944 62730 805996
rect 34514 802544 34520 802596
rect 34572 802584 34578 802596
rect 41782 802584 41788 802596
rect 34572 802556 41788 802584
rect 34572 802544 34578 802556
rect 41782 802544 41788 802556
rect 41840 802544 41846 802596
rect 32398 802408 32404 802460
rect 32456 802448 32462 802460
rect 42702 802448 42708 802460
rect 32456 802420 42708 802448
rect 32456 802408 32462 802420
rect 42702 802408 42708 802420
rect 42760 802408 42766 802460
rect 33778 801184 33784 801236
rect 33836 801224 33842 801236
rect 42610 801224 42616 801236
rect 33836 801196 42616 801224
rect 33836 801184 33842 801196
rect 42610 801184 42616 801196
rect 42668 801184 42674 801236
rect 31018 801048 31024 801100
rect 31076 801088 31082 801100
rect 43438 801088 43444 801100
rect 31076 801060 43444 801088
rect 31076 801048 31082 801060
rect 43438 801048 43444 801060
rect 43496 801048 43502 801100
rect 42426 799076 42432 799128
rect 42484 799116 42490 799128
rect 42484 799088 48314 799116
rect 42484 799076 42490 799088
rect 48286 799048 48314 799088
rect 53098 799048 53104 799060
rect 48286 799020 53104 799048
rect 53098 799008 53104 799020
rect 53156 799008 53162 799060
rect 43622 797648 43628 797700
rect 43680 797688 43686 797700
rect 57238 797688 57244 797700
rect 43680 797660 57244 797688
rect 43680 797648 43686 797660
rect 57238 797648 57244 797660
rect 57296 797648 57302 797700
rect 44634 796328 44640 796340
rect 42260 796300 44640 796328
rect 42260 795048 42288 796300
rect 44634 796288 44640 796300
rect 44692 796288 44698 796340
rect 42426 795608 42432 795660
rect 42484 795648 42490 795660
rect 43622 795648 43628 795660
rect 42484 795620 43628 795648
rect 42484 795608 42490 795620
rect 43622 795608 43628 795620
rect 43680 795608 43686 795660
rect 42242 794996 42248 795048
rect 42300 794996 42306 795048
rect 42242 793772 42248 793824
rect 42300 793812 42306 793824
rect 43162 793812 43168 793824
rect 42300 793784 43168 793812
rect 42300 793772 42306 793784
rect 43162 793772 43168 793784
rect 43220 793772 43226 793824
rect 42610 793500 42616 793552
rect 42668 793540 42674 793552
rect 43438 793540 43444 793552
rect 42668 793512 43444 793540
rect 42668 793500 42674 793512
rect 43438 793500 43444 793512
rect 43496 793500 43502 793552
rect 653398 790780 653404 790832
rect 653456 790820 653462 790832
rect 675386 790820 675392 790832
rect 653456 790792 675392 790820
rect 653456 790780 653462 790792
rect 675386 790780 675392 790792
rect 675444 790780 675450 790832
rect 53098 790712 53104 790764
rect 53156 790752 53162 790764
rect 62206 790752 62212 790764
rect 53156 790724 62212 790752
rect 53156 790712 53162 790724
rect 62206 790712 62212 790724
rect 62264 790712 62270 790764
rect 42426 790576 42432 790628
rect 42484 790576 42490 790628
rect 42150 790372 42156 790424
rect 42208 790412 42214 790424
rect 42444 790412 42472 790576
rect 42208 790384 42472 790412
rect 42208 790372 42214 790384
rect 42242 789760 42248 789812
rect 42300 789760 42306 789812
rect 42260 789540 42288 789760
rect 42242 789488 42248 789540
rect 42300 789488 42306 789540
rect 57238 789148 57244 789200
rect 57296 789188 57302 789200
rect 62114 789188 62120 789200
rect 57296 789160 62120 789188
rect 57296 789148 57302 789160
rect 62114 789148 62120 789160
rect 62172 789148 62178 789200
rect 62114 786672 62120 786684
rect 42536 786644 62120 786672
rect 42536 785664 42564 786644
rect 62114 786632 62120 786644
rect 62172 786632 62178 786684
rect 42518 785612 42524 785664
rect 42576 785612 42582 785664
rect 44818 785136 44824 785188
rect 44876 785176 44882 785188
rect 62114 785176 62120 785188
rect 44876 785148 62120 785176
rect 44876 785136 44882 785148
rect 62114 785136 62120 785148
rect 62172 785136 62178 785188
rect 670602 784252 670608 784304
rect 670660 784292 670666 784304
rect 675110 784292 675116 784304
rect 670660 784264 675116 784292
rect 670660 784252 670666 784264
rect 675110 784252 675116 784264
rect 675168 784252 675174 784304
rect 669222 784116 669228 784168
rect 669280 784156 669286 784168
rect 675386 784156 675392 784168
rect 669280 784128 675392 784156
rect 669280 784116 669286 784128
rect 675386 784116 675392 784128
rect 675444 784116 675450 784168
rect 673730 782620 673736 782672
rect 673788 782660 673794 782672
rect 675110 782660 675116 782672
rect 673788 782632 675116 782660
rect 673788 782620 673794 782632
rect 675110 782620 675116 782632
rect 675168 782620 675174 782672
rect 669038 782484 669044 782536
rect 669096 782524 669102 782536
rect 675294 782524 675300 782536
rect 669096 782496 675300 782524
rect 669096 782484 669102 782496
rect 675294 782484 675300 782496
rect 675352 782484 675358 782536
rect 655514 781056 655520 781108
rect 655572 781096 655578 781108
rect 675018 781096 675024 781108
rect 655572 781068 675024 781096
rect 655572 781056 655578 781068
rect 675018 781056 675024 781068
rect 675076 781056 675082 781108
rect 673914 779968 673920 780020
rect 673972 780008 673978 780020
rect 675110 780008 675116 780020
rect 673972 779980 675116 780008
rect 673972 779968 673978 779980
rect 675110 779968 675116 779980
rect 675168 779968 675174 780020
rect 655054 778336 655060 778388
rect 655112 778376 655118 778388
rect 674926 778376 674932 778388
rect 655112 778348 674932 778376
rect 655112 778336 655118 778348
rect 674926 778336 674932 778348
rect 674984 778336 674990 778388
rect 651466 777588 651472 777640
rect 651524 777628 651530 777640
rect 660298 777628 660304 777640
rect 651524 777600 660304 777628
rect 651524 777588 651530 777600
rect 660298 777588 660304 777600
rect 660356 777588 660362 777640
rect 670418 776976 670424 777028
rect 670476 777016 670482 777028
rect 675294 777016 675300 777028
rect 670476 776988 675300 777016
rect 670476 776976 670482 776988
rect 675294 776976 675300 776988
rect 675352 776976 675358 777028
rect 672718 775616 672724 775668
rect 672776 775656 672782 775668
rect 674926 775656 674932 775668
rect 672776 775628 674932 775656
rect 672776 775616 672782 775628
rect 674926 775616 674932 775628
rect 674984 775616 674990 775668
rect 651466 775548 651472 775600
rect 651524 775588 651530 775600
rect 669958 775588 669964 775600
rect 651524 775560 669964 775588
rect 651524 775548 651530 775560
rect 669958 775548 669964 775560
rect 670016 775548 670022 775600
rect 651374 775276 651380 775328
rect 651432 775316 651438 775328
rect 653398 775316 653404 775328
rect 651432 775288 653404 775316
rect 651432 775276 651438 775288
rect 653398 775276 653404 775288
rect 653456 775276 653462 775328
rect 35802 774188 35808 774240
rect 35860 774228 35866 774240
rect 41690 774228 41696 774240
rect 35860 774200 41696 774228
rect 35860 774188 35866 774200
rect 41690 774188 41696 774200
rect 41748 774188 41754 774240
rect 42058 774188 42064 774240
rect 42116 774228 42122 774240
rect 59998 774228 60004 774240
rect 42116 774200 60004 774228
rect 42116 774188 42122 774200
rect 59998 774188 60004 774200
rect 60056 774188 60062 774240
rect 651466 774120 651472 774172
rect 651524 774160 651530 774172
rect 655514 774160 655520 774172
rect 651524 774132 655520 774160
rect 651524 774120 651530 774132
rect 655514 774120 655520 774132
rect 655572 774120 655578 774172
rect 651466 773780 651472 773832
rect 651524 773820 651530 773832
rect 655054 773820 655060 773832
rect 651524 773792 655060 773820
rect 651524 773780 651530 773792
rect 655054 773780 655060 773792
rect 655112 773780 655118 773832
rect 671430 773372 671436 773424
rect 671488 773412 671494 773424
rect 675294 773412 675300 773424
rect 671488 773384 675300 773412
rect 671488 773372 671494 773384
rect 675294 773372 675300 773384
rect 675352 773372 675358 773424
rect 35802 773304 35808 773356
rect 35860 773344 35866 773356
rect 41690 773344 41696 773356
rect 35860 773316 41696 773344
rect 35860 773304 35866 773316
rect 41690 773304 41696 773316
rect 41748 773304 41754 773356
rect 35802 773100 35808 773152
rect 35860 773140 35866 773152
rect 40770 773140 40776 773152
rect 35860 773112 40776 773140
rect 35860 773100 35866 773112
rect 40770 773100 40776 773112
rect 40828 773100 40834 773152
rect 35526 772964 35532 773016
rect 35584 773004 35590 773016
rect 41690 773004 41696 773016
rect 35584 772976 41696 773004
rect 35584 772964 35590 772976
rect 41690 772964 41696 772976
rect 41748 772964 41754 773016
rect 42058 772964 42064 773016
rect 42116 773004 42122 773016
rect 43162 773004 43168 773016
rect 42116 772976 43168 773004
rect 42116 772964 42122 772976
rect 43162 772964 43168 772976
rect 43220 772964 43226 773016
rect 35342 772828 35348 772880
rect 35400 772868 35406 772880
rect 61378 772868 61384 772880
rect 35400 772840 41736 772868
rect 35400 772828 35406 772840
rect 41708 772744 41736 772840
rect 42076 772840 61384 772868
rect 42076 772744 42104 772840
rect 61378 772828 61384 772840
rect 61436 772828 61442 772880
rect 41690 772692 41696 772744
rect 41748 772692 41754 772744
rect 42058 772692 42064 772744
rect 42116 772692 42122 772744
rect 35802 771808 35808 771860
rect 35860 771848 35866 771860
rect 40218 771848 40224 771860
rect 35860 771820 40224 771848
rect 35860 771808 35866 771820
rect 40218 771808 40224 771820
rect 40276 771808 40282 771860
rect 41046 771644 41052 771656
rect 38626 771616 41052 771644
rect 35618 771536 35624 771588
rect 35676 771576 35682 771588
rect 38626 771576 38654 771616
rect 41046 771604 41052 771616
rect 41104 771604 41110 771656
rect 35676 771548 38654 771576
rect 35676 771536 35682 771548
rect 35802 771400 35808 771452
rect 35860 771440 35866 771452
rect 41690 771440 41696 771452
rect 35860 771412 41696 771440
rect 35860 771400 35866 771412
rect 41690 771400 41696 771412
rect 41748 771400 41754 771452
rect 42058 771400 42064 771452
rect 42116 771440 42122 771452
rect 44174 771440 44180 771452
rect 42116 771412 44180 771440
rect 42116 771400 42122 771412
rect 44174 771400 44180 771412
rect 44232 771400 44238 771452
rect 35802 770448 35808 770500
rect 35860 770488 35866 770500
rect 39850 770488 39856 770500
rect 35860 770460 39856 770488
rect 35860 770448 35866 770460
rect 39850 770448 39856 770460
rect 39908 770448 39914 770500
rect 35618 770176 35624 770228
rect 35676 770216 35682 770228
rect 41506 770216 41512 770228
rect 35676 770188 41512 770216
rect 35676 770176 35682 770188
rect 41506 770176 41512 770188
rect 41564 770176 41570 770228
rect 35802 770040 35808 770092
rect 35860 770080 35866 770092
rect 41690 770080 41696 770092
rect 35860 770052 41696 770080
rect 35860 770040 35866 770052
rect 41690 770040 41696 770052
rect 41748 770040 41754 770092
rect 42058 770040 42064 770092
rect 42116 770080 42122 770092
rect 44542 770080 44548 770092
rect 42116 770052 44548 770080
rect 42116 770040 42122 770052
rect 44542 770040 44548 770052
rect 44600 770040 44606 770092
rect 35802 769156 35808 769208
rect 35860 769196 35866 769208
rect 35860 769156 35894 769196
rect 35866 768992 35894 769156
rect 41690 768992 41696 769004
rect 35866 768964 41696 768992
rect 41690 768952 41696 768964
rect 41748 768952 41754 769004
rect 35526 768816 35532 768868
rect 35584 768856 35590 768868
rect 41230 768856 41236 768868
rect 35584 768828 41236 768856
rect 35584 768816 35590 768828
rect 41230 768816 41236 768828
rect 41288 768816 41294 768868
rect 35802 768680 35808 768732
rect 35860 768720 35866 768732
rect 40034 768720 40040 768732
rect 35860 768692 40040 768720
rect 35860 768680 35866 768692
rect 40034 768680 40040 768692
rect 40092 768680 40098 768732
rect 35802 767320 35808 767372
rect 35860 767360 35866 767372
rect 36538 767360 36544 767372
rect 35860 767332 36544 767360
rect 35860 767320 35866 767332
rect 36538 767320 36544 767332
rect 36596 767320 36602 767372
rect 35802 766028 35808 766080
rect 35860 766068 35866 766080
rect 39758 766068 39764 766080
rect 35860 766040 39764 766068
rect 35860 766028 35866 766040
rect 39758 766028 39764 766040
rect 39816 766028 39822 766080
rect 40034 765280 40040 765332
rect 40092 765320 40098 765332
rect 41690 765320 41696 765332
rect 40092 765292 41696 765320
rect 40092 765280 40098 765292
rect 41690 765280 41696 765292
rect 41748 765280 41754 765332
rect 42058 765144 42064 765196
rect 42116 765184 42122 765196
rect 42518 765184 42524 765196
rect 42116 765156 42524 765184
rect 42116 765144 42122 765156
rect 42518 765144 42524 765156
rect 42576 765144 42582 765196
rect 35802 764804 35808 764856
rect 35860 764844 35866 764856
rect 39390 764844 39396 764856
rect 35860 764816 39396 764844
rect 35860 764804 35866 764816
rect 39390 764804 39396 764816
rect 39448 764804 39454 764856
rect 41690 764640 41696 764652
rect 36004 764612 41696 764640
rect 35802 764532 35808 764584
rect 35860 764572 35866 764584
rect 36004 764572 36032 764612
rect 41690 764600 41696 764612
rect 41748 764600 41754 764652
rect 35860 764544 36032 764572
rect 35860 764532 35866 764544
rect 35618 763444 35624 763496
rect 35676 763484 35682 763496
rect 40954 763484 40960 763496
rect 35676 763456 40960 763484
rect 35676 763444 35682 763456
rect 40954 763444 40960 763456
rect 41012 763444 41018 763496
rect 40696 763252 41736 763280
rect 35802 763172 35808 763224
rect 35860 763212 35866 763224
rect 40696 763212 40724 763252
rect 35860 763184 40724 763212
rect 35860 763172 35866 763184
rect 41708 763156 41736 763252
rect 53098 763212 53104 763224
rect 41984 763184 53104 763212
rect 41690 763104 41696 763156
rect 41748 763104 41754 763156
rect 41984 763076 42012 763184
rect 53098 763172 53104 763184
rect 53156 763172 53162 763224
rect 42426 763076 42432 763088
rect 41984 763048 42432 763076
rect 42426 763036 42432 763048
rect 42484 763036 42490 763088
rect 42058 761880 42064 761932
rect 42116 761920 42122 761932
rect 48958 761920 48964 761932
rect 42116 761892 48964 761920
rect 42116 761880 42122 761892
rect 48958 761880 48964 761892
rect 49016 761880 49022 761932
rect 35802 761812 35808 761864
rect 35860 761852 35866 761864
rect 41690 761852 41696 761864
rect 35860 761824 41696 761852
rect 35860 761812 35866 761824
rect 41690 761812 41696 761824
rect 41748 761812 41754 761864
rect 35158 759772 35164 759824
rect 35216 759812 35222 759824
rect 41690 759812 41696 759824
rect 35216 759784 41696 759812
rect 35216 759772 35222 759784
rect 41690 759772 41696 759784
rect 41748 759772 41754 759824
rect 32398 759636 32404 759688
rect 32456 759676 32462 759688
rect 41598 759676 41604 759688
rect 32456 759648 41604 759676
rect 32456 759636 32462 759648
rect 41598 759636 41604 759648
rect 41656 759636 41662 759688
rect 42058 759500 42064 759552
rect 42116 759540 42122 759552
rect 42426 759540 42432 759552
rect 42116 759512 42432 759540
rect 42116 759500 42122 759512
rect 42426 759500 42432 759512
rect 42484 759500 42490 759552
rect 33778 758276 33784 758328
rect 33836 758316 33842 758328
rect 39206 758316 39212 758328
rect 33836 758288 39212 758316
rect 33836 758276 33842 758288
rect 39206 758276 39212 758288
rect 39264 758276 39270 758328
rect 42242 756032 42248 756084
rect 42300 756032 42306 756084
rect 42260 755472 42288 756032
rect 44726 755488 44732 755540
rect 44784 755528 44790 755540
rect 62942 755528 62948 755540
rect 44784 755500 62948 755528
rect 44784 755488 44790 755500
rect 62942 755488 62948 755500
rect 63000 755488 63006 755540
rect 42242 755420 42248 755472
rect 42300 755420 42306 755472
rect 43622 754876 43628 754928
rect 43680 754916 43686 754928
rect 45002 754916 45008 754928
rect 43680 754888 45008 754916
rect 43680 754876 43686 754888
rect 45002 754876 45008 754888
rect 45060 754876 45066 754928
rect 43990 753516 43996 753568
rect 44048 753556 44054 753568
rect 45370 753556 45376 753568
rect 44048 753528 45376 753556
rect 44048 753516 44054 753528
rect 45370 753516 45376 753528
rect 45428 753516 45434 753568
rect 61378 747260 61384 747312
rect 61436 747300 61442 747312
rect 63034 747300 63040 747312
rect 61436 747272 63040 747300
rect 61436 747260 61442 747272
rect 63034 747260 63040 747272
rect 63092 747260 63098 747312
rect 653398 746580 653404 746632
rect 653456 746620 653462 746632
rect 675386 746620 675392 746632
rect 653456 746592 675392 746620
rect 653456 746580 653462 746592
rect 675386 746580 675392 746592
rect 675444 746580 675450 746632
rect 44818 746512 44824 746564
rect 44876 746552 44882 746564
rect 62114 746552 62120 746564
rect 44876 746524 62120 746552
rect 44876 746512 44882 746524
rect 62114 746512 62120 746524
rect 62172 746512 62178 746564
rect 42794 744064 42800 744116
rect 42852 744104 42858 744116
rect 42852 744076 45554 744104
rect 42852 744064 42858 744076
rect 45526 743900 45554 744076
rect 62114 743900 62120 743912
rect 45526 743872 62120 743900
rect 62114 743860 62120 743872
rect 62172 743860 62178 743912
rect 46198 743724 46204 743776
rect 46256 743764 46262 743776
rect 62114 743764 62120 743776
rect 46256 743736 62120 743764
rect 46256 743724 46262 743736
rect 62114 743724 62120 743736
rect 62172 743724 62178 743776
rect 59998 742364 60004 742416
rect 60056 742404 60062 742416
rect 62114 742404 62120 742416
rect 60056 742376 62120 742404
rect 60056 742364 60062 742376
rect 62114 742364 62120 742376
rect 62172 742364 62178 742416
rect 671798 742160 671804 742212
rect 671856 742200 671862 742212
rect 675386 742200 675392 742212
rect 671856 742172 675392 742200
rect 671856 742160 671862 742172
rect 675386 742160 675392 742172
rect 675444 742160 675450 742212
rect 671614 741140 671620 741192
rect 671672 741180 671678 741192
rect 675110 741180 675116 741192
rect 671672 741152 675116 741180
rect 671672 741140 671678 741152
rect 675110 741140 675116 741152
rect 675168 741140 675174 741192
rect 673546 738624 673552 738676
rect 673604 738664 673610 738676
rect 675386 738664 675392 738676
rect 673604 738636 675392 738664
rect 673604 738624 673610 738636
rect 675386 738624 675392 738636
rect 675444 738624 675450 738676
rect 672258 738420 672264 738472
rect 672316 738460 672322 738472
rect 675110 738460 675116 738472
rect 672316 738432 675116 738460
rect 672316 738420 672322 738432
rect 675110 738420 675116 738432
rect 675168 738420 675174 738472
rect 652018 736856 652024 736908
rect 652076 736896 652082 736908
rect 656158 736896 656164 736908
rect 652076 736868 656164 736896
rect 652076 736856 652082 736868
rect 656158 736856 656164 736868
rect 656216 736856 656222 736908
rect 675294 735740 675300 735752
rect 663766 735712 675300 735740
rect 657538 735564 657544 735616
rect 657596 735604 657602 735616
rect 663766 735604 663794 735712
rect 675294 735700 675300 735712
rect 675352 735700 675358 735752
rect 657596 735576 663794 735604
rect 657596 735564 657602 735576
rect 669590 735564 669596 735616
rect 669648 735604 669654 735616
rect 675110 735604 675116 735616
rect 669648 735576 675116 735604
rect 669648 735564 669654 735576
rect 675110 735564 675116 735576
rect 675168 735564 675174 735616
rect 675110 734244 675116 734256
rect 663766 734216 675116 734244
rect 654778 734136 654784 734188
rect 654836 734176 654842 734188
rect 663766 734176 663794 734216
rect 675110 734204 675116 734216
rect 675168 734204 675174 734256
rect 654836 734148 663794 734176
rect 654836 734136 654842 734148
rect 651466 733388 651472 733440
rect 651524 733428 651530 733440
rect 668578 733428 668584 733440
rect 651524 733400 668584 733428
rect 651524 733388 651530 733400
rect 668578 733388 668584 733400
rect 668636 733388 668642 733440
rect 672074 732708 672080 732760
rect 672132 732748 672138 732760
rect 675294 732748 675300 732760
rect 672132 732720 675300 732748
rect 672132 732708 672138 732720
rect 675294 732708 675300 732720
rect 675352 732708 675358 732760
rect 651466 731416 651472 731468
rect 651524 731456 651530 731468
rect 658918 731456 658924 731468
rect 651524 731428 658924 731456
rect 651524 731416 651530 731428
rect 658918 731416 658924 731428
rect 658976 731416 658982 731468
rect 651374 731076 651380 731128
rect 651432 731116 651438 731128
rect 653398 731116 653404 731128
rect 651432 731088 653404 731116
rect 651432 731076 651438 731088
rect 653398 731076 653404 731088
rect 653456 731076 653462 731128
rect 674926 731076 674932 731128
rect 674984 731076 674990 731128
rect 674944 730912 674972 731076
rect 675110 730912 675116 730924
rect 674944 730884 675116 730912
rect 675110 730872 675116 730884
rect 675168 730872 675174 730924
rect 652662 730668 652668 730720
rect 652720 730708 652726 730720
rect 661678 730708 661684 730720
rect 652720 730680 661684 730708
rect 652720 730668 652726 730680
rect 661678 730668 661684 730680
rect 661736 730668 661742 730720
rect 43622 730260 43628 730312
rect 43680 730300 43686 730312
rect 61378 730300 61384 730312
rect 43680 730272 61384 730300
rect 43680 730260 43686 730272
rect 61378 730260 61384 730272
rect 61436 730260 61442 730312
rect 651466 729988 651472 730040
rect 651524 730028 651530 730040
rect 657538 730028 657544 730040
rect 651524 730000 657544 730028
rect 651524 729988 651530 730000
rect 657538 729988 657544 730000
rect 657596 729988 657602 730040
rect 42242 729308 42248 729360
rect 42300 729348 42306 729360
rect 62942 729348 62948 729360
rect 42300 729320 62948 729348
rect 42300 729308 42306 729320
rect 62942 729308 62948 729320
rect 63000 729308 63006 729360
rect 41690 728872 41696 728884
rect 41386 728844 41696 728872
rect 40954 728764 40960 728816
rect 41012 728804 41018 728816
rect 41386 728804 41414 728844
rect 41690 728832 41696 728844
rect 41748 728832 41754 728884
rect 42058 728832 42064 728884
rect 42116 728872 42122 728884
rect 43070 728872 43076 728884
rect 42116 728844 43076 728872
rect 42116 728832 42122 728844
rect 43070 728832 43076 728844
rect 43128 728832 43134 728884
rect 41012 728776 41414 728804
rect 41012 728764 41018 728776
rect 41138 728628 41144 728680
rect 41196 728668 41202 728680
rect 41690 728668 41696 728680
rect 41196 728640 41696 728668
rect 41196 728628 41202 728640
rect 41690 728628 41696 728640
rect 41748 728628 41754 728680
rect 42058 728628 42064 728680
rect 42116 728668 42122 728680
rect 43438 728668 43444 728680
rect 42116 728640 43444 728668
rect 42116 728628 42122 728640
rect 43438 728628 43444 728640
rect 43496 728628 43502 728680
rect 651466 728492 651472 728544
rect 651524 728532 651530 728544
rect 654778 728532 654784 728544
rect 651524 728504 654784 728532
rect 651524 728492 651530 728504
rect 654778 728492 654784 728504
rect 654836 728492 654842 728544
rect 673086 728288 673092 728340
rect 673144 728328 673150 728340
rect 673144 728300 674176 728328
rect 673144 728288 673150 728300
rect 670878 728084 670884 728136
rect 670936 728124 670942 728136
rect 670936 728096 674058 728124
rect 670936 728084 670942 728096
rect 40862 727404 40868 727456
rect 40920 727444 40926 727456
rect 41690 727444 41696 727456
rect 40920 727416 41696 727444
rect 40920 727404 40926 727416
rect 41690 727404 41696 727416
rect 41748 727404 41754 727456
rect 42058 727404 42064 727456
rect 42116 727444 42122 727456
rect 44358 727444 44364 727456
rect 42116 727416 44364 727444
rect 42116 727404 42122 727416
rect 44358 727404 44364 727416
rect 44416 727404 44422 727456
rect 41322 727268 41328 727320
rect 41380 727308 41386 727320
rect 41690 727308 41696 727320
rect 41380 727280 41696 727308
rect 41380 727268 41386 727280
rect 41690 727268 41696 727280
rect 41748 727268 41754 727320
rect 42058 727268 42064 727320
rect 42116 727308 42122 727320
rect 44634 727308 44640 727320
rect 42116 727280 44640 727308
rect 42116 727268 42122 727280
rect 44634 727268 44640 727280
rect 44692 727268 44698 727320
rect 674558 726724 674564 726776
rect 674616 726764 674622 726776
rect 683390 726764 683396 726776
rect 674616 726736 683396 726764
rect 674616 726724 674622 726736
rect 683390 726724 683396 726736
rect 683448 726724 683454 726776
rect 674742 726520 674748 726572
rect 674800 726560 674806 726572
rect 680998 726560 681004 726572
rect 674800 726532 681004 726560
rect 674800 726520 674806 726532
rect 680998 726520 681004 726532
rect 681056 726520 681062 726572
rect 674374 726384 674380 726436
rect 674432 726424 674438 726436
rect 684034 726424 684040 726436
rect 674432 726396 684040 726424
rect 674432 726384 674438 726396
rect 684034 726384 684040 726396
rect 684092 726384 684098 726436
rect 41322 726180 41328 726232
rect 41380 726220 41386 726232
rect 41690 726220 41696 726232
rect 41380 726192 41696 726220
rect 41380 726180 41386 726192
rect 41690 726180 41696 726192
rect 41748 726180 41754 726232
rect 41138 725908 41144 725960
rect 41196 725948 41202 725960
rect 41598 725948 41604 725960
rect 41196 725920 41604 725948
rect 41196 725908 41202 725920
rect 41598 725908 41604 725920
rect 41656 725908 41662 725960
rect 675294 721692 675300 721744
rect 675352 721692 675358 721744
rect 675312 721268 675340 721692
rect 675294 721216 675300 721268
rect 675352 721216 675358 721268
rect 673914 721012 673920 721064
rect 673972 721052 673978 721064
rect 673972 721024 674512 721052
rect 673972 721012 673978 721024
rect 674484 720520 674512 721024
rect 675294 720808 675300 720860
rect 675352 720808 675358 720860
rect 675312 720520 675340 720808
rect 674466 720468 674472 720520
rect 674524 720468 674530 720520
rect 675294 720468 675300 720520
rect 675352 720468 675358 720520
rect 43622 718972 43628 719024
rect 43680 719012 43686 719024
rect 55858 719012 55864 719024
rect 43680 718984 55864 719012
rect 43680 718972 43686 718984
rect 55858 718972 55864 718984
rect 55916 718972 55922 719024
rect 32398 716796 32404 716848
rect 32456 716836 32462 716848
rect 41690 716836 41696 716848
rect 32456 716808 41696 716836
rect 32456 716796 32462 716808
rect 41690 716796 41696 716808
rect 41748 716796 41754 716848
rect 674282 716456 674288 716508
rect 674340 716496 674346 716508
rect 676030 716496 676036 716508
rect 674340 716468 676036 716496
rect 674340 716456 674346 716468
rect 676030 716456 676036 716468
rect 676088 716456 676094 716508
rect 656158 716252 656164 716304
rect 656216 716292 656222 716304
rect 674006 716292 674012 716304
rect 656216 716264 674012 716292
rect 656216 716252 656222 716264
rect 674006 716252 674012 716264
rect 674064 716252 674070 716304
rect 669958 715708 669964 715760
rect 670016 715748 670022 715760
rect 674006 715748 674012 715760
rect 670016 715720 674012 715748
rect 670016 715708 670022 715720
rect 674006 715708 674012 715720
rect 674064 715708 674070 715760
rect 35158 715640 35164 715692
rect 35216 715680 35222 715692
rect 40402 715680 40408 715692
rect 35216 715652 40408 715680
rect 35216 715640 35222 715652
rect 40402 715640 40408 715652
rect 40460 715640 40466 715692
rect 31662 715436 31668 715488
rect 31720 715476 31726 715488
rect 38010 715476 38016 715488
rect 31720 715448 38016 715476
rect 31720 715436 31726 715448
rect 38010 715436 38016 715448
rect 38068 715436 38074 715488
rect 671062 715300 671068 715352
rect 671120 715340 671126 715352
rect 674006 715340 674012 715352
rect 671120 715312 674012 715340
rect 671120 715300 671126 715312
rect 674006 715300 674012 715312
rect 674064 715300 674070 715352
rect 674282 715028 674288 715080
rect 674340 715068 674346 715080
rect 676030 715068 676036 715080
rect 674340 715040 676036 715068
rect 674340 715028 674346 715040
rect 676030 715028 676036 715040
rect 676088 715028 676094 715080
rect 660298 714960 660304 715012
rect 660356 715000 660362 715012
rect 674006 715000 674012 715012
rect 660356 714972 674012 715000
rect 660356 714960 660362 714972
rect 674006 714960 674012 714972
rect 674064 714960 674070 715012
rect 674282 714892 674288 714944
rect 674340 714932 674346 714944
rect 676030 714932 676036 714944
rect 674340 714904 676036 714932
rect 674340 714892 674346 714904
rect 676030 714892 676036 714904
rect 676088 714892 676094 714944
rect 672442 714824 672448 714876
rect 672500 714864 672506 714876
rect 674006 714864 674012 714876
rect 672500 714836 674012 714864
rect 672500 714824 672506 714836
rect 674006 714824 674012 714836
rect 674064 714824 674070 714876
rect 39298 714756 39304 714808
rect 39356 714796 39362 714808
rect 41598 714796 41604 714808
rect 39356 714768 41604 714796
rect 39356 714756 39362 714768
rect 41598 714756 41604 714768
rect 41656 714756 41662 714808
rect 671890 714484 671896 714536
rect 671948 714524 671954 714536
rect 674006 714524 674012 714536
rect 671948 714496 674012 714524
rect 671948 714484 671954 714496
rect 674006 714484 674012 714496
rect 674064 714484 674070 714536
rect 42058 714008 42064 714060
rect 42116 714048 42122 714060
rect 42610 714048 42616 714060
rect 42116 714020 42616 714048
rect 42116 714008 42122 714020
rect 42610 714008 42616 714020
rect 42668 714008 42674 714060
rect 672626 713668 672632 713720
rect 672684 713708 672690 713720
rect 674006 713708 674012 713720
rect 672684 713680 674012 713708
rect 672684 713668 672690 713680
rect 674006 713668 674012 713680
rect 674064 713668 674070 713720
rect 671062 713192 671068 713244
rect 671120 713232 671126 713244
rect 674006 713232 674012 713244
rect 671120 713204 674012 713232
rect 671120 713192 671126 713204
rect 674006 713192 674012 713204
rect 674064 713192 674070 713244
rect 671890 712376 671896 712428
rect 671948 712416 671954 712428
rect 674006 712416 674012 712428
rect 671948 712388 674012 712416
rect 671948 712376 671954 712388
rect 674006 712376 674012 712388
rect 674064 712376 674070 712428
rect 51718 712144 51724 712156
rect 42260 712116 51724 712144
rect 42260 711136 42288 712116
rect 51718 712104 51724 712116
rect 51776 712104 51782 712156
rect 42242 711084 42248 711136
rect 42300 711084 42306 711136
rect 671430 709996 671436 710048
rect 671488 710036 671494 710048
rect 674006 710036 674012 710048
rect 671488 710008 674012 710036
rect 671488 709996 671494 710008
rect 674006 709996 674012 710008
rect 674064 709996 674070 710048
rect 674282 709724 674288 709776
rect 674340 709764 674346 709776
rect 676030 709764 676036 709776
rect 674340 709736 676036 709764
rect 674340 709724 674346 709736
rect 676030 709724 676036 709736
rect 676088 709724 676094 709776
rect 43622 709316 43628 709368
rect 43680 709356 43686 709368
rect 45278 709356 45284 709368
rect 43680 709328 45284 709356
rect 43680 709316 43686 709328
rect 45278 709316 45284 709328
rect 45336 709316 45342 709368
rect 669038 709316 669044 709368
rect 669096 709356 669102 709368
rect 674006 709356 674012 709368
rect 669096 709328 674012 709356
rect 669096 709316 669102 709328
rect 674006 709316 674012 709328
rect 674064 709316 674070 709368
rect 670602 709180 670608 709232
rect 670660 709220 670666 709232
rect 674006 709220 674012 709232
rect 670660 709192 674012 709220
rect 670660 709180 670666 709192
rect 674006 709180 674012 709192
rect 674064 709180 674070 709232
rect 674282 708704 674288 708756
rect 674340 708744 674346 708756
rect 676030 708744 676036 708756
rect 674340 708716 676036 708744
rect 674340 708704 674346 708716
rect 676030 708704 676036 708716
rect 676088 708704 676094 708756
rect 669222 708228 669228 708280
rect 669280 708268 669286 708280
rect 674006 708268 674012 708280
rect 669280 708240 674012 708268
rect 669280 708228 669286 708240
rect 674006 708228 674012 708240
rect 674064 708228 674070 708280
rect 674466 707140 674472 707192
rect 674524 707180 674530 707192
rect 676030 707180 676036 707192
rect 674524 707152 676036 707180
rect 674524 707140 674530 707152
rect 676030 707140 676036 707152
rect 676088 707140 676094 707192
rect 42426 705508 42432 705560
rect 42484 705548 42490 705560
rect 43438 705548 43444 705560
rect 42484 705520 43444 705548
rect 42484 705508 42490 705520
rect 43438 705508 43444 705520
rect 43496 705508 43502 705560
rect 670418 705304 670424 705356
rect 670476 705344 670482 705356
rect 674006 705344 674012 705356
rect 670476 705316 674012 705344
rect 670476 705304 670482 705316
rect 674006 705304 674012 705316
rect 674064 705304 674070 705356
rect 674282 705304 674288 705356
rect 674340 705344 674346 705356
rect 683114 705344 683120 705356
rect 674340 705316 683120 705344
rect 674340 705304 674346 705316
rect 683114 705304 683120 705316
rect 683172 705304 683178 705356
rect 667842 705168 667848 705220
rect 667900 705208 667906 705220
rect 674006 705208 674012 705220
rect 667900 705180 674012 705208
rect 667900 705168 667906 705180
rect 674006 705168 674012 705180
rect 674064 705168 674070 705220
rect 674282 705168 674288 705220
rect 674340 705208 674346 705220
rect 675846 705208 675852 705220
rect 674340 705180 675852 705208
rect 674340 705168 674346 705180
rect 675846 705168 675852 705180
rect 675904 705168 675910 705220
rect 51718 705100 51724 705152
rect 51776 705140 51782 705152
rect 62114 705140 62120 705152
rect 51776 705112 62120 705140
rect 51776 705100 51782 705112
rect 62114 705100 62120 705112
rect 62172 705100 62178 705152
rect 674282 703876 674288 703928
rect 674340 703916 674346 703928
rect 676030 703916 676036 703928
rect 674340 703888 676036 703916
rect 674340 703876 674346 703888
rect 676030 703876 676036 703888
rect 676088 703876 676094 703928
rect 667014 703808 667020 703860
rect 667072 703848 667078 703860
rect 674006 703848 674012 703860
rect 667072 703820 674012 703848
rect 667072 703808 667078 703820
rect 674006 703808 674012 703820
rect 674064 703808 674070 703860
rect 44174 703740 44180 703792
rect 44232 703780 44238 703792
rect 62114 703780 62120 703792
rect 44232 703752 62120 703780
rect 44232 703740 44238 703752
rect 62114 703740 62120 703752
rect 62172 703740 62178 703792
rect 654778 701156 654784 701208
rect 654836 701196 654842 701208
rect 673730 701196 673736 701208
rect 654836 701168 673736 701196
rect 654836 701156 654842 701168
rect 673730 701156 673736 701168
rect 673788 701156 673794 701208
rect 42702 701020 42708 701072
rect 42760 701060 42766 701072
rect 62942 701060 62948 701072
rect 42760 701032 62948 701060
rect 42760 701020 42766 701032
rect 62942 701020 62948 701032
rect 63000 701020 63006 701072
rect 42058 699184 42064 699236
rect 42116 699224 42122 699236
rect 42518 699224 42524 699236
rect 42116 699196 42524 699224
rect 42116 699184 42122 699196
rect 42518 699184 42524 699196
rect 42576 699184 42582 699236
rect 46198 698232 46204 698284
rect 46256 698272 46262 698284
rect 62206 698272 62212 698284
rect 46256 698244 62212 698272
rect 46256 698232 46262 698244
rect 62206 698232 62212 698244
rect 62264 698232 62270 698284
rect 656526 690208 656532 690260
rect 656584 690248 656590 690260
rect 674006 690248 674012 690260
rect 656584 690220 674012 690248
rect 656584 690208 656590 690220
rect 674006 690208 674012 690220
rect 674064 690208 674070 690260
rect 674466 690004 674472 690056
rect 674524 690044 674530 690056
rect 675110 690044 675116 690056
rect 674524 690016 675116 690044
rect 674524 690004 674530 690016
rect 675110 690004 675116 690016
rect 675168 690004 675174 690056
rect 674926 688984 674932 689036
rect 674984 689024 674990 689036
rect 674984 688996 675156 689024
rect 674984 688984 674990 688996
rect 675128 688832 675156 688996
rect 652754 688780 652760 688832
rect 652812 688820 652818 688832
rect 672994 688820 673000 688832
rect 652812 688792 673000 688820
rect 652812 688780 652818 688792
rect 672994 688780 673000 688792
rect 673052 688780 673058 688832
rect 675110 688780 675116 688832
rect 675168 688780 675174 688832
rect 651466 688644 651472 688696
rect 651524 688684 651530 688696
rect 657538 688684 657544 688696
rect 651524 688656 657544 688684
rect 651524 688644 651530 688656
rect 657538 688644 657544 688656
rect 657596 688644 657602 688696
rect 43438 687488 43444 687540
rect 43496 687528 43502 687540
rect 61378 687528 61384 687540
rect 43496 687500 61384 687528
rect 43496 687488 43502 687500
rect 61378 687488 61384 687500
rect 61436 687488 61442 687540
rect 651466 687216 651472 687268
rect 651524 687256 651530 687268
rect 669958 687256 669964 687268
rect 651524 687228 669964 687256
rect 651524 687216 651530 687228
rect 669958 687216 669964 687228
rect 670016 687216 670022 687268
rect 651466 687012 651472 687064
rect 651524 687052 651530 687064
rect 654778 687052 654784 687064
rect 651524 687024 654784 687052
rect 651524 687012 651530 687024
rect 654778 687012 654784 687024
rect 654836 687012 654842 687064
rect 43438 686468 43444 686520
rect 43496 686508 43502 686520
rect 62942 686508 62948 686520
rect 43496 686480 62948 686508
rect 43496 686468 43502 686480
rect 62942 686468 62948 686480
rect 63000 686468 63006 686520
rect 651650 686468 651656 686520
rect 651708 686508 651714 686520
rect 667198 686508 667204 686520
rect 651708 686480 667204 686508
rect 651708 686468 651714 686480
rect 667198 686468 667204 686480
rect 667256 686468 667262 686520
rect 41322 686264 41328 686316
rect 41380 686304 41386 686316
rect 41690 686304 41696 686316
rect 41380 686276 41696 686304
rect 41380 686264 41386 686276
rect 41690 686264 41696 686276
rect 41748 686264 41754 686316
rect 42058 686264 42064 686316
rect 42116 686304 42122 686316
rect 42794 686304 42800 686316
rect 42116 686276 42800 686304
rect 42116 686264 42122 686276
rect 42794 686264 42800 686276
rect 42852 686264 42858 686316
rect 41138 686060 41144 686112
rect 41196 686100 41202 686112
rect 41690 686100 41696 686112
rect 41196 686072 41696 686100
rect 41196 686060 41202 686072
rect 41690 686060 41696 686072
rect 41748 686060 41754 686112
rect 42058 686060 42064 686112
rect 42116 686100 42122 686112
rect 43070 686100 43076 686112
rect 42116 686072 43076 686100
rect 42116 686060 42122 686072
rect 43070 686060 43076 686072
rect 43128 686060 43134 686112
rect 40954 685856 40960 685908
rect 41012 685896 41018 685908
rect 41690 685896 41696 685908
rect 41012 685868 41696 685896
rect 41012 685856 41018 685868
rect 41690 685856 41696 685868
rect 41748 685856 41754 685908
rect 42058 685856 42064 685908
rect 42116 685896 42122 685908
rect 45094 685896 45100 685908
rect 42116 685868 45100 685896
rect 42116 685856 42122 685868
rect 45094 685856 45100 685868
rect 45152 685856 45158 685908
rect 651466 685516 651472 685568
rect 651524 685556 651530 685568
rect 656526 685556 656532 685568
rect 651524 685528 656532 685556
rect 651524 685516 651530 685528
rect 656526 685516 656532 685528
rect 656584 685516 656590 685568
rect 674282 683952 674288 684004
rect 674340 683992 674346 684004
rect 674650 683992 674656 684004
rect 674340 683964 674656 683992
rect 674340 683952 674346 683964
rect 674650 683952 674656 683964
rect 674708 683952 674714 684004
rect 41322 683408 41328 683460
rect 41380 683448 41386 683460
rect 41690 683448 41696 683460
rect 41380 683420 41696 683448
rect 41380 683408 41386 683420
rect 41690 683408 41696 683420
rect 41748 683408 41754 683460
rect 675478 682524 675484 682576
rect 675536 682564 675542 682576
rect 683206 682564 683212 682576
rect 675536 682536 683212 682564
rect 675536 682524 675542 682536
rect 683206 682524 683212 682536
rect 683264 682524 683270 682576
rect 674742 682388 674748 682440
rect 674800 682428 674806 682440
rect 683482 682428 683488 682440
rect 674800 682400 683488 682428
rect 674800 682388 674806 682400
rect 683482 682388 683488 682400
rect 683540 682388 683546 682440
rect 40770 678580 40776 678632
rect 40828 678620 40834 678632
rect 41690 678620 41696 678632
rect 40828 678592 41696 678620
rect 40828 678580 40834 678592
rect 41690 678580 41696 678592
rect 41748 678580 41754 678632
rect 40770 677696 40776 677748
rect 40828 677736 40834 677748
rect 41598 677736 41604 677748
rect 40828 677708 41604 677736
rect 40828 677696 40834 677708
rect 41598 677696 41604 677708
rect 41656 677696 41662 677748
rect 42426 676200 42432 676252
rect 42484 676240 42490 676252
rect 59998 676240 60004 676252
rect 42484 676212 60004 676240
rect 42484 676200 42490 676212
rect 59998 676200 60004 676212
rect 60056 676200 60062 676252
rect 33042 674092 33048 674144
rect 33100 674132 33106 674144
rect 41414 674132 41420 674144
rect 33100 674104 41420 674132
rect 33100 674092 33106 674104
rect 41414 674092 41420 674104
rect 41472 674092 41478 674144
rect 35158 672732 35164 672784
rect 35216 672772 35222 672784
rect 41598 672772 41604 672784
rect 35216 672744 41604 672772
rect 35216 672732 35222 672744
rect 41598 672732 41604 672744
rect 41656 672732 41662 672784
rect 42610 671304 42616 671356
rect 42668 671304 42674 671356
rect 673546 671304 673552 671356
rect 673604 671344 673610 671356
rect 673604 671316 673776 671344
rect 673604 671304 673610 671316
rect 42628 671220 42656 671304
rect 42610 671168 42616 671220
rect 42668 671168 42674 671220
rect 668578 671100 668584 671152
rect 668636 671140 668642 671152
rect 673546 671140 673552 671152
rect 668636 671112 673552 671140
rect 668636 671100 668642 671112
rect 673546 671100 673552 671112
rect 673604 671100 673610 671152
rect 36538 670964 36544 671016
rect 36596 671004 36602 671016
rect 40494 671004 40500 671016
rect 36596 670976 40500 671004
rect 36596 670964 36602 670976
rect 40494 670964 40500 670976
rect 40552 670964 40558 671016
rect 661678 670692 661684 670744
rect 661736 670732 661742 670744
rect 673748 670732 673776 671316
rect 661736 670704 673776 670732
rect 661736 670692 661742 670704
rect 672442 670556 672448 670608
rect 672500 670596 672506 670608
rect 673362 670596 673368 670608
rect 672500 670568 673368 670596
rect 672500 670556 672506 670568
rect 673362 670556 673368 670568
rect 673420 670556 673426 670608
rect 670234 669604 670240 669656
rect 670292 669644 670298 669656
rect 673362 669644 673368 669656
rect 670292 669616 673368 669644
rect 670292 669604 670298 669616
rect 673362 669604 673368 669616
rect 673420 669604 673426 669656
rect 658918 669468 658924 669520
rect 658976 669508 658982 669520
rect 673546 669508 673552 669520
rect 658976 669480 673552 669508
rect 658976 669468 658982 669480
rect 673546 669468 673552 669480
rect 673604 669468 673610 669520
rect 674834 669468 674840 669520
rect 674892 669508 674898 669520
rect 676490 669508 676496 669520
rect 674892 669480 676496 669508
rect 674892 669468 674898 669480
rect 676490 669468 676496 669480
rect 676548 669468 676554 669520
rect 42426 669332 42432 669384
rect 42484 669372 42490 669384
rect 57238 669372 57244 669384
rect 42484 669344 57244 669372
rect 42484 669332 42490 669344
rect 57238 669332 57244 669344
rect 57296 669332 57302 669384
rect 673546 668652 673552 668704
rect 673604 668692 673610 668704
rect 673604 668664 673776 668692
rect 673604 668652 673610 668664
rect 671062 668516 671068 668568
rect 671120 668556 671126 668568
rect 673546 668556 673552 668568
rect 671120 668528 673552 668556
rect 671120 668516 671126 668528
rect 673546 668516 673552 668528
rect 673604 668516 673610 668568
rect 671062 668108 671068 668160
rect 671120 668148 671126 668160
rect 673546 668148 673552 668160
rect 671120 668120 673552 668148
rect 671120 668108 671126 668120
rect 673546 668108 673552 668120
rect 673604 668108 673610 668160
rect 44542 667904 44548 667956
rect 44600 667944 44606 667956
rect 58618 667944 58624 667956
rect 44600 667916 58624 667944
rect 44600 667904 44606 667916
rect 58618 667904 58624 667916
rect 58676 667904 58682 667956
rect 671430 667904 671436 667956
rect 671488 667944 671494 667956
rect 673748 667944 673776 668664
rect 671488 667916 673776 667944
rect 671488 667904 671494 667916
rect 674834 667020 674840 667072
rect 674892 667060 674898 667072
rect 676490 667060 676496 667072
rect 674892 667032 676496 667060
rect 674892 667020 674898 667032
rect 676490 667020 676496 667032
rect 676548 667020 676554 667072
rect 671890 666884 671896 666936
rect 671948 666924 671954 666936
rect 673546 666924 673552 666936
rect 671948 666896 673552 666924
rect 671948 666884 671954 666896
rect 673546 666884 673552 666896
rect 673604 666884 673610 666936
rect 671890 666544 671896 666596
rect 671948 666584 671954 666596
rect 673546 666584 673552 666596
rect 671948 666556 673552 666584
rect 671948 666544 671954 666556
rect 673546 666544 673552 666556
rect 673604 666544 673610 666596
rect 42242 665796 42248 665848
rect 42300 665836 42306 665848
rect 44542 665836 44548 665848
rect 42300 665808 44548 665836
rect 42300 665796 42306 665808
rect 44542 665796 44548 665808
rect 44600 665796 44606 665848
rect 669590 665252 669596 665304
rect 669648 665292 669654 665304
rect 673546 665292 673552 665304
rect 669648 665264 673552 665292
rect 669648 665252 669654 665264
rect 673546 665252 673552 665264
rect 673604 665252 673610 665304
rect 672258 665116 672264 665168
rect 672316 665156 672322 665168
rect 673362 665156 673368 665168
rect 672316 665128 673368 665156
rect 672316 665116 672322 665128
rect 673362 665116 673368 665128
rect 673420 665116 673426 665168
rect 671706 664368 671712 664420
rect 671764 664408 671770 664420
rect 673546 664408 673552 664420
rect 671764 664380 673552 664408
rect 671764 664368 671770 664380
rect 673546 664368 673552 664380
rect 673604 664368 673610 664420
rect 669406 663892 669412 663944
rect 669464 663932 669470 663944
rect 673546 663932 673552 663944
rect 669464 663904 673552 663932
rect 669464 663892 669470 663904
rect 673546 663892 673552 663904
rect 673604 663892 673610 663944
rect 42610 663756 42616 663808
rect 42668 663756 42674 663808
rect 674834 663756 674840 663808
rect 674892 663796 674898 663808
rect 676030 663796 676036 663808
rect 674892 663768 676036 663796
rect 674892 663756 674898 663768
rect 676030 663756 676036 663768
rect 676088 663756 676094 663808
rect 42628 663604 42656 663756
rect 42610 663552 42616 663604
rect 42668 663552 42674 663604
rect 42242 663416 42248 663468
rect 42300 663456 42306 663468
rect 42794 663456 42800 663468
rect 42300 663428 42800 663456
rect 42300 663416 42306 663428
rect 42794 663416 42800 663428
rect 42852 663416 42858 663468
rect 673546 663348 673552 663400
rect 673604 663388 673610 663400
rect 673914 663388 673920 663400
rect 673604 663360 673920 663388
rect 673604 663348 673610 663360
rect 673914 663348 673920 663360
rect 673972 663348 673978 663400
rect 42242 663008 42248 663060
rect 42300 663048 42306 663060
rect 43990 663048 43996 663060
rect 42300 663020 43996 663048
rect 42300 663008 42306 663020
rect 43990 663008 43996 663020
rect 44048 663008 44054 663060
rect 672074 662396 672080 662448
rect 672132 662436 672138 662448
rect 673914 662436 673920 662448
rect 672132 662408 673920 662436
rect 672132 662396 672138 662408
rect 673914 662396 673920 662408
rect 673972 662396 673978 662448
rect 671246 661580 671252 661632
rect 671304 661620 671310 661632
rect 673914 661620 673920 661632
rect 671304 661592 673920 661620
rect 671304 661580 671310 661592
rect 673914 661580 673920 661592
rect 673972 661580 673978 661632
rect 669222 661104 669228 661156
rect 669280 661144 669286 661156
rect 673914 661144 673920 661156
rect 669280 661116 673920 661144
rect 669280 661104 669286 661116
rect 673914 661104 673920 661116
rect 673972 661104 673978 661156
rect 57238 660900 57244 660952
rect 57296 660940 57302 660952
rect 62114 660940 62120 660952
rect 57296 660912 62120 660940
rect 57296 660900 57302 660912
rect 62114 660900 62120 660912
rect 62172 660900 62178 660952
rect 42150 660492 42156 660544
rect 42208 660532 42214 660544
rect 43622 660532 43628 660544
rect 42208 660504 43628 660532
rect 42208 660492 42214 660504
rect 43622 660492 43628 660504
rect 43680 660492 43686 660544
rect 668854 660084 668860 660136
rect 668912 660124 668918 660136
rect 673914 660124 673920 660136
rect 668912 660096 673920 660124
rect 668912 660084 668918 660096
rect 673914 660084 673920 660096
rect 673972 660084 673978 660136
rect 674834 659812 674840 659864
rect 674892 659852 674898 659864
rect 683114 659852 683120 659864
rect 674892 659824 683120 659852
rect 674892 659812 674898 659824
rect 683114 659812 683120 659824
rect 683172 659812 683178 659864
rect 58618 659540 58624 659592
rect 58676 659580 58682 659592
rect 62114 659580 62120 659592
rect 58676 659552 62120 659580
rect 58676 659540 58682 659552
rect 62114 659540 62120 659552
rect 62172 659540 62178 659592
rect 42150 658996 42156 659048
rect 42208 659036 42214 659048
rect 42610 659036 42616 659048
rect 42208 659008 42616 659036
rect 42208 658996 42214 659008
rect 42610 658996 42616 659008
rect 42668 658996 42674 659048
rect 42518 657500 42524 657552
rect 42576 657540 42582 657552
rect 62114 657540 62120 657552
rect 42576 657512 62120 657540
rect 42576 657500 42582 657512
rect 62114 657500 62120 657512
rect 62172 657500 62178 657552
rect 653398 655528 653404 655580
rect 653456 655568 653462 655580
rect 673914 655568 673920 655580
rect 653456 655540 673920 655568
rect 653456 655528 653462 655540
rect 673914 655528 673920 655540
rect 673972 655528 673978 655580
rect 45462 655460 45468 655512
rect 45520 655500 45526 655512
rect 62114 655500 62120 655512
rect 45520 655472 62120 655500
rect 45520 655460 45526 655472
rect 62114 655460 62120 655472
rect 62172 655460 62178 655512
rect 655514 645872 655520 645924
rect 655572 645912 655578 645924
rect 674006 645912 674012 645924
rect 655572 645884 674012 645912
rect 655572 645872 655578 645884
rect 674006 645872 674012 645884
rect 674064 645872 674070 645924
rect 674558 644580 674564 644632
rect 674616 644620 674622 644632
rect 675294 644620 675300 644632
rect 674616 644592 675300 644620
rect 674616 644580 674622 644592
rect 675294 644580 675300 644592
rect 675352 644580 675358 644632
rect 35802 644444 35808 644496
rect 35860 644484 35866 644496
rect 40126 644484 40132 644496
rect 35860 644456 40132 644484
rect 35860 644444 35866 644456
rect 40126 644444 40132 644456
rect 40184 644444 40190 644496
rect 35802 643492 35808 643544
rect 35860 643532 35866 643544
rect 40586 643532 40592 643544
rect 35860 643504 40592 643532
rect 35860 643492 35866 643504
rect 40586 643492 40592 643504
rect 40644 643492 40650 643544
rect 41690 643328 41696 643340
rect 41386 643300 41696 643328
rect 35526 643220 35532 643272
rect 35584 643260 35590 643272
rect 41386 643260 41414 643300
rect 41690 643288 41696 643300
rect 41748 643288 41754 643340
rect 42058 643288 42064 643340
rect 42116 643328 42122 643340
rect 45094 643328 45100 643340
rect 42116 643300 45100 643328
rect 42116 643288 42122 643300
rect 45094 643288 45100 643300
rect 45152 643288 45158 643340
rect 35584 643232 41414 643260
rect 35584 643220 35590 643232
rect 35342 643084 35348 643136
rect 35400 643124 35406 643136
rect 41690 643124 41696 643136
rect 35400 643096 41696 643124
rect 35400 643084 35406 643096
rect 41690 643084 41696 643096
rect 41748 643084 41754 643136
rect 42058 643084 42064 643136
rect 42116 643124 42122 643136
rect 61378 643124 61384 643136
rect 42116 643096 61384 643124
rect 42116 643084 42122 643096
rect 61378 643084 61384 643096
rect 61436 643084 61442 643136
rect 655330 643084 655336 643136
rect 655388 643124 655394 643136
rect 674006 643124 674012 643136
rect 655388 643096 674012 643124
rect 655388 643084 655394 643096
rect 674006 643084 674012 643096
rect 674064 643084 674070 643136
rect 38562 642472 38568 642524
rect 38620 642512 38626 642524
rect 41690 642512 41696 642524
rect 38620 642484 41696 642512
rect 38620 642472 38626 642484
rect 41690 642472 41696 642484
rect 41748 642472 41754 642524
rect 42058 642336 42064 642388
rect 42116 642376 42122 642388
rect 62942 642376 62948 642388
rect 42116 642348 62948 642376
rect 42116 642336 42122 642348
rect 62942 642336 62948 642348
rect 63000 642336 63006 642388
rect 651466 642336 651472 642388
rect 651524 642376 651530 642388
rect 658918 642376 658924 642388
rect 651524 642348 658924 642376
rect 651524 642336 651530 642348
rect 658918 642336 658924 642348
rect 658976 642336 658982 642388
rect 35802 642132 35808 642184
rect 35860 642172 35866 642184
rect 40310 642172 40316 642184
rect 35860 642144 40316 642172
rect 35860 642132 35866 642144
rect 40310 642132 40316 642144
rect 40368 642132 40374 642184
rect 35434 641860 35440 641912
rect 35492 641900 35498 641912
rect 39942 641900 39948 641912
rect 35492 641872 39948 641900
rect 35492 641860 35498 641872
rect 39942 641860 39948 641872
rect 40000 641860 40006 641912
rect 35618 641724 35624 641776
rect 35676 641764 35682 641776
rect 41690 641764 41696 641776
rect 35676 641736 41696 641764
rect 35676 641724 35682 641736
rect 41690 641724 41696 641736
rect 41748 641724 41754 641776
rect 42058 641724 42064 641776
rect 42116 641764 42122 641776
rect 44358 641764 44364 641776
rect 42116 641736 44364 641764
rect 42116 641724 42122 641736
rect 44358 641724 44364 641736
rect 44416 641724 44422 641776
rect 674742 641044 674748 641096
rect 674800 641044 674806 641096
rect 674760 640892 674788 641044
rect 674742 640840 674748 640892
rect 674800 640840 674806 640892
rect 35802 640704 35808 640756
rect 35860 640744 35866 640756
rect 39942 640744 39948 640756
rect 35860 640716 39948 640744
rect 35860 640704 35866 640716
rect 39942 640704 39948 640716
rect 40000 640704 40006 640756
rect 42058 640500 42064 640552
rect 42116 640540 42122 640552
rect 42978 640540 42984 640552
rect 42116 640512 42984 640540
rect 42116 640500 42122 640512
rect 42978 640500 42984 640512
rect 43036 640500 43042 640552
rect 35526 640432 35532 640484
rect 35584 640472 35590 640484
rect 41690 640472 41696 640484
rect 35584 640444 41696 640472
rect 35584 640432 35590 640444
rect 41690 640432 41696 640444
rect 41748 640432 41754 640484
rect 35342 640296 35348 640348
rect 35400 640336 35406 640348
rect 41690 640336 41696 640348
rect 35400 640308 41696 640336
rect 35400 640296 35406 640308
rect 41690 640296 41696 640308
rect 41748 640296 41754 640348
rect 42058 640296 42064 640348
rect 42116 640336 42122 640348
rect 45462 640336 45468 640348
rect 42116 640308 45468 640336
rect 42116 640296 42122 640308
rect 45462 640296 45468 640308
rect 45520 640296 45526 640348
rect 651466 640296 651472 640348
rect 651524 640336 651530 640348
rect 668578 640336 668584 640348
rect 651524 640308 668584 640336
rect 651524 640296 651530 640308
rect 668578 640296 668584 640308
rect 668636 640296 668642 640348
rect 675202 640228 675208 640280
rect 675260 640228 675266 640280
rect 674834 640160 674840 640212
rect 674892 640160 674898 640212
rect 651374 640092 651380 640144
rect 651432 640132 651438 640144
rect 653398 640132 653404 640144
rect 651432 640104 653404 640132
rect 651432 640092 651438 640104
rect 653398 640092 653404 640104
rect 653456 640092 653462 640144
rect 674852 639804 674880 640160
rect 675018 639888 675024 639940
rect 675076 639928 675082 639940
rect 675220 639928 675248 640228
rect 675076 639900 675248 639928
rect 675076 639888 675082 639900
rect 674834 639752 674840 639804
rect 674892 639752 674898 639804
rect 35802 639140 35808 639192
rect 35860 639180 35866 639192
rect 35860 639140 35894 639180
rect 35866 639112 35894 639140
rect 39298 639112 39304 639124
rect 35866 639084 39304 639112
rect 39298 639072 39304 639084
rect 39356 639072 39362 639124
rect 35802 638936 35808 638988
rect 35860 638976 35866 638988
rect 40034 638976 40040 638988
rect 35860 638948 40040 638976
rect 35860 638936 35866 638948
rect 40034 638936 40040 638948
rect 40092 638936 40098 638988
rect 651650 638868 651656 638920
rect 651708 638908 651714 638920
rect 655330 638908 655336 638920
rect 651708 638880 655336 638908
rect 651708 638868 651714 638880
rect 655330 638868 655336 638880
rect 655388 638868 655394 638920
rect 651466 638732 651472 638784
rect 651524 638772 651530 638784
rect 655514 638772 655520 638784
rect 651524 638744 655520 638772
rect 651524 638732 651530 638744
rect 655514 638732 655520 638744
rect 655572 638732 655578 638784
rect 34422 638188 34428 638240
rect 34480 638228 34486 638240
rect 41690 638228 41696 638240
rect 34480 638200 41696 638228
rect 34480 638188 34486 638200
rect 41690 638188 41696 638200
rect 41748 638188 41754 638240
rect 674742 637712 674748 637764
rect 674800 637712 674806 637764
rect 674760 637628 674788 637712
rect 35802 637576 35808 637628
rect 35860 637616 35866 637628
rect 36538 637616 36544 637628
rect 35860 637588 36544 637616
rect 35860 637576 35866 637588
rect 36538 637576 36544 637588
rect 36596 637576 36602 637628
rect 674742 637576 674748 637628
rect 674800 637576 674806 637628
rect 674282 637440 674288 637492
rect 674340 637480 674346 637492
rect 675478 637480 675484 637492
rect 674340 637452 675484 637480
rect 674340 637440 674346 637452
rect 675478 637440 675484 637452
rect 675536 637440 675542 637492
rect 674742 637032 674748 637084
rect 674800 637072 674806 637084
rect 683206 637072 683212 637084
rect 674800 637044 683212 637072
rect 674800 637032 674806 637044
rect 683206 637032 683212 637044
rect 683264 637032 683270 637084
rect 35618 636828 35624 636880
rect 35676 636868 35682 636880
rect 40310 636868 40316 636880
rect 35676 636840 40316 636868
rect 35676 636828 35682 636840
rect 40310 636828 40316 636840
rect 40368 636828 40374 636880
rect 675478 636828 675484 636880
rect 675536 636868 675542 636880
rect 683390 636868 683396 636880
rect 675536 636840 683396 636868
rect 675536 636828 675542 636840
rect 683390 636828 683396 636840
rect 683448 636828 683454 636880
rect 35802 636692 35808 636744
rect 35860 636732 35866 636744
rect 35860 636692 35894 636732
rect 35866 636664 35894 636692
rect 40862 636664 40868 636676
rect 35866 636636 40868 636664
rect 40862 636624 40868 636636
rect 40920 636624 40926 636676
rect 35802 636352 35808 636404
rect 35860 636392 35866 636404
rect 40494 636392 40500 636404
rect 35860 636364 40500 636392
rect 35860 636352 35866 636364
rect 40494 636352 40500 636364
rect 40552 636352 40558 636404
rect 35526 636216 35532 636268
rect 35584 636256 35590 636268
rect 35584 636228 38654 636256
rect 35584 636216 35590 636228
rect 38626 636188 38654 636228
rect 39114 636188 39120 636200
rect 38626 636160 39120 636188
rect 39114 636148 39120 636160
rect 39172 636148 39178 636200
rect 674926 635468 674932 635520
rect 674984 635508 674990 635520
rect 675662 635508 675668 635520
rect 674984 635480 675668 635508
rect 674984 635468 674990 635480
rect 675662 635468 675668 635480
rect 675720 635468 675726 635520
rect 35802 634788 35808 634840
rect 35860 634828 35866 634840
rect 40494 634828 40500 634840
rect 35860 634800 40500 634828
rect 35860 634788 35866 634800
rect 40494 634788 40500 634800
rect 40552 634788 40558 634840
rect 652018 634040 652024 634092
rect 652076 634080 652082 634092
rect 660298 634080 660304 634092
rect 652076 634052 660304 634080
rect 652076 634040 652082 634052
rect 660298 634040 660304 634052
rect 660356 634040 660362 634092
rect 35802 633836 35808 633888
rect 35860 633876 35866 633888
rect 35860 633836 35894 633876
rect 35866 633740 35894 633836
rect 39758 633740 39764 633752
rect 35866 633712 39764 633740
rect 39758 633700 39764 633712
rect 39816 633700 39822 633752
rect 35802 633428 35808 633480
rect 35860 633468 35866 633480
rect 41506 633468 41512 633480
rect 35860 633440 41512 633468
rect 35860 633428 35866 633440
rect 41506 633428 41512 633440
rect 41564 633428 41570 633480
rect 42058 633428 42064 633480
rect 42116 633468 42122 633480
rect 60182 633468 60188 633480
rect 42116 633440 60188 633468
rect 42116 633428 42122 633440
rect 60182 633428 60188 633440
rect 60240 633428 60246 633480
rect 36538 630572 36544 630624
rect 36596 630612 36602 630624
rect 36596 630584 41414 630612
rect 36596 630572 36602 630584
rect 41386 630544 41414 630584
rect 41598 630544 41604 630556
rect 41386 630516 41604 630544
rect 41598 630504 41604 630516
rect 41656 630504 41662 630556
rect 671522 628736 671528 628788
rect 671580 628736 671586 628788
rect 35158 628532 35164 628584
rect 35216 628572 35222 628584
rect 40494 628572 40500 628584
rect 35216 628544 40500 628572
rect 35216 628532 35222 628544
rect 40494 628532 40500 628544
rect 40552 628532 40558 628584
rect 671338 628396 671344 628448
rect 671396 628436 671402 628448
rect 671540 628436 671568 628736
rect 671396 628408 671568 628436
rect 671396 628396 671402 628408
rect 669958 625948 669964 626000
rect 670016 625988 670022 626000
rect 673546 625988 673552 626000
rect 670016 625960 673552 625988
rect 670016 625948 670022 625960
rect 673546 625948 673552 625960
rect 673604 625948 673610 626000
rect 44174 625812 44180 625864
rect 44232 625852 44238 625864
rect 63126 625852 63132 625864
rect 44232 625824 63132 625852
rect 44232 625812 44238 625824
rect 63126 625812 63132 625824
rect 63184 625812 63190 625864
rect 667198 625676 667204 625728
rect 667256 625716 667262 625728
rect 674006 625716 674012 625728
rect 667256 625688 674012 625716
rect 667256 625676 667262 625688
rect 674006 625676 674012 625688
rect 674064 625676 674070 625728
rect 674742 625676 674748 625728
rect 674800 625716 674806 625728
rect 676490 625716 676496 625728
rect 674800 625688 676496 625716
rect 674800 625676 674806 625688
rect 676490 625676 676496 625688
rect 676548 625676 676554 625728
rect 657538 625132 657544 625184
rect 657596 625172 657602 625184
rect 674006 625172 674012 625184
rect 657596 625144 674012 625172
rect 657596 625132 657602 625144
rect 674006 625132 674012 625144
rect 674064 625132 674070 625184
rect 670234 624996 670240 625048
rect 670292 625036 670298 625048
rect 674006 625036 674012 625048
rect 670292 625008 674012 625036
rect 670292 624996 670298 625008
rect 674006 624996 674012 625008
rect 674064 624996 674070 625048
rect 42242 624656 42248 624708
rect 42300 624696 42306 624708
rect 44174 624696 44180 624708
rect 42300 624668 44180 624696
rect 42300 624656 42306 624668
rect 44174 624656 44180 624668
rect 44232 624656 44238 624708
rect 670234 624656 670240 624708
rect 670292 624696 670298 624708
rect 674006 624696 674012 624708
rect 670292 624668 674012 624696
rect 670292 624656 670298 624668
rect 674006 624656 674012 624668
rect 674064 624656 674070 624708
rect 671430 624316 671436 624368
rect 671488 624356 671494 624368
rect 674006 624356 674012 624368
rect 671488 624328 674012 624356
rect 671488 624316 671494 624328
rect 674006 624316 674012 624328
rect 674064 624316 674070 624368
rect 42242 624044 42248 624096
rect 42300 624084 42306 624096
rect 44358 624084 44364 624096
rect 42300 624056 44364 624084
rect 42300 624044 42306 624056
rect 44358 624044 44364 624056
rect 44416 624044 44422 624096
rect 669406 623840 669412 623892
rect 669464 623880 669470 623892
rect 674006 623880 674012 623892
rect 669464 623852 674012 623880
rect 669464 623840 669470 623852
rect 674006 623840 674012 623852
rect 674064 623840 674070 623892
rect 671062 623500 671068 623552
rect 671120 623540 671126 623552
rect 674006 623540 674012 623552
rect 671120 623512 674012 623540
rect 671120 623500 671126 623512
rect 674006 623500 674012 623512
rect 674064 623500 674070 623552
rect 670418 623024 670424 623076
rect 670476 623064 670482 623076
rect 674006 623064 674012 623076
rect 670476 623036 674012 623064
rect 670476 623024 670482 623036
rect 674006 623024 674012 623036
rect 674064 623024 674070 623076
rect 674374 623024 674380 623076
rect 674432 623064 674438 623076
rect 683390 623064 683396 623076
rect 674432 623036 683396 623064
rect 674432 623024 674438 623036
rect 683390 623024 683396 623036
rect 683448 623024 683454 623076
rect 671890 622684 671896 622736
rect 671948 622724 671954 622736
rect 674006 622724 674012 622736
rect 671948 622696 674012 622724
rect 671948 622684 671954 622696
rect 674006 622684 674012 622696
rect 674064 622684 674070 622736
rect 671430 622208 671436 622260
rect 671488 622248 671494 622260
rect 674006 622248 674012 622260
rect 671488 622220 674012 622248
rect 671488 622208 671494 622220
rect 674006 622208 674012 622220
rect 674064 622208 674070 622260
rect 42242 621664 42248 621716
rect 42300 621704 42306 621716
rect 44174 621704 44180 621716
rect 42300 621676 44180 621704
rect 42300 621664 42306 621676
rect 44174 621664 44180 621676
rect 44232 621664 44238 621716
rect 667658 621596 667664 621648
rect 667716 621636 667722 621648
rect 674006 621636 674012 621648
rect 667716 621608 674012 621636
rect 667716 621596 667722 621608
rect 674006 621596 674012 621608
rect 674064 621596 674070 621648
rect 42242 621528 42248 621580
rect 42300 621568 42306 621580
rect 43990 621568 43996 621580
rect 42300 621540 43996 621568
rect 42300 621528 42306 621540
rect 43990 621528 43996 621540
rect 44048 621528 44054 621580
rect 670878 620644 670884 620696
rect 670936 620684 670942 620696
rect 672534 620684 672540 620696
rect 670936 620656 672540 620684
rect 670936 620644 670942 620656
rect 672534 620644 672540 620656
rect 672592 620644 672598 620696
rect 42242 620372 42248 620424
rect 42300 620412 42306 620424
rect 42702 620412 42708 620424
rect 42300 620384 42708 620412
rect 42300 620372 42306 620384
rect 42702 620372 42708 620384
rect 42760 620372 42766 620424
rect 669038 620372 669044 620424
rect 669096 620412 669102 620424
rect 673638 620412 673644 620424
rect 669096 620384 673644 620412
rect 669096 620372 669102 620384
rect 673638 620372 673644 620384
rect 673696 620372 673702 620424
rect 669774 619828 669780 619880
rect 669832 619868 669838 619880
rect 673638 619868 673644 619880
rect 669832 619840 673644 619868
rect 669832 619828 669838 619840
rect 673638 619828 673644 619840
rect 673696 619828 673702 619880
rect 42242 619624 42248 619676
rect 42300 619664 42306 619676
rect 42886 619664 42892 619676
rect 42300 619636 42892 619664
rect 42300 619624 42306 619636
rect 42886 619624 42892 619636
rect 42944 619624 42950 619676
rect 668210 617924 668216 617976
rect 668268 617964 668274 617976
rect 673638 617964 673644 617976
rect 668268 617936 673644 617964
rect 668268 617924 668274 617936
rect 673638 617924 673644 617936
rect 673696 617924 673702 617976
rect 674282 617516 674288 617568
rect 674340 617556 674346 617568
rect 676214 617556 676220 617568
rect 674340 617528 676220 617556
rect 674340 617516 674346 617528
rect 676214 617516 676220 617528
rect 676272 617516 676278 617568
rect 42242 617312 42248 617364
rect 42300 617352 42306 617364
rect 43070 617352 43076 617364
rect 42300 617324 43076 617352
rect 42300 617312 42306 617324
rect 43070 617312 43076 617324
rect 43128 617312 43134 617364
rect 668394 616836 668400 616888
rect 668452 616876 668458 616888
rect 673638 616876 673644 616888
rect 668452 616848 673644 616876
rect 668452 616836 668458 616848
rect 673638 616836 673644 616848
rect 673696 616836 673702 616888
rect 44174 616768 44180 616820
rect 44232 616808 44238 616820
rect 62114 616808 62120 616820
rect 44232 616780 62120 616808
rect 44232 616768 44238 616780
rect 62114 616768 62120 616780
rect 62172 616768 62178 616820
rect 670602 615476 670608 615528
rect 670660 615516 670666 615528
rect 673638 615516 673644 615528
rect 670660 615488 673644 615516
rect 670660 615476 670666 615488
rect 673638 615476 673644 615488
rect 673696 615476 673702 615528
rect 674282 615476 674288 615528
rect 674340 615516 674346 615528
rect 683114 615516 683120 615528
rect 674340 615488 683120 615516
rect 674340 615476 674346 615488
rect 683114 615476 683120 615488
rect 683172 615476 683178 615528
rect 670602 614864 670608 614916
rect 670660 614904 670666 614916
rect 673638 614904 673644 614916
rect 670660 614876 673644 614904
rect 670660 614864 670666 614876
rect 673638 614864 673644 614876
rect 673696 614864 673702 614916
rect 42702 614116 42708 614168
rect 42760 614156 42766 614168
rect 62114 614156 62120 614168
rect 42760 614128 62120 614156
rect 42760 614116 42766 614128
rect 62114 614116 62120 614128
rect 62172 614116 62178 614168
rect 46198 613368 46204 613420
rect 46256 613408 46262 613420
rect 62114 613408 62120 613420
rect 46256 613380 62120 613408
rect 46256 613368 46262 613380
rect 62114 613368 62120 613380
rect 62172 613368 62178 613420
rect 43806 612660 43812 612672
rect 43663 612632 43812 612660
rect 42242 612348 42248 612400
rect 42300 612388 42306 612400
rect 42300 612360 43562 612388
rect 42300 612348 42306 612360
rect 43663 612306 43691 612632
rect 43806 612620 43812 612632
rect 43864 612620 43870 612672
rect 43990 612212 43996 612264
rect 44048 612252 44054 612264
rect 44726 612252 44732 612264
rect 44048 612224 44732 612252
rect 44048 612212 44054 612224
rect 44726 612212 44732 612224
rect 44784 612212 44790 612264
rect 44082 612116 44088 612128
rect 43792 612088 44088 612116
rect 44082 612076 44088 612088
rect 44140 612076 44146 612128
rect 43875 611992 43927 611998
rect 43875 611934 43927 611940
rect 44266 611708 44272 611720
rect 44022 611680 44272 611708
rect 44266 611668 44272 611680
rect 44324 611668 44330 611720
rect 44910 611572 44916 611584
rect 44114 611544 44916 611572
rect 44910 611532 44916 611544
rect 44968 611532 44974 611584
rect 653398 611328 653404 611380
rect 653456 611368 653462 611380
rect 673638 611368 673644 611380
rect 653456 611340 673644 611368
rect 653456 611328 653462 611340
rect 673638 611328 673644 611340
rect 673696 611328 673702 611380
rect 50154 611300 50160 611312
rect 44237 611272 50160 611300
rect 50154 611260 50160 611272
rect 50212 611260 50218 611312
rect 44312 611124 44318 611176
rect 44370 611124 44376 611176
rect 44461 610864 45554 610892
rect 44726 610756 44732 610768
rect 44574 610728 44732 610756
rect 44726 610716 44732 610728
rect 44784 610716 44790 610768
rect 45526 610008 45554 610864
rect 50154 610104 50160 610156
rect 50212 610144 50218 610156
rect 58618 610144 58624 610156
rect 50212 610116 58624 610144
rect 50212 610104 50218 610116
rect 58618 610104 58624 610116
rect 58676 610104 58682 610156
rect 61378 610008 61384 610020
rect 45526 609980 61384 610008
rect 61378 609968 61384 609980
rect 61436 609968 61442 610020
rect 667658 608608 667664 608660
rect 667716 608648 667722 608660
rect 673178 608648 673184 608660
rect 667716 608620 673184 608648
rect 667716 608608 667722 608620
rect 673178 608608 673184 608620
rect 673236 608608 673242 608660
rect 674282 608336 674288 608388
rect 674340 608376 674346 608388
rect 675478 608376 675484 608388
rect 674340 608348 675484 608376
rect 674340 608336 674346 608348
rect 675478 608336 675484 608348
rect 675536 608336 675542 608388
rect 674282 603236 674288 603288
rect 674340 603276 674346 603288
rect 675110 603276 675116 603288
rect 674340 603248 675116 603276
rect 674340 603236 674346 603248
rect 675110 603236 675116 603248
rect 675168 603236 675174 603288
rect 35802 601672 35808 601724
rect 35860 601712 35866 601724
rect 36538 601712 36544 601724
rect 35860 601684 36544 601712
rect 35860 601672 35866 601684
rect 36538 601672 36544 601684
rect 36596 601672 36602 601724
rect 657538 600448 657544 600500
rect 657596 600488 657602 600500
rect 657596 600460 669314 600488
rect 657596 600448 657602 600460
rect 669286 600420 669314 600460
rect 673822 600420 673828 600432
rect 669286 600392 673828 600420
rect 673822 600380 673828 600392
rect 673880 600380 673886 600432
rect 654778 598952 654784 599004
rect 654836 598992 654842 599004
rect 673178 598992 673184 599004
rect 654836 598964 673184 598992
rect 654836 598952 654842 598964
rect 673178 598952 673184 598964
rect 673236 598952 673242 599004
rect 674466 598952 674472 599004
rect 674524 598992 674530 599004
rect 675294 598992 675300 599004
rect 674524 598964 675300 598992
rect 674524 598952 674530 598964
rect 675294 598952 675300 598964
rect 675352 598952 675358 599004
rect 651466 597524 651472 597576
rect 651524 597564 651530 597576
rect 669958 597564 669964 597576
rect 651524 597536 669964 597564
rect 651524 597524 651530 597536
rect 669958 597524 669964 597536
rect 670016 597524 670022 597576
rect 43070 597388 43076 597440
rect 43128 597388 43134 597440
rect 43088 597032 43116 597388
rect 43070 596980 43076 597032
rect 43128 596980 43134 597032
rect 651466 596164 651472 596216
rect 651524 596204 651530 596216
rect 664438 596204 664444 596216
rect 651524 596176 664444 596204
rect 651524 596164 651530 596176
rect 664438 596164 664444 596176
rect 664496 596164 664502 596216
rect 40126 595756 40132 595808
rect 40184 595796 40190 595808
rect 41690 595796 41696 595808
rect 40184 595768 41696 595796
rect 40184 595756 40190 595768
rect 41690 595756 41696 595768
rect 41748 595756 41754 595808
rect 651650 595484 651656 595536
rect 651708 595524 651714 595536
rect 653398 595524 653404 595536
rect 651708 595496 653404 595524
rect 651708 595484 651714 595496
rect 653398 595484 653404 595496
rect 653456 595484 653462 595536
rect 651466 594804 651472 594856
rect 651524 594844 651530 594856
rect 661678 594844 661684 594856
rect 651524 594816 661684 594844
rect 651524 594804 651530 594816
rect 661678 594804 661684 594816
rect 661736 594804 661742 594856
rect 41322 594736 41328 594788
rect 41380 594776 41386 594788
rect 41690 594776 41696 594788
rect 41380 594748 41696 594776
rect 41380 594736 41386 594748
rect 41690 594736 41696 594748
rect 41748 594736 41754 594788
rect 651466 594668 651472 594720
rect 651524 594708 651530 594720
rect 657538 594708 657544 594720
rect 651524 594680 657544 594708
rect 651524 594668 651530 594680
rect 657538 594668 657544 594680
rect 657596 594668 657602 594720
rect 39942 594260 39948 594312
rect 40000 594300 40006 594312
rect 41598 594300 41604 594312
rect 40000 594272 41604 594300
rect 40000 594260 40006 594272
rect 41598 594260 41604 594272
rect 41656 594260 41662 594312
rect 651466 593240 651472 593292
rect 651524 593280 651530 593292
rect 654778 593280 654784 593292
rect 651524 593252 654784 593280
rect 651524 593240 651530 593252
rect 654778 593240 654784 593252
rect 654836 593240 654842 593292
rect 674282 592628 674288 592680
rect 674340 592668 674346 592680
rect 683390 592668 683396 592680
rect 674340 592640 683396 592668
rect 674340 592628 674346 592640
rect 683390 592628 683396 592640
rect 683448 592628 683454 592680
rect 674834 591472 674840 591524
rect 674892 591512 674898 591524
rect 679618 591512 679624 591524
rect 674892 591484 679624 591512
rect 674892 591472 674898 591484
rect 679618 591472 679624 591484
rect 679676 591472 679682 591524
rect 35618 590792 35624 590844
rect 35676 590832 35682 590844
rect 35676 590804 39896 590832
rect 35676 590792 35682 590804
rect 39868 590764 39896 590804
rect 41690 590764 41696 590776
rect 39868 590736 41696 590764
rect 41690 590724 41696 590736
rect 41748 590724 41754 590776
rect 35802 590656 35808 590708
rect 35860 590696 35866 590708
rect 39666 590696 39672 590708
rect 35860 590668 39672 590696
rect 35860 590656 35866 590668
rect 39666 590656 39672 590668
rect 39724 590656 39730 590708
rect 42058 590656 42064 590708
rect 42116 590696 42122 590708
rect 43254 590696 43260 590708
rect 42116 590668 43260 590696
rect 42116 590656 42122 590668
rect 43254 590656 43260 590668
rect 43312 590656 43318 590708
rect 674650 588548 674656 588600
rect 674708 588588 674714 588600
rect 684034 588588 684040 588600
rect 674708 588560 684040 588588
rect 674708 588548 674714 588560
rect 684034 588548 684040 588560
rect 684092 588548 684098 588600
rect 33042 587120 33048 587172
rect 33100 587160 33106 587172
rect 41506 587160 41512 587172
rect 33100 587132 41512 587160
rect 33100 587120 33106 587132
rect 41506 587120 41512 587132
rect 41564 587120 41570 587172
rect 42242 586236 42248 586288
rect 42300 586276 42306 586288
rect 42610 586276 42616 586288
rect 42300 586248 42616 586276
rect 42300 586236 42306 586248
rect 42610 586236 42616 586248
rect 42668 586236 42674 586288
rect 35158 586100 35164 586152
rect 35216 586140 35222 586152
rect 35216 586112 36032 586140
rect 35216 586100 35222 586112
rect 36004 586072 36032 586112
rect 39390 586072 39396 586084
rect 36004 586044 39396 586072
rect 39390 586032 39396 586044
rect 39448 586032 39454 586084
rect 33778 585896 33784 585948
rect 33836 585936 33842 585948
rect 39758 585936 39764 585948
rect 33836 585908 39764 585936
rect 33836 585896 33842 585908
rect 39758 585896 39764 585908
rect 39816 585896 39822 585948
rect 31018 585760 31024 585812
rect 31076 585800 31082 585812
rect 39206 585800 39212 585812
rect 31076 585772 39212 585800
rect 31076 585760 31082 585772
rect 39206 585760 39212 585772
rect 39264 585760 39270 585812
rect 660298 581000 660304 581052
rect 660356 581040 660362 581052
rect 673178 581040 673184 581052
rect 660356 581012 673184 581040
rect 660356 581000 660362 581012
rect 673178 581000 673184 581012
rect 673236 581000 673242 581052
rect 668578 580252 668584 580304
rect 668636 580292 668642 580304
rect 673178 580292 673184 580304
rect 668636 580264 673184 580292
rect 668636 580252 668642 580264
rect 673178 580252 673184 580264
rect 673236 580252 673242 580304
rect 670234 579980 670240 580032
rect 670292 580020 670298 580032
rect 673178 580020 673184 580032
rect 670292 579992 673184 580020
rect 670292 579980 670298 579992
rect 673178 579980 673184 579992
rect 673236 579980 673242 580032
rect 674374 579708 674380 579760
rect 674432 579748 674438 579760
rect 676214 579748 676220 579760
rect 674432 579720 676220 579748
rect 674432 579708 674438 579720
rect 676214 579708 676220 579720
rect 676272 579708 676278 579760
rect 658918 579640 658924 579692
rect 658976 579680 658982 579692
rect 673178 579680 673184 579692
rect 658976 579652 673184 579680
rect 658976 579640 658982 579652
rect 673178 579640 673184 579652
rect 673236 579640 673242 579692
rect 42242 578960 42248 579012
rect 42300 579000 42306 579012
rect 43254 579000 43260 579012
rect 42300 578972 43260 579000
rect 42300 578960 42306 578972
rect 43254 578960 43260 578972
rect 43312 578960 43318 579012
rect 669406 578892 669412 578944
rect 669464 578932 669470 578944
rect 673178 578932 673184 578944
rect 669464 578904 673184 578932
rect 669464 578892 669470 578904
rect 673178 578892 673184 578904
rect 673236 578892 673242 578944
rect 674466 578416 674472 578468
rect 674524 578456 674530 578468
rect 676214 578456 676220 578468
rect 674524 578428 676220 578456
rect 674524 578416 674530 578428
rect 676214 578416 676220 578428
rect 676272 578416 676278 578468
rect 670786 578212 670792 578264
rect 670844 578252 670850 578264
rect 673178 578252 673184 578264
rect 670844 578224 673184 578252
rect 670844 578212 670850 578224
rect 673178 578212 673184 578224
rect 673236 578212 673242 578264
rect 670234 577600 670240 577652
rect 670292 577640 670298 577652
rect 673178 577640 673184 577652
rect 670292 577612 673184 577640
rect 670292 577600 670298 577612
rect 673178 577600 673184 577612
rect 673236 577600 673242 577652
rect 674374 577532 674380 577584
rect 674432 577572 674438 577584
rect 676214 577572 676220 577584
rect 674432 577544 676220 577572
rect 674432 577532 674438 577544
rect 676214 577532 676220 577544
rect 676272 577532 676278 577584
rect 670418 577396 670424 577448
rect 670476 577436 670482 577448
rect 673178 577436 673184 577448
rect 670476 577408 673184 577436
rect 670476 577396 670482 577408
rect 673178 577396 673184 577408
rect 673236 577396 673242 577448
rect 671430 577124 671436 577176
rect 671488 577164 671494 577176
rect 673178 577164 673184 577176
rect 671488 577136 673184 577164
rect 671488 577124 671494 577136
rect 673178 577124 673184 577136
rect 673236 577124 673242 577176
rect 669406 576852 669412 576904
rect 669464 576892 669470 576904
rect 673178 576892 673184 576904
rect 669464 576864 673184 576892
rect 669464 576852 669470 576864
rect 673178 576852 673184 576864
rect 673236 576852 673242 576904
rect 45094 575424 45100 575476
rect 45152 575464 45158 575476
rect 62114 575464 62120 575476
rect 45152 575436 62120 575464
rect 45152 575424 45158 575436
rect 62114 575424 62120 575436
rect 62172 575424 62178 575476
rect 671614 574540 671620 574592
rect 671672 574580 671678 574592
rect 673914 574580 673920 574592
rect 671672 574552 673920 574580
rect 671672 574540 671678 574552
rect 673914 574540 673920 574552
rect 673972 574540 673978 574592
rect 671982 574268 671988 574320
rect 672040 574308 672046 574320
rect 673914 574308 673920 574320
rect 672040 574280 673920 574308
rect 672040 574268 672046 574280
rect 673914 574268 673920 574280
rect 673972 574268 673978 574320
rect 667474 574064 667480 574116
rect 667532 574104 667538 574116
rect 667532 574076 673960 574104
rect 667532 574064 667538 574076
rect 46934 573996 46940 574048
rect 46992 574036 46998 574048
rect 62114 574036 62120 574048
rect 46992 574008 62120 574036
rect 46992 573996 46998 574008
rect 62114 573996 62120 574008
rect 62172 573996 62178 574048
rect 673932 573912 673960 574076
rect 674374 574064 674380 574116
rect 674432 574104 674438 574116
rect 676214 574104 676220 574116
rect 674432 574076 676220 574104
rect 674432 574064 674438 574076
rect 676214 574064 676220 574076
rect 676272 574064 676278 574116
rect 673914 573860 673920 573912
rect 673972 573860 673978 573912
rect 671798 571548 671804 571600
rect 671856 571588 671862 571600
rect 673914 571588 673920 571600
rect 671856 571560 673920 571588
rect 671856 571548 671862 571560
rect 673914 571548 673920 571560
rect 673972 571548 673978 571600
rect 674558 571548 674564 571600
rect 674616 571588 674622 571600
rect 676030 571588 676036 571600
rect 674616 571560 676036 571588
rect 674616 571548 674622 571560
rect 676030 571548 676036 571560
rect 676088 571548 676094 571600
rect 674374 571412 674380 571464
rect 674432 571452 674438 571464
rect 676214 571452 676220 571464
rect 674432 571424 676220 571452
rect 674432 571412 674438 571424
rect 676214 571412 676220 571424
rect 676272 571412 676278 571464
rect 669590 571344 669596 571396
rect 669648 571384 669654 571396
rect 673914 571384 673920 571396
rect 669648 571356 673920 571384
rect 669648 571344 669654 571356
rect 673914 571344 673920 571356
rect 673972 571344 673978 571396
rect 671338 571072 671344 571124
rect 671396 571112 671402 571124
rect 673914 571112 673920 571124
rect 671396 571084 673920 571112
rect 671396 571072 671402 571084
rect 673914 571072 673920 571084
rect 673972 571072 673978 571124
rect 42058 570936 42064 570988
rect 42116 570976 42122 570988
rect 42610 570976 42616 570988
rect 42116 570948 42616 570976
rect 42116 570936 42122 570948
rect 42610 570936 42616 570948
rect 42668 570936 42674 570988
rect 674834 570460 674840 570512
rect 674892 570500 674898 570512
rect 675478 570500 675484 570512
rect 674892 570472 675484 570500
rect 674892 570460 674898 570472
rect 675478 570460 675484 570472
rect 675536 570500 675542 570512
rect 683114 570500 683120 570512
rect 675536 570472 683120 570500
rect 675536 570460 675542 570472
rect 683114 570460 683120 570472
rect 683172 570460 683178 570512
rect 671982 569916 671988 569968
rect 672040 569956 672046 569968
rect 673914 569956 673920 569968
rect 672040 569928 673920 569956
rect 672040 569916 672046 569928
rect 673914 569916 673920 569928
rect 673972 569916 673978 569968
rect 669774 568556 669780 568608
rect 669832 568596 669838 568608
rect 673914 568596 673920 568608
rect 669832 568568 673920 568596
rect 669832 568556 669838 568568
rect 673914 568556 673920 568568
rect 673972 568556 673978 568608
rect 653398 565836 653404 565888
rect 653456 565876 653462 565888
rect 673914 565876 673920 565888
rect 653456 565848 673920 565876
rect 653456 565836 653462 565848
rect 673914 565836 673920 565848
rect 673972 565836 673978 565888
rect 665082 564408 665088 564460
rect 665140 564448 665146 564460
rect 673914 564448 673920 564460
rect 665140 564420 673920 564448
rect 665140 564408 665146 564420
rect 673914 564408 673920 564420
rect 673972 564408 673978 564460
rect 657814 554752 657820 554804
rect 657872 554792 657878 554804
rect 672718 554792 672724 554804
rect 657872 554764 672724 554792
rect 657872 554752 657878 554764
rect 672718 554752 672724 554764
rect 672776 554752 672782 554804
rect 674650 553460 674656 553512
rect 674708 553500 674714 553512
rect 675294 553500 675300 553512
rect 674708 553472 675300 553500
rect 674708 553460 674714 553472
rect 675294 553460 675300 553472
rect 675352 553460 675358 553512
rect 655146 553392 655152 553444
rect 655204 553432 655210 553444
rect 669590 553432 669596 553444
rect 655204 553404 669596 553432
rect 655204 553392 655210 553404
rect 669590 553392 669596 553404
rect 669648 553392 669654 553444
rect 674926 553024 674932 553036
rect 674806 552996 674932 553024
rect 674466 552916 674472 552968
rect 674524 552956 674530 552968
rect 674806 552956 674834 552996
rect 674926 552984 674932 552996
rect 674984 552984 674990 553036
rect 674524 552928 674834 552956
rect 674524 552916 674530 552928
rect 651466 552644 651472 552696
rect 651524 552684 651530 552696
rect 665818 552684 665824 552696
rect 651524 552656 665824 552684
rect 651524 552644 651530 552656
rect 665818 552644 665824 552656
rect 665876 552644 665882 552696
rect 41322 552032 41328 552084
rect 41380 552072 41386 552084
rect 41690 552072 41696 552084
rect 41380 552044 41696 552072
rect 41380 552032 41386 552044
rect 41690 552032 41696 552044
rect 41748 552032 41754 552084
rect 674466 552032 674472 552084
rect 674524 552072 674530 552084
rect 675110 552072 675116 552084
rect 674524 552044 675116 552072
rect 674524 552032 674530 552044
rect 675110 552032 675116 552044
rect 675168 552032 675174 552084
rect 651466 550604 651472 550656
rect 651524 550644 651530 550656
rect 660298 550644 660304 550656
rect 651524 550616 660304 550644
rect 651524 550604 651530 550616
rect 660298 550604 660304 550616
rect 660356 550604 660362 550656
rect 40954 550400 40960 550452
rect 41012 550440 41018 550452
rect 41690 550440 41696 550452
rect 41012 550412 41696 550440
rect 41012 550400 41018 550412
rect 41690 550400 41696 550412
rect 41748 550400 41754 550452
rect 651374 550332 651380 550384
rect 651432 550372 651438 550384
rect 653398 550372 653404 550384
rect 651432 550344 653404 550372
rect 651432 550332 651438 550344
rect 653398 550332 653404 550344
rect 653456 550332 653462 550384
rect 651650 549856 651656 549908
rect 651708 549896 651714 549908
rect 663058 549896 663064 549908
rect 651708 549868 663064 549896
rect 651708 549856 651714 549868
rect 663058 549856 663064 549868
rect 663116 549856 663122 549908
rect 651466 549176 651472 549228
rect 651524 549216 651530 549228
rect 657814 549216 657820 549228
rect 651524 549188 657820 549216
rect 651524 549176 651530 549188
rect 657814 549176 657820 549188
rect 657872 549176 657878 549228
rect 674926 548836 674932 548888
rect 674984 548876 674990 548888
rect 675294 548876 675300 548888
rect 674984 548848 675300 548876
rect 674984 548836 674990 548848
rect 675294 548836 675300 548848
rect 675352 548836 675358 548888
rect 651466 548768 651472 548820
rect 651524 548808 651530 548820
rect 655146 548808 655152 548820
rect 651524 548780 655152 548808
rect 651524 548768 651530 548780
rect 655146 548768 655152 548780
rect 655204 548768 655210 548820
rect 41322 547884 41328 547936
rect 41380 547924 41386 547936
rect 41690 547924 41696 547936
rect 41380 547896 41696 547924
rect 41380 547884 41386 547896
rect 41690 547884 41696 547896
rect 41748 547884 41754 547936
rect 674282 547340 674288 547392
rect 674340 547380 674346 547392
rect 683206 547380 683212 547392
rect 674340 547352 683212 547380
rect 674340 547340 674346 547352
rect 683206 547340 683212 547352
rect 683264 547340 683270 547392
rect 29638 547136 29644 547188
rect 29696 547176 29702 547188
rect 41690 547176 41696 547188
rect 29696 547148 41696 547176
rect 29696 547136 29702 547148
rect 41690 547136 41696 547148
rect 41748 547136 41754 547188
rect 675570 547136 675576 547188
rect 675628 547176 675634 547188
rect 683390 547176 683396 547188
rect 675628 547148 683396 547176
rect 675628 547136 675634 547148
rect 683390 547136 683396 547148
rect 683448 547136 683454 547188
rect 675202 546592 675208 546644
rect 675260 546632 675266 546644
rect 675570 546632 675576 546644
rect 675260 546604 675576 546632
rect 675260 546592 675266 546604
rect 675570 546592 675576 546604
rect 675628 546592 675634 546644
rect 675386 546456 675392 546508
rect 675444 546496 675450 546508
rect 680998 546496 681004 546508
rect 675444 546468 681004 546496
rect 675444 546456 675450 546468
rect 680998 546456 681004 546468
rect 681056 546456 681062 546508
rect 675110 540948 675116 541000
rect 675168 540988 675174 541000
rect 675570 540988 675576 541000
rect 675168 540960 675576 540988
rect 675168 540948 675174 540960
rect 675570 540948 675576 540960
rect 675628 540948 675634 541000
rect 673546 536120 673552 536172
rect 673604 536160 673610 536172
rect 673914 536160 673920 536172
rect 673604 536132 673920 536160
rect 673604 536120 673610 536132
rect 673914 536120 673920 536132
rect 673972 536120 673978 536172
rect 669958 535916 669964 535968
rect 670016 535956 670022 535968
rect 674006 535956 674012 535968
rect 670016 535928 674012 535956
rect 670016 535916 670022 535928
rect 674006 535916 674012 535928
rect 674064 535916 674070 535968
rect 674282 535848 674288 535900
rect 674340 535888 674346 535900
rect 676030 535888 676036 535900
rect 674340 535860 676036 535888
rect 674340 535848 674346 535860
rect 676030 535848 676036 535860
rect 676088 535848 676094 535900
rect 674282 535644 674288 535696
rect 674340 535684 674346 535696
rect 676214 535684 676220 535696
rect 674340 535656 676220 535684
rect 674340 535644 674346 535656
rect 676214 535644 676220 535656
rect 676272 535644 676278 535696
rect 664438 535440 664444 535492
rect 664496 535480 664502 535492
rect 674006 535480 674012 535492
rect 664496 535452 674012 535480
rect 664496 535440 664502 535452
rect 674006 535440 674012 535452
rect 674064 535440 674070 535492
rect 670970 534964 670976 535016
rect 671028 535004 671034 535016
rect 674006 535004 674012 535016
rect 671028 534976 674012 535004
rect 671028 534964 671034 534976
rect 674006 534964 674012 534976
rect 674064 534964 674070 535016
rect 674282 534896 674288 534948
rect 674340 534936 674346 534948
rect 676030 534936 676036 534948
rect 674340 534908 676036 534936
rect 674340 534896 674346 534908
rect 676030 534896 676036 534908
rect 676088 534896 676094 534948
rect 670786 534692 670792 534744
rect 670844 534732 670850 534744
rect 674006 534732 674012 534744
rect 670844 534704 674012 534732
rect 670844 534692 670850 534704
rect 674006 534692 674012 534704
rect 674064 534692 674070 534744
rect 674282 534624 674288 534676
rect 674340 534664 674346 534676
rect 676490 534664 676496 534676
rect 674340 534636 676496 534664
rect 674340 534624 674346 534636
rect 676490 534624 676496 534636
rect 676548 534624 676554 534676
rect 674282 534488 674288 534540
rect 674340 534528 674346 534540
rect 676214 534528 676220 534540
rect 674340 534500 676220 534528
rect 674340 534488 674346 534500
rect 676214 534488 676220 534500
rect 676272 534488 676278 534540
rect 661678 534080 661684 534132
rect 661736 534120 661742 534132
rect 674006 534120 674012 534132
rect 661736 534092 674012 534120
rect 661736 534080 661742 534092
rect 674006 534080 674012 534092
rect 674064 534080 674070 534132
rect 675478 533332 675484 533384
rect 675536 533372 675542 533384
rect 683574 533372 683580 533384
rect 675536 533344 683580 533372
rect 675536 533332 675542 533344
rect 683574 533332 683580 533344
rect 683632 533332 683638 533384
rect 670234 533264 670240 533316
rect 670292 533304 670298 533316
rect 674006 533304 674012 533316
rect 670292 533276 674012 533304
rect 670292 533264 670298 533276
rect 674006 533264 674012 533276
rect 674064 533264 674070 533316
rect 674282 533196 674288 533248
rect 674340 533236 674346 533248
rect 676030 533236 676036 533248
rect 674340 533208 676036 533236
rect 674340 533196 674346 533208
rect 676030 533196 676036 533208
rect 676088 533196 676094 533248
rect 674282 532788 674288 532840
rect 674340 532828 674346 532840
rect 676030 532828 676036 532840
rect 674340 532800 676036 532828
rect 674340 532788 674346 532800
rect 676030 532788 676036 532800
rect 676088 532788 676094 532840
rect 670786 532720 670792 532772
rect 670844 532760 670850 532772
rect 674006 532760 674012 532772
rect 670844 532732 674012 532760
rect 670844 532720 670850 532732
rect 674006 532720 674012 532732
rect 674064 532720 674070 532772
rect 669406 532516 669412 532568
rect 669464 532556 669470 532568
rect 674006 532556 674012 532568
rect 669464 532528 674012 532556
rect 669464 532516 669470 532528
rect 674006 532516 674012 532528
rect 674064 532516 674070 532568
rect 674282 532448 674288 532500
rect 674340 532488 674346 532500
rect 676030 532488 676036 532500
rect 674340 532460 676036 532488
rect 674340 532448 674346 532460
rect 676030 532448 676036 532460
rect 676088 532448 676094 532500
rect 44818 531972 44824 532024
rect 44876 532012 44882 532024
rect 62114 532012 62120 532024
rect 44876 531984 62120 532012
rect 44876 531972 44882 531984
rect 62114 531972 62120 531984
rect 62172 531972 62178 532024
rect 671614 531972 671620 532024
rect 671672 532012 671678 532024
rect 674006 532012 674012 532024
rect 671672 531984 674012 532012
rect 671672 531972 671678 531984
rect 674006 531972 674012 531984
rect 674064 531972 674070 532024
rect 674282 531972 674288 532024
rect 674340 532012 674346 532024
rect 676030 532012 676036 532024
rect 674340 531984 676036 532012
rect 674340 531972 674346 531984
rect 676030 531972 676036 531984
rect 676088 531972 676094 532024
rect 667658 531836 667664 531888
rect 667716 531876 667722 531888
rect 674006 531876 674012 531888
rect 667716 531848 674012 531876
rect 667716 531836 667722 531848
rect 674006 531836 674012 531848
rect 674064 531836 674070 531888
rect 674282 531768 674288 531820
rect 674340 531808 674346 531820
rect 676214 531808 676220 531820
rect 674340 531780 676220 531808
rect 674340 531768 674346 531780
rect 676214 531768 676220 531780
rect 676272 531768 676278 531820
rect 51718 531224 51724 531276
rect 51776 531264 51782 531276
rect 62298 531264 62304 531276
rect 51776 531236 62304 531264
rect 51776 531224 51782 531236
rect 62298 531224 62304 531236
rect 62356 531224 62362 531276
rect 42702 530924 42708 530936
rect 42168 530896 42708 530924
rect 42168 530732 42196 530896
rect 42702 530884 42708 530896
rect 42760 530884 42766 530936
rect 672166 530884 672172 530936
rect 672224 530924 672230 530936
rect 674006 530924 674012 530936
rect 672224 530896 674012 530924
rect 672224 530884 672230 530896
rect 674006 530884 674012 530896
rect 674064 530884 674070 530936
rect 674282 530816 674288 530868
rect 674340 530856 674346 530868
rect 676030 530856 676036 530868
rect 674340 530828 676036 530856
rect 674340 530816 674346 530828
rect 676030 530816 676036 530828
rect 676088 530816 676094 530868
rect 42150 530680 42156 530732
rect 42208 530680 42214 530732
rect 42242 530272 42248 530324
rect 42300 530312 42306 530324
rect 42886 530312 42892 530324
rect 42300 530284 42892 530312
rect 42300 530272 42306 530284
rect 42886 530272 42892 530284
rect 42944 530272 42950 530324
rect 667290 529932 667296 529984
rect 667348 529972 667354 529984
rect 674006 529972 674012 529984
rect 667348 529944 674012 529972
rect 667348 529932 667354 529944
rect 674006 529932 674012 529944
rect 674064 529932 674070 529984
rect 674282 529932 674288 529984
rect 674340 529972 674346 529984
rect 676030 529972 676036 529984
rect 674340 529944 676036 529972
rect 674340 529932 674346 529944
rect 676030 529932 676036 529944
rect 676088 529932 676094 529984
rect 671154 529388 671160 529440
rect 671212 529428 671218 529440
rect 674006 529428 674012 529440
rect 671212 529400 674012 529428
rect 671212 529388 671218 529400
rect 674006 529388 674012 529400
rect 674064 529388 674070 529440
rect 674282 529320 674288 529372
rect 674340 529360 674346 529372
rect 676030 529360 676036 529372
rect 674340 529332 676036 529360
rect 674340 529320 674346 529332
rect 676030 529320 676036 529332
rect 676088 529320 676094 529372
rect 674282 529184 674288 529236
rect 674340 529224 674346 529236
rect 676214 529224 676220 529236
rect 674340 529196 676220 529224
rect 674340 529184 674346 529196
rect 676214 529184 676220 529196
rect 676272 529184 676278 529236
rect 668394 529116 668400 529168
rect 668452 529156 668458 529168
rect 674006 529156 674012 529168
rect 668452 529128 674012 529156
rect 668452 529116 668458 529128
rect 674006 529116 674012 529128
rect 674064 529116 674070 529168
rect 672350 528844 672356 528896
rect 672408 528884 672414 528896
rect 674006 528884 674012 528896
rect 672408 528856 674012 528884
rect 672408 528844 672414 528856
rect 674006 528844 674012 528856
rect 674064 528844 674070 528896
rect 674282 528776 674288 528828
rect 674340 528816 674346 528828
rect 676030 528816 676036 528828
rect 674340 528788 676036 528816
rect 674340 528776 674346 528788
rect 676030 528776 676036 528788
rect 676088 528776 676094 528828
rect 45186 528572 45192 528624
rect 45244 528612 45250 528624
rect 62114 528612 62120 528624
rect 45244 528584 62120 528612
rect 45244 528572 45250 528584
rect 62114 528572 62120 528584
rect 62172 528572 62178 528624
rect 672534 528028 672540 528080
rect 672592 528068 672598 528080
rect 674006 528068 674012 528080
rect 672592 528040 674012 528068
rect 672592 528028 672598 528040
rect 674006 528028 674012 528040
rect 674064 528028 674070 528080
rect 674282 527960 674288 528012
rect 674340 528000 674346 528012
rect 676030 528000 676036 528012
rect 674340 527972 676036 528000
rect 674340 527960 674346 527972
rect 676030 527960 676036 527972
rect 676088 527960 676094 528012
rect 47578 527076 47584 527128
rect 47636 527116 47642 527128
rect 62114 527116 62120 527128
rect 47636 527088 62120 527116
rect 47636 527076 47642 527088
rect 62114 527076 62120 527088
rect 62172 527076 62178 527128
rect 42058 527008 42064 527060
rect 42116 527048 42122 527060
rect 42702 527048 42708 527060
rect 42116 527020 42708 527048
rect 42116 527008 42122 527020
rect 42702 527008 42708 527020
rect 42760 527008 42766 527060
rect 669038 524560 669044 524612
rect 669096 524600 669102 524612
rect 674006 524600 674012 524612
rect 669096 524572 674012 524600
rect 669096 524560 669102 524572
rect 674006 524560 674012 524572
rect 674064 524560 674070 524612
rect 674282 524560 674288 524612
rect 674340 524600 674346 524612
rect 683114 524600 683120 524612
rect 674340 524572 683120 524600
rect 674340 524560 674346 524572
rect 683114 524560 683120 524572
rect 683172 524560 683178 524612
rect 668578 524424 668584 524476
rect 668636 524464 668642 524476
rect 669038 524464 669044 524476
rect 668636 524436 669044 524464
rect 668636 524424 668642 524436
rect 669038 524424 669044 524436
rect 669096 524424 669102 524476
rect 675478 520208 675484 520260
rect 675536 520248 675542 520260
rect 680354 520248 680360 520260
rect 675536 520220 680360 520248
rect 675536 520208 675542 520220
rect 680354 520208 680360 520220
rect 680412 520208 680418 520260
rect 675662 518780 675668 518832
rect 675720 518820 675726 518832
rect 677870 518820 677876 518832
rect 675720 518792 677876 518820
rect 675720 518780 675726 518792
rect 677870 518780 677876 518792
rect 677928 518780 677934 518832
rect 658458 518168 658464 518220
rect 658516 518208 658522 518220
rect 668578 518208 668584 518220
rect 658516 518180 668584 518208
rect 658516 518168 658522 518180
rect 668578 518168 668584 518180
rect 668636 518168 668642 518220
rect 650638 509872 650644 509924
rect 650696 509912 650702 509924
rect 658458 509912 658464 509924
rect 650696 509884 658464 509912
rect 650696 509872 650702 509884
rect 658458 509872 658464 509884
rect 658516 509872 658522 509924
rect 675110 503616 675116 503668
rect 675168 503656 675174 503668
rect 679618 503656 679624 503668
rect 675168 503628 679624 503656
rect 675168 503616 675174 503628
rect 679618 503616 679624 503628
rect 679676 503616 679682 503668
rect 675294 503480 675300 503532
rect 675352 503520 675358 503532
rect 680998 503520 681004 503532
rect 675352 503492 681004 503520
rect 675352 503480 675358 503492
rect 680998 503480 681004 503492
rect 681056 503480 681062 503532
rect 674834 500896 674840 500948
rect 674892 500936 674898 500948
rect 681182 500936 681188 500948
rect 674892 500908 681188 500936
rect 674892 500896 674898 500908
rect 681182 500896 681188 500908
rect 681240 500896 681246 500948
rect 674282 491648 674288 491700
rect 674340 491688 674346 491700
rect 676030 491688 676036 491700
rect 674340 491660 676036 491688
rect 674340 491648 674346 491660
rect 676030 491648 676036 491660
rect 676088 491648 676094 491700
rect 665818 491580 665824 491632
rect 665876 491620 665882 491632
rect 674006 491620 674012 491632
rect 665876 491592 674012 491620
rect 665876 491580 665882 491592
rect 674006 491580 674012 491592
rect 674064 491580 674070 491632
rect 663058 491444 663064 491496
rect 663116 491484 663122 491496
rect 673822 491484 673828 491496
rect 663116 491456 673828 491484
rect 663116 491444 663122 491456
rect 673822 491444 673828 491456
rect 673880 491444 673886 491496
rect 660298 491308 660304 491360
rect 660356 491348 660362 491360
rect 674006 491348 674012 491360
rect 660356 491320 674012 491348
rect 660356 491308 660362 491320
rect 674006 491308 674012 491320
rect 674064 491308 674070 491360
rect 670970 490900 670976 490952
rect 671028 490940 671034 490952
rect 674006 490940 674012 490952
rect 671028 490912 674012 490940
rect 671028 490900 671034 490912
rect 674006 490900 674012 490912
rect 674064 490900 674070 490952
rect 672534 490696 672540 490748
rect 672592 490736 672598 490748
rect 672902 490736 672908 490748
rect 672592 490708 672908 490736
rect 672592 490696 672598 490708
rect 672902 490696 672908 490708
rect 672960 490696 672966 490748
rect 672442 489608 672448 489660
rect 672500 489648 672506 489660
rect 674006 489648 674012 489660
rect 672500 489620 674012 489648
rect 672500 489608 672506 489620
rect 674006 489608 674012 489620
rect 674064 489608 674070 489660
rect 670786 489268 670792 489320
rect 670844 489308 670850 489320
rect 674006 489308 674012 489320
rect 670844 489280 674012 489308
rect 670844 489268 670850 489280
rect 674006 489268 674012 489280
rect 674064 489268 674070 489320
rect 671614 488452 671620 488504
rect 671672 488492 671678 488504
rect 674006 488492 674012 488504
rect 671672 488464 674012 488492
rect 671672 488452 671678 488464
rect 674006 488452 674012 488464
rect 674064 488452 674070 488504
rect 672626 486004 672632 486056
rect 672684 486044 672690 486056
rect 674006 486044 674012 486056
rect 672684 486016 674012 486044
rect 672684 486004 672690 486016
rect 674006 486004 674012 486016
rect 674064 486004 674070 486056
rect 674282 485868 674288 485920
rect 674340 485908 674346 485920
rect 676030 485908 676036 485920
rect 674340 485880 676036 485908
rect 674340 485868 674346 485880
rect 676030 485868 676036 485880
rect 676088 485868 676094 485920
rect 665082 485800 665088 485852
rect 665140 485840 665146 485852
rect 674006 485840 674012 485852
rect 665140 485812 674012 485840
rect 665140 485800 665146 485812
rect 674006 485800 674012 485812
rect 674064 485800 674070 485852
rect 674282 485120 674288 485172
rect 674340 485160 674346 485172
rect 676030 485160 676036 485172
rect 674340 485132 676036 485160
rect 674340 485120 674346 485132
rect 676030 485120 676036 485132
rect 676088 485120 676094 485172
rect 668762 484372 668768 484424
rect 668820 484412 668826 484424
rect 674006 484412 674012 484424
rect 668820 484384 674012 484412
rect 668820 484372 668826 484384
rect 674006 484372 674012 484384
rect 674064 484372 674070 484424
rect 674466 483964 674472 484016
rect 674524 484004 674530 484016
rect 676030 484004 676036 484016
rect 674524 483976 676036 484004
rect 674524 483964 674530 483976
rect 676030 483964 676036 483976
rect 676088 483964 676094 484016
rect 671798 483148 671804 483200
rect 671856 483188 671862 483200
rect 674006 483188 674012 483200
rect 671856 483160 674012 483188
rect 671856 483148 671862 483160
rect 674006 483148 674012 483160
rect 674064 483148 674070 483200
rect 676214 482944 676220 482996
rect 676272 482984 676278 482996
rect 677410 482984 677416 482996
rect 676272 482956 677416 482984
rect 676272 482944 676278 482956
rect 677410 482944 677416 482956
rect 677468 482944 677474 482996
rect 674650 482332 674656 482384
rect 674708 482372 674714 482384
rect 676030 482372 676036 482384
rect 674708 482344 676036 482372
rect 674708 482332 674714 482344
rect 676030 482332 676036 482344
rect 676088 482332 676094 482384
rect 665174 480360 665180 480412
rect 665232 480400 665238 480412
rect 670418 480400 670424 480412
rect 665232 480372 670424 480400
rect 665232 480360 665238 480372
rect 670418 480360 670424 480372
rect 670476 480400 670482 480412
rect 674006 480400 674012 480412
rect 670476 480372 674012 480400
rect 670476 480360 670482 480372
rect 674006 480360 674012 480372
rect 674064 480360 674070 480412
rect 674282 480360 674288 480412
rect 674340 480400 674346 480412
rect 683114 480400 683120 480412
rect 674340 480372 683120 480400
rect 674340 480360 674346 480372
rect 683114 480360 683120 480372
rect 683172 480360 683178 480412
rect 659654 476144 659660 476196
rect 659712 476184 659718 476196
rect 665174 476184 665180 476196
rect 659712 476156 665180 476184
rect 659712 476144 659718 476156
rect 665174 476144 665180 476156
rect 665232 476144 665238 476196
rect 676030 475124 676036 475176
rect 676088 475164 676094 475176
rect 680354 475164 680360 475176
rect 676088 475136 680360 475164
rect 676088 475124 676094 475136
rect 680354 475124 680360 475136
rect 680412 475124 680418 475176
rect 656158 473424 656164 473476
rect 656216 473464 656222 473476
rect 659654 473464 659660 473476
rect 656216 473436 659660 473464
rect 656216 473424 656222 473436
rect 659654 473424 659660 473436
rect 659712 473424 659718 473476
rect 650822 470568 650828 470620
rect 650880 470608 650886 470620
rect 656158 470608 656164 470620
rect 650880 470580 656164 470608
rect 650880 470568 650886 470580
rect 656158 470568 656164 470580
rect 656216 470568 656222 470620
rect 667014 456560 667020 456612
rect 667072 456600 667078 456612
rect 667072 456572 673988 456600
rect 667072 456560 667078 456572
rect 673960 456246 673988 456572
rect 667842 455948 667848 456000
rect 667900 455988 667906 456000
rect 667900 455960 673854 455988
rect 667900 455948 667906 455960
rect 673362 455812 673368 455864
rect 673420 455852 673426 455864
rect 673420 455824 673762 455852
rect 673420 455812 673426 455824
rect 669222 455608 669228 455660
rect 669280 455648 669286 455660
rect 669280 455620 673624 455648
rect 669280 455608 669286 455620
rect 673270 455336 673276 455388
rect 673328 455336 673334 455388
rect 673288 455022 673316 455336
rect 673388 455252 673440 455258
rect 673388 455194 673440 455200
rect 673506 455252 673558 455258
rect 673506 455194 673558 455200
rect 674282 454860 674288 454912
rect 674340 454900 674346 454912
rect 675846 454900 675852 454912
rect 674340 454872 675852 454900
rect 674340 454860 674346 454872
rect 675846 454860 675852 454872
rect 675904 454860 675910 454912
rect 672074 454792 672080 454844
rect 672132 454832 672138 454844
rect 672132 454804 673190 454832
rect 672132 454792 672138 454804
rect 673046 454640 673098 454646
rect 674282 454588 674288 454640
rect 674340 454628 674346 454640
rect 675478 454628 675484 454640
rect 674340 454600 675484 454628
rect 674340 454588 674346 454600
rect 675478 454588 675484 454600
rect 675536 454588 675542 454640
rect 673046 454582 673098 454588
rect 672810 454452 672816 454504
rect 672868 454452 672874 454504
rect 672828 454206 672856 454452
rect 672954 454368 673006 454374
rect 674282 454316 674288 454368
rect 674340 454356 674346 454368
rect 675662 454356 675668 454368
rect 674340 454328 675668 454356
rect 674340 454316 674346 454328
rect 675662 454316 675668 454328
rect 675720 454316 675726 454368
rect 672954 454310 673006 454316
rect 672258 453908 672264 453960
rect 672316 453948 672322 453960
rect 672316 453920 672750 453948
rect 672316 453908 672322 453920
rect 674282 453908 674288 453960
rect 674340 453948 674346 453960
rect 676030 453948 676036 453960
rect 674340 453920 676036 453948
rect 674340 453908 674346 453920
rect 676030 453908 676036 453920
rect 676088 453908 676094 453960
rect 35802 429156 35808 429208
rect 35860 429196 35866 429208
rect 41690 429196 41696 429208
rect 35860 429168 41696 429196
rect 35860 429156 35866 429168
rect 41690 429156 41696 429168
rect 41748 429156 41754 429208
rect 35802 427932 35808 427984
rect 35860 427972 35866 427984
rect 41690 427972 41696 427984
rect 35860 427944 41696 427972
rect 35860 427932 35866 427944
rect 41690 427932 41696 427944
rect 41748 427932 41754 427984
rect 40954 424328 40960 424380
rect 41012 424368 41018 424380
rect 41690 424368 41696 424380
rect 41012 424340 41696 424368
rect 41012 424328 41018 424340
rect 41690 424328 41696 424340
rect 41748 424328 41754 424380
rect 41138 422356 41144 422408
rect 41196 422396 41202 422408
rect 41598 422396 41604 422408
rect 41196 422368 41604 422396
rect 41196 422356 41202 422368
rect 41598 422356 41604 422368
rect 41656 422356 41662 422408
rect 32030 417392 32036 417444
rect 32088 417432 32094 417444
rect 41690 417432 41696 417444
rect 32088 417404 41696 417432
rect 32088 417392 32094 417404
rect 41690 417392 41696 417404
rect 41748 417392 41754 417444
rect 42058 417256 42064 417308
rect 42116 417296 42122 417308
rect 42610 417296 42616 417308
rect 42116 417268 42616 417296
rect 42116 417256 42122 417268
rect 42610 417256 42616 417268
rect 42668 417256 42674 417308
rect 34514 416032 34520 416084
rect 34572 416072 34578 416084
rect 41690 416072 41696 416084
rect 34572 416044 41696 416072
rect 34572 416032 34578 416044
rect 41690 416032 41696 416044
rect 41748 416032 41754 416084
rect 42242 409776 42248 409828
rect 42300 409816 42306 409828
rect 43162 409816 43168 409828
rect 42300 409788 43168 409816
rect 42300 409776 42306 409788
rect 43162 409776 43168 409788
rect 43220 409776 43226 409828
rect 42242 406988 42248 407040
rect 42300 407028 42306 407040
rect 42610 407028 42616 407040
rect 42300 407000 42616 407028
rect 42300 406988 42306 407000
rect 42610 406988 42616 407000
rect 42668 406988 42674 407040
rect 44726 404268 44732 404320
rect 44784 404308 44790 404320
rect 62114 404308 62120 404320
rect 44784 404280 62120 404308
rect 44784 404268 44790 404280
rect 62114 404268 62120 404280
rect 62172 404268 62178 404320
rect 674558 403248 674564 403300
rect 674616 403288 674622 403300
rect 676214 403288 676220 403300
rect 674616 403260 676220 403288
rect 674616 403248 674622 403260
rect 676214 403248 676220 403260
rect 676272 403248 676278 403300
rect 51442 402908 51448 402960
rect 51500 402948 51506 402960
rect 62114 402948 62120 402960
rect 51500 402920 62120 402948
rect 51500 402908 51506 402920
rect 62114 402908 62120 402920
rect 62172 402908 62178 402960
rect 42426 402228 42432 402280
rect 42484 402268 42490 402280
rect 42978 402268 42984 402280
rect 42484 402240 42984 402268
rect 42484 402228 42490 402240
rect 42978 402228 42984 402240
rect 43036 402228 43042 402280
rect 45186 400256 45192 400308
rect 45244 400256 45250 400308
rect 45204 400092 45232 400256
rect 51074 400188 51080 400240
rect 51132 400228 51138 400240
rect 62114 400228 62120 400240
rect 51132 400200 62120 400228
rect 51132 400188 51138 400200
rect 62114 400188 62120 400200
rect 62172 400188 62178 400240
rect 62114 400092 62120 400104
rect 45204 400064 62120 400092
rect 62114 400052 62120 400064
rect 62172 400052 62178 400104
rect 46382 399440 46388 399492
rect 46440 399480 46446 399492
rect 56042 399480 56048 399492
rect 46440 399452 56048 399480
rect 46440 399440 46446 399452
rect 56042 399440 56048 399452
rect 56100 399440 56106 399492
rect 674926 398828 674932 398880
rect 674984 398868 674990 398880
rect 676030 398868 676036 398880
rect 674984 398840 676036 398868
rect 674984 398828 674990 398840
rect 676030 398828 676036 398840
rect 676088 398828 676094 398880
rect 47762 398760 47768 398812
rect 47820 398800 47826 398812
rect 62114 398800 62120 398812
rect 47820 398772 62120 398800
rect 47820 398760 47826 398772
rect 62114 398760 62120 398772
rect 62172 398760 62178 398812
rect 674558 396040 674564 396092
rect 674616 396080 674622 396092
rect 676030 396080 676036 396092
rect 674616 396052 676036 396080
rect 674616 396040 674622 396052
rect 676030 396040 676036 396052
rect 676088 396040 676094 396092
rect 675202 395700 675208 395752
rect 675260 395740 675266 395752
rect 676214 395740 676220 395752
rect 675260 395712 676220 395740
rect 675260 395700 675266 395712
rect 676214 395700 676220 395712
rect 676272 395700 676278 395752
rect 674374 394272 674380 394324
rect 674432 394312 674438 394324
rect 676214 394312 676220 394324
rect 674432 394284 676220 394312
rect 674432 394272 674438 394284
rect 676214 394272 676220 394284
rect 676272 394272 676278 394324
rect 679618 386764 679624 386776
rect 675588 386736 679624 386764
rect 41322 386384 41328 386436
rect 41380 386424 41386 386436
rect 41690 386424 41696 386436
rect 41380 386396 41696 386424
rect 41380 386384 41386 386396
rect 41690 386384 41696 386396
rect 41748 386384 41754 386436
rect 675588 386424 675616 386736
rect 679618 386724 679624 386736
rect 679676 386724 679682 386776
rect 675496 386396 675616 386424
rect 675496 386028 675524 386396
rect 675478 385976 675484 386028
rect 675536 385976 675542 386028
rect 674834 384752 674840 384804
rect 674892 384792 674898 384804
rect 675386 384792 675392 384804
rect 674892 384764 675392 384792
rect 674892 384752 674898 384764
rect 675386 384752 675392 384764
rect 675444 384752 675450 384804
rect 41322 382236 41328 382288
rect 41380 382276 41386 382288
rect 41690 382276 41696 382288
rect 41380 382248 41696 382276
rect 41380 382236 41386 382248
rect 41690 382236 41696 382248
rect 41748 382236 41754 382288
rect 674374 382168 674380 382220
rect 674432 382208 674438 382220
rect 675110 382208 675116 382220
rect 674432 382180 675116 382208
rect 674432 382168 674438 382180
rect 675110 382168 675116 382180
rect 675168 382168 675174 382220
rect 41322 379720 41328 379772
rect 41380 379760 41386 379772
rect 41506 379760 41512 379772
rect 41380 379732 41512 379760
rect 41380 379720 41386 379732
rect 41506 379720 41512 379732
rect 41564 379720 41570 379772
rect 40402 379624 40408 379636
rect 36096 379596 40408 379624
rect 35802 379516 35808 379568
rect 35860 379556 35866 379568
rect 35860 379528 36032 379556
rect 35860 379516 35866 379528
rect 36004 379488 36032 379528
rect 36096 379488 36124 379596
rect 40402 379584 40408 379596
rect 40460 379584 40466 379636
rect 36004 379460 36124 379488
rect 35802 378156 35808 378208
rect 35860 378196 35866 378208
rect 41690 378196 41696 378208
rect 35860 378168 41696 378196
rect 35860 378156 35866 378168
rect 41690 378156 41696 378168
rect 41748 378156 41754 378208
rect 674374 378088 674380 378140
rect 674432 378128 674438 378140
rect 675110 378128 675116 378140
rect 674432 378100 675116 378128
rect 674432 378088 674438 378100
rect 675110 378088 675116 378100
rect 675168 378088 675174 378140
rect 651466 373940 651472 373992
rect 651524 373980 651530 373992
rect 657538 373980 657544 373992
rect 651524 373952 657544 373980
rect 651524 373940 651530 373952
rect 657538 373940 657544 373952
rect 657596 373940 657602 373992
rect 33962 373260 33968 373312
rect 34020 373300 34026 373312
rect 41690 373300 41696 373312
rect 34020 373272 41696 373300
rect 34020 373260 34026 373272
rect 41690 373260 41696 373272
rect 41748 373260 41754 373312
rect 674650 372512 674656 372564
rect 674708 372552 674714 372564
rect 675294 372552 675300 372564
rect 674708 372524 675300 372552
rect 674708 372512 674714 372524
rect 675294 372512 675300 372524
rect 675352 372512 675358 372564
rect 39298 372036 39304 372088
rect 39356 372076 39362 372088
rect 41690 372076 41696 372088
rect 39356 372048 41696 372076
rect 39356 372036 39362 372048
rect 41690 372036 41696 372048
rect 41748 372036 41754 372088
rect 42058 371900 42064 371952
rect 42116 371940 42122 371952
rect 42702 371940 42708 371952
rect 42116 371912 42708 371940
rect 42116 371900 42122 371912
rect 42702 371900 42708 371912
rect 42760 371900 42766 371952
rect 651466 370948 651472 371000
rect 651524 370988 651530 371000
rect 654778 370988 654784 371000
rect 651524 370960 654784 370988
rect 651524 370948 651530 370960
rect 654778 370948 654784 370960
rect 654836 370948 654842 371000
rect 42426 366800 42432 366852
rect 42484 366840 42490 366852
rect 43070 366840 43076 366852
rect 42484 366812 43076 366840
rect 42484 366800 42490 366812
rect 43070 366800 43076 366812
rect 43128 366800 43134 366852
rect 42242 365848 42248 365900
rect 42300 365888 42306 365900
rect 42702 365888 42708 365900
rect 42300 365860 42708 365888
rect 42300 365848 42306 365860
rect 42702 365848 42708 365860
rect 42760 365848 42766 365900
rect 655514 364964 655520 365016
rect 655572 365004 655578 365016
rect 668578 365004 668584 365016
rect 655572 364976 668584 365004
rect 655572 364964 655578 364976
rect 668578 364964 668584 364976
rect 668636 364964 668642 365016
rect 42334 362856 42340 362908
rect 42392 362896 42398 362908
rect 42702 362896 42708 362908
rect 42392 362868 42708 362896
rect 42392 362856 42398 362868
rect 42702 362856 42708 362868
rect 42760 362856 42766 362908
rect 651006 361564 651012 361616
rect 651064 361604 651070 361616
rect 655514 361604 655520 361616
rect 651064 361576 655520 361604
rect 651064 361564 651070 361576
rect 655514 361564 655520 361576
rect 655572 361564 655578 361616
rect 44634 361496 44640 361548
rect 44692 361536 44698 361548
rect 62114 361536 62120 361548
rect 44692 361508 62120 361536
rect 44692 361496 44698 361508
rect 62114 361496 62120 361508
rect 62172 361496 62178 361548
rect 51074 360136 51080 360188
rect 51132 360176 51138 360188
rect 62114 360176 62120 360188
rect 51132 360148 62120 360176
rect 51132 360136 51138 360148
rect 62114 360136 62120 360148
rect 62172 360136 62178 360188
rect 44634 357416 44640 357468
rect 44692 357456 44698 357468
rect 62114 357456 62120 357468
rect 44692 357428 62120 357456
rect 44692 357416 44698 357428
rect 62114 357416 62120 357428
rect 62172 357416 62178 357468
rect 42242 355988 42248 356040
rect 42300 356028 42306 356040
rect 42886 356028 42892 356040
rect 42300 356000 42892 356028
rect 42300 355988 42306 356000
rect 42886 355988 42892 356000
rect 42944 355988 42950 356040
rect 47762 355988 47768 356040
rect 47820 356028 47826 356040
rect 62114 356028 62120 356040
rect 47820 356000 62120 356028
rect 47820 355988 47826 356000
rect 62114 355988 62120 356000
rect 62172 355988 62178 356040
rect 45462 354600 45468 354612
rect 44867 354572 45468 354600
rect 44640 354544 44692 354550
rect 44640 354486 44692 354492
rect 44732 354340 44784 354346
rect 44867 354314 44895 354572
rect 45462 354560 45468 354572
rect 45520 354560 45526 354612
rect 44732 354282 44784 354288
rect 45462 354124 45468 354136
rect 44988 354096 45468 354124
rect 45462 354084 45468 354096
rect 45520 354084 45526 354136
rect 45462 353852 45468 353864
rect 45105 353824 45468 353852
rect 45462 353812 45468 353824
rect 45520 353812 45526 353864
rect 45297 353716 45303 353728
rect 45218 353688 45303 353716
rect 45297 353676 45303 353688
rect 45355 353676 45361 353728
rect 47946 353444 47952 353456
rect 45329 353416 47952 353444
rect 47946 353404 47952 353416
rect 48004 353404 48010 353456
rect 45422 353184 45474 353190
rect 45422 353126 45474 353132
rect 35802 344564 35808 344616
rect 35860 344604 35866 344616
rect 40034 344604 40040 344616
rect 35860 344576 40040 344604
rect 35860 344564 35866 344576
rect 40034 344564 40040 344576
rect 40092 344564 40098 344616
rect 35526 343748 35532 343800
rect 35584 343788 35590 343800
rect 40034 343788 40040 343800
rect 35584 343760 40040 343788
rect 35584 343748 35590 343760
rect 40034 343748 40040 343760
rect 40092 343748 40098 343800
rect 35802 342252 35808 342304
rect 35860 342292 35866 342304
rect 40218 342292 40224 342304
rect 35860 342264 40224 342292
rect 35860 342252 35866 342264
rect 40218 342252 40224 342264
rect 40276 342252 40282 342304
rect 33042 341368 33048 341420
rect 33100 341408 33106 341420
rect 40218 341408 40224 341420
rect 33100 341380 40224 341408
rect 33100 341368 33106 341380
rect 40218 341368 40224 341380
rect 40276 341368 40282 341420
rect 45462 341368 45468 341420
rect 45520 341408 45526 341420
rect 62206 341408 62212 341420
rect 45520 341380 62212 341408
rect 45520 341368 45526 341380
rect 62206 341368 62212 341380
rect 62264 341368 62270 341420
rect 35802 341164 35808 341216
rect 35860 341204 35866 341216
rect 40218 341204 40224 341216
rect 35860 341176 40224 341204
rect 35860 341164 35866 341176
rect 40218 341164 40224 341176
rect 40276 341164 40282 341216
rect 35618 341028 35624 341080
rect 35676 341068 35682 341080
rect 40034 341068 40040 341080
rect 35676 341040 40040 341068
rect 35676 341028 35682 341040
rect 40034 341028 40040 341040
rect 40092 341028 40098 341080
rect 35526 339600 35532 339652
rect 35584 339640 35590 339652
rect 36538 339640 36544 339652
rect 35584 339612 36544 339640
rect 35584 339600 35590 339612
rect 36538 339600 36544 339612
rect 36596 339600 36602 339652
rect 35802 339464 35808 339516
rect 35860 339504 35866 339516
rect 38838 339504 38844 339516
rect 35860 339476 38844 339504
rect 35860 339464 35866 339476
rect 38838 339464 38844 339476
rect 38896 339464 38902 339516
rect 35802 335316 35808 335368
rect 35860 335356 35866 335368
rect 40218 335356 40224 335368
rect 35860 335328 40224 335356
rect 35860 335316 35866 335328
rect 40218 335316 40224 335328
rect 40276 335316 40282 335368
rect 35618 334228 35624 334280
rect 35676 334268 35682 334280
rect 39390 334268 39396 334280
rect 35676 334240 39396 334268
rect 35676 334228 35682 334240
rect 39390 334228 39396 334240
rect 39448 334228 39454 334280
rect 35802 333956 35808 334008
rect 35860 333996 35866 334008
rect 41690 333996 41696 334008
rect 35860 333968 41696 333996
rect 35860 333956 35866 333968
rect 41690 333956 41696 333968
rect 41748 333956 41754 334008
rect 42058 333956 42064 334008
rect 42116 333996 42122 334008
rect 42978 333996 42984 334008
rect 42116 333968 42984 333996
rect 42116 333956 42122 333968
rect 42978 333956 42984 333968
rect 43036 333956 43042 334008
rect 674466 333888 674472 333940
rect 674524 333928 674530 333940
rect 675110 333928 675116 333940
rect 674524 333900 675116 333928
rect 674524 333888 674530 333900
rect 675110 333888 675116 333900
rect 675168 333888 675174 333940
rect 651374 328244 651380 328296
rect 651432 328284 651438 328296
rect 654778 328284 654784 328296
rect 651432 328256 654784 328284
rect 651432 328244 651438 328256
rect 654778 328244 654784 328256
rect 654836 328244 654842 328296
rect 651374 325592 651380 325644
rect 651432 325632 651438 325644
rect 653398 325632 653404 325644
rect 651432 325604 653404 325632
rect 651432 325592 651438 325604
rect 653398 325592 653404 325604
rect 653456 325592 653462 325644
rect 42242 322872 42248 322924
rect 42300 322912 42306 322924
rect 43162 322912 43168 322924
rect 42300 322884 43168 322912
rect 42300 322872 42306 322884
rect 43162 322872 43168 322884
rect 43220 322872 43226 322924
rect 42242 320220 42248 320272
rect 42300 320220 42306 320272
rect 42260 320124 42288 320220
rect 42260 320096 42656 320124
rect 42628 320000 42656 320096
rect 42610 319948 42616 320000
rect 42668 319948 42674 320000
rect 60366 315936 60372 315988
rect 60424 315976 60430 315988
rect 62114 315976 62120 315988
rect 60424 315948 62120 315976
rect 60424 315936 60430 315948
rect 62114 315936 62120 315948
rect 62172 315936 62178 315988
rect 51074 314712 51080 314764
rect 51132 314752 51138 314764
rect 62114 314752 62120 314764
rect 51132 314724 62120 314752
rect 51132 314712 51138 314724
rect 62114 314712 62120 314724
rect 62172 314712 62178 314764
rect 46382 309068 46388 309120
rect 46440 309108 46446 309120
rect 47762 309108 47768 309120
rect 46440 309080 47768 309108
rect 46440 309068 46446 309080
rect 47762 309068 47768 309080
rect 47820 309068 47826 309120
rect 676214 306348 676220 306400
rect 676272 306388 676278 306400
rect 676858 306388 676864 306400
rect 676272 306360 676864 306388
rect 676272 306348 676278 306360
rect 676858 306348 676864 306360
rect 676916 306348 676922 306400
rect 675846 304920 675852 304972
rect 675904 304960 675910 304972
rect 676398 304960 676404 304972
rect 675904 304932 676404 304960
rect 675904 304920 675910 304932
rect 676398 304920 676404 304932
rect 676456 304920 676462 304972
rect 651374 303492 651380 303544
rect 651432 303532 651438 303544
rect 653398 303532 653404 303544
rect 651432 303504 653404 303532
rect 651432 303492 651438 303504
rect 653398 303492 653404 303504
rect 653456 303492 653462 303544
rect 651466 300772 651472 300824
rect 651524 300812 651530 300824
rect 660298 300812 660304 300824
rect 651524 300784 660304 300812
rect 651524 300772 651530 300784
rect 660298 300772 660304 300784
rect 660356 300772 660362 300824
rect 41138 299616 41144 299668
rect 41196 299656 41202 299668
rect 41598 299656 41604 299668
rect 41196 299628 41604 299656
rect 41196 299616 41202 299628
rect 41598 299616 41604 299628
rect 41656 299616 41662 299668
rect 675846 297032 675852 297084
rect 675904 297072 675910 297084
rect 679618 297072 679624 297084
rect 675904 297044 679624 297072
rect 675904 297032 675910 297044
rect 679618 297032 679624 297044
rect 679676 297032 679682 297084
rect 651926 296760 651932 296812
rect 651984 296800 651990 296812
rect 651984 296772 654134 296800
rect 651984 296760 651990 296772
rect 654106 296732 654134 296772
rect 665818 296732 665824 296744
rect 654106 296704 665824 296732
rect 665818 296692 665824 296704
rect 665876 296692 665882 296744
rect 675478 296352 675484 296404
rect 675536 296352 675542 296404
rect 41322 295604 41328 295656
rect 41380 295644 41386 295656
rect 41690 295644 41696 295656
rect 41380 295616 41696 295644
rect 41380 295604 41386 295616
rect 41690 295604 41696 295616
rect 41748 295604 41754 295656
rect 50522 295332 50528 295384
rect 50580 295372 50586 295384
rect 62114 295372 62120 295384
rect 50580 295344 62120 295372
rect 50580 295332 50586 295344
rect 62114 295332 62120 295344
rect 62172 295332 62178 295384
rect 675496 295248 675524 296352
rect 675478 295196 675484 295248
rect 675536 295196 675542 295248
rect 57238 294040 57244 294092
rect 57296 294080 57302 294092
rect 62114 294080 62120 294092
rect 57296 294052 62120 294080
rect 57296 294040 57302 294052
rect 62114 294040 62120 294052
rect 62172 294040 62178 294092
rect 651466 293972 651472 294024
rect 651524 294012 651530 294024
rect 664438 294012 664444 294024
rect 651524 293984 664444 294012
rect 651524 293972 651530 293984
rect 664438 293972 664444 293984
rect 664496 293972 664502 294024
rect 51902 292544 51908 292596
rect 51960 292584 51966 292596
rect 62114 292584 62120 292596
rect 51960 292556 62120 292584
rect 51960 292544 51966 292556
rect 62114 292544 62120 292556
rect 62172 292544 62178 292596
rect 41138 292204 41144 292256
rect 41196 292244 41202 292256
rect 41598 292244 41604 292256
rect 41196 292216 41604 292244
rect 41196 292204 41202 292216
rect 41598 292204 41604 292216
rect 41656 292204 41662 292256
rect 47578 292136 47584 292188
rect 47636 292176 47642 292188
rect 53466 292176 53472 292188
rect 47636 292148 53472 292176
rect 47636 292136 47642 292148
rect 53466 292136 53472 292148
rect 53524 292136 53530 292188
rect 47762 292000 47768 292052
rect 47820 292040 47826 292052
rect 53650 292040 53656 292052
rect 47820 292012 53656 292040
rect 47820 292000 47826 292012
rect 53650 292000 53656 292012
rect 53708 292000 53714 292052
rect 41230 291252 41236 291304
rect 41288 291292 41294 291304
rect 41690 291292 41696 291304
rect 41288 291264 41696 291292
rect 41288 291252 41294 291264
rect 41690 291252 41696 291264
rect 41748 291252 41754 291304
rect 651466 291184 651472 291236
rect 651524 291224 651530 291236
rect 663058 291224 663064 291236
rect 651524 291196 663064 291224
rect 651524 291184 651530 291196
rect 663058 291184 663064 291196
rect 663116 291184 663122 291236
rect 53282 291116 53288 291168
rect 53340 291156 53346 291168
rect 62114 291156 62120 291168
rect 53340 291128 62120 291156
rect 53340 291116 53346 291128
rect 62114 291116 62120 291128
rect 62172 291116 62178 291168
rect 651374 290368 651380 290420
rect 651432 290408 651438 290420
rect 653398 290408 653404 290420
rect 651432 290380 653404 290408
rect 651432 290368 651438 290380
rect 653398 290368 653404 290380
rect 653456 290368 653462 290420
rect 651466 288396 651472 288448
rect 651524 288436 651530 288448
rect 672166 288436 672172 288448
rect 651524 288408 672172 288436
rect 651524 288396 651530 288408
rect 672166 288396 672172 288408
rect 672224 288396 672230 288448
rect 651466 287036 651472 287088
rect 651524 287076 651530 287088
rect 667566 287076 667572 287088
rect 651524 287048 667572 287076
rect 651524 287036 651530 287048
rect 667566 287036 667572 287048
rect 667624 287036 667630 287088
rect 33778 286288 33784 286340
rect 33836 286328 33842 286340
rect 41690 286328 41696 286340
rect 33836 286300 41696 286328
rect 33836 286288 33842 286300
rect 41690 286288 41696 286300
rect 41748 286288 41754 286340
rect 46382 285676 46388 285728
rect 46440 285716 46446 285728
rect 63034 285716 63040 285728
rect 46440 285688 63040 285716
rect 46440 285676 46446 285688
rect 63034 285676 63040 285688
rect 63092 285676 63098 285728
rect 651466 285676 651472 285728
rect 651524 285716 651530 285728
rect 667382 285716 667388 285728
rect 651524 285688 667388 285716
rect 651524 285676 651530 285688
rect 667382 285676 667388 285688
rect 667440 285676 667446 285728
rect 674466 285608 674472 285660
rect 674524 285648 674530 285660
rect 675110 285648 675116 285660
rect 674524 285620 675116 285648
rect 674524 285608 674530 285620
rect 675110 285608 675116 285620
rect 675168 285608 675174 285660
rect 53650 284928 53656 284980
rect 53708 284968 53714 284980
rect 56318 284968 56324 284980
rect 53708 284940 56324 284968
rect 53708 284928 53714 284940
rect 56318 284928 56324 284940
rect 56376 284928 56382 284980
rect 39298 284724 39304 284776
rect 39356 284764 39362 284776
rect 41690 284764 41696 284776
rect 39356 284736 41696 284764
rect 39356 284724 39362 284736
rect 41690 284724 41696 284736
rect 41748 284724 41754 284776
rect 42058 284656 42064 284708
rect 42116 284696 42122 284708
rect 42610 284696 42616 284708
rect 42116 284668 42616 284696
rect 42116 284656 42122 284668
rect 42610 284656 42616 284668
rect 42668 284656 42674 284708
rect 60366 284384 60372 284436
rect 60424 284424 60430 284436
rect 62114 284424 62120 284436
rect 60424 284396 62120 284424
rect 60424 284384 60430 284396
rect 62114 284384 62120 284396
rect 62172 284384 62178 284436
rect 651466 284316 651472 284368
rect 651524 284356 651530 284368
rect 672350 284356 672356 284368
rect 651524 284328 672356 284356
rect 651524 284316 651530 284328
rect 672350 284316 672356 284328
rect 672408 284316 672414 284368
rect 47762 282888 47768 282940
rect 47820 282928 47826 282940
rect 62114 282928 62120 282940
rect 47820 282900 62120 282928
rect 47820 282888 47826 282900
rect 62114 282888 62120 282900
rect 62172 282888 62178 282940
rect 651466 282140 651472 282192
rect 651524 282180 651530 282192
rect 666554 282180 666560 282192
rect 651524 282152 666560 282180
rect 651524 282140 651530 282152
rect 666554 282140 666560 282152
rect 666612 282140 666618 282192
rect 53282 281528 53288 281580
rect 53340 281568 53346 281580
rect 62114 281568 62120 281580
rect 53340 281540 62120 281568
rect 53340 281528 53346 281540
rect 62114 281528 62120 281540
rect 62172 281528 62178 281580
rect 58802 280168 58808 280220
rect 58860 280208 58866 280220
rect 62114 280208 62120 280220
rect 58860 280180 62120 280208
rect 58860 280168 58866 280180
rect 62114 280168 62120 280180
rect 62172 280168 62178 280220
rect 651466 280168 651472 280220
rect 651524 280208 651530 280220
rect 667198 280208 667204 280220
rect 651524 280180 667204 280208
rect 651524 280168 651530 280180
rect 667198 280168 667204 280180
rect 667256 280168 667262 280220
rect 62574 278672 62580 278724
rect 62632 278712 62638 278724
rect 671338 278712 671344 278724
rect 62632 278684 671344 278712
rect 62632 278672 62638 278684
rect 671338 278672 671344 278684
rect 671396 278672 671402 278724
rect 63402 278536 63408 278588
rect 63460 278576 63466 278588
rect 671706 278576 671712 278588
rect 63460 278548 671712 278576
rect 63460 278536 63466 278548
rect 671706 278536 671712 278548
rect 671764 278536 671770 278588
rect 56042 278400 56048 278452
rect 56100 278440 56106 278452
rect 651006 278440 651012 278452
rect 56100 278412 651012 278440
rect 56100 278400 56106 278412
rect 651006 278400 651012 278412
rect 651064 278400 651070 278452
rect 51718 278264 51724 278316
rect 51776 278304 51782 278316
rect 634998 278304 635004 278316
rect 51776 278276 635004 278304
rect 51776 278264 51782 278276
rect 634998 278264 635004 278276
rect 635056 278264 635062 278316
rect 47946 278128 47952 278180
rect 48004 278168 48010 278180
rect 637758 278168 637764 278180
rect 48004 278140 637764 278168
rect 48004 278128 48010 278140
rect 637758 278128 637764 278140
rect 637816 278128 637822 278180
rect 64138 277992 64144 278044
rect 64196 278032 64202 278044
rect 667934 278032 667940 278044
rect 64196 278004 667940 278032
rect 64196 277992 64202 278004
rect 667934 277992 667940 278004
rect 667992 277992 667998 278044
rect 53466 277856 53472 277908
rect 53524 277896 53530 277908
rect 53524 277868 68784 277896
rect 53524 277856 53530 277868
rect 56318 277720 56324 277772
rect 56376 277760 56382 277772
rect 68756 277760 68784 277868
rect 69658 277856 69664 277908
rect 69716 277896 69722 277908
rect 629478 277896 629484 277908
rect 69716 277868 629484 277896
rect 69716 277856 69722 277868
rect 629478 277856 629484 277868
rect 629536 277856 629542 277908
rect 650822 277896 650828 277908
rect 629956 277868 650828 277896
rect 629956 277760 629984 277868
rect 650822 277856 650828 277868
rect 650880 277856 650886 277908
rect 650638 277760 650644 277772
rect 56376 277732 68692 277760
rect 68756 277732 629984 277760
rect 630048 277732 650644 277760
rect 56376 277720 56382 277732
rect 64322 277584 64328 277636
rect 64380 277624 64386 277636
rect 68664 277624 68692 277732
rect 630048 277624 630076 277732
rect 650638 277720 650644 277732
rect 650696 277720 650702 277772
rect 636194 277624 636200 277636
rect 64380 277596 64874 277624
rect 68664 277596 630076 277624
rect 634786 277596 636200 277624
rect 64380 277584 64386 277596
rect 64846 277488 64874 277596
rect 69658 277488 69664 277500
rect 64846 277460 69664 277488
rect 69658 277448 69664 277460
rect 69716 277448 69722 277500
rect 629478 277448 629484 277500
rect 629536 277488 629542 277500
rect 634786 277488 634814 277596
rect 636194 277584 636200 277596
rect 636252 277584 636258 277636
rect 629536 277460 634814 277488
rect 629536 277448 629542 277460
rect 42242 277312 42248 277364
rect 42300 277352 42306 277364
rect 42794 277352 42800 277364
rect 42300 277324 42800 277352
rect 42300 277312 42306 277324
rect 42794 277312 42800 277324
rect 42852 277312 42858 277364
rect 482830 277312 482836 277364
rect 482888 277352 482894 277364
rect 557534 277352 557540 277364
rect 482888 277324 557540 277352
rect 482888 277312 482894 277324
rect 557534 277312 557540 277324
rect 557592 277312 557598 277364
rect 487982 277176 487988 277228
rect 488040 277216 488046 277228
rect 565814 277216 565820 277228
rect 488040 277188 565820 277216
rect 488040 277176 488046 277188
rect 565814 277176 565820 277188
rect 565872 277176 565878 277228
rect 497918 277040 497924 277092
rect 497976 277080 497982 277092
rect 579982 277080 579988 277092
rect 497976 277052 579988 277080
rect 497976 277040 497982 277052
rect 579982 277040 579988 277052
rect 580040 277040 580046 277092
rect 511626 276904 511632 276956
rect 511684 276944 511690 276956
rect 600130 276944 600136 276956
rect 511684 276916 600136 276944
rect 511684 276904 511690 276916
rect 600130 276904 600136 276916
rect 600188 276904 600194 276956
rect 514478 276768 514484 276820
rect 514536 276808 514542 276820
rect 603626 276808 603632 276820
rect 514536 276780 603632 276808
rect 514536 276768 514542 276780
rect 603626 276768 603632 276780
rect 603684 276768 603690 276820
rect 518710 276632 518716 276684
rect 518768 276672 518774 276684
rect 609606 276672 609612 276684
rect 518768 276644 609612 276672
rect 518768 276632 518774 276644
rect 609606 276632 609612 276644
rect 609664 276632 609670 276684
rect 479978 276496 479984 276548
rect 480036 276536 480042 276548
rect 555234 276536 555240 276548
rect 480036 276508 555240 276536
rect 480036 276496 480042 276508
rect 555234 276496 555240 276508
rect 555292 276496 555298 276548
rect 477034 276360 477040 276412
rect 477092 276400 477098 276412
rect 550450 276400 550456 276412
rect 477092 276372 550456 276400
rect 477092 276360 477098 276372
rect 550450 276360 550456 276372
rect 550508 276360 550514 276412
rect 471606 276224 471612 276276
rect 471664 276264 471670 276276
rect 543366 276264 543372 276276
rect 471664 276236 543372 276264
rect 471664 276224 471670 276236
rect 543366 276224 543372 276236
rect 543424 276224 543430 276276
rect 107194 275952 107200 276004
rect 107252 275992 107258 276004
rect 163498 275992 163504 276004
rect 107252 275964 163504 275992
rect 107252 275952 107258 275964
rect 163498 275952 163504 275964
rect 163556 275952 163562 276004
rect 167546 275952 167552 276004
rect 167604 275992 167610 276004
rect 178862 275992 178868 276004
rect 167604 275964 178868 275992
rect 167604 275952 167610 275964
rect 178862 275952 178868 275964
rect 178920 275952 178926 276004
rect 185210 275952 185216 276004
rect 185268 275992 185274 276004
rect 221274 275992 221280 276004
rect 185268 275964 221280 275992
rect 185268 275952 185274 275964
rect 221274 275952 221280 275964
rect 221332 275952 221338 276004
rect 232498 275952 232504 276004
rect 232556 275992 232562 276004
rect 239214 275992 239220 276004
rect 232556 275964 239220 275992
rect 232556 275952 232562 275964
rect 239214 275952 239220 275964
rect 239272 275952 239278 276004
rect 410794 275952 410800 276004
rect 410852 275992 410858 276004
rect 455874 275992 455880 276004
rect 410852 275964 455880 275992
rect 410852 275952 410858 275964
rect 455874 275952 455880 275964
rect 455932 275952 455938 276004
rect 456058 275952 456064 276004
rect 456116 275992 456122 276004
rect 509050 275992 509056 276004
rect 456116 275964 509056 275992
rect 456116 275952 456122 275964
rect 509050 275952 509056 275964
rect 509108 275952 509114 276004
rect 513190 275952 513196 276004
rect 513248 275992 513254 276004
rect 601326 275992 601332 276004
rect 513248 275964 601332 275992
rect 513248 275952 513254 275964
rect 601326 275952 601332 275964
rect 601384 275952 601390 276004
rect 139118 275816 139124 275868
rect 139176 275856 139182 275868
rect 174262 275856 174268 275868
rect 139176 275828 174268 275856
rect 139176 275816 139182 275828
rect 174262 275816 174268 275828
rect 174320 275816 174326 275868
rect 178126 275816 178132 275868
rect 178184 275856 178190 275868
rect 216674 275856 216680 275868
rect 178184 275828 216680 275856
rect 178184 275816 178190 275828
rect 216674 275816 216680 275828
rect 216732 275816 216738 275868
rect 224218 275816 224224 275868
rect 224276 275856 224282 275868
rect 232682 275856 232688 275868
rect 224276 275828 232688 275856
rect 224276 275816 224282 275828
rect 232682 275816 232688 275828
rect 232740 275816 232746 275868
rect 236086 275816 236092 275868
rect 236144 275856 236150 275868
rect 250438 275856 250444 275868
rect 236144 275828 250444 275856
rect 236144 275816 236150 275828
rect 250438 275816 250444 275828
rect 250496 275816 250502 275868
rect 286870 275816 286876 275868
rect 286928 275856 286934 275868
rect 291838 275856 291844 275868
rect 286928 275828 291844 275856
rect 286928 275816 286934 275828
rect 291838 275816 291844 275828
rect 291896 275816 291902 275868
rect 430206 275816 430212 275868
rect 430264 275856 430270 275868
rect 484302 275856 484308 275868
rect 430264 275828 484308 275856
rect 430264 275816 430270 275828
rect 484302 275816 484308 275828
rect 484360 275816 484366 275868
rect 490558 275816 490564 275868
rect 490616 275856 490622 275868
rect 505554 275856 505560 275868
rect 490616 275828 505560 275856
rect 490616 275816 490622 275828
rect 505554 275816 505560 275828
rect 505612 275816 505618 275868
rect 522758 275816 522764 275868
rect 522816 275856 522822 275868
rect 615494 275856 615500 275868
rect 522816 275828 615500 275856
rect 522816 275816 522822 275828
rect 615494 275816 615500 275828
rect 615552 275816 615558 275868
rect 260926 275748 260932 275800
rect 260984 275788 260990 275800
rect 266354 275788 266360 275800
rect 260984 275760 266360 275788
rect 260984 275748 260990 275760
rect 266354 275748 266360 275760
rect 266412 275748 266418 275800
rect 93026 275680 93032 275732
rect 93084 275720 93090 275732
rect 152826 275720 152832 275732
rect 93084 275692 152832 275720
rect 93084 275680 93090 275692
rect 152826 275680 152832 275692
rect 152884 275680 152890 275732
rect 160462 275680 160468 275732
rect 160520 275720 160526 275732
rect 199562 275720 199568 275732
rect 160520 275692 199568 275720
rect 160520 275680 160526 275692
rect 199562 275680 199568 275692
rect 199620 275680 199626 275732
rect 217134 275680 217140 275732
rect 217192 275720 217198 275732
rect 224218 275720 224224 275732
rect 217192 275692 224224 275720
rect 217192 275680 217198 275692
rect 224218 275680 224224 275692
rect 224276 275680 224282 275732
rect 229002 275680 229008 275732
rect 229060 275720 229066 275732
rect 243538 275720 243544 275732
rect 229060 275692 243544 275720
rect 229060 275680 229066 275692
rect 243538 275680 243544 275692
rect 243596 275680 243602 275732
rect 250254 275680 250260 275732
rect 250312 275720 250318 275732
rect 259362 275720 259368 275732
rect 250312 275692 259368 275720
rect 250312 275680 250318 275692
rect 259362 275680 259368 275692
rect 259420 275680 259426 275732
rect 284570 275680 284576 275732
rect 284628 275720 284634 275732
rect 290090 275720 290096 275732
rect 284628 275692 290096 275720
rect 284628 275680 284634 275692
rect 290090 275680 290096 275692
rect 290148 275680 290154 275732
rect 416406 275680 416412 275732
rect 416464 275720 416470 275732
rect 462958 275720 462964 275732
rect 416464 275692 462964 275720
rect 416464 275680 416470 275692
rect 462958 275680 462964 275692
rect 463016 275680 463022 275732
rect 463142 275680 463148 275732
rect 463200 275720 463206 275732
rect 516226 275720 516232 275732
rect 463200 275692 516232 275720
rect 463200 275680 463206 275692
rect 516226 275680 516232 275692
rect 516284 275680 516290 275732
rect 528186 275680 528192 275732
rect 528244 275720 528250 275732
rect 622578 275720 622584 275732
rect 528244 275692 622584 275720
rect 528244 275680 528250 275692
rect 622578 275680 622584 275692
rect 622636 275680 622642 275732
rect 76466 275544 76472 275596
rect 76524 275584 76530 275596
rect 86218 275584 86224 275596
rect 76524 275556 86224 275584
rect 76524 275544 76530 275556
rect 86218 275544 86224 275556
rect 86276 275544 86282 275596
rect 90726 275544 90732 275596
rect 90784 275584 90790 275596
rect 154758 275584 154764 275596
rect 90784 275556 154764 275584
rect 90784 275544 90790 275556
rect 154758 275544 154764 275556
rect 154816 275544 154822 275596
rect 171042 275544 171048 275596
rect 171100 275584 171106 275596
rect 211614 275584 211620 275596
rect 171100 275556 211620 275584
rect 171100 275544 171106 275556
rect 211614 275544 211620 275556
rect 211672 275544 211678 275596
rect 218330 275544 218336 275596
rect 218388 275584 218394 275596
rect 233878 275584 233884 275596
rect 218388 275556 233884 275584
rect 218388 275544 218394 275556
rect 233878 275544 233884 275556
rect 233936 275544 233942 275596
rect 239582 275544 239588 275596
rect 239640 275584 239646 275596
rect 255958 275584 255964 275596
rect 239640 275556 255964 275584
rect 239640 275544 239646 275556
rect 255958 275544 255964 275556
rect 256016 275544 256022 275596
rect 257338 275544 257344 275596
rect 257396 275584 257402 275596
rect 262306 275584 262312 275596
rect 257396 275556 262312 275584
rect 257396 275544 257402 275556
rect 262306 275544 262312 275556
rect 262364 275544 262370 275596
rect 266814 275544 266820 275596
rect 266872 275584 266878 275596
rect 276474 275584 276480 275596
rect 266872 275556 276480 275584
rect 266872 275544 266878 275556
rect 276474 275544 276480 275556
rect 276532 275544 276538 275596
rect 363874 275544 363880 275596
rect 363932 275584 363938 275596
rect 388530 275584 388536 275596
rect 363932 275556 388536 275584
rect 363932 275544 363938 275556
rect 388530 275544 388536 275556
rect 388588 275544 388594 275596
rect 445018 275544 445024 275596
rect 445076 275584 445082 275596
rect 498470 275584 498476 275596
rect 445076 275556 498476 275584
rect 445076 275544 445082 275556
rect 498470 275544 498476 275556
rect 498528 275544 498534 275596
rect 498838 275544 498844 275596
rect 498896 275584 498902 275596
rect 512638 275584 512644 275596
rect 498896 275556 512644 275584
rect 498896 275544 498902 275556
rect 512638 275544 512644 275556
rect 512696 275544 512702 275596
rect 516778 275544 516784 275596
rect 516836 275584 516842 275596
rect 526806 275584 526812 275596
rect 516836 275556 526812 275584
rect 516836 275544 516842 275556
rect 526806 275544 526812 275556
rect 526864 275544 526870 275596
rect 532326 275544 532332 275596
rect 532384 275584 532390 275596
rect 629662 275584 629668 275596
rect 532384 275556 629668 275584
rect 532384 275544 532390 275556
rect 629662 275544 629668 275556
rect 629720 275544 629726 275596
rect 277486 275476 277492 275528
rect 277544 275516 277550 275528
rect 285122 275516 285128 275528
rect 277544 275488 285128 275516
rect 277544 275476 277550 275488
rect 285122 275476 285128 275488
rect 285180 275476 285186 275528
rect 100110 275408 100116 275460
rect 100168 275448 100174 275460
rect 100168 275420 142154 275448
rect 100168 275408 100174 275420
rect 71774 275272 71780 275324
rect 71832 275312 71838 275324
rect 141050 275312 141056 275324
rect 71832 275284 141056 275312
rect 71832 275272 71838 275284
rect 141050 275272 141056 275284
rect 141108 275272 141114 275324
rect 142126 275312 142154 275420
rect 156874 275408 156880 275460
rect 156932 275448 156938 275460
rect 156932 275420 161474 275448
rect 156932 275408 156938 275420
rect 159450 275312 159456 275324
rect 142126 275284 159456 275312
rect 159450 275272 159456 275284
rect 159508 275272 159514 275324
rect 161446 275312 161474 275420
rect 163958 275408 163964 275460
rect 164016 275448 164022 275460
rect 206370 275448 206376 275460
rect 164016 275420 206376 275448
rect 164016 275408 164022 275420
rect 206370 275408 206376 275420
rect 206428 275408 206434 275460
rect 221918 275408 221924 275460
rect 221976 275448 221982 275460
rect 243722 275448 243728 275460
rect 221976 275420 243728 275448
rect 221976 275408 221982 275420
rect 243722 275408 243728 275420
rect 243780 275408 243786 275460
rect 256142 275408 256148 275460
rect 256200 275448 256206 275460
rect 256200 275420 269068 275448
rect 256200 275408 256206 275420
rect 200758 275312 200764 275324
rect 161446 275284 200764 275312
rect 200758 275272 200764 275284
rect 200816 275272 200822 275324
rect 214834 275272 214840 275324
rect 214892 275312 214898 275324
rect 239398 275312 239404 275324
rect 214892 275284 239404 275312
rect 214892 275272 214898 275284
rect 239398 275272 239404 275284
rect 239456 275272 239462 275324
rect 243170 275272 243176 275324
rect 243228 275312 243234 275324
rect 256694 275312 256700 275324
rect 243228 275284 256700 275312
rect 243228 275272 243234 275284
rect 256694 275272 256700 275284
rect 256752 275272 256758 275324
rect 269040 275244 269068 275420
rect 358630 275408 358636 275460
rect 358688 275448 358694 275460
rect 381446 275448 381452 275460
rect 358688 275420 381452 275448
rect 358688 275408 358694 275420
rect 381446 275408 381452 275420
rect 381504 275408 381510 275460
rect 386046 275408 386052 275460
rect 386104 275448 386110 275460
rect 420454 275448 420460 275460
rect 386104 275420 420460 275448
rect 386104 275408 386110 275420
rect 420454 275408 420460 275420
rect 420512 275408 420518 275460
rect 435634 275408 435640 275460
rect 435692 275448 435698 275460
rect 485038 275448 485044 275460
rect 435692 275420 485044 275448
rect 435692 275408 435698 275420
rect 485038 275408 485044 275420
rect 485096 275408 485102 275460
rect 485222 275408 485228 275460
rect 485280 275448 485286 275460
rect 530394 275448 530400 275460
rect 485280 275420 530400 275448
rect 485280 275408 485286 275420
rect 530394 275408 530400 275420
rect 530452 275408 530458 275460
rect 537662 275408 537668 275460
rect 537720 275448 537726 275460
rect 636746 275448 636752 275460
rect 537720 275420 636752 275448
rect 537720 275408 537726 275420
rect 636746 275408 636752 275420
rect 636804 275408 636810 275460
rect 269206 275340 269212 275392
rect 269264 275380 269270 275392
rect 274634 275380 274640 275392
rect 269264 275352 274640 275380
rect 269264 275340 269270 275352
rect 274634 275340 274640 275352
rect 274692 275340 274698 275392
rect 276290 275272 276296 275324
rect 276348 275312 276354 275324
rect 283098 275312 283104 275324
rect 276348 275284 283104 275312
rect 276348 275272 276354 275284
rect 283098 275272 283104 275284
rect 283156 275272 283162 275324
rect 285674 275272 285680 275324
rect 285732 275312 285738 275324
rect 291286 275312 291292 275324
rect 285732 275284 291292 275312
rect 285732 275272 285738 275284
rect 291286 275272 291292 275284
rect 291344 275272 291350 275324
rect 291654 275272 291660 275324
rect 291712 275312 291718 275324
rect 295334 275312 295340 275324
rect 291712 275284 295340 275312
rect 291712 275272 291718 275284
rect 295334 275272 295340 275284
rect 295392 275272 295398 275324
rect 299934 275272 299940 275324
rect 299992 275312 299998 275324
rect 301130 275312 301136 275324
rect 299992 275284 301136 275312
rect 299992 275272 299998 275284
rect 301130 275272 301136 275284
rect 301188 275272 301194 275324
rect 326430 275272 326436 275324
rect 326488 275312 326494 275324
rect 335354 275312 335360 275324
rect 326488 275284 335360 275312
rect 326488 275272 326494 275284
rect 335354 275272 335360 275284
rect 335412 275272 335418 275324
rect 371050 275272 371056 275324
rect 371108 275312 371114 275324
rect 399202 275312 399208 275324
rect 371108 275284 399208 275312
rect 371108 275272 371114 275284
rect 399202 275272 399208 275284
rect 399260 275272 399266 275324
rect 418798 275272 418804 275324
rect 418856 275312 418862 275324
rect 466546 275312 466552 275324
rect 418856 275284 466552 275312
rect 418856 275272 418862 275284
rect 466546 275272 466552 275284
rect 466604 275272 466610 275324
rect 467558 275272 467564 275324
rect 467616 275312 467622 275324
rect 537478 275312 537484 275324
rect 467616 275284 537484 275312
rect 467616 275272 467622 275284
rect 537478 275272 537484 275284
rect 537536 275272 537542 275324
rect 542262 275272 542268 275324
rect 542320 275312 542326 275324
rect 643830 275312 643836 275324
rect 542320 275284 643836 275312
rect 542320 275272 542326 275284
rect 643830 275272 643836 275284
rect 643888 275272 643894 275324
rect 270126 275244 270132 275256
rect 269040 275216 270132 275244
rect 270126 275204 270132 275216
rect 270184 275204 270190 275256
rect 96614 275136 96620 275188
rect 96672 275176 96678 275188
rect 149606 275176 149612 275188
rect 96672 275148 149612 275176
rect 96672 275136 96678 275148
rect 149606 275136 149612 275148
rect 149664 275136 149670 275188
rect 153378 275136 153384 275188
rect 153436 275176 153442 275188
rect 169018 275176 169024 275188
rect 153436 275148 169024 275176
rect 153436 275136 153442 275148
rect 169018 275136 169024 275148
rect 169076 275136 169082 275188
rect 189994 275136 190000 275188
rect 190052 275176 190058 275188
rect 222930 275176 222936 275188
rect 190052 275148 222936 275176
rect 190052 275136 190058 275148
rect 222930 275136 222936 275148
rect 222988 275136 222994 275188
rect 292850 275136 292856 275188
rect 292908 275176 292914 275188
rect 295794 275176 295800 275188
rect 292908 275148 295800 275176
rect 292908 275136 292914 275148
rect 295794 275136 295800 275148
rect 295852 275136 295858 275188
rect 298738 275136 298744 275188
rect 298796 275176 298802 275188
rect 300026 275176 300032 275188
rect 298796 275148 300032 275176
rect 298796 275136 298802 275148
rect 300026 275136 300032 275148
rect 300084 275136 300090 275188
rect 427078 275136 427084 275188
rect 427136 275176 427142 275188
rect 477218 275176 477224 275188
rect 427136 275148 477224 275176
rect 427136 275136 427142 275148
rect 477218 275136 477224 275148
rect 477276 275136 477282 275188
rect 485038 275136 485044 275188
rect 485096 275176 485102 275188
rect 491386 275176 491392 275188
rect 485096 275148 491392 275176
rect 485096 275136 485102 275148
rect 491386 275136 491392 275148
rect 491444 275136 491450 275188
rect 507486 275136 507492 275188
rect 507544 275176 507550 275188
rect 594242 275176 594248 275188
rect 507544 275148 594248 275176
rect 507544 275136 507550 275148
rect 594242 275136 594248 275148
rect 594300 275136 594306 275188
rect 263226 275068 263232 275120
rect 263284 275108 263290 275120
rect 273254 275108 273260 275120
rect 263284 275080 273260 275108
rect 263284 275068 263290 275080
rect 273254 275068 273260 275080
rect 273312 275068 273318 275120
rect 136818 275000 136824 275052
rect 136876 275040 136882 275052
rect 137646 275040 137652 275052
rect 136876 275012 137652 275040
rect 136876 275000 136882 275012
rect 137646 275000 137652 275012
rect 137704 275000 137710 275052
rect 146202 275000 146208 275052
rect 146260 275040 146266 275052
rect 185302 275040 185308 275052
rect 146260 275012 185308 275040
rect 146260 275000 146266 275012
rect 185302 275000 185308 275012
rect 185360 275000 185366 275052
rect 288066 275000 288072 275052
rect 288124 275040 288130 275052
rect 292850 275040 292856 275052
rect 288124 275012 292856 275040
rect 288124 275000 288130 275012
rect 292850 275000 292856 275012
rect 292908 275000 292914 275052
rect 420546 275000 420552 275052
rect 420604 275040 420610 275052
rect 470134 275040 470140 275052
rect 420604 275012 470140 275040
rect 420604 275000 420610 275012
rect 470134 275000 470140 275012
rect 470192 275000 470198 275052
rect 484302 275000 484308 275052
rect 484360 275040 484366 275052
rect 485222 275040 485228 275052
rect 484360 275012 485228 275040
rect 484360 275000 484366 275012
rect 485222 275000 485228 275012
rect 485280 275000 485286 275052
rect 503438 275000 503444 275052
rect 503496 275040 503502 275052
rect 587066 275040 587072 275052
rect 503496 275012 587072 275040
rect 503496 275000 503502 275012
rect 587066 275000 587072 275012
rect 587124 275000 587130 275052
rect 81250 274932 81256 274984
rect 81308 274972 81314 274984
rect 81308 274944 84194 274972
rect 81308 274932 81314 274944
rect 84166 274904 84194 274944
rect 293954 274932 293960 274984
rect 294012 274972 294018 274984
rect 297174 274972 297180 274984
rect 294012 274944 297180 274972
rect 294012 274932 294018 274944
rect 297174 274932 297180 274944
rect 297232 274932 297238 274984
rect 145282 274904 145288 274916
rect 84166 274876 145288 274904
rect 145282 274864 145288 274876
rect 145340 274864 145346 274916
rect 149790 274864 149796 274916
rect 149848 274904 149854 274916
rect 189074 274904 189080 274916
rect 149848 274876 189080 274904
rect 149848 274864 149854 274876
rect 189074 274864 189080 274876
rect 189132 274864 189138 274916
rect 289262 274864 289268 274916
rect 289320 274904 289326 274916
rect 292666 274904 292672 274916
rect 289320 274876 292672 274904
rect 289320 274864 289326 274876
rect 292666 274864 292672 274876
rect 292724 274864 292730 274916
rect 473078 274864 473084 274916
rect 473136 274904 473142 274916
rect 544562 274904 544568 274916
rect 473136 274876 544568 274904
rect 473136 274864 473142 274876
rect 544562 274864 544568 274876
rect 544620 274864 544626 274916
rect 296346 274796 296352 274848
rect 296404 274836 296410 274848
rect 298370 274836 298376 274848
rect 296404 274808 298376 274836
rect 296404 274796 296410 274808
rect 298370 274796 298376 274808
rect 298428 274796 298434 274848
rect 128538 274728 128544 274780
rect 128596 274768 128602 274780
rect 168282 274768 168288 274780
rect 128596 274740 168288 274768
rect 128596 274728 128602 274740
rect 168282 274728 168288 274740
rect 168340 274728 168346 274780
rect 207750 274728 207756 274780
rect 207808 274768 207814 274780
rect 210694 274768 210700 274780
rect 207808 274740 210700 274768
rect 207808 274728 207814 274740
rect 210694 274728 210700 274740
rect 210752 274728 210758 274780
rect 476758 274728 476764 274780
rect 476816 274768 476822 274780
rect 523310 274768 523316 274780
rect 476816 274740 523316 274768
rect 476816 274728 476822 274740
rect 523310 274728 523316 274740
rect 523368 274728 523374 274780
rect 523678 274728 523684 274780
rect 523736 274768 523742 274780
rect 533890 274768 533896 274780
rect 523736 274740 533896 274768
rect 523736 274728 523742 274740
rect 533890 274728 533896 274740
rect 533948 274728 533954 274780
rect 534718 274728 534724 274780
rect 534776 274768 534782 274780
rect 540974 274768 540980 274780
rect 534776 274740 540980 274768
rect 534776 274728 534782 274740
rect 540974 274728 540980 274740
rect 541032 274728 541038 274780
rect 74166 274660 74172 274712
rect 74224 274700 74230 274712
rect 76834 274700 76840 274712
rect 74224 274672 76840 274700
rect 74224 274660 74230 274672
rect 76834 274660 76840 274672
rect 76892 274660 76898 274712
rect 85942 274660 85948 274712
rect 86000 274700 86006 274712
rect 90358 274700 90364 274712
rect 86000 274672 90364 274700
rect 86000 274660 86006 274672
rect 90358 274660 90364 274672
rect 90416 274660 90422 274712
rect 103698 274660 103704 274712
rect 103756 274700 103762 274712
rect 104802 274700 104808 274712
rect 103756 274672 104808 274700
rect 103756 274660 103762 274672
rect 104802 274660 104808 274672
rect 104860 274660 104866 274712
rect 110782 274660 110788 274712
rect 110840 274700 110846 274712
rect 111702 274700 111708 274712
rect 110840 274672 111708 274700
rect 110840 274660 110846 274672
rect 111702 274660 111708 274672
rect 111760 274660 111766 274712
rect 253842 274660 253848 274712
rect 253900 274700 253906 274712
rect 256878 274700 256884 274712
rect 253900 274672 256884 274700
rect 253900 274660 253906 274672
rect 256878 274660 256884 274672
rect 256936 274660 256942 274712
rect 275094 274660 275100 274712
rect 275152 274700 275158 274712
rect 278314 274700 278320 274712
rect 275152 274672 278320 274700
rect 275152 274660 275158 274672
rect 278314 274660 278320 274672
rect 278372 274660 278378 274712
rect 283374 274660 283380 274712
rect 283432 274700 283438 274712
rect 289170 274700 289176 274712
rect 283432 274672 289176 274700
rect 283432 274660 283438 274672
rect 289170 274660 289176 274672
rect 289228 274660 289234 274712
rect 290458 274660 290464 274712
rect 290516 274700 290522 274712
rect 294138 274700 294144 274712
rect 290516 274672 294144 274700
rect 290516 274660 290522 274672
rect 294138 274660 294144 274672
rect 294196 274660 294202 274712
rect 295150 274660 295156 274712
rect 295208 274700 295214 274712
rect 296806 274700 296812 274712
rect 295208 274672 296812 274700
rect 295208 274660 295214 274672
rect 296806 274660 296812 274672
rect 296864 274660 296870 274712
rect 297542 274660 297548 274712
rect 297600 274700 297606 274712
rect 299474 274700 299480 274712
rect 297600 274672 299480 274700
rect 297600 274660 297606 274672
rect 299474 274660 299480 274672
rect 299532 274660 299538 274712
rect 303430 274660 303436 274712
rect 303488 274700 303494 274712
rect 303982 274700 303988 274712
rect 303488 274672 303988 274700
rect 303488 274660 303494 274672
rect 303982 274660 303988 274672
rect 304040 274660 304046 274712
rect 321186 274660 321192 274712
rect 321244 274700 321250 274712
rect 328270 274700 328276 274712
rect 321244 274672 328276 274700
rect 321244 274660 321250 274672
rect 328270 274660 328276 274672
rect 328328 274660 328334 274712
rect 114370 274592 114376 274644
rect 114428 274632 114434 274644
rect 171594 274632 171600 274644
rect 114428 274604 171600 274632
rect 114428 274592 114434 274604
rect 171594 274592 171600 274604
rect 171652 274592 171658 274644
rect 179322 274592 179328 274644
rect 179380 274632 179386 274644
rect 214558 274632 214564 274644
rect 179380 274604 214564 274632
rect 179380 274592 179386 274604
rect 214558 274592 214564 274604
rect 214616 274592 214622 274644
rect 409782 274592 409788 274644
rect 409840 274632 409846 274644
rect 453574 274632 453580 274644
rect 409840 274604 453580 274632
rect 409840 274592 409846 274604
rect 453574 274592 453580 274604
rect 453632 274592 453638 274644
rect 457438 274592 457444 274644
rect 457496 274632 457502 274644
rect 480714 274632 480720 274644
rect 457496 274604 480720 274632
rect 457496 274592 457502 274604
rect 480714 274592 480720 274604
rect 480772 274592 480778 274644
rect 486786 274592 486792 274644
rect 486844 274632 486850 274644
rect 563422 274632 563428 274644
rect 486844 274604 563428 274632
rect 486844 274592 486850 274604
rect 563422 274592 563428 274604
rect 563480 274592 563486 274644
rect 101306 274456 101312 274508
rect 101364 274496 101370 274508
rect 160922 274496 160928 274508
rect 101364 274468 160928 274496
rect 101364 274456 101370 274468
rect 160922 274456 160928 274468
rect 160980 274456 160986 274508
rect 168742 274456 168748 274508
rect 168800 274496 168806 274508
rect 208394 274496 208400 274508
rect 168800 274468 208400 274496
rect 168800 274456 168806 274468
rect 208394 274456 208400 274468
rect 208452 274456 208458 274508
rect 381538 274456 381544 274508
rect 381596 274496 381602 274508
rect 392118 274496 392124 274508
rect 381596 274468 392124 274496
rect 381596 274456 381602 274468
rect 392118 274456 392124 274468
rect 392176 274456 392182 274508
rect 413830 274456 413836 274508
rect 413888 274496 413894 274508
rect 460658 274496 460664 274508
rect 413888 274468 460664 274496
rect 413888 274456 413894 274468
rect 460658 274456 460664 274468
rect 460716 274456 460722 274508
rect 463234 274456 463240 274508
rect 463292 274496 463298 274508
rect 484302 274496 484308 274508
rect 463292 274468 484308 274496
rect 463292 274456 463298 274468
rect 484302 274456 484308 274468
rect 484360 274456 484366 274508
rect 488350 274456 488356 274508
rect 488408 274496 488414 274508
rect 567010 274496 567016 274508
rect 488408 274468 567016 274496
rect 488408 274456 488414 274468
rect 567010 274456 567016 274468
rect 567068 274456 567074 274508
rect 95418 274320 95424 274372
rect 95476 274360 95482 274372
rect 157610 274360 157616 274372
rect 95476 274332 157616 274360
rect 95476 274320 95482 274332
rect 157610 274320 157616 274332
rect 157668 274320 157674 274372
rect 159266 274320 159272 274372
rect 159324 274360 159330 274372
rect 202322 274360 202328 274372
rect 159324 274332 202328 274360
rect 159324 274320 159330 274332
rect 202322 274320 202328 274332
rect 202380 274320 202386 274372
rect 223114 274320 223120 274372
rect 223172 274360 223178 274372
rect 247218 274360 247224 274372
rect 223172 274332 247224 274360
rect 223172 274320 223178 274332
rect 247218 274320 247224 274332
rect 247276 274320 247282 274372
rect 369118 274320 369124 274372
rect 369176 274360 369182 274372
rect 387334 274360 387340 274372
rect 369176 274332 387340 274360
rect 369176 274320 369182 274332
rect 387334 274320 387340 274332
rect 387392 274320 387398 274372
rect 419074 274320 419080 274372
rect 419132 274360 419138 274372
rect 467742 274360 467748 274372
rect 419132 274332 467748 274360
rect 419132 274320 419138 274332
rect 467742 274320 467748 274332
rect 467800 274320 467806 274372
rect 506198 274320 506204 274372
rect 506256 274360 506262 274372
rect 591850 274360 591856 274372
rect 506256 274332 591856 274360
rect 506256 274320 506262 274332
rect 591850 274320 591856 274332
rect 591908 274320 591914 274372
rect 331858 274252 331864 274304
rect 331916 274292 331922 274304
rect 337746 274292 337752 274304
rect 331916 274264 337752 274292
rect 331916 274252 331922 274264
rect 337746 274252 337752 274264
rect 337804 274252 337810 274304
rect 67082 274184 67088 274236
rect 67140 274224 67146 274236
rect 130378 274224 130384 274236
rect 67140 274196 130384 274224
rect 67140 274184 67146 274196
rect 130378 274184 130384 274196
rect 130436 274184 130442 274236
rect 130838 274184 130844 274236
rect 130896 274224 130902 274236
rect 182450 274224 182456 274236
rect 130896 274196 182456 274224
rect 130896 274184 130902 274196
rect 182450 274184 182456 274196
rect 182508 274184 182514 274236
rect 193490 274184 193496 274236
rect 193548 274224 193554 274236
rect 226426 274224 226432 274236
rect 193548 274196 226432 274224
rect 193548 274184 193554 274196
rect 226426 274184 226432 274196
rect 226484 274184 226490 274236
rect 239214 274184 239220 274236
rect 239272 274224 239278 274236
rect 253934 274224 253940 274236
rect 239272 274196 253940 274224
rect 239272 274184 239278 274196
rect 253934 274184 253940 274196
rect 253992 274184 253998 274236
rect 359458 274184 359464 274236
rect 359516 274224 359522 274236
rect 380250 274224 380256 274236
rect 359516 274196 380256 274224
rect 359516 274184 359522 274196
rect 380250 274184 380256 274196
rect 380308 274184 380314 274236
rect 388990 274184 388996 274236
rect 389048 274224 389054 274236
rect 425146 274224 425152 274236
rect 389048 274196 425152 274224
rect 389048 274184 389054 274196
rect 425146 274184 425152 274196
rect 425204 274184 425210 274236
rect 425698 274184 425704 274236
rect 425756 274224 425762 274236
rect 474826 274224 474832 274236
rect 425756 274196 474832 274224
rect 425756 274184 425762 274196
rect 474826 274184 474832 274196
rect 474884 274184 474890 274236
rect 511810 274184 511816 274236
rect 511868 274224 511874 274236
rect 598934 274224 598940 274236
rect 511868 274196 598940 274224
rect 511868 274184 511874 274196
rect 598934 274184 598940 274196
rect 598992 274184 598998 274236
rect 77662 274048 77668 274100
rect 77720 274088 77726 274100
rect 144914 274088 144920 274100
rect 77720 274060 144920 274088
rect 77720 274048 77726 274060
rect 144914 274048 144920 274060
rect 144972 274048 144978 274100
rect 154482 274048 154488 274100
rect 154540 274088 154546 274100
rect 198090 274088 198096 274100
rect 154540 274060 198096 274088
rect 154540 274048 154546 274060
rect 198090 274048 198096 274060
rect 198148 274048 198154 274100
rect 210050 274048 210056 274100
rect 210108 274088 210114 274100
rect 237834 274088 237840 274100
rect 210108 274060 237840 274088
rect 210108 274048 210114 274060
rect 237834 274048 237840 274060
rect 237892 274048 237898 274100
rect 249058 274048 249064 274100
rect 249116 274088 249122 274100
rect 265250 274088 265256 274100
rect 249116 274060 265256 274088
rect 249116 274048 249122 274060
rect 265250 274048 265256 274060
rect 265308 274048 265314 274100
rect 266354 274048 266360 274100
rect 266412 274088 266418 274100
rect 273530 274088 273536 274100
rect 266412 274060 273536 274088
rect 266412 274048 266418 274060
rect 273530 274048 273536 274060
rect 273588 274048 273594 274100
rect 278590 274048 278596 274100
rect 278648 274088 278654 274100
rect 285858 274088 285864 274100
rect 278648 274060 285864 274088
rect 278648 274048 278654 274060
rect 285858 274048 285864 274060
rect 285916 274048 285922 274100
rect 337746 274048 337752 274100
rect 337804 274088 337810 274100
rect 351914 274088 351920 274100
rect 337804 274060 351920 274088
rect 337804 274048 337810 274060
rect 351914 274048 351920 274060
rect 351972 274048 351978 274100
rect 353938 274048 353944 274100
rect 353996 274088 354002 274100
rect 369578 274088 369584 274100
rect 353996 274060 369584 274088
rect 353996 274048 354002 274060
rect 369578 274048 369584 274060
rect 369636 274048 369642 274100
rect 373258 274048 373264 274100
rect 373316 274088 373322 274100
rect 400306 274088 400312 274100
rect 373316 274060 400312 274088
rect 373316 274048 373322 274060
rect 400306 274048 400312 274060
rect 400364 274048 400370 274100
rect 401502 274048 401508 274100
rect 401560 274088 401566 274100
rect 442902 274088 442908 274100
rect 401560 274060 442908 274088
rect 401560 274048 401566 274060
rect 442902 274048 442908 274060
rect 442960 274048 442966 274100
rect 451182 274048 451188 274100
rect 451240 274088 451246 274100
rect 513834 274088 513840 274100
rect 451240 274060 513840 274088
rect 451240 274048 451246 274060
rect 513834 274048 513840 274060
rect 513892 274048 513898 274100
rect 536742 274048 536748 274100
rect 536800 274088 536806 274100
rect 634354 274088 634360 274100
rect 536800 274060 634360 274088
rect 536800 274048 536806 274060
rect 634354 274048 634360 274060
rect 634412 274048 634418 274100
rect 69382 273912 69388 273964
rect 69440 273952 69446 273964
rect 139394 273952 139400 273964
rect 69440 273924 139400 273952
rect 69440 273912 69446 273924
rect 139394 273912 139400 273924
rect 139452 273912 139458 273964
rect 148594 273912 148600 273964
rect 148652 273952 148658 273964
rect 194778 273952 194784 273964
rect 148652 273924 194784 273952
rect 148652 273912 148658 273924
rect 194778 273912 194784 273924
rect 194836 273912 194842 273964
rect 208854 273912 208860 273964
rect 208912 273952 208918 273964
rect 237466 273952 237472 273964
rect 208912 273924 237472 273952
rect 208912 273912 208918 273924
rect 237466 273912 237472 273924
rect 237524 273912 237530 273964
rect 238478 273912 238484 273964
rect 238536 273952 238542 273964
rect 238536 273924 238754 273952
rect 238536 273912 238542 273924
rect 88334 273776 88340 273828
rect 88392 273816 88398 273828
rect 119338 273816 119344 273828
rect 88392 273788 119344 273816
rect 88392 273776 88398 273788
rect 119338 273776 119344 273788
rect 119396 273776 119402 273828
rect 120258 273776 120264 273828
rect 120316 273816 120322 273828
rect 175274 273816 175280 273828
rect 120316 273788 175280 273816
rect 120316 273776 120322 273788
rect 175274 273776 175280 273788
rect 175332 273776 175338 273828
rect 192386 273776 192392 273828
rect 192444 273816 192450 273828
rect 224954 273816 224960 273828
rect 192444 273788 224960 273816
rect 192444 273776 192450 273788
rect 224954 273776 224960 273788
rect 225012 273776 225018 273828
rect 238726 273816 238754 273924
rect 271506 273912 271512 273964
rect 271564 273952 271570 273964
rect 280338 273952 280344 273964
rect 271564 273924 280344 273952
rect 271564 273912 271570 273924
rect 280338 273912 280344 273924
rect 280396 273912 280402 273964
rect 322750 273912 322756 273964
rect 322808 273952 322814 273964
rect 330570 273952 330576 273964
rect 322808 273924 330576 273952
rect 322808 273912 322814 273924
rect 330570 273912 330576 273924
rect 330628 273912 330634 273964
rect 335262 273912 335268 273964
rect 335320 273952 335326 273964
rect 348326 273952 348332 273964
rect 335320 273924 348332 273952
rect 335320 273912 335326 273924
rect 348326 273912 348332 273924
rect 348384 273912 348390 273964
rect 350350 273912 350356 273964
rect 350408 273952 350414 273964
rect 368474 273952 368480 273964
rect 350408 273924 368480 273952
rect 350408 273912 350414 273924
rect 368474 273912 368480 273924
rect 368532 273912 368538 273964
rect 377766 273912 377772 273964
rect 377824 273952 377830 273964
rect 408586 273952 408592 273964
rect 377824 273924 408592 273952
rect 377824 273912 377830 273924
rect 408586 273912 408592 273924
rect 408644 273912 408650 273964
rect 422110 273912 422116 273964
rect 422168 273952 422174 273964
rect 472434 273952 472440 273964
rect 422168 273924 472440 273952
rect 422168 273912 422174 273924
rect 472434 273912 472440 273924
rect 472492 273912 472498 273964
rect 474642 273912 474648 273964
rect 474700 273952 474706 273964
rect 545758 273952 545764 273964
rect 474700 273924 545764 273952
rect 474700 273912 474706 273924
rect 545758 273912 545764 273924
rect 545816 273912 545822 273964
rect 545942 273912 545948 273964
rect 546000 273952 546006 273964
rect 639138 273952 639144 273964
rect 546000 273924 639144 273952
rect 546000 273912 546006 273924
rect 639138 273912 639144 273924
rect 639196 273912 639202 273964
rect 258074 273816 258080 273828
rect 238726 273788 258080 273816
rect 258074 273776 258080 273788
rect 258132 273776 258138 273828
rect 259362 273776 259368 273828
rect 259420 273816 259426 273828
rect 266354 273816 266360 273828
rect 259420 273788 266360 273816
rect 259420 273776 259426 273788
rect 266354 273776 266360 273788
rect 266412 273776 266418 273828
rect 396994 273776 397000 273828
rect 397052 273816 397058 273828
rect 435818 273816 435824 273828
rect 397052 273788 435824 273816
rect 397052 273776 397058 273788
rect 435818 273776 435824 273788
rect 435876 273776 435882 273828
rect 438118 273776 438124 273828
rect 438176 273816 438182 273828
rect 473630 273816 473636 273828
rect 438176 273788 473636 273816
rect 438176 273776 438182 273788
rect 473630 273776 473636 273788
rect 473688 273776 473694 273828
rect 481358 273776 481364 273828
rect 481416 273816 481422 273828
rect 556338 273816 556344 273828
rect 481416 273788 556344 273816
rect 481416 273776 481422 273788
rect 556338 273776 556344 273788
rect 556396 273776 556402 273828
rect 556798 273776 556804 273828
rect 556856 273816 556862 273828
rect 590654 273816 590660 273828
rect 556856 273788 590660 273816
rect 556856 273776 556862 273788
rect 590654 273776 590660 273788
rect 590712 273776 590718 273828
rect 119062 273640 119068 273692
rect 119120 273680 119126 273692
rect 173250 273680 173256 273692
rect 119120 273652 173256 273680
rect 119120 273640 119126 273652
rect 173250 273640 173256 273652
rect 173308 273640 173314 273692
rect 447594 273640 447600 273692
rect 447652 273680 447658 273692
rect 481910 273680 481916 273692
rect 447652 273652 481916 273680
rect 447652 273640 447658 273652
rect 481910 273640 481916 273652
rect 481968 273640 481974 273692
rect 484210 273640 484216 273692
rect 484268 273680 484274 273692
rect 559926 273680 559932 273692
rect 484268 273652 559932 273680
rect 484268 273640 484274 273652
rect 559926 273640 559932 273652
rect 559984 273640 559990 273692
rect 132034 273504 132040 273556
rect 132092 273544 132098 273556
rect 153838 273544 153844 273556
rect 132092 273516 153844 273544
rect 132092 273504 132098 273516
rect 153838 273504 153844 273516
rect 153896 273504 153902 273556
rect 440878 273504 440884 273556
rect 440936 273544 440942 273556
rect 471238 273544 471244 273556
rect 440936 273516 471244 273544
rect 440936 273504 440942 273516
rect 471238 273504 471244 273516
rect 471296 273504 471302 273556
rect 476022 273504 476028 273556
rect 476080 273544 476086 273556
rect 549254 273544 549260 273556
rect 476080 273516 549260 273544
rect 476080 273504 476086 273516
rect 549254 273504 549260 273516
rect 549312 273504 549318 273556
rect 549898 273504 549904 273556
rect 549956 273544 549962 273556
rect 583570 273544 583576 273556
rect 549956 273516 583576 273544
rect 549956 273504 549962 273516
rect 583570 273504 583576 273516
rect 583628 273504 583634 273556
rect 145282 273368 145288 273420
rect 145340 273408 145346 273420
rect 147858 273408 147864 273420
rect 145340 273380 147864 273408
rect 145340 273368 145346 273380
rect 147858 273368 147864 273380
rect 147916 273368 147922 273420
rect 478690 273368 478696 273420
rect 478748 273408 478754 273420
rect 552842 273408 552848 273420
rect 478748 273380 552848 273408
rect 478748 273368 478754 273380
rect 552842 273368 552848 273380
rect 552900 273368 552906 273420
rect 327718 273232 327724 273284
rect 327776 273272 327782 273284
rect 329466 273272 329472 273284
rect 327776 273244 329472 273272
rect 327776 273232 327782 273244
rect 329466 273232 329472 273244
rect 329524 273232 329530 273284
rect 42426 273164 42432 273216
rect 42484 273204 42490 273216
rect 43254 273204 43260 273216
rect 42484 273176 43260 273204
rect 42484 273164 42490 273176
rect 43254 273164 43260 273176
rect 43312 273164 43318 273216
rect 108390 273164 108396 273216
rect 108448 273204 108454 273216
rect 165890 273204 165896 273216
rect 108448 273176 165896 273204
rect 108448 273164 108454 273176
rect 165890 273164 165896 273176
rect 165948 273164 165954 273216
rect 186406 273164 186412 273216
rect 186464 273204 186470 273216
rect 218698 273204 218704 273216
rect 186464 273176 218704 273204
rect 186464 273164 186470 273176
rect 218698 273164 218704 273176
rect 218756 273164 218762 273216
rect 362770 273164 362776 273216
rect 362828 273204 362834 273216
rect 385862 273204 385868 273216
rect 362828 273176 385868 273204
rect 362828 273164 362834 273176
rect 385862 273164 385868 273176
rect 385920 273164 385926 273216
rect 400030 273164 400036 273216
rect 400088 273204 400094 273216
rect 439314 273204 439320 273216
rect 400088 273176 439320 273204
rect 400088 273164 400094 273176
rect 439314 273164 439320 273176
rect 439372 273164 439378 273216
rect 444006 273164 444012 273216
rect 444064 273204 444070 273216
rect 503162 273204 503168 273216
rect 444064 273176 503168 273204
rect 444064 273164 444070 273176
rect 503162 273164 503168 273176
rect 503220 273164 503226 273216
rect 504174 273164 504180 273216
rect 504232 273204 504238 273216
rect 511442 273204 511448 273216
rect 504232 273176 511448 273204
rect 504232 273164 504238 273176
rect 511442 273164 511448 273176
rect 511500 273164 511506 273216
rect 515214 273204 515220 273216
rect 511644 273176 515220 273204
rect 102502 273028 102508 273080
rect 102560 273068 102566 273080
rect 162854 273068 162860 273080
rect 102560 273040 162860 273068
rect 102560 273028 102566 273040
rect 162854 273028 162860 273040
rect 162912 273028 162918 273080
rect 172238 273028 172244 273080
rect 172296 273068 172302 273080
rect 209774 273068 209780 273080
rect 172296 273040 209780 273068
rect 172296 273028 172302 273040
rect 209774 273028 209780 273040
rect 209832 273028 209838 273080
rect 219526 273028 219532 273080
rect 219584 273068 219590 273080
rect 244550 273068 244556 273080
rect 219584 273040 244556 273068
rect 219584 273028 219590 273040
rect 244550 273028 244556 273040
rect 244608 273028 244614 273080
rect 280982 273028 280988 273080
rect 281040 273068 281046 273080
rect 286318 273068 286324 273080
rect 281040 273040 286324 273068
rect 281040 273028 281046 273040
rect 286318 273028 286324 273040
rect 286376 273028 286382 273080
rect 361206 273028 361212 273080
rect 361264 273068 361270 273080
rect 384942 273068 384948 273080
rect 361264 273040 384948 273068
rect 361264 273028 361270 273040
rect 384942 273028 384948 273040
rect 385000 273028 385006 273080
rect 385678 273028 385684 273080
rect 385736 273068 385742 273080
rect 395614 273068 395620 273080
rect 385736 273040 395620 273068
rect 385736 273028 385742 273040
rect 395614 273028 395620 273040
rect 395672 273028 395678 273080
rect 404170 273028 404176 273080
rect 404228 273068 404234 273080
rect 446490 273068 446496 273080
rect 404228 273040 446496 273068
rect 404228 273028 404234 273040
rect 446490 273028 446496 273040
rect 446548 273028 446554 273080
rect 446858 273028 446864 273080
rect 446916 273068 446922 273080
rect 507946 273068 507952 273080
rect 446916 273040 507952 273068
rect 446916 273028 446922 273040
rect 507946 273028 507952 273040
rect 508004 273028 508010 273080
rect 509694 273028 509700 273080
rect 509752 273068 509758 273080
rect 511644 273068 511672 273176
rect 515214 273164 515220 273176
rect 515272 273164 515278 273216
rect 515398 273164 515404 273216
rect 515456 273204 515462 273216
rect 519722 273204 519728 273216
rect 515456 273176 519728 273204
rect 515456 273164 515462 273176
rect 519722 273164 519728 273176
rect 519780 273164 519786 273216
rect 521470 273164 521476 273216
rect 521528 273204 521534 273216
rect 614298 273204 614304 273216
rect 521528 273176 614304 273204
rect 521528 273164 521534 273176
rect 614298 273164 614304 273176
rect 614356 273164 614362 273216
rect 509752 273040 511672 273068
rect 509752 273028 509758 273040
rect 513834 273028 513840 273080
rect 513892 273068 513898 273080
rect 518526 273068 518532 273080
rect 513892 273040 518532 273068
rect 513892 273028 513898 273040
rect 518526 273028 518532 273040
rect 518584 273028 518590 273080
rect 569402 273068 569408 273080
rect 518866 273040 569408 273068
rect 94222 272892 94228 272944
rect 94280 272932 94286 272944
rect 155954 272932 155960 272944
rect 94280 272904 155960 272932
rect 94280 272892 94286 272904
rect 155954 272892 155960 272904
rect 156012 272892 156018 272944
rect 166350 272892 166356 272944
rect 166408 272932 166414 272944
rect 207290 272932 207296 272944
rect 166408 272904 207296 272932
rect 166408 272892 166414 272904
rect 207290 272892 207296 272904
rect 207348 272892 207354 272944
rect 211246 272892 211252 272944
rect 211304 272932 211310 272944
rect 220078 272932 220084 272944
rect 211304 272904 220084 272932
rect 211304 272892 211310 272904
rect 220078 272892 220084 272904
rect 220136 272892 220142 272944
rect 220722 272892 220728 272944
rect 220780 272932 220786 272944
rect 245746 272932 245752 272944
rect 220780 272904 245752 272932
rect 220780 272892 220786 272904
rect 245746 272892 245752 272904
rect 245804 272892 245810 272944
rect 247862 272892 247868 272944
rect 247920 272932 247926 272944
rect 264238 272932 264244 272944
rect 247920 272904 264244 272932
rect 247920 272892 247926 272904
rect 264238 272892 264244 272904
rect 264296 272892 264302 272944
rect 333790 272892 333796 272944
rect 333848 272932 333854 272944
rect 345934 272932 345940 272944
rect 333848 272904 345940 272932
rect 333848 272892 333854 272904
rect 345934 272892 345940 272904
rect 345992 272892 345998 272944
rect 348418 272892 348424 272944
rect 348476 272932 348482 272944
rect 362494 272932 362500 272944
rect 348476 272904 362500 272932
rect 348476 272892 348482 272904
rect 362494 272892 362500 272904
rect 362552 272892 362558 272944
rect 365438 272892 365444 272944
rect 365496 272932 365502 272944
rect 390922 272932 390928 272944
rect 365496 272904 390928 272932
rect 365496 272892 365502 272904
rect 390922 272892 390928 272904
rect 390980 272892 390986 272944
rect 405550 272892 405556 272944
rect 405608 272932 405614 272944
rect 448790 272932 448796 272944
rect 405608 272904 448796 272932
rect 405608 272892 405614 272904
rect 448790 272892 448796 272904
rect 448848 272892 448854 272944
rect 455322 272892 455328 272944
rect 455380 272932 455386 272944
rect 461394 272932 461400 272944
rect 455380 272904 461400 272932
rect 455380 272892 455386 272904
rect 461394 272892 461400 272904
rect 461452 272892 461458 272944
rect 515030 272932 515036 272944
rect 461596 272904 515036 272932
rect 82446 272756 82452 272808
rect 82504 272796 82510 272808
rect 148410 272796 148416 272808
rect 82504 272768 148416 272796
rect 82504 272756 82510 272768
rect 148410 272756 148416 272768
rect 148468 272756 148474 272808
rect 155678 272756 155684 272808
rect 155736 272796 155742 272808
rect 200114 272796 200120 272808
rect 155736 272768 200120 272796
rect 155736 272756 155742 272768
rect 200114 272756 200120 272768
rect 200172 272756 200178 272808
rect 205358 272756 205364 272808
rect 205416 272796 205422 272808
rect 234798 272796 234804 272808
rect 205416 272768 234804 272796
rect 205416 272756 205422 272768
rect 234798 272756 234804 272768
rect 234856 272756 234862 272808
rect 245378 272756 245384 272808
rect 245436 272796 245442 272808
rect 245436 272768 258074 272796
rect 245436 272756 245442 272768
rect 72970 272620 72976 272672
rect 73028 272660 73034 272672
rect 142154 272660 142160 272672
rect 73028 272632 142160 272660
rect 73028 272620 73034 272632
rect 142154 272620 142160 272632
rect 142212 272620 142218 272672
rect 142706 272620 142712 272672
rect 142764 272660 142770 272672
rect 145558 272660 145564 272672
rect 142764 272632 145564 272660
rect 142764 272620 142770 272632
rect 145558 272620 145564 272632
rect 145616 272620 145622 272672
rect 147398 272620 147404 272672
rect 147456 272660 147462 272672
rect 193214 272660 193220 272672
rect 147456 272632 193220 272660
rect 147456 272620 147462 272632
rect 193214 272620 193220 272632
rect 193272 272620 193278 272672
rect 197078 272620 197084 272672
rect 197136 272660 197142 272672
rect 229094 272660 229100 272672
rect 197136 272632 229100 272660
rect 197136 272620 197142 272632
rect 229094 272620 229100 272632
rect 229152 272620 229158 272672
rect 233694 272620 233700 272672
rect 233752 272660 233758 272672
rect 254394 272660 254400 272672
rect 233752 272632 254400 272660
rect 233752 272620 233758 272632
rect 254394 272620 254400 272632
rect 254452 272620 254458 272672
rect 258046 272660 258074 272768
rect 262306 272756 262312 272808
rect 262364 272796 262370 272808
rect 270954 272796 270960 272808
rect 262364 272768 270960 272796
rect 262364 272756 262370 272768
rect 270954 272756 270960 272768
rect 271012 272756 271018 272808
rect 274266 272756 274272 272808
rect 274324 272796 274330 272808
rect 282914 272796 282920 272808
rect 274324 272768 282920 272796
rect 274324 272756 274330 272768
rect 282914 272756 282920 272768
rect 282972 272756 282978 272808
rect 325326 272756 325332 272808
rect 325384 272796 325390 272808
rect 332962 272796 332968 272808
rect 325384 272768 332968 272796
rect 325384 272756 325390 272768
rect 332962 272756 332968 272768
rect 333020 272756 333026 272808
rect 344646 272756 344652 272808
rect 344704 272796 344710 272808
rect 361390 272796 361396 272808
rect 344704 272768 361396 272796
rect 344704 272756 344710 272768
rect 361390 272756 361396 272768
rect 361448 272756 361454 272808
rect 362218 272756 362224 272808
rect 362276 272796 362282 272808
rect 370314 272796 370320 272808
rect 362276 272768 370320 272796
rect 362276 272756 362282 272768
rect 370314 272756 370320 272768
rect 370372 272756 370378 272808
rect 370498 272756 370504 272808
rect 370556 272796 370562 272808
rect 396810 272796 396816 272808
rect 370556 272768 396816 272796
rect 370556 272756 370562 272768
rect 396810 272756 396816 272768
rect 396868 272756 396874 272808
rect 406838 272756 406844 272808
rect 406896 272796 406902 272808
rect 449986 272796 449992 272808
rect 406896 272768 449992 272796
rect 406896 272756 406902 272768
rect 449986 272756 449992 272768
rect 450044 272756 450050 272808
rect 452286 272756 452292 272808
rect 452344 272796 452350 272808
rect 461596 272796 461624 272904
rect 515030 272892 515036 272904
rect 515088 272892 515094 272944
rect 515214 272892 515220 272944
rect 515272 272932 515278 272944
rect 518866 272932 518894 273040
rect 569402 273028 569408 273040
rect 569460 273028 569466 273080
rect 515272 272904 518894 272932
rect 515272 272892 515278 272904
rect 532510 272892 532516 272944
rect 532568 272932 532574 272944
rect 532568 272904 538904 272932
rect 532568 272892 532574 272904
rect 513834 272796 513840 272808
rect 452344 272768 461624 272796
rect 461688 272768 513840 272796
rect 452344 272756 452350 272768
rect 262674 272660 262680 272672
rect 258046 272632 262680 272660
rect 262674 272620 262680 272632
rect 262732 272620 262738 272672
rect 264422 272620 264428 272672
rect 264480 272660 264486 272672
rect 276014 272660 276020 272672
rect 264480 272632 276020 272660
rect 264480 272620 264486 272632
rect 276014 272620 276020 272632
rect 276072 272620 276078 272672
rect 324038 272620 324044 272672
rect 324096 272660 324102 272672
rect 331398 272660 331404 272672
rect 324096 272632 331404 272660
rect 324096 272620 324102 272632
rect 331398 272620 331404 272632
rect 331456 272620 331462 272672
rect 332318 272620 332324 272672
rect 332376 272660 332382 272672
rect 343634 272660 343640 272672
rect 332376 272632 343640 272660
rect 332376 272620 332382 272632
rect 343634 272620 343640 272632
rect 343692 272620 343698 272672
rect 346210 272620 346216 272672
rect 346268 272660 346274 272672
rect 363690 272660 363696 272672
rect 346268 272632 363696 272660
rect 346268 272620 346274 272632
rect 363690 272620 363696 272632
rect 363748 272620 363754 272672
rect 376110 272620 376116 272672
rect 376168 272660 376174 272672
rect 406286 272660 406292 272672
rect 376168 272632 406292 272660
rect 376168 272620 376174 272632
rect 406286 272620 406292 272632
rect 406344 272620 406350 272672
rect 412266 272620 412272 272672
rect 412324 272660 412330 272672
rect 456794 272660 456800 272672
rect 412324 272632 456800 272660
rect 412324 272620 412330 272632
rect 456794 272620 456800 272632
rect 456852 272620 456858 272672
rect 457162 272620 457168 272672
rect 457220 272660 457226 272672
rect 461026 272660 461032 272672
rect 457220 272632 461032 272660
rect 457220 272620 457226 272632
rect 461026 272620 461032 272632
rect 461084 272620 461090 272672
rect 461394 272620 461400 272672
rect 461452 272660 461458 272672
rect 461688 272660 461716 272768
rect 513834 272756 513840 272768
rect 513892 272756 513898 272808
rect 514018 272756 514024 272808
rect 514076 272796 514082 272808
rect 525610 272796 525616 272808
rect 514076 272768 525616 272796
rect 514076 272756 514082 272768
rect 525610 272756 525616 272768
rect 525668 272756 525674 272808
rect 529842 272756 529848 272808
rect 529900 272796 529906 272808
rect 532878 272796 532884 272808
rect 529900 272768 532884 272796
rect 529900 272756 529906 272768
rect 532878 272756 532884 272768
rect 532936 272756 532942 272808
rect 533706 272756 533712 272808
rect 533764 272796 533770 272808
rect 538674 272796 538680 272808
rect 533764 272768 538680 272796
rect 533764 272756 533770 272768
rect 538674 272756 538680 272768
rect 538732 272756 538738 272808
rect 538876 272796 538904 272904
rect 539042 272892 539048 272944
rect 539100 272932 539106 272944
rect 624970 272932 624976 272944
rect 539100 272904 624976 272932
rect 539100 272892 539106 272904
rect 624970 272892 624976 272904
rect 625028 272892 625034 272944
rect 632054 272932 632060 272944
rect 628668 272904 632060 272932
rect 628466 272796 628472 272808
rect 538876 272768 628472 272796
rect 628466 272756 628472 272768
rect 628524 272756 628530 272808
rect 461452 272632 461716 272660
rect 461452 272620 461458 272632
rect 461854 272620 461860 272672
rect 461912 272660 461918 272672
rect 461912 272632 463924 272660
rect 461912 272620 461918 272632
rect 463896 272592 463924 272632
rect 466408 272620 466414 272672
rect 466466 272660 466472 272672
rect 522114 272660 522120 272672
rect 466466 272632 522120 272660
rect 466466 272620 466472 272632
rect 522114 272620 522120 272632
rect 522172 272620 522178 272672
rect 526806 272620 526812 272672
rect 526864 272660 526870 272672
rect 621382 272660 621388 272672
rect 526864 272632 621388 272660
rect 526864 272620 526870 272632
rect 621382 272620 621388 272632
rect 621440 272620 621446 272672
rect 463896 272564 466316 272592
rect 65886 272484 65892 272536
rect 65944 272524 65950 272536
rect 136818 272524 136824 272536
rect 65944 272496 136824 272524
rect 65944 272484 65950 272496
rect 136818 272484 136824 272496
rect 136876 272484 136882 272536
rect 137922 272484 137928 272536
rect 137980 272524 137986 272536
rect 137980 272496 180794 272524
rect 137980 272484 137986 272496
rect 116670 272348 116676 272400
rect 116728 272388 116734 272400
rect 172514 272388 172520 272400
rect 116728 272360 172520 272388
rect 116728 272348 116734 272360
rect 172514 272348 172520 272360
rect 172572 272348 172578 272400
rect 180766 272388 180794 272496
rect 181714 272484 181720 272536
rect 181772 272524 181778 272536
rect 186958 272524 186964 272536
rect 181772 272496 186964 272524
rect 181772 272484 181778 272496
rect 186958 272484 186964 272496
rect 187016 272484 187022 272536
rect 195882 272484 195888 272536
rect 195940 272524 195946 272536
rect 227898 272524 227904 272536
rect 195940 272496 227904 272524
rect 195940 272484 195946 272496
rect 227898 272484 227904 272496
rect 227956 272484 227962 272536
rect 228082 272484 228088 272536
rect 228140 272524 228146 272536
rect 249058 272524 249064 272536
rect 228140 272496 249064 272524
rect 228140 272484 228146 272496
rect 249058 272484 249064 272496
rect 249116 272484 249122 272536
rect 254946 272484 254952 272536
rect 255004 272524 255010 272536
rect 269298 272524 269304 272536
rect 255004 272496 269304 272524
rect 255004 272484 255010 272496
rect 269298 272484 269304 272496
rect 269356 272484 269362 272536
rect 270310 272484 270316 272536
rect 270368 272524 270374 272536
rect 280522 272524 280528 272536
rect 270368 272496 280528 272524
rect 270368 272484 270374 272496
rect 280522 272484 280528 272496
rect 280580 272484 280586 272536
rect 329742 272484 329748 272536
rect 329800 272524 329806 272536
rect 338850 272524 338856 272536
rect 329800 272496 338856 272524
rect 329800 272484 329806 272496
rect 338850 272484 338856 272496
rect 338908 272484 338914 272536
rect 339218 272484 339224 272536
rect 339276 272524 339282 272536
rect 354214 272524 354220 272536
rect 339276 272496 354220 272524
rect 339276 272484 339282 272496
rect 354214 272484 354220 272496
rect 354272 272484 354278 272536
rect 354490 272484 354496 272536
rect 354548 272524 354554 272536
rect 375558 272524 375564 272536
rect 354548 272496 375564 272524
rect 354548 272484 354554 272496
rect 375558 272484 375564 272496
rect 375616 272484 375622 272536
rect 379422 272484 379428 272536
rect 379480 272524 379486 272536
rect 410978 272524 410984 272536
rect 379480 272496 410984 272524
rect 379480 272484 379486 272496
rect 410978 272484 410984 272496
rect 411036 272484 411042 272536
rect 416590 272484 416596 272536
rect 416648 272524 416654 272536
rect 463694 272524 463700 272536
rect 416648 272496 463700 272524
rect 416648 272484 416654 272496
rect 463694 272484 463700 272496
rect 463752 272484 463758 272536
rect 466288 272524 466316 272564
rect 470548 272524 470554 272536
rect 466288 272496 470554 272524
rect 470548 272484 470554 272496
rect 470606 272484 470612 272536
rect 470686 272484 470692 272536
rect 470744 272524 470750 272536
rect 532694 272524 532700 272536
rect 470744 272496 532700 272524
rect 470744 272484 470750 272496
rect 532694 272484 532700 272496
rect 532752 272484 532758 272536
rect 532878 272484 532884 272536
rect 532936 272524 532942 272536
rect 538490 272524 538496 272536
rect 532936 272496 538496 272524
rect 532936 272484 532942 272496
rect 538490 272484 538496 272496
rect 538548 272484 538554 272536
rect 538674 272484 538680 272536
rect 538732 272524 538738 272536
rect 628668 272524 628696 272904
rect 632054 272892 632060 272904
rect 632112 272892 632118 272944
rect 635550 272796 635556 272808
rect 538732 272496 628696 272524
rect 629956 272768 635556 272796
rect 538732 272484 538738 272496
rect 187694 272388 187700 272400
rect 180766 272360 187700 272388
rect 187694 272348 187700 272360
rect 187752 272348 187758 272400
rect 194962 272348 194968 272400
rect 195020 272388 195026 272400
rect 227162 272388 227168 272400
rect 195020 272360 227168 272388
rect 195020 272348 195026 272360
rect 227162 272348 227168 272360
rect 227220 272348 227226 272400
rect 318702 272348 318708 272400
rect 318760 272388 318766 272400
rect 324682 272388 324688 272400
rect 318760 272360 324688 272388
rect 318760 272348 318766 272360
rect 324682 272348 324688 272360
rect 324740 272348 324746 272400
rect 395982 272348 395988 272400
rect 396040 272388 396046 272400
rect 434622 272388 434628 272400
rect 396040 272360 434628 272388
rect 396040 272348 396046 272360
rect 434622 272348 434628 272360
rect 434680 272348 434686 272400
rect 449710 272348 449716 272400
rect 449768 272388 449774 272400
rect 504174 272388 504180 272400
rect 449768 272360 504180 272388
rect 449768 272348 449774 272360
rect 504174 272348 504180 272360
rect 504232 272348 504238 272400
rect 504358 272348 504364 272400
rect 504416 272388 504422 272400
rect 514018 272388 514024 272400
rect 504416 272360 514024 272388
rect 504416 272348 504422 272360
rect 514018 272348 514024 272360
rect 514076 272348 514082 272400
rect 517422 272348 517428 272400
rect 517480 272388 517486 272400
rect 600958 272388 600964 272400
rect 517480 272360 600964 272388
rect 517480 272348 517486 272360
rect 600958 272348 600964 272360
rect 601016 272348 601022 272400
rect 601142 272348 601148 272400
rect 601200 272388 601206 272400
rect 629956 272388 629984 272768
rect 635550 272756 635556 272768
rect 635608 272756 635614 272808
rect 634078 272620 634084 272672
rect 634136 272660 634142 272672
rect 640334 272660 640340 272672
rect 634136 272632 640340 272660
rect 634136 272620 634142 272632
rect 640334 272620 640340 272632
rect 640392 272620 640398 272672
rect 601200 272360 629984 272388
rect 601200 272348 601206 272360
rect 127342 272212 127348 272264
rect 127400 272252 127406 272264
rect 179874 272252 179880 272264
rect 127400 272224 179880 272252
rect 127400 272212 127406 272224
rect 179874 272212 179880 272224
rect 179932 272212 179938 272264
rect 189074 272212 189080 272264
rect 189132 272252 189138 272264
rect 196434 272252 196440 272264
rect 189132 272224 196440 272252
rect 189132 272212 189138 272224
rect 196434 272212 196440 272224
rect 196492 272212 196498 272264
rect 391842 272212 391848 272264
rect 391900 272252 391906 272264
rect 428734 272252 428740 272264
rect 391900 272224 428740 272252
rect 391900 272212 391906 272224
rect 428734 272212 428740 272224
rect 428792 272212 428798 272264
rect 450538 272212 450544 272264
rect 450596 272252 450602 272264
rect 510246 272252 510252 272264
rect 450596 272224 510252 272252
rect 450596 272212 450602 272224
rect 510246 272212 510252 272224
rect 510304 272212 510310 272264
rect 520090 272212 520096 272264
rect 520148 272252 520154 272264
rect 610710 272252 610716 272264
rect 520148 272224 610716 272252
rect 520148 272212 520154 272224
rect 610710 272212 610716 272224
rect 610768 272212 610774 272264
rect 145098 272076 145104 272128
rect 145156 272116 145162 272128
rect 192386 272116 192392 272128
rect 145156 272088 192392 272116
rect 145156 272076 145162 272088
rect 192386 272076 192392 272088
rect 192444 272076 192450 272128
rect 384942 272076 384948 272128
rect 385000 272116 385006 272128
rect 418062 272116 418068 272128
rect 385000 272088 418068 272116
rect 385000 272076 385006 272088
rect 418062 272076 418068 272088
rect 418120 272076 418126 272128
rect 428458 272076 428464 272128
rect 428516 272116 428522 272128
rect 470548 272116 470554 272128
rect 428516 272088 470554 272116
rect 428516 272076 428522 272088
rect 470548 272076 470554 272088
rect 470606 272076 470612 272128
rect 470778 272076 470784 272128
rect 470836 272116 470842 272128
rect 470836 272088 480392 272116
rect 470836 272076 470842 272088
rect 124950 271940 124956 271992
rect 125008 271980 125014 271992
rect 151078 271980 151084 271992
rect 125008 271952 151084 271980
rect 125008 271940 125014 271952
rect 151078 271940 151084 271952
rect 151136 271940 151142 271992
rect 431678 271940 431684 271992
rect 431736 271980 431742 271992
rect 480162 271980 480168 271992
rect 431736 271952 480168 271980
rect 431736 271940 431742 271952
rect 480162 271940 480168 271952
rect 480220 271940 480226 271992
rect 480364 271980 480392 272088
rect 480530 272076 480536 272128
rect 480588 272116 480594 272128
rect 547506 272116 547512 272128
rect 480588 272088 547512 272116
rect 480588 272076 480594 272088
rect 547506 272076 547512 272088
rect 547564 272076 547570 272128
rect 547690 272076 547696 272128
rect 547748 272116 547754 272128
rect 547748 272088 586514 272116
rect 547748 272076 547754 272088
rect 504358 271980 504364 271992
rect 480364 271952 504364 271980
rect 504358 271940 504364 271952
rect 504416 271940 504422 271992
rect 504542 271940 504548 271992
rect 504600 271980 504606 271992
rect 562318 271980 562324 271992
rect 504600 271952 562324 271980
rect 504600 271940 504606 271952
rect 562318 271940 562324 271952
rect 562376 271940 562382 271992
rect 586486 271980 586514 272088
rect 600958 272076 600964 272128
rect 601016 272116 601022 272128
rect 607214 272116 607220 272128
rect 601016 272088 607220 272116
rect 601016 272076 601022 272088
rect 607214 272076 607220 272088
rect 607272 272076 607278 272128
rect 601142 271980 601148 271992
rect 586486 271952 601148 271980
rect 601142 271940 601148 271952
rect 601200 271940 601206 271992
rect 105998 271804 106004 271856
rect 106056 271844 106062 271856
rect 164970 271844 164976 271856
rect 106056 271816 164976 271844
rect 106056 271804 106062 271816
rect 164970 271804 164976 271816
rect 165028 271804 165034 271856
rect 174262 271804 174268 271856
rect 174320 271844 174326 271856
rect 189258 271844 189264 271856
rect 174320 271816 189264 271844
rect 174320 271804 174326 271816
rect 189258 271804 189264 271816
rect 189316 271804 189322 271856
rect 202966 271804 202972 271856
rect 203024 271844 203030 271856
rect 233234 271844 233240 271856
rect 203024 271816 233240 271844
rect 203024 271804 203030 271816
rect 233234 271804 233240 271816
rect 233292 271804 233298 271856
rect 274634 271804 274640 271856
rect 274692 271844 274698 271856
rect 279234 271844 279240 271856
rect 274692 271816 279240 271844
rect 274692 271804 274698 271816
rect 279234 271804 279240 271816
rect 279292 271804 279298 271856
rect 355318 271804 355324 271856
rect 355376 271844 355382 271856
rect 356606 271844 356612 271856
rect 355376 271816 356612 271844
rect 355376 271804 355382 271816
rect 356606 271804 356612 271816
rect 356664 271804 356670 271856
rect 375282 271804 375288 271856
rect 375340 271844 375346 271856
rect 403894 271844 403900 271856
rect 375340 271816 403900 271844
rect 375340 271804 375346 271816
rect 403894 271804 403900 271816
rect 403952 271804 403958 271856
rect 433150 271804 433156 271856
rect 433208 271844 433214 271856
rect 480162 271844 480168 271856
rect 433208 271816 480168 271844
rect 433208 271804 433214 271816
rect 480162 271804 480168 271816
rect 480220 271804 480226 271856
rect 480438 271804 480444 271856
rect 480496 271844 480502 271856
rect 484854 271844 484860 271856
rect 480496 271816 484860 271844
rect 480496 271804 480502 271816
rect 484854 271804 484860 271816
rect 484912 271804 484918 271856
rect 501414 271844 501420 271856
rect 489886 271816 501420 271844
rect 97810 271668 97816 271720
rect 97868 271708 97874 271720
rect 158806 271708 158812 271720
rect 97868 271680 158812 271708
rect 97868 271668 97874 271680
rect 158806 271668 158812 271680
rect 158864 271668 158870 271720
rect 169846 271668 169852 271720
rect 169904 271708 169910 271720
rect 209958 271708 209964 271720
rect 169904 271680 209964 271708
rect 169904 271668 169910 271680
rect 209958 271668 209964 271680
rect 210016 271668 210022 271720
rect 225414 271668 225420 271720
rect 225472 271708 225478 271720
rect 228358 271708 228364 271720
rect 225472 271680 228364 271708
rect 225472 271668 225478 271680
rect 228358 271668 228364 271680
rect 228416 271668 228422 271720
rect 351178 271668 351184 271720
rect 351236 271708 351242 271720
rect 366082 271708 366088 271720
rect 351236 271680 366088 271708
rect 351236 271668 351242 271680
rect 366082 271668 366088 271680
rect 366140 271668 366146 271720
rect 381998 271668 382004 271720
rect 382056 271708 382062 271720
rect 414566 271708 414572 271720
rect 382056 271680 414572 271708
rect 382056 271668 382062 271680
rect 414566 271668 414572 271680
rect 414624 271668 414630 271720
rect 430390 271668 430396 271720
rect 430448 271708 430454 271720
rect 483566 271708 483572 271720
rect 430448 271680 483572 271708
rect 430448 271668 430454 271680
rect 483566 271668 483572 271680
rect 483624 271668 483630 271720
rect 485038 271668 485044 271720
rect 485096 271708 485102 271720
rect 489886 271708 489914 271816
rect 501414 271804 501420 271816
rect 501472 271804 501478 271856
rect 578510 271844 578516 271856
rect 504376 271816 578516 271844
rect 485096 271680 489914 271708
rect 485096 271668 485102 271680
rect 496538 271668 496544 271720
rect 496596 271708 496602 271720
rect 504376 271708 504404 271816
rect 578510 271804 578516 271816
rect 578568 271804 578574 271856
rect 578878 271804 578884 271856
rect 578936 271844 578942 271856
rect 604822 271844 604828 271856
rect 578936 271816 604828 271844
rect 578936 271804 578942 271816
rect 604822 271804 604828 271816
rect 604880 271804 604886 271856
rect 496596 271680 504404 271708
rect 496596 271668 496602 271680
rect 504542 271668 504548 271720
rect 504600 271708 504606 271720
rect 585962 271708 585968 271720
rect 504600 271680 585968 271708
rect 504600 271668 504606 271680
rect 585962 271668 585968 271680
rect 586020 271668 586026 271720
rect 87138 271532 87144 271584
rect 87196 271572 87202 271584
rect 151998 271572 152004 271584
rect 87196 271544 152004 271572
rect 87196 271532 87202 271544
rect 151998 271532 152004 271544
rect 152056 271532 152062 271584
rect 165154 271532 165160 271584
rect 165212 271572 165218 271584
rect 205634 271572 205640 271584
rect 165212 271544 205640 271572
rect 165212 271532 165218 271544
rect 205634 271532 205640 271544
rect 205692 271532 205698 271584
rect 215938 271532 215944 271584
rect 215996 271572 216002 271584
rect 242066 271572 242072 271584
rect 215996 271544 242072 271572
rect 215996 271532 216002 271544
rect 242066 271532 242072 271544
rect 242124 271532 242130 271584
rect 337930 271532 337936 271584
rect 337988 271572 337994 271584
rect 350718 271572 350724 271584
rect 337988 271544 350724 271572
rect 337988 271532 337994 271544
rect 350718 271532 350724 271544
rect 350776 271532 350782 271584
rect 360838 271532 360844 271584
rect 360896 271572 360902 271584
rect 377582 271572 377588 271584
rect 360896 271544 377588 271572
rect 360896 271532 360902 271544
rect 377582 271532 377588 271544
rect 377640 271532 377646 271584
rect 387702 271532 387708 271584
rect 387760 271572 387766 271584
rect 421650 271572 421656 271584
rect 387760 271544 421656 271572
rect 387760 271532 387766 271544
rect 421650 271532 421656 271544
rect 421708 271532 421714 271584
rect 437198 271532 437204 271584
rect 437256 271572 437262 271584
rect 493686 271572 493692 271584
rect 437256 271544 493692 271572
rect 437256 271532 437262 271544
rect 493686 271532 493692 271544
rect 493744 271532 493750 271584
rect 499298 271532 499304 271584
rect 499356 271572 499362 271584
rect 582374 271572 582380 271584
rect 499356 271544 582380 271572
rect 499356 271532 499362 271544
rect 582374 271532 582380 271544
rect 582432 271532 582438 271584
rect 583018 271532 583024 271584
rect 583076 271572 583082 271584
rect 611630 271572 611636 271584
rect 583076 271544 611636 271572
rect 583076 271532 583082 271544
rect 611630 271532 611636 271544
rect 611688 271532 611694 271584
rect 611998 271532 612004 271584
rect 612056 271572 612062 271584
rect 618990 271572 618996 271584
rect 612056 271544 618996 271572
rect 612056 271532 612062 271544
rect 618990 271532 618996 271544
rect 619048 271532 619054 271584
rect 75362 271396 75368 271448
rect 75420 271436 75426 271448
rect 142706 271436 142712 271448
rect 75420 271408 142712 271436
rect 75420 271396 75426 271408
rect 142706 271396 142712 271408
rect 142764 271396 142770 271448
rect 162670 271396 162676 271448
rect 162728 271436 162734 271448
rect 204714 271436 204720 271448
rect 162728 271408 204720 271436
rect 162728 271396 162734 271408
rect 204714 271396 204720 271408
rect 204772 271396 204778 271448
rect 213638 271396 213644 271448
rect 213696 271436 213702 271448
rect 240410 271436 240416 271448
rect 213696 271408 240416 271436
rect 213696 271396 213702 271408
rect 240410 271396 240416 271408
rect 240468 271396 240474 271448
rect 240778 271396 240784 271448
rect 240836 271436 240842 271448
rect 259638 271436 259644 271448
rect 240836 271408 259644 271436
rect 240836 271396 240842 271408
rect 259638 271396 259644 271408
rect 259696 271396 259702 271448
rect 260098 271396 260104 271448
rect 260156 271436 260162 271448
rect 272610 271436 272616 271448
rect 260156 271408 272616 271436
rect 260156 271396 260162 271408
rect 272610 271396 272616 271408
rect 272668 271396 272674 271448
rect 325510 271396 325516 271448
rect 325568 271436 325574 271448
rect 334158 271436 334164 271448
rect 325568 271408 334164 271436
rect 325568 271396 325574 271408
rect 334158 271396 334164 271408
rect 334216 271396 334222 271448
rect 347682 271396 347688 271448
rect 347740 271436 347746 271448
rect 364886 271436 364892 271448
rect 347740 271408 364892 271436
rect 347740 271396 347746 271408
rect 364886 271396 364892 271408
rect 364944 271396 364950 271448
rect 366358 271396 366364 271448
rect 366416 271436 366422 271448
rect 383838 271436 383844 271448
rect 366416 271408 383844 271436
rect 366416 271396 366422 271408
rect 383838 271396 383844 271408
rect 383896 271396 383902 271448
rect 384758 271396 384764 271448
rect 384816 271436 384822 271448
rect 419258 271436 419264 271448
rect 384816 271408 419264 271436
rect 384816 271396 384822 271408
rect 419258 271396 419264 271408
rect 419316 271396 419322 271448
rect 420178 271396 420184 271448
rect 420236 271436 420242 271448
rect 431126 271436 431132 271448
rect 420236 271408 431132 271436
rect 420236 271396 420242 271408
rect 431126 271396 431132 271408
rect 431184 271396 431190 271448
rect 439958 271396 439964 271448
rect 440016 271436 440022 271448
rect 497274 271436 497280 271448
rect 440016 271408 497280 271436
rect 440016 271396 440022 271408
rect 497274 271396 497280 271408
rect 497332 271396 497338 271448
rect 501966 271396 501972 271448
rect 502024 271436 502030 271448
rect 504542 271436 504548 271448
rect 502024 271408 504548 271436
rect 502024 271396 502030 271408
rect 504542 271396 504548 271408
rect 504600 271396 504606 271448
rect 505002 271396 505008 271448
rect 505060 271436 505066 271448
rect 589458 271436 589464 271448
rect 505060 271408 589464 271436
rect 505060 271396 505066 271408
rect 589458 271396 589464 271408
rect 589516 271396 589522 271448
rect 589918 271396 589924 271448
rect 589976 271436 589982 271448
rect 633250 271436 633256 271448
rect 589976 271408 633256 271436
rect 589976 271396 589982 271408
rect 633250 271396 633256 271408
rect 633308 271396 633314 271448
rect 76834 271260 76840 271312
rect 76892 271300 76898 271312
rect 143534 271300 143540 271312
rect 76892 271272 143540 271300
rect 76892 271260 76898 271272
rect 143534 271260 143540 271272
rect 143592 271260 143598 271312
rect 152182 271260 152188 271312
rect 152240 271300 152246 271312
rect 197354 271300 197360 271312
rect 152240 271272 197360 271300
rect 152240 271260 152246 271272
rect 197354 271260 197360 271272
rect 197412 271260 197418 271312
rect 198274 271260 198280 271312
rect 198332 271300 198338 271312
rect 229554 271300 229560 271312
rect 198332 271272 229560 271300
rect 198332 271260 198338 271272
rect 229554 271260 229560 271272
rect 229612 271260 229618 271312
rect 235258 271260 235264 271312
rect 235316 271300 235322 271312
rect 255314 271300 255320 271312
rect 235316 271272 255320 271300
rect 235316 271260 235322 271272
rect 255314 271260 255320 271272
rect 255372 271260 255378 271312
rect 256694 271260 256700 271312
rect 256752 271300 256758 271312
rect 261018 271300 261024 271312
rect 256752 271272 261024 271300
rect 256752 271260 256758 271272
rect 261018 271260 261024 271272
rect 261076 271260 261082 271312
rect 262030 271260 262036 271312
rect 262088 271300 262094 271312
rect 274634 271300 274640 271312
rect 262088 271272 274640 271300
rect 262088 271260 262094 271272
rect 274634 271260 274640 271272
rect 274692 271260 274698 271312
rect 329558 271260 329564 271312
rect 329616 271300 329622 271312
rect 340046 271300 340052 271312
rect 329616 271272 340052 271300
rect 329616 271260 329622 271272
rect 340046 271260 340052 271272
rect 340104 271260 340110 271312
rect 340598 271260 340604 271312
rect 340656 271300 340662 271312
rect 355134 271300 355140 271312
rect 340656 271272 355140 271300
rect 340656 271260 340662 271272
rect 355134 271260 355140 271272
rect 355192 271260 355198 271312
rect 357158 271260 357164 271312
rect 357216 271300 357222 271312
rect 379054 271300 379060 271312
rect 357216 271272 379060 271300
rect 357216 271260 357222 271272
rect 379054 271260 379060 271272
rect 379112 271260 379118 271312
rect 390278 271260 390284 271312
rect 390336 271300 390342 271312
rect 426342 271300 426348 271312
rect 390336 271272 426348 271300
rect 390336 271260 390342 271272
rect 426342 271260 426348 271272
rect 426400 271260 426406 271312
rect 432230 271300 432236 271312
rect 427096 271272 432236 271300
rect 68186 271124 68192 271176
rect 68244 271164 68250 271176
rect 138474 271164 138480 271176
rect 68244 271136 138480 271164
rect 68244 271124 68250 271136
rect 138474 271124 138480 271136
rect 138532 271124 138538 271176
rect 141510 271124 141516 271176
rect 141568 271164 141574 271176
rect 189074 271164 189080 271176
rect 141568 271136 189080 271164
rect 141568 271124 141574 271136
rect 189074 271124 189080 271136
rect 189132 271124 189138 271176
rect 191190 271124 191196 271176
rect 191248 271164 191254 271176
rect 225138 271164 225144 271176
rect 191248 271136 225144 271164
rect 191248 271124 191254 271136
rect 225138 271124 225144 271136
rect 225196 271124 225202 271176
rect 230198 271124 230204 271176
rect 230256 271164 230262 271176
rect 252002 271164 252008 271176
rect 230256 271136 252008 271164
rect 230256 271124 230262 271136
rect 252002 271124 252008 271136
rect 252060 271124 252066 271176
rect 268010 271124 268016 271176
rect 268068 271164 268074 271176
rect 278774 271164 278780 271176
rect 268068 271136 278780 271164
rect 268068 271124 268074 271136
rect 278774 271124 278780 271136
rect 278832 271124 278838 271176
rect 279786 271124 279792 271176
rect 279844 271164 279850 271176
rect 287054 271164 287060 271176
rect 279844 271136 287060 271164
rect 279844 271124 279850 271136
rect 287054 271124 287060 271136
rect 287112 271124 287118 271176
rect 331122 271124 331128 271176
rect 331180 271164 331186 271176
rect 342438 271164 342444 271176
rect 331180 271136 342444 271164
rect 331180 271124 331186 271136
rect 342438 271124 342444 271136
rect 342496 271124 342502 271176
rect 343542 271124 343548 271176
rect 343600 271164 343606 271176
rect 360194 271164 360200 271176
rect 343600 271136 360200 271164
rect 343600 271124 343606 271136
rect 360194 271124 360200 271136
rect 360252 271124 360258 271176
rect 364150 271124 364156 271176
rect 364208 271164 364214 271176
rect 389726 271164 389732 271176
rect 364208 271136 389732 271164
rect 364208 271124 364214 271136
rect 389726 271124 389732 271136
rect 389784 271124 389790 271176
rect 394326 271124 394332 271176
rect 394384 271164 394390 271176
rect 427096 271164 427124 271272
rect 432230 271260 432236 271272
rect 432288 271260 432294 271312
rect 442902 271260 442908 271312
rect 442960 271300 442966 271312
rect 500862 271300 500868 271312
rect 442960 271272 500868 271300
rect 442960 271260 442966 271272
rect 500862 271260 500868 271272
rect 500920 271260 500926 271312
rect 507670 271260 507676 271312
rect 507728 271300 507734 271312
rect 593046 271300 593052 271312
rect 507728 271272 593052 271300
rect 507728 271260 507734 271272
rect 593046 271260 593052 271272
rect 593104 271260 593110 271312
rect 598198 271260 598204 271312
rect 598256 271300 598262 271312
rect 645026 271300 645032 271312
rect 598256 271272 645032 271300
rect 598256 271260 598262 271272
rect 645026 271260 645032 271272
rect 645084 271260 645090 271312
rect 437934 271164 437940 271176
rect 394384 271136 427124 271164
rect 427188 271136 437940 271164
rect 394384 271124 394390 271136
rect 113450 270988 113456 271040
rect 113508 271028 113514 271040
rect 169938 271028 169944 271040
rect 113508 271000 169944 271028
rect 113508 270988 113514 271000
rect 169938 270988 169944 271000
rect 169996 270988 170002 271040
rect 187418 270988 187424 271040
rect 187476 271028 187482 271040
rect 215938 271028 215944 271040
rect 187476 271000 215944 271028
rect 187476 270988 187482 271000
rect 215938 270988 215944 271000
rect 215996 270988 216002 271040
rect 251450 270988 251456 271040
rect 251508 271028 251514 271040
rect 266906 271028 266912 271040
rect 251508 271000 266912 271028
rect 251508 270988 251514 271000
rect 266906 270988 266912 271000
rect 266964 270988 266970 271040
rect 417418 270988 417424 271040
rect 417476 271028 417482 271040
rect 427188 271028 427216 271136
rect 437934 271124 437940 271136
rect 437992 271124 437998 271176
rect 441338 271124 441344 271176
rect 441396 271164 441402 271176
rect 445018 271164 445024 271176
rect 441396 271136 445024 271164
rect 441396 271124 441402 271136
rect 445018 271124 445024 271136
rect 445076 271124 445082 271176
rect 445662 271124 445668 271176
rect 445720 271164 445726 271176
rect 503990 271164 503996 271176
rect 445720 271136 503996 271164
rect 445720 271124 445726 271136
rect 503990 271124 503996 271136
rect 504048 271124 504054 271176
rect 524046 271124 524052 271176
rect 524104 271164 524110 271176
rect 617334 271164 617340 271176
rect 524104 271136 617340 271164
rect 524104 271124 524110 271136
rect 617334 271124 617340 271136
rect 617392 271124 617398 271176
rect 617518 271124 617524 271176
rect 617576 271164 617582 271176
rect 626074 271164 626080 271176
rect 617576 271136 626080 271164
rect 617576 271124 617582 271136
rect 626074 271124 626080 271136
rect 626132 271124 626138 271176
rect 417476 271000 427216 271028
rect 417476 270988 417482 271000
rect 427446 270988 427452 271040
rect 427504 271028 427510 271040
rect 479150 271028 479156 271040
rect 427504 271000 479156 271028
rect 427504 270988 427510 271000
rect 479150 270988 479156 271000
rect 479208 270988 479214 271040
rect 480254 270988 480260 271040
rect 480312 271028 480318 271040
rect 486602 271028 486608 271040
rect 480312 271000 486608 271028
rect 480312 270988 480318 271000
rect 486602 270988 486608 271000
rect 486660 270988 486666 271040
rect 495066 270988 495072 271040
rect 495124 271028 495130 271040
rect 575290 271028 575296 271040
rect 495124 271000 575296 271028
rect 495124 270988 495130 271000
rect 575290 270988 575296 271000
rect 575348 270988 575354 271040
rect 123754 270852 123760 270904
rect 123812 270892 123818 270904
rect 177482 270892 177488 270904
rect 123812 270864 177488 270892
rect 123812 270852 123818 270864
rect 177482 270852 177488 270864
rect 177540 270852 177546 270904
rect 407758 270852 407764 270904
rect 407816 270892 407822 270904
rect 440510 270892 440516 270904
rect 407816 270864 440516 270892
rect 407816 270852 407822 270864
rect 440510 270852 440516 270864
rect 440568 270852 440574 270904
rect 449158 270852 449164 270904
rect 449216 270892 449222 270904
rect 490190 270892 490196 270904
rect 449216 270864 490196 270892
rect 449216 270852 449222 270864
rect 490190 270852 490196 270864
rect 490248 270852 490254 270904
rect 492582 270852 492588 270904
rect 492640 270892 492646 270904
rect 571702 270892 571708 270904
rect 492640 270864 571708 270892
rect 492640 270852 492646 270864
rect 571702 270852 571708 270864
rect 571760 270852 571766 270904
rect 134426 270716 134432 270768
rect 134484 270756 134490 270768
rect 185118 270756 185124 270768
rect 134484 270728 185124 270756
rect 134484 270716 134490 270728
rect 185118 270716 185124 270728
rect 185176 270716 185182 270768
rect 321370 270716 321376 270768
rect 321428 270756 321434 270768
rect 327074 270756 327080 270768
rect 321428 270728 327080 270756
rect 321428 270716 321434 270728
rect 327074 270716 327080 270728
rect 327132 270716 327138 270768
rect 414658 270716 414664 270768
rect 414716 270756 414722 270768
rect 450814 270756 450820 270768
rect 414716 270728 450820 270756
rect 414716 270716 414722 270728
rect 450814 270716 450820 270728
rect 450872 270716 450878 270768
rect 486970 270716 486976 270768
rect 487028 270756 487034 270768
rect 564618 270756 564624 270768
rect 487028 270728 564624 270756
rect 487028 270716 487034 270728
rect 564618 270716 564624 270728
rect 564676 270716 564682 270768
rect 567838 270716 567844 270768
rect 567896 270756 567902 270768
rect 597738 270756 597744 270768
rect 567896 270728 597744 270756
rect 567896 270716 567902 270728
rect 597738 270716 597744 270728
rect 597796 270716 597802 270768
rect 121454 270580 121460 270632
rect 121512 270620 121518 270632
rect 168098 270620 168104 270632
rect 121512 270592 168104 270620
rect 121512 270580 121518 270592
rect 168098 270580 168104 270592
rect 168156 270580 168162 270632
rect 403618 270580 403624 270632
rect 403676 270620 403682 270632
rect 433426 270620 433432 270632
rect 403676 270592 433432 270620
rect 403676 270580 403682 270592
rect 433426 270580 433432 270592
rect 433484 270580 433490 270632
rect 453298 270580 453304 270632
rect 453356 270620 453362 270632
rect 487798 270620 487804 270632
rect 453356 270592 487804 270620
rect 453356 270580 453362 270592
rect 487798 270580 487804 270592
rect 487856 270580 487862 270632
rect 489638 270580 489644 270632
rect 489696 270620 489702 270632
rect 568206 270620 568212 270632
rect 489696 270592 568212 270620
rect 489696 270580 489702 270592
rect 568206 270580 568212 270592
rect 568264 270580 568270 270632
rect 84102 270444 84108 270496
rect 84160 270484 84166 270496
rect 137462 270484 137468 270496
rect 84160 270456 137468 270484
rect 84160 270444 84166 270456
rect 137462 270444 137468 270456
rect 137520 270444 137526 270496
rect 137646 270444 137652 270496
rect 137704 270484 137710 270496
rect 186130 270484 186136 270496
rect 137704 270456 186136 270484
rect 137704 270444 137710 270456
rect 186130 270444 186136 270456
rect 186188 270444 186194 270496
rect 200758 270444 200764 270496
rect 200816 270484 200822 270496
rect 201862 270484 201868 270496
rect 200816 270456 201868 270484
rect 200816 270444 200822 270456
rect 201862 270444 201868 270456
rect 201920 270444 201926 270496
rect 206830 270444 206836 270496
rect 206888 270484 206894 270496
rect 235810 270484 235816 270496
rect 206888 270456 235816 270484
rect 206888 270444 206894 270456
rect 235810 270444 235816 270456
rect 235868 270444 235874 270496
rect 278314 270444 278320 270496
rect 278372 270484 278378 270496
rect 283834 270484 283840 270496
rect 278372 270456 283840 270484
rect 278372 270444 278378 270456
rect 283834 270444 283840 270456
rect 283892 270444 283898 270496
rect 400858 270444 400864 270496
rect 400916 270484 400922 270496
rect 441614 270484 441620 270496
rect 400916 270456 441620 270484
rect 400916 270444 400922 270456
rect 441614 270444 441620 270456
rect 441672 270444 441678 270496
rect 456426 270444 456432 270496
rect 456484 270484 456490 270496
rect 520274 270484 520280 270496
rect 456484 270456 520280 270484
rect 456484 270444 456490 270456
rect 520274 270444 520280 270456
rect 520332 270444 520338 270496
rect 523126 270444 523132 270496
rect 523184 270484 523190 270496
rect 532878 270484 532884 270496
rect 523184 270456 532884 270484
rect 523184 270444 523190 270456
rect 532878 270444 532884 270456
rect 532936 270444 532942 270496
rect 619634 270484 619640 270496
rect 533356 270456 619640 270484
rect 78858 270308 78864 270360
rect 78916 270348 78922 270360
rect 132494 270348 132500 270360
rect 78916 270320 132500 270348
rect 78916 270308 78922 270320
rect 132494 270308 132500 270320
rect 132552 270308 132558 270360
rect 133782 270308 133788 270360
rect 133840 270348 133846 270360
rect 183646 270348 183652 270360
rect 133840 270320 183652 270348
rect 133840 270308 133846 270320
rect 183646 270308 183652 270320
rect 183704 270308 183710 270360
rect 185302 270308 185308 270360
rect 185360 270348 185366 270360
rect 194410 270348 194416 270360
rect 185360 270320 194416 270348
rect 185360 270308 185366 270320
rect 194410 270308 194416 270320
rect 194468 270308 194474 270360
rect 199930 270308 199936 270360
rect 199988 270348 199994 270360
rect 230842 270348 230848 270360
rect 199988 270320 230848 270348
rect 199988 270308 199994 270320
rect 230842 270308 230848 270320
rect 230900 270308 230906 270360
rect 232682 270308 232688 270360
rect 232740 270348 232746 270360
rect 248230 270348 248236 270360
rect 232740 270320 248236 270348
rect 232740 270308 232746 270320
rect 248230 270308 248236 270320
rect 248288 270308 248294 270360
rect 283098 270308 283104 270360
rect 283156 270348 283162 270360
rect 284662 270348 284668 270360
rect 283156 270320 284668 270348
rect 283156 270308 283162 270320
rect 284662 270308 284668 270320
rect 284720 270308 284726 270360
rect 355042 270308 355048 270360
rect 355100 270348 355106 270360
rect 376938 270348 376944 270360
rect 355100 270320 376944 270348
rect 355100 270308 355106 270320
rect 376938 270308 376944 270320
rect 376996 270308 377002 270360
rect 379698 270308 379704 270360
rect 379756 270348 379762 270360
rect 404354 270348 404360 270360
rect 379756 270320 404360 270348
rect 379756 270308 379762 270320
rect 404354 270308 404360 270320
rect 404412 270308 404418 270360
rect 415026 270308 415032 270360
rect 415084 270348 415090 270360
rect 461210 270348 461216 270360
rect 415084 270320 461216 270348
rect 415084 270308 415090 270320
rect 461210 270308 461216 270320
rect 461268 270308 461274 270360
rect 461394 270308 461400 270360
rect 461452 270348 461458 270360
rect 461452 270320 524644 270348
rect 461452 270308 461458 270320
rect 111978 270172 111984 270224
rect 112036 270212 112042 270224
rect 168742 270212 168748 270224
rect 112036 270184 168748 270212
rect 112036 270172 112042 270184
rect 168742 270172 168748 270184
rect 168800 270172 168806 270224
rect 184842 270172 184848 270224
rect 184900 270212 184906 270224
rect 219342 270212 219348 270224
rect 184900 270184 219348 270212
rect 184900 270172 184906 270184
rect 219342 270172 219348 270184
rect 219400 270172 219406 270224
rect 244366 270172 244372 270224
rect 244424 270212 244430 270224
rect 262306 270212 262312 270224
rect 244424 270184 262312 270212
rect 244424 270172 244430 270184
rect 262306 270172 262312 270184
rect 262364 270172 262370 270224
rect 334342 270172 334348 270224
rect 334400 270212 334406 270224
rect 346394 270212 346400 270224
rect 334400 270184 346400 270212
rect 334400 270172 334406 270184
rect 346394 270172 346400 270184
rect 346452 270172 346458 270224
rect 372246 270172 372252 270224
rect 372304 270212 372310 270224
rect 397454 270212 397460 270224
rect 372304 270184 397460 270212
rect 372304 270172 372310 270184
rect 397454 270172 397460 270184
rect 397512 270172 397518 270224
rect 409598 270172 409604 270224
rect 409656 270212 409662 270224
rect 454034 270212 454040 270224
rect 409656 270184 454040 270212
rect 409656 270172 409662 270184
rect 454034 270172 454040 270184
rect 454092 270172 454098 270224
rect 458818 270172 458824 270224
rect 458876 270212 458882 270224
rect 524414 270212 524420 270224
rect 458876 270184 524420 270212
rect 458876 270172 458882 270184
rect 524414 270172 524420 270184
rect 524472 270172 524478 270224
rect 524616 270212 524644 270320
rect 525610 270308 525616 270360
rect 525668 270348 525674 270360
rect 533356 270348 533384 270456
rect 619634 270444 619640 270456
rect 619692 270444 619698 270496
rect 525668 270320 533384 270348
rect 525668 270308 525674 270320
rect 533522 270308 533528 270360
rect 533580 270348 533586 270360
rect 626534 270348 626540 270360
rect 533580 270320 626540 270348
rect 533580 270308 533586 270320
rect 626534 270308 626540 270320
rect 626592 270308 626598 270360
rect 527174 270212 527180 270224
rect 524616 270184 527180 270212
rect 527174 270172 527180 270184
rect 527232 270172 527238 270224
rect 528370 270172 528376 270224
rect 528428 270212 528434 270224
rect 623958 270212 623964 270224
rect 528428 270184 623964 270212
rect 528428 270172 528434 270184
rect 623958 270172 623964 270184
rect 624016 270172 624022 270224
rect 89622 270036 89628 270088
rect 89680 270076 89686 270088
rect 153010 270076 153016 270088
rect 89680 270048 153016 270076
rect 89680 270036 89686 270048
rect 153010 270036 153016 270048
rect 153068 270036 153074 270088
rect 176562 270036 176568 270088
rect 176620 270076 176626 270088
rect 211154 270076 211160 270088
rect 176620 270048 211160 270076
rect 176620 270036 176626 270048
rect 211154 270036 211160 270048
rect 211212 270036 211218 270088
rect 212442 270036 212448 270088
rect 212500 270076 212506 270088
rect 239950 270076 239956 270088
rect 212500 270048 239956 270076
rect 212500 270036 212506 270048
rect 239950 270036 239956 270048
rect 240008 270036 240014 270088
rect 241882 270036 241888 270088
rect 241940 270076 241946 270088
rect 260650 270076 260656 270088
rect 241940 270048 260656 270076
rect 241940 270036 241946 270048
rect 260650 270036 260656 270048
rect 260708 270036 260714 270088
rect 266170 270036 266176 270088
rect 266228 270076 266234 270088
rect 277210 270076 277216 270088
rect 266228 270048 277216 270076
rect 266228 270036 266234 270048
rect 277210 270036 277216 270048
rect 277268 270036 277274 270088
rect 345290 270036 345296 270088
rect 345348 270076 345354 270088
rect 358814 270076 358820 270088
rect 345348 270048 358820 270076
rect 345348 270036 345354 270048
rect 358814 270036 358820 270048
rect 358872 270036 358878 270088
rect 366634 270036 366640 270088
rect 366692 270076 366698 270088
rect 393314 270076 393320 270088
rect 366692 270048 393320 270076
rect 366692 270036 366698 270048
rect 393314 270036 393320 270048
rect 393372 270036 393378 270088
rect 394694 270036 394700 270088
rect 394752 270076 394758 270088
rect 408770 270076 408776 270088
rect 394752 270048 408776 270076
rect 394752 270036 394758 270048
rect 408770 270036 408776 270048
rect 408828 270036 408834 270088
rect 412450 270036 412456 270088
rect 412508 270076 412514 270088
rect 458174 270076 458180 270088
rect 412508 270048 458180 270076
rect 412508 270036 412514 270048
rect 458174 270036 458180 270048
rect 458232 270036 458238 270088
rect 463510 270036 463516 270088
rect 463568 270076 463574 270088
rect 530762 270076 530768 270088
rect 463568 270048 530768 270076
rect 463568 270036 463574 270048
rect 530762 270036 530768 270048
rect 530820 270036 530826 270088
rect 530946 270036 530952 270088
rect 531004 270076 531010 270088
rect 533154 270076 533160 270088
rect 531004 270048 533160 270076
rect 531004 270036 531010 270048
rect 533154 270036 533160 270048
rect 533212 270036 533218 270088
rect 538306 270076 538312 270088
rect 533356 270048 538312 270076
rect 85482 269900 85488 269952
rect 85540 269940 85546 269952
rect 149422 269940 149428 269952
rect 85540 269912 149428 269940
rect 85540 269900 85546 269912
rect 149422 269900 149428 269912
rect 149480 269900 149486 269952
rect 152826 269900 152832 269952
rect 152884 269940 152890 269952
rect 157150 269940 157156 269952
rect 152884 269912 157156 269940
rect 152884 269900 152890 269912
rect 157150 269900 157156 269912
rect 157208 269900 157214 269952
rect 173802 269900 173808 269952
rect 173860 269940 173866 269952
rect 212626 269940 212632 269952
rect 173860 269912 212632 269940
rect 173860 269900 173866 269912
rect 212626 269900 212632 269912
rect 212684 269900 212690 269952
rect 226610 269900 226616 269952
rect 226668 269940 226674 269952
rect 249886 269940 249892 269952
rect 226668 269912 249892 269940
rect 226668 269900 226674 269912
rect 249886 269900 249892 269912
rect 249944 269900 249950 269952
rect 256878 269900 256884 269952
rect 256936 269940 256942 269952
rect 268930 269940 268936 269952
rect 256936 269912 268936 269940
rect 256936 269900 256942 269912
rect 268930 269900 268936 269912
rect 268988 269900 268994 269952
rect 330202 269900 330208 269952
rect 330260 269940 330266 269952
rect 340874 269940 340880 269952
rect 330260 269912 340880 269940
rect 330260 269900 330266 269912
rect 340874 269900 340880 269912
rect 340932 269900 340938 269952
rect 341794 269900 341800 269952
rect 341852 269940 341858 269952
rect 357434 269940 357440 269952
rect 341852 269912 357440 269940
rect 341852 269900 341858 269912
rect 357434 269900 357440 269912
rect 357492 269900 357498 269952
rect 359182 269900 359188 269952
rect 359240 269940 359246 269952
rect 382274 269940 382280 269952
rect 359240 269912 382280 269940
rect 359240 269900 359246 269912
rect 382274 269900 382280 269912
rect 382332 269900 382338 269952
rect 383010 269900 383016 269952
rect 383068 269940 383074 269952
rect 411254 269940 411260 269952
rect 383068 269912 411260 269940
rect 383068 269900 383074 269912
rect 411254 269900 411260 269912
rect 411312 269900 411318 269952
rect 419626 269900 419632 269952
rect 419684 269940 419690 269952
rect 467926 269940 467932 269952
rect 419684 269912 467932 269940
rect 419684 269900 419690 269912
rect 467926 269900 467932 269912
rect 467984 269900 467990 269952
rect 468478 269900 468484 269952
rect 468536 269940 468542 269952
rect 533356 269940 533384 270048
rect 538306 270036 538312 270048
rect 538364 270036 538370 270088
rect 630674 270076 630680 270088
rect 538876 270048 630680 270076
rect 468536 269912 533384 269940
rect 468536 269900 468542 269912
rect 533982 269900 533988 269952
rect 534040 269940 534046 269952
rect 538876 269940 538904 270048
rect 630674 270036 630680 270048
rect 630732 270036 630738 270088
rect 534040 269912 538904 269940
rect 534040 269900 534046 269912
rect 540514 269900 540520 269952
rect 540572 269940 540578 269952
rect 640518 269940 640524 269952
rect 540572 269912 640524 269940
rect 540572 269900 540578 269912
rect 640518 269900 640524 269912
rect 640576 269900 640582 269952
rect 70578 269764 70584 269816
rect 70636 269804 70642 269816
rect 79318 269804 79324 269816
rect 70636 269776 79324 269804
rect 70636 269764 70642 269776
rect 79318 269764 79324 269776
rect 79376 269764 79382 269816
rect 80054 269764 80060 269816
rect 80112 269804 80118 269816
rect 146386 269804 146392 269816
rect 80112 269776 146392 269804
rect 80112 269764 80118 269776
rect 146386 269764 146392 269776
rect 146444 269764 146450 269816
rect 158622 269764 158628 269816
rect 158680 269804 158686 269816
rect 201034 269804 201040 269816
rect 158680 269776 201040 269804
rect 158680 269764 158686 269776
rect 201034 269764 201040 269776
rect 201092 269764 201098 269816
rect 201678 269764 201684 269816
rect 201736 269804 201742 269816
rect 232498 269804 232504 269816
rect 201736 269776 232504 269804
rect 201736 269764 201742 269776
rect 232498 269764 232504 269776
rect 232556 269764 232562 269816
rect 237282 269764 237288 269816
rect 237340 269804 237346 269816
rect 257338 269804 257344 269816
rect 237340 269776 257344 269804
rect 237340 269764 237346 269776
rect 257338 269764 257344 269776
rect 257396 269764 257402 269816
rect 258534 269764 258540 269816
rect 258592 269804 258598 269816
rect 272242 269804 272248 269816
rect 258592 269776 272248 269804
rect 258592 269764 258598 269776
rect 272242 269764 272248 269776
rect 272300 269764 272306 269816
rect 273070 269764 273076 269816
rect 273128 269804 273134 269816
rect 282178 269804 282184 269816
rect 273128 269776 282184 269804
rect 273128 269764 273134 269776
rect 282178 269764 282184 269776
rect 282236 269764 282242 269816
rect 326890 269764 326896 269816
rect 326948 269804 326954 269816
rect 335538 269804 335544 269816
rect 326948 269776 335544 269804
rect 326948 269764 326954 269776
rect 335538 269764 335544 269776
rect 335596 269764 335602 269816
rect 335998 269764 336004 269816
rect 336056 269804 336062 269816
rect 349154 269804 349160 269816
rect 336056 269776 349160 269804
rect 336056 269764 336062 269776
rect 349154 269764 349160 269776
rect 349212 269764 349218 269816
rect 351730 269764 351736 269816
rect 351788 269804 351794 269816
rect 371234 269804 371240 269816
rect 351788 269776 371240 269804
rect 351788 269764 351794 269776
rect 371234 269764 371240 269776
rect 371292 269764 371298 269816
rect 376570 269764 376576 269816
rect 376628 269804 376634 269816
rect 407114 269804 407120 269816
rect 376628 269776 407120 269804
rect 376628 269764 376634 269776
rect 407114 269764 407120 269776
rect 407172 269764 407178 269816
rect 417142 269764 417148 269816
rect 417200 269804 417206 269816
rect 465074 269804 465080 269816
rect 417200 269776 465080 269804
rect 417200 269764 417206 269776
rect 465074 269764 465080 269776
rect 465132 269764 465138 269816
rect 465994 269764 466000 269816
rect 466052 269804 466058 269816
rect 530394 269804 530400 269816
rect 466052 269776 530400 269804
rect 466052 269764 466058 269776
rect 530394 269764 530400 269776
rect 530452 269764 530458 269816
rect 538490 269804 538496 269816
rect 530596 269776 538496 269804
rect 122742 269628 122748 269680
rect 122800 269668 122806 269680
rect 176194 269668 176200 269680
rect 122800 269640 176200 269668
rect 122800 269628 122806 269640
rect 176194 269628 176200 269640
rect 176252 269628 176258 269680
rect 183462 269628 183468 269680
rect 183520 269668 183526 269680
rect 205450 269668 205456 269680
rect 183520 269640 205456 269668
rect 183520 269628 183526 269640
rect 205450 269628 205456 269640
rect 205508 269628 205514 269680
rect 392026 269628 392032 269680
rect 392084 269668 392090 269680
rect 401686 269668 401692 269680
rect 392084 269640 401692 269668
rect 392084 269628 392090 269640
rect 401686 269628 401692 269640
rect 401744 269628 401750 269680
rect 404354 269628 404360 269680
rect 404412 269668 404418 269680
rect 423674 269668 423680 269680
rect 404412 269640 423680 269668
rect 404412 269628 404418 269640
rect 423674 269628 423680 269640
rect 423732 269628 423738 269680
rect 423858 269628 423864 269680
rect 423916 269668 423922 269680
rect 451366 269668 451372 269680
rect 423916 269640 451372 269668
rect 423916 269628 423922 269640
rect 451366 269628 451372 269640
rect 451424 269628 451430 269680
rect 453574 269628 453580 269680
rect 453632 269668 453638 269680
rect 509234 269668 509240 269680
rect 453632 269640 509240 269668
rect 453632 269628 453638 269640
rect 509234 269628 509240 269640
rect 509292 269628 509298 269680
rect 530596 269668 530624 269776
rect 538490 269764 538496 269776
rect 538548 269764 538554 269816
rect 538674 269764 538680 269816
rect 538732 269804 538738 269816
rect 541158 269804 541164 269816
rect 538732 269776 541164 269804
rect 538732 269764 538738 269776
rect 541158 269764 541164 269776
rect 541216 269764 541222 269816
rect 541342 269764 541348 269816
rect 541400 269804 541406 269816
rect 637574 269804 637580 269816
rect 541400 269776 637580 269804
rect 541400 269764 541406 269776
rect 637574 269764 637580 269776
rect 637632 269764 637638 269816
rect 509712 269640 530624 269668
rect 129642 269492 129648 269544
rect 129700 269532 129706 269544
rect 181162 269532 181168 269544
rect 129700 269504 181168 269532
rect 129700 269492 129706 269504
rect 181162 269492 181168 269504
rect 181220 269492 181226 269544
rect 204162 269492 204168 269544
rect 204220 269532 204226 269544
rect 223482 269532 223488 269544
rect 204220 269504 223488 269532
rect 204220 269492 204226 269504
rect 223482 269492 223488 269504
rect 223540 269492 223546 269544
rect 398742 269492 398748 269544
rect 398800 269532 398806 269544
rect 412634 269532 412640 269544
rect 398800 269504 412640 269532
rect 398800 269492 398806 269504
rect 412634 269492 412640 269504
rect 412692 269492 412698 269544
rect 424594 269492 424600 269544
rect 424652 269532 424658 269544
rect 475010 269532 475016 269544
rect 424652 269504 475016 269532
rect 424652 269492 424658 269504
rect 475010 269492 475016 269504
rect 475068 269492 475074 269544
rect 495250 269492 495256 269544
rect 495308 269532 495314 269544
rect 509712 269532 509740 269640
rect 532878 269628 532884 269680
rect 532936 269668 532942 269680
rect 616414 269668 616420 269680
rect 532936 269640 616420 269668
rect 532936 269628 532942 269640
rect 616414 269628 616420 269640
rect 616472 269628 616478 269680
rect 495308 269504 509740 269532
rect 495308 269492 495314 269504
rect 509878 269492 509884 269544
rect 509936 269532 509942 269544
rect 596174 269532 596180 269544
rect 509936 269504 596180 269532
rect 509936 269492 509942 269504
rect 596174 269492 596180 269504
rect 596232 269492 596238 269544
rect 126882 269356 126888 269408
rect 126940 269396 126946 269408
rect 178678 269396 178684 269408
rect 126940 269368 178684 269396
rect 126940 269356 126946 269368
rect 178678 269356 178684 269368
rect 178736 269356 178742 269408
rect 408402 269356 408408 269408
rect 408460 269396 408466 269408
rect 426526 269396 426532 269408
rect 408460 269368 426532 269396
rect 408460 269356 408466 269368
rect 426526 269356 426532 269368
rect 426584 269356 426590 269408
rect 441614 269356 441620 269408
rect 441672 269396 441678 269408
rect 458450 269396 458456 269408
rect 441672 269368 458456 269396
rect 441672 269356 441678 269368
rect 458450 269356 458456 269368
rect 458508 269356 458514 269408
rect 470962 269356 470968 269408
rect 471020 269396 471026 269408
rect 538306 269396 538312 269408
rect 471020 269368 538312 269396
rect 471020 269356 471026 269368
rect 538306 269356 538312 269368
rect 538364 269356 538370 269408
rect 538490 269356 538496 269408
rect 538548 269396 538554 269408
rect 575474 269396 575480 269408
rect 538548 269368 575480 269396
rect 538548 269356 538554 269368
rect 575474 269356 575480 269368
rect 575532 269356 575538 269408
rect 143902 269220 143908 269272
rect 143960 269260 143966 269272
rect 191098 269260 191104 269272
rect 143960 269232 191104 269260
rect 143960 269220 143966 269232
rect 191098 269220 191104 269232
rect 191156 269220 191162 269272
rect 282730 269220 282736 269272
rect 282788 269260 282794 269272
rect 288802 269260 288808 269272
rect 282788 269232 288808 269260
rect 282788 269220 282794 269232
rect 288802 269220 288808 269232
rect 288860 269220 288866 269272
rect 401686 269220 401692 269272
rect 401744 269260 401750 269272
rect 416774 269260 416780 269272
rect 401744 269232 416780 269260
rect 401744 269220 401750 269232
rect 416774 269220 416780 269232
rect 416832 269220 416838 269272
rect 474274 269220 474280 269272
rect 474332 269260 474338 269272
rect 474332 269232 534074 269260
rect 474332 269220 474338 269232
rect 534046 269192 534074 269232
rect 546494 269192 546500 269204
rect 534046 269164 546500 269192
rect 546494 269152 546500 269164
rect 546552 269152 546558 269204
rect 319438 269084 319444 269136
rect 319496 269124 319502 269136
rect 325694 269124 325700 269136
rect 319496 269096 325700 269124
rect 319496 269084 319502 269096
rect 325694 269084 325700 269096
rect 325752 269084 325758 269136
rect 118602 269016 118608 269068
rect 118660 269056 118666 269068
rect 174538 269056 174544 269068
rect 118660 269028 174544 269056
rect 118660 269016 118666 269028
rect 174538 269016 174544 269028
rect 174596 269016 174602 269068
rect 175090 269016 175096 269068
rect 175148 269056 175154 269068
rect 177666 269056 177672 269068
rect 175148 269028 177672 269056
rect 175148 269016 175154 269028
rect 177666 269016 177672 269028
rect 177724 269016 177730 269068
rect 273254 269016 273260 269068
rect 273312 269056 273318 269068
rect 275554 269056 275560 269068
rect 273312 269028 275560 269056
rect 273312 269016 273318 269028
rect 275554 269016 275560 269028
rect 275612 269016 275618 269068
rect 433702 269016 433708 269068
rect 433760 269056 433766 269068
rect 488534 269056 488540 269068
rect 433760 269028 488540 269056
rect 433760 269016 433766 269028
rect 488534 269016 488540 269028
rect 488592 269016 488598 269068
rect 493318 269016 493324 269068
rect 493376 269056 493382 269068
rect 574094 269056 574100 269068
rect 493376 269028 574100 269056
rect 493376 269016 493382 269028
rect 574094 269016 574100 269028
rect 574152 269016 574158 269068
rect 115842 268880 115848 268932
rect 115900 268920 115906 268932
rect 171226 268920 171232 268932
rect 115900 268892 171232 268920
rect 115900 268880 115906 268892
rect 171226 268880 171232 268892
rect 171284 268880 171290 268932
rect 382366 268880 382372 268932
rect 382424 268920 382430 268932
rect 415394 268920 415400 268932
rect 382424 268892 415400 268920
rect 382424 268880 382430 268892
rect 415394 268880 415400 268892
rect 415452 268880 415458 268932
rect 436554 268880 436560 268932
rect 436612 268920 436618 268932
rect 491662 268920 491668 268932
rect 436612 268892 491668 268920
rect 436612 268880 436618 268892
rect 491662 268880 491668 268892
rect 491720 268880 491726 268932
rect 498286 268880 498292 268932
rect 498344 268920 498350 268932
rect 580994 268920 581000 268932
rect 498344 268892 581000 268920
rect 498344 268880 498350 268892
rect 580994 268880 581000 268892
rect 581052 268880 581058 268932
rect 110322 268744 110328 268796
rect 110380 268784 110386 268796
rect 167914 268784 167920 268796
rect 110380 268756 167920 268784
rect 110380 268744 110386 268756
rect 167914 268744 167920 268756
rect 167972 268744 167978 268796
rect 168282 268744 168288 268796
rect 168340 268784 168346 268796
rect 181990 268784 181996 268796
rect 168340 268756 181996 268784
rect 168340 268744 168346 268756
rect 181990 268744 181996 268756
rect 182048 268744 182054 268796
rect 188890 268744 188896 268796
rect 188948 268784 188954 268796
rect 190454 268784 190460 268796
rect 188948 268756 190460 268784
rect 188948 268744 188954 268756
rect 190454 268744 190460 268756
rect 190512 268744 190518 268796
rect 200574 268744 200580 268796
rect 200632 268784 200638 268796
rect 231302 268784 231308 268796
rect 200632 268756 231308 268784
rect 200632 268744 200638 268756
rect 231302 268744 231308 268756
rect 231360 268744 231366 268796
rect 387334 268744 387340 268796
rect 387392 268784 387398 268796
rect 422294 268784 422300 268796
rect 387392 268756 422300 268784
rect 387392 268744 387398 268756
rect 422294 268744 422300 268756
rect 422352 268744 422358 268796
rect 438670 268744 438676 268796
rect 438728 268784 438734 268796
rect 495434 268784 495440 268796
rect 438728 268756 495440 268784
rect 438728 268744 438734 268756
rect 495434 268744 495440 268756
rect 495492 268744 495498 268796
rect 500770 268744 500776 268796
rect 500828 268784 500834 268796
rect 583754 268784 583760 268796
rect 500828 268756 583760 268784
rect 500828 268744 500834 268756
rect 583754 268744 583760 268756
rect 583812 268744 583818 268796
rect 104986 268608 104992 268660
rect 105044 268648 105050 268660
rect 163774 268648 163780 268660
rect 105044 268620 163780 268648
rect 105044 268608 105050 268620
rect 163774 268608 163780 268620
rect 163832 268608 163838 268660
rect 176930 268608 176936 268660
rect 176988 268648 176994 268660
rect 215110 268648 215116 268660
rect 176988 268620 215116 268648
rect 176988 268608 176994 268620
rect 215110 268608 215116 268620
rect 215168 268608 215174 268660
rect 224218 268608 224224 268660
rect 224276 268648 224282 268660
rect 243262 268648 243268 268660
rect 224276 268620 243268 268648
rect 224276 268608 224282 268620
rect 243262 268608 243268 268620
rect 243320 268608 243326 268660
rect 352558 268608 352564 268660
rect 352616 268648 352622 268660
rect 372614 268648 372620 268660
rect 352616 268620 372620 268648
rect 352616 268608 352622 268620
rect 372614 268608 372620 268620
rect 372672 268608 372678 268660
rect 393682 268608 393688 268660
rect 393740 268648 393746 268660
rect 429194 268648 429200 268660
rect 393740 268620 429200 268648
rect 393740 268608 393746 268620
rect 429194 268608 429200 268620
rect 429252 268608 429258 268660
rect 441154 268608 441160 268660
rect 441212 268648 441218 268660
rect 499574 268648 499580 268660
rect 441212 268620 499580 268648
rect 441212 268608 441218 268620
rect 499574 268608 499580 268620
rect 499632 268608 499638 268660
rect 503254 268608 503260 268660
rect 503312 268648 503318 268660
rect 587894 268648 587900 268660
rect 503312 268620 587900 268648
rect 503312 268608 503318 268620
rect 587894 268608 587900 268620
rect 587952 268608 587958 268660
rect 99282 268472 99288 268524
rect 99340 268512 99346 268524
rect 160462 268512 160468 268524
rect 99340 268484 160468 268512
rect 99340 268472 99346 268484
rect 160462 268472 160468 268484
rect 160520 268472 160526 268524
rect 180610 268472 180616 268524
rect 180668 268512 180674 268524
rect 217594 268512 217600 268524
rect 180668 268484 217600 268512
rect 180668 268472 180674 268484
rect 217594 268472 217600 268484
rect 217652 268472 217658 268524
rect 231670 268472 231676 268524
rect 231728 268512 231734 268524
rect 253198 268512 253204 268524
rect 231728 268484 253204 268512
rect 231728 268472 231734 268484
rect 253198 268472 253204 268484
rect 253256 268472 253262 268524
rect 338482 268472 338488 268524
rect 338540 268512 338546 268524
rect 352098 268512 352104 268524
rect 338540 268484 352104 268512
rect 338540 268472 338546 268484
rect 352098 268472 352104 268484
rect 352156 268472 352162 268524
rect 367462 268472 367468 268524
rect 367520 268512 367526 268524
rect 393498 268512 393504 268524
rect 367520 268484 393504 268512
rect 367520 268472 367526 268484
rect 393498 268472 393504 268484
rect 393556 268472 393562 268524
rect 397270 268472 397276 268524
rect 397328 268512 397334 268524
rect 436094 268512 436100 268524
rect 397328 268484 436100 268512
rect 397328 268472 397334 268484
rect 436094 268472 436100 268484
rect 436152 268472 436158 268524
rect 446122 268472 446128 268524
rect 446180 268512 446186 268524
rect 506474 268512 506480 268524
rect 446180 268484 506480 268512
rect 446180 268472 446186 268484
rect 506474 268472 506480 268484
rect 506532 268472 506538 268524
rect 508222 268472 508228 268524
rect 508280 268512 508286 268524
rect 594794 268512 594800 268524
rect 508280 268484 594800 268512
rect 508280 268472 508286 268484
rect 594794 268472 594800 268484
rect 594852 268472 594858 268524
rect 92382 268336 92388 268388
rect 92440 268376 92446 268388
rect 155494 268376 155500 268388
rect 92440 268348 155500 268376
rect 92440 268336 92446 268348
rect 155494 268336 155500 268348
rect 155552 268336 155558 268388
rect 161566 268336 161572 268388
rect 161624 268376 161630 268388
rect 203518 268376 203524 268388
rect 161624 268348 203524 268376
rect 161624 268336 161630 268348
rect 203518 268336 203524 268348
rect 203576 268336 203582 268388
rect 210694 268336 210700 268388
rect 210752 268376 210758 268388
rect 236638 268376 236644 268388
rect 210752 268348 236644 268376
rect 210752 268336 210758 268348
rect 236638 268336 236644 268348
rect 236696 268336 236702 268388
rect 252646 268336 252652 268388
rect 252704 268376 252710 268388
rect 268102 268376 268108 268388
rect 252704 268348 268108 268376
rect 252704 268336 252710 268348
rect 268102 268336 268108 268348
rect 268160 268336 268166 268388
rect 348786 268336 348792 268388
rect 348844 268376 348850 268388
rect 367094 268376 367100 268388
rect 348844 268348 367100 268376
rect 348844 268336 348850 268348
rect 367094 268336 367100 268348
rect 367152 268336 367158 268388
rect 372430 268336 372436 268388
rect 372488 268376 372494 268388
rect 400490 268376 400496 268388
rect 372488 268348 400496 268376
rect 372488 268336 372494 268348
rect 400490 268336 400496 268348
rect 400548 268336 400554 268388
rect 402238 268336 402244 268388
rect 402296 268376 402302 268388
rect 443086 268376 443092 268388
rect 402296 268348 443092 268376
rect 402296 268336 402302 268348
rect 443086 268336 443092 268348
rect 443144 268336 443150 268388
rect 461854 268336 461860 268388
rect 461912 268376 461918 268388
rect 528554 268376 528560 268388
rect 461912 268348 528560 268376
rect 461912 268336 461918 268348
rect 528554 268336 528560 268348
rect 528612 268336 528618 268388
rect 541342 268336 541348 268388
rect 541400 268376 541406 268388
rect 641714 268376 641720 268388
rect 541400 268348 641720 268376
rect 541400 268336 541406 268348
rect 641714 268336 641720 268348
rect 641772 268336 641778 268388
rect 135622 268200 135628 268252
rect 135680 268240 135686 268252
rect 140130 268240 140136 268252
rect 135680 268212 140136 268240
rect 135680 268200 135686 268212
rect 140130 268200 140136 268212
rect 140188 268200 140194 268252
rect 140682 268200 140688 268252
rect 140740 268240 140746 268252
rect 188614 268240 188620 268252
rect 140740 268212 188620 268240
rect 140740 268200 140746 268212
rect 188614 268200 188620 268212
rect 188672 268200 188678 268252
rect 416222 268200 416228 268252
rect 416280 268240 416286 268252
rect 447134 268240 447140 268252
rect 416280 268212 447140 268240
rect 416280 268200 416286 268212
rect 447134 268200 447140 268212
rect 447192 268200 447198 268252
rect 448422 268200 448428 268252
rect 448480 268240 448486 268252
rect 494054 268240 494060 268252
rect 448480 268212 494060 268240
rect 448480 268200 448486 268212
rect 494054 268200 494060 268212
rect 494112 268200 494118 268252
rect 495802 268200 495808 268252
rect 495860 268240 495866 268252
rect 576854 268240 576860 268252
rect 495860 268212 576860 268240
rect 495860 268200 495866 268212
rect 576854 268200 576860 268212
rect 576912 268200 576918 268252
rect 151722 268064 151728 268116
rect 151780 268104 151786 268116
rect 196066 268104 196072 268116
rect 151780 268076 196072 268104
rect 151780 268064 151786 268076
rect 196066 268064 196072 268076
rect 196124 268064 196130 268116
rect 422294 268064 422300 268116
rect 422352 268104 422358 268116
rect 444374 268104 444380 268116
rect 422352 268076 444380 268104
rect 422352 268064 422358 268076
rect 444374 268064 444380 268076
rect 444432 268064 444438 268116
rect 527174 268064 527180 268116
rect 527232 268104 527238 268116
rect 607398 268104 607404 268116
rect 527232 268076 607404 268104
rect 527232 268064 527238 268076
rect 607398 268064 607404 268076
rect 607456 268064 607462 268116
rect 490834 267928 490840 267980
rect 490892 267968 490898 267980
rect 569954 267968 569960 267980
rect 490892 267940 569960 267968
rect 490892 267928 490898 267940
rect 569954 267928 569960 267940
rect 570012 267928 570018 267980
rect 276474 267724 276480 267776
rect 276532 267764 276538 267776
rect 278038 267764 278044 267776
rect 276532 267736 278044 267764
rect 276532 267724 276538 267736
rect 278038 267724 278044 267736
rect 278096 267724 278102 267776
rect 119338 267656 119344 267708
rect 119396 267696 119402 267708
rect 153470 267696 153476 267708
rect 119396 267668 153476 267696
rect 119396 267656 119402 267668
rect 153470 267656 153476 267668
rect 153528 267656 153534 267708
rect 153838 267656 153844 267708
rect 153896 267696 153902 267708
rect 184474 267696 184480 267708
rect 153896 267668 184480 267696
rect 153896 267656 153902 267668
rect 184474 267656 184480 267668
rect 184532 267656 184538 267708
rect 365806 267656 365812 267708
rect 365864 267696 365870 267708
rect 381538 267696 381544 267708
rect 365864 267668 381544 267696
rect 365864 267656 365870 267668
rect 381538 267656 381544 267668
rect 381596 267656 381602 267708
rect 388162 267656 388168 267708
rect 388220 267696 388226 267708
rect 404354 267696 404360 267708
rect 388220 267668 404360 267696
rect 388220 267656 388226 267668
rect 404354 267656 404360 267668
rect 404412 267656 404418 267708
rect 408034 267656 408040 267708
rect 408092 267696 408098 267708
rect 423858 267696 423864 267708
rect 408092 267668 423864 267696
rect 408092 267656 408098 267668
rect 423858 267656 423864 267668
rect 423916 267656 423922 267708
rect 445294 267656 445300 267708
rect 445352 267696 445358 267708
rect 490558 267696 490564 267708
rect 445352 267668 490564 267696
rect 445352 267656 445358 267668
rect 490558 267656 490564 267668
rect 490616 267656 490622 267708
rect 509878 267656 509884 267708
rect 509936 267696 509942 267708
rect 567838 267696 567844 267708
rect 509936 267668 567844 267696
rect 509936 267656 509942 267668
rect 567838 267656 567844 267668
rect 567896 267656 567902 267708
rect 111702 267520 111708 267572
rect 111760 267560 111766 267572
rect 168558 267560 168564 267572
rect 111760 267532 168564 267560
rect 111760 267520 111766 267532
rect 168558 267520 168564 267532
rect 168616 267520 168622 267572
rect 169018 267520 169024 267572
rect 169076 267560 169082 267572
rect 199378 267560 199384 267572
rect 169076 267532 199384 267560
rect 169076 267520 169082 267532
rect 199378 267520 199384 267532
rect 199436 267520 199442 267572
rect 215938 267520 215944 267572
rect 215996 267560 216002 267572
rect 222562 267560 222568 267572
rect 215996 267532 222568 267560
rect 215996 267520 216002 267532
rect 222562 267520 222568 267532
rect 222620 267520 222626 267572
rect 371602 267520 371608 267572
rect 371660 267560 371666 267572
rect 373258 267560 373264 267572
rect 371660 267532 373264 267560
rect 371660 267520 371666 267532
rect 373258 267520 373264 267532
rect 373316 267520 373322 267572
rect 390646 267520 390652 267572
rect 390704 267560 390710 267572
rect 408402 267560 408408 267572
rect 390704 267532 408408 267560
rect 390704 267520 390710 267532
rect 408402 267520 408408 267532
rect 408460 267520 408466 267572
rect 421282 267520 421288 267572
rect 421340 267560 421346 267572
rect 440878 267560 440884 267572
rect 421340 267532 440884 267560
rect 421340 267520 421346 267532
rect 440878 267520 440884 267532
rect 440936 267520 440942 267572
rect 447778 267520 447784 267572
rect 447836 267560 447842 267572
rect 456058 267560 456064 267572
rect 447836 267532 456064 267560
rect 447836 267520 447842 267532
rect 456058 267520 456064 267532
rect 456116 267520 456122 267572
rect 460198 267520 460204 267572
rect 460256 267560 460262 267572
rect 516778 267560 516784 267572
rect 460256 267532 516784 267560
rect 460256 267520 460262 267532
rect 516778 267520 516784 267532
rect 516836 267520 516842 267572
rect 519814 267520 519820 267572
rect 519872 267560 519878 267572
rect 583018 267560 583024 267572
rect 519872 267532 583024 267560
rect 519872 267520 519878 267532
rect 583018 267520 583024 267532
rect 583076 267520 583082 267572
rect 86218 267384 86224 267436
rect 86276 267424 86282 267436
rect 144730 267424 144736 267436
rect 86276 267396 144736 267424
rect 86276 267384 86282 267396
rect 144730 267384 144736 267396
rect 144788 267384 144794 267436
rect 145558 267384 145564 267436
rect 145616 267424 145622 267436
rect 191926 267424 191932 267436
rect 145616 267396 191932 267424
rect 145616 267384 145622 267396
rect 191926 267384 191932 267396
rect 191984 267384 191990 267436
rect 199562 267384 199568 267436
rect 199620 267424 199626 267436
rect 204346 267424 204352 267436
rect 199620 267396 204352 267424
rect 199620 267384 199626 267396
rect 204346 267384 204352 267396
rect 204404 267384 204410 267436
rect 205450 267384 205456 267436
rect 205508 267424 205514 267436
rect 218422 267424 218428 267436
rect 205508 267396 218428 267424
rect 205508 267384 205514 267396
rect 218422 267384 218428 267396
rect 218480 267384 218486 267436
rect 233878 267384 233884 267436
rect 233936 267424 233942 267436
rect 233936 267396 238754 267424
rect 233936 267384 233942 267396
rect 104802 267248 104808 267300
rect 104860 267288 104866 267300
rect 164602 267288 164608 267300
rect 104860 267260 164608 267288
rect 104860 267248 104866 267260
rect 164602 267248 164608 267260
rect 164660 267248 164666 267300
rect 186958 267248 186964 267300
rect 187016 267288 187022 267300
rect 219250 267288 219256 267300
rect 187016 267260 219256 267288
rect 187016 267248 187022 267260
rect 219250 267248 219256 267260
rect 219308 267248 219314 267300
rect 223482 267248 223488 267300
rect 223540 267288 223546 267300
rect 234154 267288 234160 267300
rect 223540 267260 234160 267288
rect 223540 267248 223546 267260
rect 234154 267248 234160 267260
rect 234212 267248 234218 267300
rect 238726 267288 238754 267396
rect 243538 267384 243544 267436
rect 243596 267424 243602 267436
rect 251542 267424 251548 267436
rect 243596 267396 251548 267424
rect 243596 267384 243602 267396
rect 251542 267384 251548 267396
rect 251600 267384 251606 267436
rect 315298 267384 315304 267436
rect 315356 267424 315362 267436
rect 319162 267424 319168 267436
rect 315356 267396 319168 267424
rect 315356 267384 315362 267396
rect 319162 267384 319168 267396
rect 319220 267384 319226 267436
rect 340966 267384 340972 267436
rect 341024 267424 341030 267436
rect 355318 267424 355324 267436
rect 341024 267396 355324 267424
rect 341024 267384 341030 267396
rect 355318 267384 355324 267396
rect 355376 267384 355382 267436
rect 362494 267384 362500 267436
rect 362552 267424 362558 267436
rect 369118 267424 369124 267436
rect 362552 267396 369124 267424
rect 362552 267384 362558 267396
rect 369118 267384 369124 267396
rect 369176 267384 369182 267436
rect 374454 267424 374460 267436
rect 369320 267396 374460 267424
rect 244090 267288 244096 267300
rect 238726 267260 244096 267288
rect 244090 267248 244096 267260
rect 244148 267248 244154 267300
rect 321922 267248 321928 267300
rect 321980 267288 321986 267300
rect 327718 267288 327724 267300
rect 321980 267260 327724 267288
rect 321980 267248 321986 267260
rect 327718 267248 327724 267260
rect 327776 267248 327782 267300
rect 350902 267248 350908 267300
rect 350960 267288 350966 267300
rect 362218 267288 362224 267300
rect 350960 267260 362224 267288
rect 350960 267248 350966 267260
rect 362218 267248 362224 267260
rect 362276 267248 362282 267300
rect 90358 267112 90364 267164
rect 90416 267152 90422 267164
rect 151354 267152 151360 267164
rect 90416 267124 151360 267152
rect 90416 267112 90422 267124
rect 151354 267112 151360 267124
rect 151412 267112 151418 267164
rect 168098 267112 168104 267164
rect 168156 267152 168162 267164
rect 177022 267152 177028 267164
rect 168156 267124 177028 267152
rect 168156 267112 168162 267124
rect 177022 267112 177028 267124
rect 177080 267112 177086 267164
rect 177666 267112 177672 267164
rect 177724 267152 177730 267164
rect 214282 267152 214288 267164
rect 177724 267124 214288 267152
rect 177724 267112 177730 267124
rect 214282 267112 214288 267124
rect 214340 267112 214346 267164
rect 220078 267112 220084 267164
rect 220136 267152 220142 267164
rect 239122 267152 239128 267164
rect 220136 267124 239128 267152
rect 220136 267112 220142 267124
rect 239122 267112 239128 267124
rect 239180 267112 239186 267164
rect 246942 267112 246948 267164
rect 247000 267152 247006 267164
rect 263962 267152 263968 267164
rect 247000 267124 263968 267152
rect 247000 267112 247006 267124
rect 263962 267112 263968 267124
rect 264020 267112 264026 267164
rect 312814 267112 312820 267164
rect 312872 267152 312878 267164
rect 316034 267152 316040 267164
rect 312872 267124 316040 267152
rect 312872 267112 312878 267124
rect 316034 267112 316040 267124
rect 316092 267112 316098 267164
rect 360010 267112 360016 267164
rect 360068 267152 360074 267164
rect 366358 267152 366364 267164
rect 360068 267124 366364 267152
rect 360068 267112 360074 267124
rect 366358 267112 366364 267124
rect 366416 267112 366422 267164
rect 79318 266976 79324 267028
rect 79376 267016 79382 267028
rect 79376 266988 122834 267016
rect 79376 266976 79382 266988
rect 122806 266880 122834 266988
rect 140130 266976 140136 267028
rect 140188 267016 140194 267028
rect 186958 267016 186964 267028
rect 140188 266988 186964 267016
rect 140188 266976 140194 266988
rect 186958 266976 186964 266988
rect 187016 266976 187022 267028
rect 190454 266976 190460 267028
rect 190512 267016 190518 267028
rect 224218 267016 224224 267028
rect 190512 266988 224224 267016
rect 190512 266976 190518 266988
rect 224218 266976 224224 266988
rect 224276 266976 224282 267028
rect 228358 266976 228364 267028
rect 228416 267016 228422 267028
rect 228416 266988 238754 267016
rect 228416 266976 228422 266988
rect 140590 266880 140596 266892
rect 122806 266852 140596 266880
rect 140590 266840 140596 266852
rect 140648 266840 140654 266892
rect 150526 266880 150532 266892
rect 140792 266852 150532 266880
rect 137462 266704 137468 266756
rect 137520 266744 137526 266756
rect 140792 266744 140820 266852
rect 150526 266840 150532 266852
rect 150584 266840 150590 266892
rect 159450 266840 159456 266892
rect 159508 266880 159514 266892
rect 162118 266880 162124 266892
rect 159508 266852 162124 266880
rect 159508 266840 159514 266852
rect 162118 266840 162124 266852
rect 162176 266840 162182 266892
rect 178862 266840 178868 266892
rect 178920 266880 178926 266892
rect 209314 266880 209320 266892
rect 178920 266852 209320 266880
rect 178920 266840 178926 266852
rect 209314 266840 209320 266852
rect 209372 266840 209378 266892
rect 218698 266840 218704 266892
rect 218756 266880 218762 266892
rect 220906 266880 220912 266892
rect 218756 266852 220912 266880
rect 218756 266840 218762 266852
rect 220906 266840 220912 266852
rect 220964 266840 220970 266892
rect 238726 266880 238754 266988
rect 249058 266976 249064 267028
rect 249116 267016 249122 267028
rect 250714 267016 250720 267028
rect 249116 266988 250720 267016
rect 249116 266976 249122 266988
rect 250714 266976 250720 266988
rect 250772 266976 250778 267028
rect 255958 266976 255964 267028
rect 256016 267016 256022 267028
rect 258994 267016 259000 267028
rect 256016 266988 259000 267016
rect 256016 266976 256022 266988
rect 258994 266976 259000 266988
rect 259052 266976 259058 267028
rect 286318 266976 286324 267028
rect 286376 267016 286382 267028
rect 287974 267016 287980 267028
rect 286376 266988 287980 267016
rect 286376 266976 286382 266988
rect 287974 266976 287980 266988
rect 288032 266976 288038 267028
rect 314470 266976 314476 267028
rect 314528 267016 314534 267028
rect 318978 267016 318984 267028
rect 314528 266988 318984 267016
rect 314528 266976 314534 266988
rect 318978 266976 318984 266988
rect 319036 266976 319042 267028
rect 353386 266976 353392 267028
rect 353444 267016 353450 267028
rect 369320 267016 369348 267396
rect 374454 267384 374460 267396
rect 374512 267384 374518 267436
rect 380710 267384 380716 267436
rect 380768 267424 380774 267436
rect 398742 267424 398748 267436
rect 380768 267396 398748 267424
rect 380768 267384 380774 267396
rect 398742 267384 398748 267396
rect 398800 267384 398806 267436
rect 403066 267384 403072 267436
rect 403124 267424 403130 267436
rect 422294 267424 422300 267436
rect 403124 267396 422300 267424
rect 403124 267384 403130 267396
rect 422294 267384 422300 267396
rect 422352 267384 422358 267436
rect 428734 267384 428740 267436
rect 428792 267424 428798 267436
rect 447594 267424 447600 267436
rect 428792 267396 447600 267424
rect 428792 267384 428798 267396
rect 447594 267384 447600 267396
rect 447652 267384 447658 267436
rect 450262 267384 450268 267436
rect 450320 267424 450326 267436
rect 498838 267424 498844 267436
rect 450320 267396 498844 267424
rect 450320 267384 450326 267396
rect 498838 267384 498844 267396
rect 498896 267384 498902 267436
rect 514846 267384 514852 267436
rect 514904 267424 514910 267436
rect 578878 267424 578884 267436
rect 514904 267396 578884 267424
rect 514904 267384 514910 267396
rect 578878 267384 578884 267396
rect 578936 267384 578942 267436
rect 373258 267248 373264 267300
rect 373316 267288 373322 267300
rect 392026 267288 392032 267300
rect 373316 267260 392032 267288
rect 373316 267248 373322 267260
rect 392026 267248 392032 267260
rect 392084 267248 392090 267300
rect 398098 267248 398104 267300
rect 398156 267288 398162 267300
rect 417418 267288 417424 267300
rect 398156 267260 417424 267288
rect 398156 267248 398162 267260
rect 417418 267248 417424 267260
rect 417476 267248 417482 267300
rect 436738 267248 436744 267300
rect 436796 267288 436802 267300
rect 457438 267288 457444 267300
rect 436796 267260 457444 267288
rect 436796 267248 436802 267260
rect 457438 267248 457444 267260
rect 457496 267248 457502 267300
rect 459370 267248 459376 267300
rect 459428 267288 459434 267300
rect 460842 267288 460848 267300
rect 459428 267260 460848 267288
rect 459428 267248 459434 267260
rect 460842 267248 460848 267260
rect 460900 267248 460906 267300
rect 465166 267248 465172 267300
rect 465224 267288 465230 267300
rect 523678 267288 523684 267300
rect 465224 267260 523684 267288
rect 465224 267248 465230 267260
rect 523678 267248 523684 267260
rect 523736 267248 523742 267300
rect 524782 267248 524788 267300
rect 524840 267288 524846 267300
rect 611998 267288 612004 267300
rect 524840 267260 612004 267288
rect 524840 267248 524846 267260
rect 611998 267248 612004 267260
rect 612056 267248 612062 267300
rect 385678 267152 385684 267164
rect 353444 266988 369348 267016
rect 373966 267124 385684 267152
rect 353444 266976 353450 266988
rect 249058 266880 249064 266892
rect 238726 266852 249064 266880
rect 249058 266840 249064 266852
rect 249116 266840 249122 266892
rect 332686 266840 332692 266892
rect 332744 266880 332750 266892
rect 343818 266880 343824 266892
rect 332744 266852 343824 266880
rect 332744 266840 332750 266852
rect 343818 266840 343824 266852
rect 343876 266840 343882 266892
rect 368290 266840 368296 266892
rect 368348 266880 368354 266892
rect 373966 266880 373994 267124
rect 385678 267112 385684 267124
rect 385736 267112 385742 267164
rect 393130 267112 393136 267164
rect 393188 267152 393194 267164
rect 420178 267152 420184 267164
rect 393188 267124 420184 267152
rect 393188 267112 393194 267124
rect 420178 267112 420184 267124
rect 420236 267112 420242 267164
rect 432874 267112 432880 267164
rect 432932 267152 432938 267164
rect 453298 267152 453304 267164
rect 432932 267124 453304 267152
rect 432932 267112 432938 267124
rect 453298 267112 453304 267124
rect 453356 267112 453362 267164
rect 455138 267112 455144 267164
rect 455196 267152 455202 267164
rect 515398 267152 515404 267164
rect 455196 267124 515404 267152
rect 455196 267112 455202 267124
rect 515398 267112 515404 267124
rect 515456 267112 515462 267164
rect 517238 267112 517244 267164
rect 517296 267152 517302 267164
rect 527174 267152 527180 267164
rect 517296 267124 527180 267152
rect 517296 267112 517302 267124
rect 527174 267112 527180 267124
rect 527232 267112 527238 267164
rect 529658 267112 529664 267164
rect 529716 267152 529722 267164
rect 617518 267152 617524 267164
rect 529716 267124 617524 267152
rect 529716 267112 529722 267124
rect 617518 267112 617524 267124
rect 617576 267112 617582 267164
rect 383194 266976 383200 267028
rect 383252 267016 383258 267028
rect 401686 267016 401692 267028
rect 383252 266988 401692 267016
rect 383252 266976 383258 266988
rect 401686 266976 401692 266988
rect 401744 266976 401750 267028
rect 413002 266976 413008 267028
rect 413060 267016 413066 267028
rect 413060 266988 441614 267016
rect 413060 266976 413066 266988
rect 441586 266892 441614 266988
rect 470134 266976 470140 267028
rect 470192 267016 470198 267028
rect 534718 267016 534724 267028
rect 470192 266988 534724 267016
rect 470192 266976 470198 266988
rect 534718 266976 534724 266988
rect 534776 266976 534782 267028
rect 535546 266976 535552 267028
rect 535604 267016 535610 267028
rect 536742 267016 536748 267028
rect 535604 266988 536748 267016
rect 535604 266976 535610 266988
rect 536742 266976 536748 266988
rect 536800 266976 536806 267028
rect 539686 266976 539692 267028
rect 539744 267016 539750 267028
rect 634078 267016 634084 267028
rect 539744 266988 634084 267016
rect 539744 266976 539750 266988
rect 634078 266976 634084 266988
rect 634136 266976 634142 267028
rect 368348 266852 373994 266880
rect 368348 266840 368354 266852
rect 378226 266840 378232 266892
rect 378284 266880 378290 266892
rect 394694 266880 394700 266892
rect 378284 266852 394700 266880
rect 378284 266840 378290 266852
rect 394694 266840 394700 266852
rect 394752 266840 394758 266892
rect 404722 266840 404728 266892
rect 404780 266880 404786 266892
rect 416222 266880 416228 266892
rect 404780 266852 416228 266880
rect 404780 266840 404786 266852
rect 416222 266840 416228 266852
rect 416280 266840 416286 266892
rect 422938 266840 422944 266892
rect 422996 266880 423002 266892
rect 438118 266880 438124 266892
rect 422996 266852 438124 266880
rect 422996 266840 423002 266852
rect 438118 266840 438124 266852
rect 438176 266840 438182 266892
rect 441586 266852 441620 266892
rect 441614 266840 441620 266852
rect 441672 266840 441678 266892
rect 442718 266840 442724 266892
rect 442776 266880 442782 266892
rect 485038 266880 485044 266892
rect 442776 266852 485044 266880
rect 442776 266840 442782 266852
rect 485038 266840 485044 266852
rect 485096 266840 485102 266892
rect 499942 266840 499948 266892
rect 500000 266880 500006 266892
rect 507854 266880 507860 266892
rect 500000 266852 507860 266880
rect 500000 266840 500006 266852
rect 507854 266840 507860 266852
rect 507912 266840 507918 266892
rect 534718 266840 534724 266892
rect 534776 266880 534782 266892
rect 589918 266880 589924 266892
rect 534776 266852 589924 266880
rect 534776 266840 534782 266852
rect 589918 266840 589924 266852
rect 589976 266840 589982 266892
rect 316954 266772 316960 266824
rect 317012 266812 317018 266824
rect 321554 266812 321560 266824
rect 317012 266784 321560 266812
rect 317012 266772 317018 266784
rect 321554 266772 321560 266784
rect 321612 266772 321618 266824
rect 137520 266716 140820 266744
rect 137520 266704 137526 266716
rect 151078 266704 151084 266756
rect 151136 266744 151142 266756
rect 179506 266744 179512 266756
rect 151136 266716 179512 266744
rect 151136 266704 151142 266716
rect 179506 266704 179512 266716
rect 179564 266704 179570 266756
rect 394786 266704 394792 266756
rect 394844 266744 394850 266756
rect 403618 266744 403624 266756
rect 394844 266716 403624 266744
rect 394844 266704 394850 266716
rect 403618 266704 403624 266716
rect 403676 266704 403682 266756
rect 407206 266704 407212 266756
rect 407264 266744 407270 266756
rect 414658 266744 414664 266756
rect 407264 266716 414664 266744
rect 407264 266704 407270 266716
rect 414658 266704 414664 266716
rect 414716 266704 414722 266756
rect 449158 266744 449164 266756
rect 441586 266716 449164 266744
rect 308674 266636 308680 266688
rect 308732 266676 308738 266688
rect 310514 266676 310520 266688
rect 308732 266648 310520 266676
rect 308732 266636 308738 266648
rect 310514 266636 310520 266648
rect 310572 266636 310578 266688
rect 313642 266636 313648 266688
rect 313700 266676 313706 266688
rect 317414 266676 317420 266688
rect 313700 266648 317420 266676
rect 313700 266636 313706 266648
rect 317414 266636 317420 266648
rect 317472 266636 317478 266688
rect 317782 266636 317788 266688
rect 317840 266676 317846 266688
rect 322934 266676 322940 266688
rect 317840 266648 322940 266676
rect 317840 266636 317846 266648
rect 322934 266636 322940 266648
rect 322992 266636 322998 266688
rect 347498 266636 347504 266688
rect 347556 266676 347562 266688
rect 351178 266676 351184 266688
rect 347556 266648 351184 266676
rect 347556 266636 347562 266648
rect 351178 266636 351184 266648
rect 351236 266636 351242 266688
rect 427906 266636 427912 266688
rect 427964 266676 427970 266688
rect 436738 266676 436744 266688
rect 427964 266648 436744 266676
rect 427964 266636 427970 266648
rect 436738 266636 436744 266648
rect 436796 266636 436802 266688
rect 441586 266676 441614 266716
rect 449158 266704 449164 266716
rect 449216 266704 449222 266756
rect 457714 266704 457720 266756
rect 457772 266744 457778 266756
rect 476758 266744 476764 266756
rect 457772 266716 476764 266744
rect 457772 266704 457778 266716
rect 476758 266704 476764 266716
rect 476816 266704 476822 266756
rect 485038 266704 485044 266756
rect 485096 266744 485102 266756
rect 485096 266716 489914 266744
rect 485096 266704 485102 266716
rect 436940 266648 441614 266676
rect 130378 266568 130384 266620
rect 130436 266608 130442 266620
rect 138106 266608 138112 266620
rect 130436 266580 138112 266608
rect 130436 266568 130442 266580
rect 138106 266568 138112 266580
rect 138164 266568 138170 266620
rect 149606 266568 149612 266620
rect 149664 266608 149670 266620
rect 159634 266608 159640 266620
rect 149664 266580 159640 266608
rect 149664 266568 149670 266580
rect 159634 266568 159640 266580
rect 159692 266568 159698 266620
rect 399754 266568 399760 266620
rect 399812 266608 399818 266620
rect 407758 266608 407764 266620
rect 399812 266580 407764 266608
rect 399812 266568 399818 266580
rect 407758 266568 407764 266580
rect 407816 266568 407822 266620
rect 310330 266500 310336 266552
rect 310388 266540 310394 266552
rect 311894 266540 311900 266552
rect 310388 266512 311900 266540
rect 310388 266500 310394 266512
rect 311894 266500 311900 266512
rect 311952 266500 311958 266552
rect 312262 266500 312268 266552
rect 312320 266540 312326 266552
rect 314654 266540 314660 266552
rect 312320 266512 314660 266540
rect 312320 266500 312326 266512
rect 314654 266500 314660 266512
rect 314712 266500 314718 266552
rect 316126 266500 316132 266552
rect 316184 266540 316190 266552
rect 320174 266540 320180 266552
rect 316184 266512 320180 266540
rect 316184 266500 316190 266512
rect 320174 266500 320180 266512
rect 320232 266500 320238 266552
rect 327718 266500 327724 266552
rect 327776 266540 327782 266552
rect 331858 266540 331864 266552
rect 327776 266512 331864 266540
rect 327776 266500 327782 266512
rect 331858 266500 331864 266512
rect 331916 266500 331922 266552
rect 345106 266500 345112 266552
rect 345164 266540 345170 266552
rect 348418 266540 348424 266552
rect 345164 266512 348424 266540
rect 345164 266500 345170 266512
rect 348418 266500 348424 266512
rect 348476 266500 348482 266552
rect 350074 266500 350080 266552
rect 350132 266540 350138 266552
rect 353938 266540 353944 266552
rect 350132 266512 353944 266540
rect 350132 266500 350138 266512
rect 353938 266500 353944 266512
rect 353996 266500 354002 266552
rect 355870 266500 355876 266552
rect 355928 266540 355934 266552
rect 360838 266540 360844 266552
rect 355928 266512 360844 266540
rect 355928 266500 355934 266512
rect 360838 266500 360844 266512
rect 360896 266500 360902 266552
rect 369946 266500 369952 266552
rect 370004 266540 370010 266552
rect 372246 266540 372252 266552
rect 370004 266512 372252 266540
rect 370004 266500 370010 266512
rect 372246 266500 372252 266512
rect 372304 266500 372310 266552
rect 374914 266500 374920 266552
rect 374972 266540 374978 266552
rect 379698 266540 379704 266552
rect 374972 266512 379704 266540
rect 374972 266500 374978 266512
rect 379698 266500 379704 266512
rect 379756 266500 379762 266552
rect 423766 266500 423772 266552
rect 423824 266540 423830 266552
rect 425698 266540 425704 266552
rect 423824 266512 425704 266540
rect 423824 266500 423830 266512
rect 425698 266500 425704 266512
rect 425756 266500 425762 266552
rect 426250 266500 426256 266552
rect 426308 266540 426314 266552
rect 428458 266540 428464 266552
rect 426308 266512 428464 266540
rect 426308 266500 426314 266512
rect 428458 266500 428464 266512
rect 428516 266500 428522 266552
rect 434530 266500 434536 266552
rect 434588 266540 434594 266552
rect 436940 266540 436968 266648
rect 452746 266568 452752 266620
rect 452804 266608 452810 266620
rect 462958 266608 462964 266620
rect 452804 266580 462964 266608
rect 452804 266568 452810 266580
rect 462958 266568 462964 266580
rect 463016 266568 463022 266620
rect 489886 266608 489914 266716
rect 490006 266704 490012 266756
rect 490064 266744 490070 266756
rect 509694 266744 509700 266756
rect 490064 266716 509700 266744
rect 490064 266704 490070 266716
rect 509694 266704 509700 266716
rect 509752 266704 509758 266756
rect 510706 266704 510712 266756
rect 510764 266744 510770 266756
rect 511810 266744 511816 266756
rect 510764 266716 511816 266744
rect 510764 266704 510770 266716
rect 511810 266704 511816 266716
rect 511868 266704 511874 266756
rect 512362 266704 512368 266756
rect 512420 266744 512426 266756
rect 513190 266744 513196 266756
rect 512420 266716 513196 266744
rect 512420 266704 512426 266716
rect 513190 266704 513196 266716
rect 513248 266704 513254 266756
rect 516502 266704 516508 266756
rect 516560 266744 516566 266756
rect 517422 266744 517428 266756
rect 516560 266716 517428 266744
rect 516560 266704 516566 266716
rect 517422 266704 517428 266716
rect 517480 266704 517486 266756
rect 518986 266704 518992 266756
rect 519044 266744 519050 266756
rect 520090 266744 520096 266756
rect 519044 266716 520096 266744
rect 519044 266704 519050 266716
rect 520090 266704 520096 266716
rect 520148 266704 520154 266756
rect 527266 266704 527272 266756
rect 527324 266744 527330 266756
rect 528186 266744 528192 266756
rect 527324 266716 528192 266744
rect 527324 266704 527330 266716
rect 528186 266704 528192 266716
rect 528244 266704 528250 266756
rect 528922 266704 528928 266756
rect 528980 266744 528986 266756
rect 529842 266744 529848 266756
rect 528980 266716 529848 266744
rect 528980 266704 528986 266716
rect 529842 266704 529848 266716
rect 529900 266704 529906 266756
rect 531406 266704 531412 266756
rect 531464 266744 531470 266756
rect 532510 266744 532516 266756
rect 531464 266716 532516 266744
rect 531464 266704 531470 266716
rect 532510 266704 532516 266716
rect 532568 266704 532574 266756
rect 533062 266704 533068 266756
rect 533120 266744 533126 266756
rect 533982 266744 533988 266756
rect 533120 266716 533988 266744
rect 533120 266704 533126 266716
rect 533982 266704 533988 266716
rect 534040 266704 534046 266756
rect 542998 266704 543004 266756
rect 543056 266744 543062 266756
rect 598198 266744 598204 266756
rect 543056 266716 598204 266744
rect 543056 266704 543062 266716
rect 598198 266704 598204 266716
rect 598256 266704 598262 266756
rect 501598 266608 501604 266620
rect 489886 266580 501604 266608
rect 501598 266568 501604 266580
rect 501656 266568 501662 266620
rect 504818 266568 504824 266620
rect 504876 266608 504882 266620
rect 556798 266608 556804 266620
rect 504876 266580 556804 266608
rect 504876 266568 504882 266580
rect 556798 266568 556804 266580
rect 556856 266568 556862 266620
rect 434588 266512 436968 266540
rect 434588 266500 434594 266512
rect 437842 266500 437848 266552
rect 437900 266540 437906 266552
rect 448422 266540 448428 266552
rect 437900 266512 448428 266540
rect 437900 266500 437906 266512
rect 448422 266500 448428 266512
rect 448480 266500 448486 266552
rect 132494 266432 132500 266484
rect 132552 266472 132558 266484
rect 147214 266472 147220 266484
rect 132552 266444 147220 266472
rect 132552 266432 132558 266444
rect 147214 266432 147220 266444
rect 147272 266432 147278 266484
rect 491662 266432 491668 266484
rect 491720 266472 491726 266484
rect 492582 266472 492588 266484
rect 491720 266444 492588 266472
rect 491720 266432 491726 266444
rect 492582 266432 492588 266444
rect 492640 266432 492646 266484
rect 494146 266432 494152 266484
rect 494204 266472 494210 266484
rect 495066 266472 495072 266484
rect 494204 266444 495072 266472
rect 494204 266432 494210 266444
rect 495066 266432 495072 266444
rect 495124 266432 495130 266484
rect 502426 266432 502432 266484
rect 502484 266472 502490 266484
rect 503438 266472 503444 266484
rect 502484 266444 503444 266472
rect 502484 266432 502490 266444
rect 503438 266432 503444 266444
rect 503496 266432 503502 266484
rect 504082 266432 504088 266484
rect 504140 266472 504146 266484
rect 505002 266472 505008 266484
rect 504140 266444 505008 266472
rect 504140 266432 504146 266444
rect 505002 266432 505008 266444
rect 505060 266432 505066 266484
rect 506566 266432 506572 266484
rect 506624 266472 506630 266484
rect 507670 266472 507676 266484
rect 506624 266444 507676 266472
rect 506624 266432 506630 266444
rect 507670 266432 507676 266444
rect 507728 266432 507734 266484
rect 507854 266432 507860 266484
rect 507912 266472 507918 266484
rect 549898 266472 549904 266484
rect 507912 266444 549904 266472
rect 507912 266432 507918 266444
rect 549898 266432 549904 266444
rect 549956 266432 549962 266484
rect 163498 266364 163504 266416
rect 163556 266404 163562 266416
rect 167086 266404 167092 266416
rect 163556 266376 167092 266404
rect 163556 266364 163562 266376
rect 167086 266364 167092 266376
rect 167144 266364 167150 266416
rect 168558 266364 168564 266416
rect 168616 266404 168622 266416
rect 169570 266404 169576 266416
rect 168616 266376 169576 266404
rect 168616 266364 168622 266376
rect 169570 266364 169576 266376
rect 169628 266364 169634 266416
rect 211154 266364 211160 266416
rect 211212 266404 211218 266416
rect 213454 266404 213460 266416
rect 211212 266376 213460 266404
rect 211212 266364 211218 266376
rect 213454 266364 213460 266376
rect 213512 266364 213518 266416
rect 214558 266364 214564 266416
rect 214616 266404 214622 266416
rect 215938 266404 215944 266416
rect 214616 266376 215944 266404
rect 214616 266364 214622 266376
rect 215938 266364 215944 266376
rect 215996 266364 216002 266416
rect 239398 266364 239404 266416
rect 239456 266404 239462 266416
rect 241606 266404 241612 266416
rect 239456 266376 241612 266404
rect 239456 266364 239462 266376
rect 241606 266364 241612 266376
rect 241664 266364 241670 266416
rect 243722 266364 243728 266416
rect 243780 266404 243786 266416
rect 246574 266404 246580 266416
rect 243780 266376 246580 266404
rect 243780 266364 243786 266376
rect 246574 266364 246580 266376
rect 246632 266364 246638 266416
rect 250438 266364 250444 266416
rect 250496 266404 250502 266416
rect 256510 266404 256516 266416
rect 250496 266376 256516 266404
rect 250496 266364 250502 266376
rect 256510 266364 256516 266376
rect 256568 266364 256574 266416
rect 300946 266364 300952 266416
rect 301004 266404 301010 266416
rect 302050 266404 302056 266416
rect 301004 266376 302056 266404
rect 301004 266364 301010 266376
rect 302050 266364 302056 266376
rect 302108 266364 302114 266416
rect 303706 266364 303712 266416
rect 303764 266404 303770 266416
rect 304534 266404 304540 266416
rect 303764 266376 304540 266404
rect 303764 266364 303770 266376
rect 304534 266364 304540 266376
rect 304592 266364 304598 266416
rect 307846 266364 307852 266416
rect 307904 266404 307910 266416
rect 309134 266404 309140 266416
rect 307904 266376 309140 266404
rect 307904 266364 307910 266376
rect 309134 266364 309140 266376
rect 309192 266364 309198 266416
rect 309502 266364 309508 266416
rect 309560 266404 309566 266416
rect 310698 266404 310704 266416
rect 309560 266376 310704 266404
rect 309560 266364 309566 266376
rect 310698 266364 310704 266376
rect 310756 266364 310762 266416
rect 311158 266364 311164 266416
rect 311216 266404 311222 266416
rect 313274 266404 313280 266416
rect 311216 266376 313280 266404
rect 311216 266364 311222 266376
rect 313274 266364 313280 266376
rect 313332 266364 313338 266416
rect 320266 266364 320272 266416
rect 320324 266404 320330 266416
rect 321370 266404 321376 266416
rect 320324 266376 321376 266404
rect 320324 266364 320330 266376
rect 321370 266364 321376 266376
rect 321428 266364 321434 266416
rect 324406 266364 324412 266416
rect 324464 266404 324470 266416
rect 325326 266404 325332 266416
rect 324464 266376 325332 266404
rect 324464 266364 324470 266376
rect 325326 266364 325332 266376
rect 325384 266364 325390 266416
rect 328546 266364 328552 266416
rect 328604 266404 328610 266416
rect 329742 266404 329748 266416
rect 328604 266376 329748 266404
rect 328604 266364 328610 266376
rect 329742 266364 329748 266376
rect 329800 266364 329806 266416
rect 336826 266364 336832 266416
rect 336884 266404 336890 266416
rect 337930 266404 337936 266416
rect 336884 266376 337936 266404
rect 336884 266364 336890 266376
rect 337930 266364 337936 266376
rect 337988 266364 337994 266416
rect 342622 266364 342628 266416
rect 342680 266404 342686 266416
rect 345290 266404 345296 266416
rect 342680 266376 345296 266404
rect 342680 266364 342686 266376
rect 345290 266364 345296 266376
rect 345348 266364 345354 266416
rect 346762 266364 346768 266416
rect 346820 266404 346826 266416
rect 347682 266404 347688 266416
rect 346820 266376 347688 266404
rect 346820 266364 346826 266376
rect 347682 266364 347688 266376
rect 347740 266364 347746 266416
rect 349246 266364 349252 266416
rect 349304 266404 349310 266416
rect 350350 266404 350356 266416
rect 349304 266376 350356 266404
rect 349304 266364 349310 266376
rect 350350 266364 350356 266376
rect 350408 266364 350414 266416
rect 357526 266364 357532 266416
rect 357584 266404 357590 266416
rect 359458 266404 359464 266416
rect 357584 266376 359464 266404
rect 357584 266364 357590 266376
rect 359458 266364 359464 266376
rect 359516 266364 359522 266416
rect 361666 266364 361672 266416
rect 361724 266404 361730 266416
rect 362770 266404 362776 266416
rect 361724 266376 362776 266404
rect 361724 266364 361730 266376
rect 362770 266364 362776 266376
rect 362828 266364 362834 266416
rect 369118 266364 369124 266416
rect 369176 266404 369182 266416
rect 370498 266404 370504 266416
rect 369176 266376 370504 266404
rect 369176 266364 369182 266376
rect 370498 266364 370504 266376
rect 370556 266364 370562 266416
rect 374086 266364 374092 266416
rect 374144 266404 374150 266416
rect 375282 266404 375288 266416
rect 374144 266376 375288 266404
rect 374144 266364 374150 266376
rect 375282 266364 375288 266376
rect 375340 266364 375346 266416
rect 379882 266364 379888 266416
rect 379940 266404 379946 266416
rect 383010 266404 383016 266416
rect 379940 266376 383016 266404
rect 379940 266364 379946 266376
rect 383010 266364 383016 266376
rect 383068 266364 383074 266416
rect 384022 266364 384028 266416
rect 384080 266404 384086 266416
rect 384942 266404 384948 266416
rect 384080 266376 384948 266404
rect 384080 266364 384086 266376
rect 384942 266364 384948 266376
rect 385000 266364 385006 266416
rect 386506 266364 386512 266416
rect 386564 266404 386570 266416
rect 387702 266404 387708 266416
rect 386564 266376 387708 266404
rect 386564 266364 386570 266376
rect 387702 266364 387708 266376
rect 387760 266364 387766 266416
rect 392302 266364 392308 266416
rect 392360 266404 392366 266416
rect 393682 266404 393688 266416
rect 392360 266376 393688 266404
rect 392360 266364 392366 266376
rect 393682 266364 393688 266376
rect 393740 266364 393746 266416
rect 398926 266364 398932 266416
rect 398984 266404 398990 266416
rect 400030 266404 400036 266416
rect 398984 266376 400036 266404
rect 398984 266364 398990 266376
rect 400030 266364 400036 266376
rect 400088 266364 400094 266416
rect 408862 266364 408868 266416
rect 408920 266404 408926 266416
rect 409782 266404 409788 266416
rect 408920 266376 409788 266404
rect 408920 266364 408926 266376
rect 409782 266364 409788 266376
rect 409840 266364 409846 266416
rect 411346 266364 411352 266416
rect 411404 266404 411410 266416
rect 412266 266404 412272 266416
rect 411404 266376 412272 266404
rect 411404 266364 411410 266376
rect 412266 266364 412272 266376
rect 412324 266364 412330 266416
rect 415486 266364 415492 266416
rect 415544 266404 415550 266416
rect 416406 266404 416412 266416
rect 415544 266376 416412 266404
rect 415544 266364 415550 266376
rect 416406 266364 416412 266376
rect 416464 266364 416470 266416
rect 417970 266364 417976 266416
rect 418028 266404 418034 266416
rect 418798 266404 418804 266416
rect 418028 266376 418804 266404
rect 418028 266364 418034 266376
rect 418798 266364 418804 266376
rect 418856 266364 418862 266416
rect 425422 266364 425428 266416
rect 425480 266404 425486 266416
rect 427078 266404 427084 266416
rect 425480 266376 427084 266404
rect 425480 266364 425486 266376
rect 427078 266364 427084 266376
rect 427136 266364 427142 266416
rect 429562 266364 429568 266416
rect 429620 266404 429626 266416
rect 430390 266404 430396 266416
rect 429620 266376 430396 266404
rect 429620 266364 429626 266376
rect 430390 266364 430396 266376
rect 430448 266364 430454 266416
rect 432046 266364 432052 266416
rect 432104 266404 432110 266416
rect 433150 266404 433156 266416
rect 432104 266376 433156 266404
rect 432104 266364 432110 266376
rect 433150 266364 433156 266376
rect 433208 266364 433214 266416
rect 440326 266364 440332 266416
rect 440384 266404 440390 266416
rect 441338 266404 441344 266416
rect 440384 266376 441344 266404
rect 440384 266364 440390 266376
rect 441338 266364 441344 266376
rect 441396 266364 441402 266416
rect 441982 266364 441988 266416
rect 442040 266404 442046 266416
rect 442902 266404 442908 266416
rect 442040 266376 442908 266404
rect 442040 266364 442046 266376
rect 442902 266364 442908 266376
rect 442960 266364 442966 266416
rect 444466 266364 444472 266416
rect 444524 266404 444530 266416
rect 445662 266404 445668 266416
rect 444524 266376 445668 266404
rect 444524 266364 444530 266376
rect 445662 266364 445668 266376
rect 445720 266364 445726 266416
rect 448606 266364 448612 266416
rect 448664 266404 448670 266416
rect 450538 266404 450544 266416
rect 448664 266376 450544 266404
rect 448664 266364 448670 266376
rect 450538 266364 450544 266376
rect 450596 266364 450602 266416
rect 454402 266364 454408 266416
rect 454460 266404 454466 266416
rect 455322 266404 455328 266416
rect 454460 266376 455328 266404
rect 454460 266364 454466 266376
rect 455322 266364 455328 266376
rect 455380 266364 455386 266416
rect 473446 266364 473452 266416
rect 473504 266404 473510 266416
rect 474642 266404 474648 266416
rect 473504 266376 474648 266404
rect 473504 266364 473510 266376
rect 474642 266364 474648 266376
rect 474700 266364 474706 266416
rect 475102 266364 475108 266416
rect 475160 266404 475166 266416
rect 479518 266404 479524 266416
rect 475160 266376 479524 266404
rect 475160 266364 475166 266376
rect 479518 266364 479524 266376
rect 479576 266364 479582 266416
rect 481726 266364 481732 266416
rect 481784 266404 481790 266416
rect 482830 266404 482836 266416
rect 481784 266376 482836 266404
rect 481784 266364 481790 266376
rect 482830 266364 482836 266376
rect 482888 266364 482894 266416
rect 483382 266364 483388 266416
rect 483440 266404 483446 266416
rect 484210 266404 484216 266416
rect 483440 266376 484216 266404
rect 483440 266364 483446 266376
rect 484210 266364 484216 266376
rect 484268 266364 484274 266416
rect 485866 266364 485872 266416
rect 485924 266404 485930 266416
rect 486786 266404 486792 266416
rect 485924 266376 486792 266404
rect 485924 266364 485930 266376
rect 486786 266364 486792 266376
rect 486844 266364 486850 266416
rect 487154 266296 487160 266348
rect 487212 266336 487218 266348
rect 557718 266336 557724 266348
rect 487212 266308 557724 266336
rect 487212 266296 487218 266308
rect 557718 266296 557724 266308
rect 557776 266296 557782 266348
rect 484210 266160 484216 266212
rect 484268 266200 484274 266212
rect 560294 266200 560300 266212
rect 484268 266172 560300 266200
rect 484268 266160 484274 266172
rect 560294 266160 560300 266172
rect 560352 266160 560358 266212
rect 482554 266024 482560 266076
rect 482612 266064 482618 266076
rect 487154 266064 487160 266076
rect 482612 266036 487160 266064
rect 482612 266024 482618 266036
rect 487154 266024 487160 266036
rect 487212 266024 487218 266076
rect 492490 266024 492496 266076
rect 492548 266064 492554 266076
rect 572714 266064 572720 266076
rect 492548 266036 572720 266064
rect 492548 266024 492554 266036
rect 572714 266024 572720 266036
rect 572772 266024 572778 266076
rect 513190 265888 513196 265940
rect 513248 265928 513254 265940
rect 601694 265928 601700 265940
rect 513248 265900 601700 265928
rect 513248 265888 513254 265900
rect 601694 265888 601700 265900
rect 601752 265888 601758 265940
rect 515674 265752 515680 265804
rect 515732 265792 515738 265804
rect 605834 265792 605840 265804
rect 515732 265764 605840 265792
rect 515732 265752 515738 265764
rect 605834 265752 605840 265764
rect 605892 265752 605898 265804
rect 189074 265616 189080 265668
rect 189132 265656 189138 265668
rect 189902 265656 189908 265668
rect 189132 265628 189908 265656
rect 189132 265616 189138 265628
rect 189902 265616 189908 265628
rect 189960 265616 189966 265668
rect 209774 265616 209780 265668
rect 209832 265656 209838 265668
rect 210694 265656 210700 265668
rect 209832 265628 210700 265656
rect 209832 265616 209838 265628
rect 210694 265616 210700 265628
rect 210752 265616 210758 265668
rect 224954 265616 224960 265668
rect 225012 265656 225018 265668
rect 225598 265656 225604 265668
rect 225012 265628 225604 265656
rect 225012 265616 225018 265628
rect 225598 265616 225604 265628
rect 225656 265616 225662 265668
rect 280338 265616 280344 265668
rect 280396 265656 280402 265668
rect 280982 265656 280988 265668
rect 280396 265628 280988 265656
rect 280396 265616 280402 265628
rect 280982 265616 280988 265628
rect 281040 265616 281046 265668
rect 292666 265616 292672 265668
rect 292724 265656 292730 265668
rect 293494 265656 293500 265668
rect 292724 265628 293500 265656
rect 292724 265616 292730 265628
rect 293494 265616 293500 265628
rect 293552 265616 293558 265668
rect 296806 265616 296812 265668
rect 296864 265656 296870 265668
rect 297542 265656 297548 265668
rect 296864 265628 297548 265656
rect 296864 265616 296870 265628
rect 297542 265616 297548 265628
rect 297600 265616 297606 265668
rect 520642 265616 520648 265668
rect 520700 265656 520706 265668
rect 612734 265656 612740 265668
rect 520700 265628 612740 265656
rect 520700 265616 520706 265628
rect 612734 265616 612740 265628
rect 612792 265616 612798 265668
rect 479242 265480 479248 265532
rect 479300 265520 479306 265532
rect 553394 265520 553400 265532
rect 479300 265492 553400 265520
rect 479300 265480 479306 265492
rect 553394 265480 553400 265492
rect 553452 265480 553458 265532
rect 477586 265344 477592 265396
rect 477644 265384 477650 265396
rect 550634 265384 550640 265396
rect 477644 265356 550640 265384
rect 477644 265344 477650 265356
rect 550634 265344 550640 265356
rect 550692 265344 550698 265396
rect 469306 265208 469312 265260
rect 469364 265248 469370 265260
rect 539962 265248 539968 265260
rect 469364 265220 539968 265248
rect 469364 265208 469370 265220
rect 539962 265208 539968 265220
rect 540020 265208 540026 265260
rect 466822 265072 466828 265124
rect 466880 265112 466886 265124
rect 535730 265112 535736 265124
rect 466880 265084 535736 265112
rect 466880 265072 466886 265084
rect 535730 265072 535736 265084
rect 535788 265072 535794 265124
rect 58618 264324 58624 264376
rect 58676 264364 58682 264376
rect 668118 264364 668124 264376
rect 58676 264336 668124 264364
rect 58676 264324 58682 264336
rect 668118 264324 668124 264336
rect 668176 264324 668182 264376
rect 46198 264188 46204 264240
rect 46256 264228 46262 264240
rect 669222 264228 669228 264240
rect 46256 264200 669228 264228
rect 46256 264188 46262 264200
rect 669222 264188 669228 264200
rect 669280 264188 669286 264240
rect 570598 261468 570604 261520
rect 570656 261508 570662 261520
rect 645854 261508 645860 261520
rect 570656 261480 645860 261508
rect 570656 261468 570662 261480
rect 645854 261468 645860 261480
rect 645912 261468 645918 261520
rect 554406 260856 554412 260908
rect 554464 260896 554470 260908
rect 568574 260896 568580 260908
rect 554464 260868 568580 260896
rect 554464 260856 554470 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 554314 259428 554320 259480
rect 554372 259468 554378 259480
rect 563698 259468 563704 259480
rect 554372 259440 563704 259468
rect 554372 259428 554378 259440
rect 563698 259428 563704 259440
rect 563756 259428 563762 259480
rect 675846 258748 675852 258800
rect 675904 258788 675910 258800
rect 676398 258788 676404 258800
rect 675904 258760 676404 258788
rect 675904 258748 675910 258760
rect 676398 258748 676404 258760
rect 676456 258748 676462 258800
rect 35802 256912 35808 256964
rect 35860 256952 35866 256964
rect 39482 256952 39488 256964
rect 35860 256924 39488 256952
rect 35860 256912 35866 256924
rect 39482 256912 39488 256924
rect 39540 256912 39546 256964
rect 35618 256708 35624 256760
rect 35676 256748 35682 256760
rect 41690 256748 41696 256760
rect 35676 256720 41696 256748
rect 35676 256708 35682 256720
rect 41690 256708 41696 256720
rect 41748 256708 41754 256760
rect 42058 256708 42064 256760
rect 42116 256748 42122 256760
rect 43346 256748 43352 256760
rect 42116 256720 43352 256748
rect 42116 256708 42122 256720
rect 43346 256708 43352 256720
rect 43404 256708 43410 256760
rect 553946 256708 553952 256760
rect 554004 256748 554010 256760
rect 560938 256748 560944 256760
rect 554004 256720 560944 256748
rect 554004 256708 554010 256720
rect 560938 256708 560944 256720
rect 560996 256708 561002 256760
rect 554498 255552 554504 255604
rect 554556 255592 554562 255604
rect 558178 255592 558184 255604
rect 554556 255564 558184 255592
rect 554556 255552 554562 255564
rect 558178 255552 558184 255564
rect 558236 255552 558242 255604
rect 35802 255416 35808 255468
rect 35860 255456 35866 255468
rect 40218 255456 40224 255468
rect 35860 255428 40224 255456
rect 35860 255416 35866 255428
rect 40218 255416 40224 255428
rect 40276 255416 40282 255468
rect 51718 254532 51724 254584
rect 51776 254572 51782 254584
rect 62390 254572 62396 254584
rect 51776 254544 62396 254572
rect 51776 254532 51782 254544
rect 62390 254532 62396 254544
rect 62448 254532 62454 254584
rect 35618 252696 35624 252748
rect 35676 252736 35682 252748
rect 40678 252736 40684 252748
rect 35676 252708 40684 252736
rect 35676 252696 35682 252708
rect 40678 252696 40684 252708
rect 40736 252696 40742 252748
rect 35802 252560 35808 252612
rect 35860 252600 35866 252612
rect 41322 252600 41328 252612
rect 35860 252572 41328 252600
rect 35860 252560 35866 252572
rect 41322 252560 41328 252572
rect 41380 252560 41386 252612
rect 554406 252560 554412 252612
rect 554464 252600 554470 252612
rect 562318 252600 562324 252612
rect 554464 252572 562324 252600
rect 554464 252560 554470 252572
rect 562318 252560 562324 252572
rect 562376 252560 562382 252612
rect 35802 251200 35808 251252
rect 35860 251240 35866 251252
rect 39298 251240 39304 251252
rect 35860 251212 39304 251240
rect 35860 251200 35866 251212
rect 39298 251200 39304 251212
rect 39356 251200 39362 251252
rect 554130 251200 554136 251252
rect 554188 251240 554194 251252
rect 556798 251240 556804 251252
rect 554188 251212 556804 251240
rect 554188 251200 554194 251212
rect 556798 251200 556804 251212
rect 556856 251200 556862 251252
rect 35618 250044 35624 250096
rect 35676 250084 35682 250096
rect 40126 250084 40132 250096
rect 35676 250056 40132 250084
rect 35676 250044 35682 250056
rect 40126 250044 40132 250056
rect 40184 250044 40190 250096
rect 35802 249772 35808 249824
rect 35860 249812 35866 249824
rect 41690 249812 41696 249824
rect 35860 249784 41696 249812
rect 35860 249772 35866 249784
rect 41690 249772 41696 249784
rect 41748 249772 41754 249824
rect 42058 249772 42064 249824
rect 42116 249812 42122 249824
rect 42978 249812 42984 249824
rect 42116 249784 42984 249812
rect 42116 249772 42122 249784
rect 42978 249772 42984 249784
rect 43036 249772 43042 249824
rect 674926 249704 674932 249756
rect 674984 249744 674990 249756
rect 675478 249744 675484 249756
rect 674984 249716 675484 249744
rect 674984 249704 674990 249716
rect 675478 249704 675484 249716
rect 675536 249704 675542 249756
rect 674926 249160 674932 249212
rect 674984 249160 674990 249212
rect 674944 249076 674972 249160
rect 674926 249024 674932 249076
rect 674984 249024 674990 249076
rect 35802 247256 35808 247308
rect 35860 247296 35866 247308
rect 39850 247296 39856 247308
rect 35860 247268 39856 247296
rect 35860 247256 35866 247268
rect 39850 247256 39856 247268
rect 39908 247256 39914 247308
rect 559558 246304 559564 246356
rect 559616 246344 559622 246356
rect 647234 246344 647240 246356
rect 559616 246316 647240 246344
rect 559616 246304 559622 246316
rect 647234 246304 647240 246316
rect 647292 246304 647298 246356
rect 553854 245624 553860 245676
rect 553912 245664 553918 245676
rect 596818 245664 596824 245676
rect 553912 245636 596824 245664
rect 553912 245624 553918 245636
rect 596818 245624 596824 245636
rect 596876 245624 596882 245676
rect 674834 245420 674840 245472
rect 674892 245460 674898 245472
rect 675202 245460 675208 245472
rect 674892 245432 675208 245460
rect 674892 245420 674898 245432
rect 675202 245420 675208 245432
rect 675260 245420 675266 245472
rect 553486 244264 553492 244316
rect 553544 244304 553550 244316
rect 555418 244304 555424 244316
rect 553544 244276 555424 244304
rect 553544 244264 553550 244276
rect 555418 244264 555424 244276
rect 555476 244264 555482 244316
rect 39298 242700 39304 242752
rect 39356 242740 39362 242752
rect 41690 242740 41696 242752
rect 39356 242712 41696 242740
rect 39356 242700 39362 242712
rect 41690 242700 41696 242712
rect 41748 242700 41754 242752
rect 42058 242632 42064 242684
rect 42116 242672 42122 242684
rect 42518 242672 42524 242684
rect 42116 242644 42524 242672
rect 42116 242632 42122 242644
rect 42518 242632 42524 242644
rect 42576 242632 42582 242684
rect 34422 242156 34428 242208
rect 34480 242196 34486 242208
rect 41690 242196 41696 242208
rect 34480 242168 41696 242196
rect 34480 242156 34486 242168
rect 41690 242156 41696 242168
rect 41748 242156 41754 242208
rect 576118 242156 576124 242208
rect 576176 242196 576182 242208
rect 648614 242196 648620 242208
rect 576176 242168 648620 242196
rect 576176 242156 576182 242168
rect 648614 242156 648620 242168
rect 648672 242156 648678 242208
rect 553670 241476 553676 241528
rect 553728 241516 553734 241528
rect 629938 241516 629944 241528
rect 553728 241488 629944 241516
rect 553728 241476 553734 241488
rect 629938 241476 629944 241488
rect 629996 241476 630002 241528
rect 554498 240116 554504 240168
rect 554556 240156 554562 240168
rect 577498 240156 577504 240168
rect 554556 240128 577504 240156
rect 554556 240116 554562 240128
rect 577498 240116 577504 240128
rect 577556 240116 577562 240168
rect 554314 238688 554320 238740
rect 554372 238728 554378 238740
rect 576118 238728 576124 238740
rect 554372 238700 576124 238728
rect 554372 238688 554378 238700
rect 576118 238688 576124 238700
rect 576176 238688 576182 238740
rect 672258 236988 672264 237040
rect 672316 237028 672322 237040
rect 672756 237028 672784 237082
rect 672316 237000 672784 237028
rect 672316 236988 672322 237000
rect 671246 236852 671252 236904
rect 671304 236892 671310 236904
rect 671304 236864 672888 236892
rect 671304 236852 671310 236864
rect 553762 236784 553768 236836
rect 553820 236824 553826 236836
rect 559558 236824 559564 236836
rect 553820 236796 559564 236824
rect 553820 236784 553826 236796
rect 559558 236784 559564 236796
rect 559616 236784 559622 236836
rect 672954 236700 673006 236706
rect 672954 236642 673006 236648
rect 672966 236524 673118 236552
rect 671706 236444 671712 236496
rect 671764 236484 671770 236496
rect 672966 236484 672994 236524
rect 671764 236456 672994 236484
rect 673184 236496 673236 236502
rect 671764 236444 671770 236456
rect 673184 236438 673236 236444
rect 671540 236048 673330 236076
rect 671062 235900 671068 235952
rect 671120 235940 671126 235952
rect 671540 235940 671568 236048
rect 671120 235912 671568 235940
rect 671120 235900 671126 235912
rect 673408 235832 673414 235884
rect 673466 235832 673472 235884
rect 672074 235696 672080 235748
rect 672132 235736 672138 235748
rect 672132 235708 673554 235736
rect 672132 235696 672138 235708
rect 673178 235492 673184 235544
rect 673236 235532 673242 235544
rect 673236 235504 673670 235532
rect 673236 235492 673242 235504
rect 672994 235016 673000 235068
rect 673052 235056 673058 235068
rect 673764 235056 673792 235314
rect 673052 235028 673792 235056
rect 673052 235016 673058 235028
rect 673454 234812 673460 234864
rect 673512 234852 673518 234864
rect 673886 234852 673914 235110
rect 673512 234824 673914 234852
rect 673512 234812 673518 234824
rect 673978 234648 674006 234906
rect 674088 234728 674140 234734
rect 674088 234670 674140 234676
rect 673316 234620 674006 234648
rect 554406 234540 554412 234592
rect 554464 234580 554470 234592
rect 570598 234580 570604 234592
rect 554464 234552 570604 234580
rect 554464 234540 554470 234552
rect 570598 234540 570604 234552
rect 570656 234540 570662 234592
rect 669774 234540 669780 234592
rect 669832 234580 669838 234592
rect 673316 234580 673344 234620
rect 669832 234552 673344 234580
rect 669832 234540 669838 234552
rect 669590 234132 669596 234184
rect 669648 234172 669654 234184
rect 674208 234172 674236 234498
rect 669648 234144 674236 234172
rect 669648 234132 669654 234144
rect 675846 233996 675852 234048
rect 675904 234036 675910 234048
rect 678238 234036 678244 234048
rect 675904 234008 678244 234036
rect 675904 233996 675910 234008
rect 678238 233996 678244 234008
rect 678296 233996 678302 234048
rect 670878 233968 670884 233980
rect 663766 233940 670884 233968
rect 652386 233860 652392 233912
rect 652444 233900 652450 233912
rect 663766 233900 663794 233940
rect 670878 233928 670884 233940
rect 670936 233928 670942 233980
rect 652444 233872 663794 233900
rect 652444 233860 652450 233872
rect 671366 233724 671372 233776
rect 671424 233764 671430 233776
rect 674098 233764 674104 233776
rect 671424 233736 674104 233764
rect 671424 233724 671430 233736
rect 674098 233724 674104 233736
rect 674156 233724 674162 233776
rect 672258 233248 672264 233300
rect 672316 233288 672322 233300
rect 673178 233288 673184 233300
rect 672316 233260 673184 233288
rect 672316 233248 672322 233260
rect 673178 233248 673184 233260
rect 673236 233248 673242 233300
rect 670878 233180 670884 233232
rect 670936 233220 670942 233232
rect 672074 233220 672080 233232
rect 670936 233192 672080 233220
rect 670936 233180 670942 233192
rect 672074 233180 672080 233192
rect 672132 233180 672138 233232
rect 673454 233180 673460 233232
rect 673512 233220 673518 233232
rect 674282 233220 674288 233232
rect 673512 233192 674288 233220
rect 673512 233180 673518 233192
rect 674282 233180 674288 233192
rect 674340 233180 674346 233232
rect 670326 233044 670332 233096
rect 670384 233084 670390 233096
rect 672994 233084 673000 233096
rect 670384 233056 673000 233084
rect 670384 233044 670390 233056
rect 672994 233044 673000 233056
rect 673052 233044 673058 233096
rect 663058 232636 663064 232688
rect 663116 232676 663122 232688
rect 674098 232676 674104 232688
rect 663116 232648 674104 232676
rect 663116 232636 663122 232648
rect 674098 232636 674104 232648
rect 674156 232636 674162 232688
rect 675846 232636 675852 232688
rect 675904 232676 675910 232688
rect 683206 232676 683212 232688
rect 675904 232648 683212 232676
rect 675904 232636 675910 232648
rect 683206 232636 683212 232648
rect 683264 232636 683270 232688
rect 653398 232500 653404 232552
rect 653456 232540 653462 232552
rect 653456 232512 663794 232540
rect 653456 232500 653462 232512
rect 663766 232472 663794 232512
rect 676030 232500 676036 232552
rect 676088 232540 676094 232552
rect 683390 232540 683396 232552
rect 676088 232512 683396 232540
rect 676088 232500 676094 232512
rect 683390 232500 683396 232512
rect 683448 232500 683454 232552
rect 663766 232444 666554 232472
rect 666526 232404 666554 232444
rect 674098 232404 674104 232416
rect 666526 232376 674104 232404
rect 674098 232364 674104 232376
rect 674156 232364 674162 232416
rect 666278 231548 666284 231600
rect 666336 231588 666342 231600
rect 674834 231588 674840 231600
rect 666336 231560 674840 231588
rect 666336 231548 666342 231560
rect 674834 231548 674840 231560
rect 674892 231548 674898 231600
rect 134978 231412 134984 231464
rect 135036 231452 135042 231464
rect 137646 231452 137652 231464
rect 135036 231424 137652 231452
rect 135036 231412 135042 231424
rect 137646 231412 137652 231424
rect 137704 231412 137710 231464
rect 61378 231276 61384 231328
rect 61436 231316 61442 231328
rect 668854 231316 668860 231328
rect 61436 231288 668860 231316
rect 61436 231276 61442 231288
rect 668854 231276 668860 231288
rect 668912 231276 668918 231328
rect 92382 231140 92388 231192
rect 92440 231180 92446 231192
rect 170766 231180 170772 231192
rect 92440 231152 170772 231180
rect 92440 231140 92446 231152
rect 170766 231140 170772 231152
rect 170824 231140 170830 231192
rect 665082 231140 665088 231192
rect 665140 231180 665146 231192
rect 665140 231152 675326 231180
rect 665140 231140 665146 231152
rect 128262 231004 128268 231056
rect 128320 231044 128326 231056
rect 195882 231044 195888 231056
rect 128320 231016 195888 231044
rect 128320 231004 128326 231016
rect 195882 231004 195888 231016
rect 195940 231004 195946 231056
rect 666462 230936 666468 230988
rect 666520 230976 666526 230988
rect 666520 230948 675142 230976
rect 666520 230936 666526 230948
rect 104802 230868 104808 230920
rect 104860 230908 104866 230920
rect 179138 230908 179144 230920
rect 104860 230880 179144 230908
rect 104860 230868 104866 230880
rect 179138 230868 179144 230880
rect 179196 230868 179202 230920
rect 674834 230800 674840 230852
rect 674892 230840 674898 230852
rect 674892 230812 674982 230840
rect 674892 230800 674898 230812
rect 118602 230732 118608 230784
rect 118660 230772 118666 230784
rect 188154 230772 188160 230784
rect 118660 230744 188160 230772
rect 118660 230732 118666 230744
rect 188154 230732 188160 230744
rect 188212 230732 188218 230784
rect 94498 230596 94504 230648
rect 94556 230636 94562 230648
rect 171410 230636 171416 230648
rect 94556 230608 171416 230636
rect 94556 230596 94562 230608
rect 171410 230596 171416 230608
rect 171468 230596 171474 230648
rect 194410 230596 194416 230648
rect 194468 230636 194474 230648
rect 196894 230636 196900 230648
rect 194468 230608 196900 230636
rect 194468 230596 194474 230608
rect 196894 230596 196900 230608
rect 196952 230596 196958 230648
rect 672074 230596 672080 230648
rect 672132 230636 672138 230648
rect 672132 230608 674820 230636
rect 672132 230596 672138 230608
rect 439314 230528 439320 230580
rect 439372 230568 439378 230580
rect 439372 230540 439544 230568
rect 439372 230528 439378 230540
rect 137646 230460 137652 230512
rect 137704 230500 137710 230512
rect 201034 230500 201040 230512
rect 137704 230472 201040 230500
rect 137704 230460 137710 230472
rect 201034 230460 201040 230472
rect 201092 230460 201098 230512
rect 42150 230392 42156 230444
rect 42208 230432 42214 230444
rect 43254 230432 43260 230444
rect 42208 230404 43260 230432
rect 42208 230392 42214 230404
rect 43254 230392 43260 230404
rect 43312 230392 43318 230444
rect 133782 230392 133788 230444
rect 133840 230432 133846 230444
rect 137462 230432 137468 230444
rect 133840 230404 137468 230432
rect 133840 230392 133846 230404
rect 137462 230392 137468 230404
rect 137520 230392 137526 230444
rect 213086 230392 213092 230444
rect 213144 230432 213150 230444
rect 261570 230432 261576 230444
rect 213144 230404 261576 230432
rect 213144 230392 213150 230404
rect 261570 230392 261576 230404
rect 261628 230392 261634 230444
rect 311986 230392 311992 230444
rect 312044 230432 312050 230444
rect 313090 230432 313096 230444
rect 312044 230404 313096 230432
rect 312044 230392 312050 230404
rect 313090 230392 313096 230404
rect 313148 230392 313154 230444
rect 374638 230392 374644 230444
rect 374696 230432 374702 230444
rect 376202 230432 376208 230444
rect 374696 230404 376208 230432
rect 374696 230392 374702 230404
rect 376202 230392 376208 230404
rect 376260 230392 376266 230444
rect 433426 230392 433432 230444
rect 433484 230432 433490 230444
rect 434162 230432 434168 230444
rect 433484 230404 434168 230432
rect 433484 230392 433490 230404
rect 434162 230392 434168 230404
rect 434220 230392 434226 230444
rect 439516 230432 439544 230540
rect 440694 230432 440700 230444
rect 439516 230404 440700 230432
rect 440694 230392 440700 230404
rect 440752 230392 440758 230444
rect 441890 230392 441896 230444
rect 441948 230432 441954 230444
rect 443454 230432 443460 230444
rect 441948 230404 443460 230432
rect 441948 230392 441954 230404
rect 443454 230392 443460 230404
rect 443512 230392 443518 230444
rect 451550 230392 451556 230444
rect 451608 230432 451614 230444
rect 453298 230432 453304 230444
rect 451608 230404 453304 230432
rect 451608 230392 451614 230404
rect 453298 230392 453304 230404
rect 453356 230392 453362 230444
rect 532510 230392 532516 230444
rect 532568 230432 532574 230444
rect 538306 230432 538312 230444
rect 532568 230404 538312 230432
rect 532568 230392 532574 230404
rect 538306 230392 538312 230404
rect 538364 230392 538370 230444
rect 673270 230392 673276 230444
rect 673328 230432 673334 230444
rect 673328 230404 674702 230432
rect 673328 230392 673334 230404
rect 387426 230324 387432 230376
rect 387484 230364 387490 230376
rect 388438 230364 388444 230376
rect 387484 230336 388444 230364
rect 387484 230324 387490 230336
rect 388438 230324 388444 230336
rect 388496 230324 388502 230376
rect 398098 230324 398104 230376
rect 398156 230364 398162 230376
rect 399386 230364 399392 230376
rect 398156 230336 399392 230364
rect 398156 230324 398162 230336
rect 399386 230324 399392 230336
rect 399444 230324 399450 230376
rect 436094 230324 436100 230376
rect 436152 230364 436158 230376
rect 436738 230364 436744 230376
rect 436152 230336 436744 230364
rect 436152 230324 436158 230336
rect 436738 230324 436744 230336
rect 436796 230324 436802 230376
rect 438670 230324 438676 230376
rect 438728 230364 438734 230376
rect 439314 230364 439320 230376
rect 438728 230336 439320 230364
rect 438728 230324 438734 230336
rect 439314 230324 439320 230336
rect 439372 230324 439378 230376
rect 443822 230324 443828 230376
rect 443880 230364 443886 230376
rect 444926 230364 444932 230376
rect 443880 230336 444932 230364
rect 443880 230324 443886 230336
rect 444926 230324 444932 230336
rect 444984 230324 444990 230376
rect 455414 230324 455420 230376
rect 455472 230364 455478 230376
rect 457162 230364 457168 230376
rect 455472 230336 457168 230364
rect 455472 230324 455478 230336
rect 457162 230324 457168 230336
rect 457220 230324 457226 230376
rect 463786 230324 463792 230376
rect 463844 230364 463850 230376
rect 465718 230364 465724 230376
rect 463844 230336 465724 230364
rect 463844 230324 463850 230336
rect 465718 230324 465724 230336
rect 465776 230324 465782 230376
rect 470870 230324 470876 230376
rect 470928 230364 470934 230376
rect 471882 230364 471888 230376
rect 470928 230336 471888 230364
rect 470928 230324 470934 230336
rect 471882 230324 471888 230336
rect 471940 230324 471946 230376
rect 476022 230324 476028 230376
rect 476080 230364 476086 230376
rect 478598 230364 478604 230376
rect 476080 230336 478604 230364
rect 476080 230324 476086 230336
rect 478598 230324 478604 230336
rect 478656 230324 478662 230376
rect 493410 230324 493416 230376
rect 493468 230364 493474 230376
rect 496354 230364 496360 230376
rect 493468 230336 496360 230364
rect 493468 230324 493474 230336
rect 496354 230324 496360 230336
rect 496412 230324 496418 230376
rect 497274 230324 497280 230376
rect 497332 230364 497338 230376
rect 498102 230364 498108 230376
rect 497332 230336 498108 230364
rect 497332 230324 497338 230336
rect 498102 230324 498108 230336
rect 498160 230324 498166 230376
rect 510798 230324 510804 230376
rect 510856 230364 510862 230376
rect 511902 230364 511908 230376
rect 510856 230336 511908 230364
rect 510856 230324 510862 230336
rect 511902 230324 511908 230336
rect 511960 230324 511966 230376
rect 521102 230324 521108 230376
rect 521160 230364 521166 230376
rect 526438 230364 526444 230376
rect 521160 230336 526444 230364
rect 521160 230324 521166 230336
rect 526438 230324 526444 230336
rect 526496 230324 526502 230376
rect 530118 230324 530124 230376
rect 530176 230364 530182 230376
rect 531130 230364 531136 230376
rect 530176 230336 531136 230364
rect 530176 230324 530182 230336
rect 531130 230324 531136 230336
rect 531188 230324 531194 230376
rect 126882 230256 126888 230308
rect 126940 230296 126946 230308
rect 194410 230296 194416 230308
rect 126940 230268 194416 230296
rect 126940 230256 126946 230268
rect 194410 230256 194416 230268
rect 194468 230256 194474 230308
rect 194870 230256 194876 230308
rect 194928 230296 194934 230308
rect 195422 230296 195428 230308
rect 194928 230268 195428 230296
rect 194928 230256 194934 230268
rect 195422 230256 195428 230268
rect 195480 230256 195486 230308
rect 195606 230256 195612 230308
rect 195664 230296 195670 230308
rect 204898 230296 204904 230308
rect 195664 230268 204904 230296
rect 195664 230256 195670 230268
rect 204898 230256 204904 230268
rect 204956 230256 204962 230308
rect 206278 230256 206284 230308
rect 206336 230296 206342 230308
rect 256418 230296 256424 230308
rect 206336 230268 256424 230296
rect 206336 230256 206342 230268
rect 256418 230256 256424 230268
rect 256476 230256 256482 230308
rect 256602 230256 256608 230308
rect 256660 230296 256666 230308
rect 297634 230296 297640 230308
rect 256660 230268 297640 230296
rect 256660 230256 256666 230268
rect 297634 230256 297640 230268
rect 297692 230256 297698 230308
rect 297818 230256 297824 230308
rect 297876 230296 297882 230308
rect 323394 230296 323400 230308
rect 297876 230268 323400 230296
rect 297876 230256 297882 230268
rect 323394 230256 323400 230268
rect 323452 230256 323458 230308
rect 539594 230296 539600 230308
rect 532528 230268 539600 230296
rect 444466 230188 444472 230240
rect 444524 230228 444530 230240
rect 447594 230228 447600 230240
rect 444524 230200 447600 230228
rect 444524 230188 444530 230200
rect 447594 230188 447600 230200
rect 447652 230188 447658 230240
rect 452838 230188 452844 230240
rect 452896 230228 452902 230240
rect 454310 230228 454316 230240
rect 452896 230200 454316 230228
rect 452896 230188 452902 230200
rect 454310 230188 454316 230200
rect 454368 230188 454374 230240
rect 468294 230188 468300 230240
rect 468352 230228 468358 230240
rect 469122 230228 469128 230240
rect 468352 230200 469128 230228
rect 468352 230188 468358 230200
rect 469122 230188 469128 230200
rect 469180 230188 469186 230240
rect 487614 230188 487620 230240
rect 487672 230228 487678 230240
rect 488442 230228 488448 230240
rect 487672 230200 488448 230228
rect 487672 230188 487678 230200
rect 488442 230188 488448 230200
rect 488500 230188 488506 230240
rect 495158 230228 495164 230240
rect 489886 230200 495164 230228
rect 95234 230120 95240 230172
rect 95292 230160 95298 230172
rect 165982 230160 165988 230172
rect 95292 230132 165988 230160
rect 95292 230120 95298 230132
rect 165982 230120 165988 230132
rect 166040 230120 166046 230172
rect 166258 230120 166264 230172
rect 166316 230160 166322 230172
rect 185578 230160 185584 230172
rect 166316 230132 185584 230160
rect 166316 230120 166322 230132
rect 185578 230120 185584 230132
rect 185636 230120 185642 230172
rect 186038 230120 186044 230172
rect 186096 230160 186102 230172
rect 235810 230160 235816 230172
rect 186096 230132 235816 230160
rect 186096 230120 186102 230132
rect 235810 230120 235816 230132
rect 235868 230120 235874 230172
rect 240318 230120 240324 230172
rect 240376 230160 240382 230172
rect 282178 230160 282184 230172
rect 240376 230132 282184 230160
rect 240376 230120 240382 230132
rect 282178 230120 282184 230132
rect 282236 230120 282242 230172
rect 282638 230120 282644 230172
rect 282696 230160 282702 230172
rect 307938 230160 307944 230172
rect 282696 230132 307944 230160
rect 282696 230120 282702 230132
rect 307938 230120 307944 230132
rect 307996 230120 308002 230172
rect 308122 230120 308128 230172
rect 308180 230160 308186 230172
rect 334986 230160 334992 230172
rect 308180 230132 334992 230160
rect 308180 230120 308186 230132
rect 334986 230120 334992 230132
rect 335044 230120 335050 230172
rect 335170 230120 335176 230172
rect 335228 230160 335234 230172
rect 350442 230160 350448 230172
rect 335228 230132 350448 230160
rect 335228 230120 335234 230132
rect 350442 230120 350448 230132
rect 350500 230120 350506 230172
rect 454126 230052 454132 230104
rect 454184 230092 454190 230104
rect 455322 230092 455328 230104
rect 454184 230064 455328 230092
rect 454184 230052 454190 230064
rect 455322 230052 455328 230064
rect 455380 230052 455386 230104
rect 82078 229984 82084 230036
rect 82136 230024 82142 230036
rect 82136 229996 84194 230024
rect 82136 229984 82142 229996
rect 84166 229888 84194 229996
rect 86218 229984 86224 230036
rect 86276 230024 86282 230036
rect 137278 230024 137284 230036
rect 86276 229996 137284 230024
rect 86276 229984 86282 229996
rect 137278 229984 137284 229996
rect 137336 229984 137342 230036
rect 137462 229984 137468 230036
rect 137520 230024 137526 230036
rect 195054 230024 195060 230036
rect 137520 229996 195060 230024
rect 137520 229984 137526 229996
rect 195054 229984 195060 229996
rect 195112 229984 195118 230036
rect 195422 229984 195428 230036
rect 195480 230024 195486 230036
rect 215202 230024 215208 230036
rect 195480 229996 215208 230024
rect 195480 229984 195486 229996
rect 215202 229984 215208 229996
rect 215260 229984 215266 230036
rect 230474 229984 230480 230036
rect 230532 230024 230538 230036
rect 277026 230024 277032 230036
rect 230532 229996 277032 230024
rect 230532 229984 230538 229996
rect 277026 229984 277032 229996
rect 277084 229984 277090 230036
rect 277210 229984 277216 230036
rect 277268 230024 277274 230036
rect 302786 230024 302792 230036
rect 277268 229996 302792 230024
rect 277268 229984 277274 229996
rect 302786 229984 302792 229996
rect 302844 229984 302850 230036
rect 303246 229984 303252 230036
rect 303304 230024 303310 230036
rect 329834 230024 329840 230036
rect 303304 229996 329840 230024
rect 303304 229984 303310 229996
rect 329834 229984 329840 229996
rect 329892 229984 329898 230036
rect 330938 229984 330944 230036
rect 330996 230024 331002 230036
rect 355594 230024 355600 230036
rect 330996 229996 355600 230024
rect 330996 229984 331002 229996
rect 355594 229984 355600 229996
rect 355652 229984 355658 230036
rect 448330 229984 448336 230036
rect 448388 230024 448394 230036
rect 448974 230024 448980 230036
rect 448388 229996 448980 230024
rect 448388 229984 448394 229996
rect 448974 229984 448980 229996
rect 449032 229984 449038 230036
rect 484394 229984 484400 230036
rect 484452 230024 484458 230036
rect 489886 230024 489914 230200
rect 495158 230188 495164 230200
rect 495216 230188 495222 230240
rect 511442 230188 511448 230240
rect 511500 230228 511506 230240
rect 517514 230228 517520 230240
rect 511500 230200 517520 230228
rect 511500 230188 511506 230200
rect 517514 230188 517520 230200
rect 517572 230188 517578 230240
rect 530762 230188 530768 230240
rect 530820 230228 530826 230240
rect 532528 230228 532556 230268
rect 539594 230256 539600 230268
rect 539652 230256 539658 230308
rect 530820 230200 532556 230228
rect 530820 230188 530826 230200
rect 673454 230188 673460 230240
rect 673512 230228 673518 230240
rect 673512 230200 674590 230228
rect 673512 230188 673518 230200
rect 532694 230120 532700 230172
rect 532752 230160 532758 230172
rect 547138 230160 547144 230172
rect 532752 230132 547144 230160
rect 532752 230120 532758 230132
rect 547138 230120 547144 230132
rect 547196 230120 547202 230172
rect 491478 230052 491484 230104
rect 491536 230092 491542 230104
rect 492490 230092 492496 230104
rect 491536 230064 492496 230092
rect 491536 230052 491542 230064
rect 492490 230052 492496 230064
rect 492548 230052 492554 230104
rect 528830 230052 528836 230104
rect 528888 230092 528894 230104
rect 532510 230092 532516 230104
rect 528888 230064 532516 230092
rect 528888 230052 528894 230064
rect 532510 230052 532516 230064
rect 532568 230052 532574 230104
rect 560938 230052 560944 230104
rect 560996 230092 561002 230104
rect 568114 230092 568120 230104
rect 560996 230064 568120 230092
rect 560996 230052 561002 230064
rect 568114 230052 568120 230064
rect 568172 230052 568178 230104
rect 484452 229996 489914 230024
rect 484452 229984 484458 229996
rect 517238 229984 517244 230036
rect 517296 230024 517302 230036
rect 524598 230024 524604 230036
rect 517296 229996 524604 230024
rect 517296 229984 517302 229996
rect 524598 229984 524604 229996
rect 524656 229984 524662 230036
rect 534626 229984 534632 230036
rect 534684 230024 534690 230036
rect 550542 230024 550548 230036
rect 534684 229996 550548 230024
rect 534684 229984 534690 229996
rect 550542 229984 550548 229996
rect 550600 229984 550606 230036
rect 674098 229984 674104 230036
rect 674156 230024 674162 230036
rect 674156 229996 674478 230024
rect 674156 229984 674162 229996
rect 453482 229916 453488 229968
rect 453540 229956 453546 229968
rect 455782 229956 455788 229968
rect 453540 229928 455788 229956
rect 453540 229916 453546 229928
rect 455782 229916 455788 229928
rect 455840 229916 455846 229968
rect 151722 229888 151728 229900
rect 84166 229860 151728 229888
rect 151722 229848 151728 229860
rect 151780 229848 151786 229900
rect 151906 229848 151912 229900
rect 151964 229888 151970 229900
rect 166258 229888 166264 229900
rect 151964 229860 166264 229888
rect 151964 229848 151970 229860
rect 166258 229848 166264 229860
rect 166316 229848 166322 229900
rect 225506 229888 225512 229900
rect 171106 229860 225512 229888
rect 68278 229712 68284 229764
rect 68336 229752 68342 229764
rect 144454 229752 144460 229764
rect 68336 229724 144460 229752
rect 68336 229712 68342 229724
rect 144454 229712 144460 229724
rect 144512 229712 144518 229764
rect 144822 229712 144828 229764
rect 144880 229752 144886 229764
rect 146294 229752 146300 229764
rect 144880 229724 146300 229752
rect 144880 229712 144886 229724
rect 146294 229712 146300 229724
rect 146352 229712 146358 229764
rect 154022 229752 154028 229764
rect 146956 229724 154028 229752
rect 137278 229576 137284 229628
rect 137336 229616 137342 229628
rect 146956 229616 146984 229724
rect 154022 229712 154028 229724
rect 154080 229712 154086 229764
rect 154206 229712 154212 229764
rect 154264 229752 154270 229764
rect 161382 229752 161388 229764
rect 154264 229724 161388 229752
rect 154264 229712 154270 229724
rect 161382 229712 161388 229724
rect 161440 229712 161446 229764
rect 161750 229752 161756 229764
rect 161584 229724 161756 229752
rect 137336 229588 146984 229616
rect 137336 229576 137342 229588
rect 151170 229576 151176 229628
rect 151228 229616 151234 229628
rect 161584 229616 161612 229724
rect 161750 229712 161756 229724
rect 161808 229712 161814 229764
rect 163958 229712 163964 229764
rect 164016 229752 164022 229764
rect 171106 229752 171134 229860
rect 225506 229848 225512 229860
rect 225564 229848 225570 229900
rect 225690 229848 225696 229900
rect 225748 229888 225754 229900
rect 271874 229888 271880 229900
rect 225748 229860 271880 229888
rect 225748 229848 225754 229860
rect 271874 229848 271880 229860
rect 271932 229848 271938 229900
rect 275646 229848 275652 229900
rect 275704 229888 275710 229900
rect 311986 229888 311992 229900
rect 275704 229860 311992 229888
rect 275704 229848 275710 229860
rect 311986 229848 311992 229860
rect 312044 229848 312050 229900
rect 312630 229848 312636 229900
rect 312688 229888 312694 229900
rect 340138 229888 340144 229900
rect 312688 229860 340144 229888
rect 312688 229848 312694 229860
rect 340138 229848 340144 229860
rect 340196 229848 340202 229900
rect 345658 229848 345664 229900
rect 345716 229888 345722 229900
rect 360746 229888 360752 229900
rect 345716 229860 360752 229888
rect 345716 229848 345722 229860
rect 360746 229848 360752 229860
rect 360804 229848 360810 229900
rect 361206 229848 361212 229900
rect 361264 229888 361270 229900
rect 378778 229888 378784 229900
rect 361264 229860 378784 229888
rect 361264 229848 361270 229860
rect 378778 229848 378784 229860
rect 378836 229848 378842 229900
rect 449618 229848 449624 229900
rect 449676 229888 449682 229900
rect 450538 229888 450544 229900
rect 449676 229860 450544 229888
rect 449676 229848 449682 229860
rect 450538 229848 450544 229860
rect 450596 229848 450602 229900
rect 467006 229848 467012 229900
rect 467064 229888 467070 229900
rect 473998 229888 474004 229900
rect 467064 229860 474004 229888
rect 467064 229848 467070 229860
rect 473998 229848 474004 229860
rect 474056 229848 474062 229900
rect 476666 229848 476672 229900
rect 476724 229888 476730 229900
rect 481634 229888 481640 229900
rect 476724 229860 481640 229888
rect 476724 229848 476730 229860
rect 481634 229848 481640 229860
rect 481692 229848 481698 229900
rect 481818 229848 481824 229900
rect 481876 229888 481882 229900
rect 493594 229888 493600 229900
rect 481876 229860 493600 229888
rect 481876 229848 481882 229860
rect 493594 229848 493600 229860
rect 493652 229848 493658 229900
rect 495986 229848 495992 229900
rect 496044 229888 496050 229900
rect 506382 229888 506388 229900
rect 496044 229860 506388 229888
rect 496044 229848 496050 229860
rect 506382 229848 506388 229860
rect 506440 229848 506446 229900
rect 507578 229848 507584 229900
rect 507636 229888 507642 229900
rect 516778 229888 516784 229900
rect 507636 229860 516784 229888
rect 507636 229848 507642 229860
rect 516778 229848 516784 229860
rect 516836 229848 516842 229900
rect 519170 229848 519176 229900
rect 519228 229888 519234 229900
rect 528554 229888 528560 229900
rect 519228 229860 528560 229888
rect 519228 229848 519234 229860
rect 528554 229848 528560 229860
rect 528612 229848 528618 229900
rect 536558 229848 536564 229900
rect 536616 229888 536622 229900
rect 559558 229888 559564 229900
rect 536616 229860 559564 229888
rect 536616 229848 536622 229860
rect 559558 229848 559564 229860
rect 559616 229848 559622 229900
rect 674098 229780 674104 229832
rect 674156 229820 674162 229832
rect 674156 229792 674360 229820
rect 674156 229780 674162 229792
rect 164016 229724 171134 229752
rect 164016 229712 164022 229724
rect 173710 229712 173716 229764
rect 173768 229752 173774 229764
rect 175918 229752 175924 229764
rect 173768 229724 175924 229752
rect 173768 229712 173774 229724
rect 175918 229712 175924 229724
rect 175976 229712 175982 229764
rect 176378 229712 176384 229764
rect 176436 229752 176442 229764
rect 185394 229752 185400 229764
rect 176436 229724 185400 229752
rect 176436 229712 176442 229724
rect 185394 229712 185400 229724
rect 185452 229712 185458 229764
rect 185578 229712 185584 229764
rect 185636 229752 185642 229764
rect 194870 229752 194876 229764
rect 185636 229724 194876 229752
rect 185636 229712 185642 229724
rect 194870 229712 194876 229724
rect 194928 229712 194934 229764
rect 195054 229712 195060 229764
rect 195112 229752 195118 229764
rect 202322 229752 202328 229764
rect 195112 229724 202328 229752
rect 195112 229712 195118 229724
rect 202322 229712 202328 229724
rect 202380 229712 202386 229764
rect 204898 229712 204904 229764
rect 204956 229752 204962 229764
rect 246114 229752 246120 229764
rect 204956 229724 246120 229752
rect 204956 229712 204962 229724
rect 246114 229712 246120 229724
rect 246172 229712 246178 229764
rect 246482 229712 246488 229764
rect 246540 229752 246546 229764
rect 287330 229752 287336 229764
rect 246540 229724 287336 229752
rect 246540 229712 246546 229724
rect 287330 229712 287336 229724
rect 287388 229712 287394 229764
rect 287698 229712 287704 229764
rect 287756 229752 287762 229764
rect 318242 229752 318248 229764
rect 287756 229724 318248 229752
rect 287756 229712 287762 229724
rect 318242 229712 318248 229724
rect 318300 229712 318306 229764
rect 345290 229752 345296 229764
rect 325666 229724 345296 229752
rect 151228 229588 161612 229616
rect 151228 229576 151234 229588
rect 161750 229576 161756 229628
rect 161808 229616 161814 229628
rect 220354 229616 220360 229628
rect 161808 229588 220360 229616
rect 161808 229576 161814 229588
rect 220354 229576 220360 229588
rect 220412 229576 220418 229628
rect 251266 229616 251272 229628
rect 229066 229588 251272 229616
rect 150986 229548 150992 229560
rect 147048 229520 150992 229548
rect 102134 229440 102140 229492
rect 102192 229480 102198 229492
rect 145650 229480 145656 229492
rect 102192 229452 145656 229480
rect 102192 229440 102198 229452
rect 145650 229440 145656 229452
rect 145708 229440 145714 229492
rect 146018 229372 146024 229424
rect 146076 229412 146082 229424
rect 147048 229412 147076 229520
rect 150986 229508 150992 229520
rect 151044 229508 151050 229560
rect 151768 229440 151774 229492
rect 151826 229480 151832 229492
rect 210050 229480 210056 229492
rect 151826 229452 210056 229480
rect 151826 229440 151832 229452
rect 210050 229440 210056 229452
rect 210108 229440 210114 229492
rect 220446 229440 220452 229492
rect 220504 229480 220510 229492
rect 229066 229480 229094 229588
rect 251266 229576 251272 229588
rect 251324 229576 251330 229628
rect 251726 229576 251732 229628
rect 251784 229616 251790 229628
rect 292482 229616 292488 229628
rect 251784 229588 292488 229616
rect 251784 229576 251790 229588
rect 292482 229576 292488 229588
rect 292540 229576 292546 229628
rect 318058 229576 318064 229628
rect 318116 229616 318122 229628
rect 325666 229616 325694 229724
rect 345290 229712 345296 229724
rect 345348 229712 345354 229764
rect 351730 229712 351736 229764
rect 351788 229752 351794 229764
rect 371050 229752 371056 229764
rect 351788 229724 371056 229752
rect 351788 229712 351794 229724
rect 371050 229712 371056 229724
rect 371108 229712 371114 229764
rect 377674 229712 377680 229764
rect 377732 229752 377738 229764
rect 389082 229752 389088 229764
rect 377732 229724 389088 229752
rect 377732 229712 377738 229724
rect 389082 229712 389088 229724
rect 389140 229712 389146 229764
rect 399846 229712 399852 229764
rect 399904 229752 399910 229764
rect 409690 229752 409696 229764
rect 399904 229724 409696 229752
rect 399904 229712 399910 229724
rect 409690 229712 409696 229724
rect 409748 229712 409754 229764
rect 410886 229712 410892 229764
rect 410944 229752 410950 229764
rect 417418 229752 417424 229764
rect 410944 229724 417424 229752
rect 410944 229712 410950 229724
rect 417418 229712 417424 229724
rect 417476 229712 417482 229764
rect 457346 229712 457352 229764
rect 457404 229752 457410 229764
rect 463878 229752 463884 229764
rect 457404 229724 463884 229752
rect 457404 229712 457410 229724
rect 463878 229712 463884 229724
rect 463936 229712 463942 229764
rect 465442 229712 465448 229764
rect 465500 229752 465506 229764
rect 467466 229752 467472 229764
rect 465500 229724 467472 229752
rect 465500 229712 465506 229724
rect 467466 229712 467472 229724
rect 467524 229712 467530 229764
rect 469582 229712 469588 229764
rect 469640 229752 469646 229764
rect 476758 229752 476764 229764
rect 469640 229724 476764 229752
rect 469640 229712 469646 229724
rect 476758 229712 476764 229724
rect 476816 229712 476822 229764
rect 479242 229712 479248 229764
rect 479300 229752 479306 229764
rect 489914 229752 489920 229764
rect 479300 229724 489920 229752
rect 479300 229712 479306 229724
rect 489914 229712 489920 229724
rect 489972 229712 489978 229764
rect 492122 229712 492128 229764
rect 492180 229752 492186 229764
rect 507118 229752 507124 229764
rect 492180 229724 507124 229752
rect 492180 229712 492186 229724
rect 507118 229712 507124 229724
rect 507176 229712 507182 229764
rect 523034 229712 523040 229764
rect 523092 229752 523098 229764
rect 534718 229752 534724 229764
rect 523092 229724 534724 229752
rect 523092 229712 523098 229724
rect 534718 229712 534724 229724
rect 534776 229712 534782 229764
rect 538490 229712 538496 229764
rect 538548 229752 538554 229764
rect 566826 229752 566832 229764
rect 538548 229724 566832 229752
rect 538548 229712 538554 229724
rect 566826 229712 566832 229724
rect 566884 229712 566890 229764
rect 663702 229712 663708 229764
rect 663760 229752 663766 229764
rect 672074 229752 672080 229764
rect 663760 229724 672080 229752
rect 663760 229712 663766 229724
rect 672074 229712 672080 229724
rect 672132 229712 672138 229764
rect 509510 229644 509516 229696
rect 509568 229684 509574 229696
rect 515490 229684 515496 229696
rect 509568 229656 515496 229684
rect 509568 229644 509574 229656
rect 515490 229644 515496 229656
rect 515548 229644 515554 229696
rect 318116 229588 325694 229616
rect 318116 229576 318122 229588
rect 388622 229576 388628 229628
rect 388680 229616 388686 229628
rect 398742 229616 398748 229628
rect 388680 229588 398748 229616
rect 388680 229576 388686 229588
rect 398742 229576 398748 229588
rect 398800 229576 398806 229628
rect 526898 229576 526904 229628
rect 526956 229616 526962 229628
rect 536098 229616 536104 229628
rect 526956 229588 536104 229616
rect 526956 229576 526962 229588
rect 536098 229576 536104 229588
rect 536156 229576 536162 229628
rect 673362 229576 673368 229628
rect 673420 229616 673426 229628
rect 673420 229588 674268 229616
rect 673420 229576 673426 229588
rect 449250 229508 449256 229560
rect 449308 229548 449314 229560
rect 451918 229548 451924 229560
rect 449308 229520 451924 229548
rect 449308 229508 449314 229520
rect 451918 229508 451924 229520
rect 451976 229508 451982 229560
rect 220504 229452 229094 229480
rect 220504 229440 220510 229452
rect 146076 229384 147076 229412
rect 146076 229372 146082 229384
rect 148318 229372 148324 229424
rect 148376 229412 148382 229424
rect 151630 229412 151636 229424
rect 148376 229384 151636 229412
rect 148376 229372 148382 229384
rect 151630 229372 151636 229384
rect 151688 229372 151694 229424
rect 674104 229356 674156 229362
rect 110322 229304 110328 229356
rect 110380 229344 110386 229356
rect 145834 229344 145840 229356
rect 110380 229316 145840 229344
rect 110380 229304 110386 229316
rect 145834 229304 145840 229316
rect 145892 229304 145898 229356
rect 153378 229344 153384 229356
rect 151786 229316 153384 229344
rect 123478 229168 123484 229220
rect 123536 229208 123542 229220
rect 151786 229208 151814 229316
rect 153378 229304 153384 229316
rect 153436 229304 153442 229356
rect 153838 229304 153844 229356
rect 153896 229344 153902 229356
rect 157794 229344 157800 229356
rect 153896 229316 157800 229344
rect 153896 229304 153902 229316
rect 157794 229304 157800 229316
rect 157852 229304 157858 229356
rect 157978 229304 157984 229356
rect 158036 229344 158042 229356
rect 163682 229344 163688 229356
rect 158036 229316 163688 229344
rect 158036 229304 158042 229316
rect 163682 229304 163688 229316
rect 163740 229304 163746 229356
rect 164234 229304 164240 229356
rect 164292 229344 164298 229356
rect 169110 229344 169116 229356
rect 164292 229316 169116 229344
rect 164292 229304 164298 229316
rect 169110 229304 169116 229316
rect 169168 229304 169174 229356
rect 170950 229304 170956 229356
rect 171008 229344 171014 229356
rect 230658 229344 230664 229356
rect 171008 229316 230664 229344
rect 171008 229304 171014 229316
rect 230658 229304 230664 229316
rect 230716 229304 230722 229356
rect 413830 229304 413836 229356
rect 413888 229344 413894 229356
rect 419994 229344 420000 229356
rect 413888 229316 420000 229344
rect 413888 229304 413894 229316
rect 419994 229304 420000 229316
rect 420052 229304 420058 229356
rect 472158 229304 472164 229356
rect 472216 229344 472222 229356
rect 472986 229344 472992 229356
rect 472216 229316 472992 229344
rect 472216 229304 472222 229316
rect 472986 229304 472992 229316
rect 473044 229304 473050 229356
rect 674104 229298 674156 229304
rect 446398 229236 446404 229288
rect 446456 229276 446462 229288
rect 448606 229276 448612 229288
rect 446456 229248 448612 229276
rect 446456 229236 446462 229248
rect 448606 229236 448612 229248
rect 448664 229236 448670 229288
rect 450262 229236 450268 229288
rect 450320 229276 450326 229288
rect 451734 229276 451740 229288
rect 450320 229248 451740 229276
rect 450320 229236 450326 229248
rect 451734 229236 451740 229248
rect 451792 229236 451798 229288
rect 495342 229236 495348 229288
rect 495400 229276 495406 229288
rect 500218 229276 500224 229288
rect 495400 229248 500224 229276
rect 495400 229236 495406 229248
rect 500218 229236 500224 229248
rect 500276 229236 500282 229288
rect 505646 229236 505652 229288
rect 505704 229276 505710 229288
rect 510614 229276 510620 229288
rect 505704 229248 510620 229276
rect 505704 229236 505710 229248
rect 510614 229236 510620 229248
rect 510672 229236 510678 229288
rect 513374 229236 513380 229288
rect 513432 229276 513438 229288
rect 519170 229276 519176 229288
rect 513432 229248 519176 229276
rect 513432 229236 513438 229248
rect 519170 229236 519176 229248
rect 519228 229236 519234 229288
rect 660942 229236 660948 229288
rect 661000 229276 661006 229288
rect 666278 229276 666284 229288
rect 661000 229248 666284 229276
rect 661000 229236 661006 229248
rect 666278 229236 666284 229248
rect 666336 229236 666342 229288
rect 123536 229180 151814 229208
rect 123536 229168 123542 229180
rect 151906 229168 151912 229220
rect 151964 229208 151970 229220
rect 155954 229208 155960 229220
rect 151964 229180 155960 229208
rect 151964 229168 151970 229180
rect 155954 229168 155960 229180
rect 156012 229168 156018 229220
rect 157242 229168 157248 229220
rect 157300 229208 157306 229220
rect 161290 229208 161296 229220
rect 157300 229180 161296 229208
rect 157300 229168 157306 229180
rect 161290 229168 161296 229180
rect 161348 229168 161354 229220
rect 161474 229168 161480 229220
rect 161532 229208 161538 229220
rect 173710 229208 173716 229220
rect 161532 229180 173716 229208
rect 161532 229168 161538 229180
rect 173710 229168 173716 229180
rect 173768 229168 173774 229220
rect 173894 229168 173900 229220
rect 173952 229208 173958 229220
rect 174814 229208 174820 229220
rect 173952 229180 174820 229208
rect 173952 229168 173958 229180
rect 174814 229168 174820 229180
rect 174872 229168 174878 229220
rect 175918 229168 175924 229220
rect 175976 229208 175982 229220
rect 180426 229208 180432 229220
rect 175976 229180 180432 229208
rect 175976 229168 175982 229180
rect 180426 229168 180432 229180
rect 180484 229168 180490 229220
rect 183370 229168 183376 229220
rect 183428 229208 183434 229220
rect 240962 229208 240968 229220
rect 183428 229180 240968 229208
rect 183428 229168 183434 229180
rect 240962 229168 240968 229180
rect 241020 229168 241026 229220
rect 423490 229100 423496 229152
rect 423548 229140 423554 229152
rect 427722 229140 427728 229152
rect 423548 229112 427728 229140
rect 423548 229100 423554 229112
rect 427722 229100 427728 229112
rect 427780 229100 427786 229152
rect 441246 229100 441252 229152
rect 441304 229140 441310 229152
rect 442074 229140 442080 229152
rect 441304 229112 442080 229140
rect 441304 229100 441310 229112
rect 442074 229100 442080 229112
rect 442132 229100 442138 229152
rect 450906 229100 450912 229152
rect 450964 229140 450970 229152
rect 452746 229140 452752 229152
rect 450964 229112 452752 229140
rect 450964 229100 450970 229112
rect 452746 229100 452752 229112
rect 452804 229100 452810 229152
rect 503714 229100 503720 229152
rect 503772 229140 503778 229152
rect 509878 229140 509884 229152
rect 503772 229112 509884 229140
rect 503772 229100 503778 229112
rect 509878 229100 509884 229112
rect 509936 229100 509942 229152
rect 515306 229100 515312 229152
rect 515364 229140 515370 229152
rect 520918 229140 520924 229152
rect 515364 229112 520924 229140
rect 515364 229100 515370 229112
rect 520918 229100 520924 229112
rect 520976 229100 520982 229152
rect 524966 229100 524972 229152
rect 525024 229140 525030 229152
rect 529934 229140 529940 229152
rect 525024 229112 529940 229140
rect 525024 229100 525030 229112
rect 529934 229100 529940 229112
rect 529992 229100 529998 229152
rect 662322 229100 662328 229152
rect 662380 229140 662386 229152
rect 666462 229140 666468 229152
rect 662380 229112 666468 229140
rect 662380 229100 662386 229112
rect 666462 229100 666468 229112
rect 666520 229100 666526 229152
rect 673546 229100 673552 229152
rect 673604 229140 673610 229152
rect 673604 229112 674038 229140
rect 673604 229100 673610 229112
rect 100662 229032 100668 229084
rect 100720 229072 100726 229084
rect 174630 229072 174636 229084
rect 100720 229044 174636 229072
rect 100720 229032 100726 229044
rect 174630 229032 174636 229044
rect 174688 229032 174694 229084
rect 174814 229032 174820 229084
rect 174872 229072 174878 229084
rect 179782 229072 179788 229084
rect 174872 229044 179788 229072
rect 174872 229032 174878 229044
rect 179782 229032 179788 229044
rect 179840 229032 179846 229084
rect 180058 229032 180064 229084
rect 180116 229072 180122 229084
rect 185578 229072 185584 229084
rect 180116 229044 185584 229072
rect 180116 229032 180122 229044
rect 185578 229032 185584 229044
rect 185636 229032 185642 229084
rect 189718 229032 189724 229084
rect 189776 229072 189782 229084
rect 189776 229044 190454 229072
rect 189776 229032 189782 229044
rect 106182 228896 106188 228948
rect 106240 228936 106246 228948
rect 173894 228936 173900 228948
rect 106240 228908 173900 228936
rect 106240 228896 106246 228908
rect 173894 228896 173900 228908
rect 173952 228896 173958 228948
rect 184934 228936 184940 228948
rect 175936 228908 184940 228936
rect 93578 228760 93584 228812
rect 93636 228800 93642 228812
rect 161428 228800 161434 228812
rect 93636 228772 161434 228800
rect 93636 228760 93642 228772
rect 161428 228760 161434 228772
rect 161486 228760 161492 228812
rect 161566 228760 161572 228812
rect 161624 228800 161630 228812
rect 161624 228772 166212 228800
rect 161624 228760 161630 228772
rect 166184 228732 166212 228772
rect 166534 228760 166540 228812
rect 166592 228800 166598 228812
rect 175936 228800 175964 228908
rect 184934 228896 184940 228908
rect 184992 228896 184998 228948
rect 185394 228896 185400 228948
rect 185452 228936 185458 228948
rect 190086 228936 190092 228948
rect 185452 228908 190092 228936
rect 185452 228896 185458 228908
rect 190086 228896 190092 228908
rect 190144 228896 190150 228948
rect 190426 228936 190454 229044
rect 192846 229032 192852 229084
rect 192904 229072 192910 229084
rect 195238 229072 195244 229084
rect 192904 229044 195244 229072
rect 192904 229032 192910 229044
rect 195238 229032 195244 229044
rect 195296 229032 195302 229084
rect 201402 229032 201408 229084
rect 201460 229072 201466 229084
rect 252554 229072 252560 229084
rect 201460 229044 252560 229072
rect 201460 229032 201466 229044
rect 252554 229032 252560 229044
rect 252612 229032 252618 229084
rect 255222 229032 255228 229084
rect 255280 229072 255286 229084
rect 295702 229072 295708 229084
rect 255280 229044 295708 229072
rect 255280 229032 255286 229044
rect 295702 229032 295708 229044
rect 295760 229032 295766 229084
rect 305546 229032 305552 229084
rect 305604 229072 305610 229084
rect 315666 229072 315672 229084
rect 305604 229044 315672 229072
rect 305604 229032 305610 229044
rect 315666 229032 315672 229044
rect 315724 229032 315730 229084
rect 326890 229032 326896 229084
rect 326948 229072 326954 229084
rect 351086 229072 351092 229084
rect 326948 229044 351092 229072
rect 326948 229032 326954 229044
rect 351086 229032 351092 229044
rect 351144 229032 351150 229084
rect 195238 228936 195244 228948
rect 190426 228908 195244 228936
rect 195238 228896 195244 228908
rect 195296 228896 195302 228948
rect 195422 228896 195428 228948
rect 195480 228936 195486 228948
rect 246758 228936 246764 228948
rect 195480 228908 246764 228936
rect 195480 228896 195486 228908
rect 246758 228896 246764 228908
rect 246816 228896 246822 228948
rect 248230 228896 248236 228948
rect 248288 228936 248294 228948
rect 291838 228936 291844 228948
rect 248288 228908 291844 228936
rect 248288 228896 248294 228908
rect 291838 228896 291844 228908
rect 291896 228896 291902 228948
rect 302142 228896 302148 228948
rect 302200 228936 302206 228948
rect 331214 228936 331220 228948
rect 302200 228908 331220 228936
rect 302200 228896 302206 228908
rect 331214 228896 331220 228908
rect 331272 228896 331278 228948
rect 506382 228896 506388 228948
rect 506440 228936 506446 228948
rect 512730 228936 512736 228948
rect 506440 228908 512736 228936
rect 506440 228896 506446 228908
rect 512730 228896 512736 228908
rect 512788 228896 512794 228948
rect 526438 228896 526444 228948
rect 526496 228936 526502 228948
rect 544010 228936 544016 228948
rect 526496 228908 544016 228936
rect 526496 228896 526502 228908
rect 544010 228896 544016 228908
rect 544068 228896 544074 228948
rect 166592 228772 175964 228800
rect 166592 228760 166598 228772
rect 176102 228760 176108 228812
rect 176160 228800 176166 228812
rect 231302 228800 231308 228812
rect 176160 228772 231308 228800
rect 176160 228760 176166 228772
rect 231302 228760 231308 228772
rect 231360 228760 231366 228812
rect 238570 228760 238576 228812
rect 238628 228800 238634 228812
rect 282822 228800 282828 228812
rect 238628 228772 282828 228800
rect 238628 228760 238634 228772
rect 282822 228760 282828 228772
rect 282880 228760 282886 228812
rect 291838 228760 291844 228812
rect 291896 228800 291902 228812
rect 300210 228800 300216 228812
rect 291896 228772 300216 228800
rect 291896 228760 291902 228772
rect 300210 228760 300216 228772
rect 300268 228760 300274 228812
rect 300670 228760 300676 228812
rect 300728 228800 300734 228812
rect 330478 228800 330484 228812
rect 300728 228772 330484 228800
rect 300728 228760 300734 228772
rect 330478 228760 330484 228772
rect 330536 228760 330542 228812
rect 376018 228760 376024 228812
rect 376076 228800 376082 228812
rect 387794 228800 387800 228812
rect 376076 228772 387800 228800
rect 376076 228760 376082 228772
rect 387794 228760 387800 228772
rect 387852 228760 387858 228812
rect 478874 228760 478880 228812
rect 478932 228800 478938 228812
rect 490374 228800 490380 228812
rect 478932 228772 490380 228800
rect 478932 228760 478938 228772
rect 490374 228760 490380 228772
rect 490432 228760 490438 228812
rect 499850 228760 499856 228812
rect 499908 228800 499914 228812
rect 518158 228800 518164 228812
rect 499908 228772 518164 228800
rect 499908 228760 499914 228772
rect 518158 228760 518164 228772
rect 518216 228760 518222 228812
rect 518526 228760 518532 228812
rect 518584 228800 518590 228812
rect 541526 228800 541532 228812
rect 518584 228772 541532 228800
rect 518584 228760 518590 228772
rect 541526 228760 541532 228772
rect 541584 228760 541590 228812
rect 166184 228704 166396 228732
rect 67542 228624 67548 228676
rect 67600 228664 67606 228676
rect 146202 228664 146208 228676
rect 67600 228636 146208 228664
rect 67600 228624 67606 228636
rect 146202 228624 146208 228636
rect 146260 228624 146266 228676
rect 165982 228664 165988 228676
rect 146956 228636 165988 228664
rect 61378 228488 61384 228540
rect 61436 228528 61442 228540
rect 61436 228500 137232 228528
rect 61436 228488 61442 228500
rect 57238 228352 57244 228404
rect 57296 228392 57302 228404
rect 136818 228392 136824 228404
rect 57296 228364 136824 228392
rect 57296 228352 57302 228364
rect 136818 228352 136824 228364
rect 136876 228352 136882 228404
rect 137204 228392 137232 228500
rect 137370 228488 137376 228540
rect 137428 228528 137434 228540
rect 146956 228528 146984 228636
rect 165982 228624 165988 228636
rect 166040 228624 166046 228676
rect 166368 228664 166396 228704
rect 181438 228664 181444 228676
rect 166368 228636 181444 228664
rect 181438 228624 181444 228636
rect 181496 228624 181502 228676
rect 181622 228624 181628 228676
rect 181680 228664 181686 228676
rect 185394 228664 185400 228676
rect 181680 228636 185400 228664
rect 181680 228624 181686 228636
rect 185394 228624 185400 228636
rect 185452 228624 185458 228676
rect 185578 228624 185584 228676
rect 185636 228664 185642 228676
rect 226150 228664 226156 228676
rect 185636 228636 226156 228664
rect 185636 228624 185642 228636
rect 226150 228624 226156 228636
rect 226208 228624 226214 228676
rect 226334 228624 226340 228676
rect 226392 228664 226398 228676
rect 272518 228664 272524 228676
rect 226392 228636 272524 228664
rect 226392 228624 226398 228636
rect 272518 228624 272524 228636
rect 272576 228624 272582 228676
rect 296622 228624 296628 228676
rect 296680 228664 296686 228676
rect 329190 228664 329196 228676
rect 296680 228636 329196 228664
rect 296680 228624 296686 228636
rect 329190 228624 329196 228636
rect 329248 228624 329254 228676
rect 336458 228624 336464 228676
rect 336516 228664 336522 228676
rect 358814 228664 358820 228676
rect 336516 228636 358820 228664
rect 336516 228624 336522 228636
rect 358814 228624 358820 228636
rect 358872 228624 358878 228676
rect 359918 228624 359924 228676
rect 359976 228664 359982 228676
rect 376846 228664 376852 228676
rect 359976 228636 376852 228664
rect 359976 228624 359982 228636
rect 376846 228624 376852 228636
rect 376904 228624 376910 228676
rect 485682 228624 485688 228676
rect 485740 228664 485746 228676
rect 498286 228664 498292 228676
rect 485740 228636 498292 228664
rect 485740 228624 485746 228636
rect 498286 228624 498292 228636
rect 498344 228624 498350 228676
rect 498562 228624 498568 228676
rect 498620 228664 498626 228676
rect 515766 228664 515772 228676
rect 498620 228636 515772 228664
rect 498620 228624 498626 228636
rect 515766 228624 515772 228636
rect 515824 228624 515830 228676
rect 517882 228624 517888 228676
rect 517940 228664 517946 228676
rect 539410 228664 539416 228676
rect 517940 228636 539416 228664
rect 517940 228624 517946 228636
rect 539410 228624 539416 228636
rect 539468 228624 539474 228676
rect 539594 228624 539600 228676
rect 539652 228664 539658 228676
rect 556982 228664 556988 228676
rect 539652 228636 556988 228664
rect 539652 228624 539658 228636
rect 556982 228624 556988 228636
rect 557040 228624 557046 228676
rect 137428 228500 146984 228528
rect 137428 228488 137434 228500
rect 147122 228488 147128 228540
rect 147180 228528 147186 228540
rect 200114 228528 200120 228540
rect 147180 228500 200120 228528
rect 147180 228488 147186 228500
rect 200114 228488 200120 228500
rect 200172 228488 200178 228540
rect 200298 228488 200304 228540
rect 200356 228528 200362 228540
rect 220998 228528 221004 228540
rect 200356 228500 221004 228528
rect 200356 228488 200362 228500
rect 220998 228488 221004 228500
rect 221056 228488 221062 228540
rect 264790 228528 264796 228540
rect 221200 228500 264796 228528
rect 137204 228364 137416 228392
rect 112990 228216 112996 228268
rect 113048 228256 113054 228268
rect 137186 228256 137192 228268
rect 113048 228228 137192 228256
rect 113048 228216 113054 228228
rect 137186 228216 137192 228228
rect 137244 228216 137250 228268
rect 137388 228256 137416 228364
rect 139302 228352 139308 228404
rect 139360 228392 139366 228404
rect 139360 228364 151814 228392
rect 139360 228352 139366 228364
rect 143074 228256 143080 228268
rect 137388 228228 143080 228256
rect 143074 228216 143080 228228
rect 143132 228216 143138 228268
rect 143442 228216 143448 228268
rect 143500 228256 143506 228268
rect 146018 228256 146024 228268
rect 143500 228228 146024 228256
rect 143500 228216 143506 228228
rect 146018 228216 146024 228228
rect 146076 228216 146082 228268
rect 146202 228216 146208 228268
rect 146260 228256 146266 228268
rect 148870 228256 148876 228268
rect 146260 228228 148876 228256
rect 146260 228216 146266 228228
rect 148870 228216 148876 228228
rect 148928 228216 148934 228268
rect 151786 228256 151814 228364
rect 153470 228352 153476 228404
rect 153528 228392 153534 228404
rect 154206 228392 154212 228404
rect 153528 228364 154212 228392
rect 153528 228352 153534 228364
rect 154206 228352 154212 228364
rect 154264 228352 154270 228404
rect 154390 228352 154396 228404
rect 154448 228392 154454 228404
rect 215846 228392 215852 228404
rect 154448 228364 215852 228392
rect 154448 228352 154454 228364
rect 215846 228352 215852 228364
rect 215904 228352 215910 228404
rect 216398 228352 216404 228404
rect 216456 228392 216462 228404
rect 221200 228392 221228 228500
rect 264790 228488 264796 228500
rect 264848 228488 264854 228540
rect 272518 228488 272524 228540
rect 272576 228528 272582 228540
rect 309870 228528 309876 228540
rect 272576 228500 309876 228528
rect 272576 228488 272582 228500
rect 309870 228488 309876 228500
rect 309928 228488 309934 228540
rect 313826 228488 313832 228540
rect 313884 228528 313890 228540
rect 320818 228528 320824 228540
rect 313884 228500 320824 228528
rect 313884 228488 313890 228500
rect 320818 228488 320824 228500
rect 320876 228488 320882 228540
rect 325418 228488 325424 228540
rect 325476 228528 325482 228540
rect 349154 228528 349160 228540
rect 325476 228500 349160 228528
rect 325476 228488 325482 228500
rect 349154 228488 349160 228500
rect 349212 228488 349218 228540
rect 350442 228488 350448 228540
rect 350500 228528 350506 228540
rect 369118 228528 369124 228540
rect 350500 228500 369124 228528
rect 350500 228488 350506 228500
rect 369118 228488 369124 228500
rect 369176 228488 369182 228540
rect 371050 228488 371056 228540
rect 371108 228528 371114 228540
rect 385218 228528 385224 228540
rect 371108 228500 385224 228528
rect 371108 228488 371114 228500
rect 385218 228488 385224 228500
rect 385276 228488 385282 228540
rect 386046 228488 386052 228540
rect 386104 228528 386110 228540
rect 397454 228528 397460 228540
rect 386104 228500 397460 228528
rect 386104 228488 386110 228500
rect 397454 228488 397460 228500
rect 397512 228488 397518 228540
rect 407758 228528 407764 228540
rect 400232 228500 407764 228528
rect 216456 228364 221228 228392
rect 216456 228352 216462 228364
rect 224770 228352 224776 228404
rect 224828 228392 224834 228404
rect 273806 228392 273812 228404
rect 224828 228364 273812 228392
rect 224828 228352 224834 228364
rect 273806 228352 273812 228364
rect 273864 228352 273870 228404
rect 285582 228352 285588 228404
rect 285640 228392 285646 228404
rect 318886 228392 318892 228404
rect 285640 228364 318892 228392
rect 285640 228352 285646 228364
rect 318886 228352 318892 228364
rect 318944 228352 318950 228404
rect 330478 228352 330484 228404
rect 330536 228392 330542 228404
rect 354950 228392 354956 228404
rect 330536 228364 354956 228392
rect 330536 228352 330542 228364
rect 354950 228352 354956 228364
rect 355008 228352 355014 228404
rect 355318 228352 355324 228404
rect 355376 228392 355382 228404
rect 372982 228392 372988 228404
rect 355376 228364 372988 228392
rect 355376 228352 355382 228364
rect 372982 228352 372988 228364
rect 373040 228352 373046 228404
rect 373442 228352 373448 228404
rect 373500 228392 373506 228404
rect 387150 228392 387156 228404
rect 373500 228364 387156 228392
rect 373500 228352 373506 228364
rect 387150 228352 387156 228364
rect 387208 228352 387214 228404
rect 390002 228352 390008 228404
rect 390060 228392 390066 228404
rect 400030 228392 400036 228404
rect 390060 228364 400036 228392
rect 390060 228352 390066 228364
rect 400030 228352 400036 228364
rect 400088 228352 400094 228404
rect 205542 228256 205548 228268
rect 151786 228228 205548 228256
rect 205542 228216 205548 228228
rect 205600 228216 205606 228268
rect 205726 228216 205732 228268
rect 205784 228256 205790 228268
rect 257062 228256 257068 228268
rect 205784 228228 257068 228256
rect 205784 228216 205790 228228
rect 257062 228216 257068 228228
rect 257120 228216 257126 228268
rect 257614 228216 257620 228268
rect 257672 228256 257678 228268
rect 296346 228256 296352 228268
rect 257672 228228 296352 228256
rect 257672 228216 257678 228228
rect 296346 228216 296352 228228
rect 296404 228216 296410 228268
rect 400232 228256 400260 228500
rect 407758 228488 407764 228500
rect 407816 228488 407822 228540
rect 409782 228488 409788 228540
rect 409840 228528 409846 228540
rect 415486 228528 415492 228540
rect 409840 228500 415492 228528
rect 409840 228488 409846 228500
rect 415486 228488 415492 228500
rect 415544 228488 415550 228540
rect 485038 228488 485044 228540
rect 485096 228528 485102 228540
rect 498654 228528 498660 228540
rect 485096 228500 498660 228528
rect 485096 228488 485102 228500
rect 498654 228488 498660 228500
rect 498712 228488 498718 228540
rect 502426 228488 502432 228540
rect 502484 228528 502490 228540
rect 521102 228528 521108 228540
rect 502484 228500 521108 228528
rect 502484 228488 502490 228500
rect 521102 228488 521108 228500
rect 521160 228488 521166 228540
rect 527542 228488 527548 228540
rect 527600 228528 527606 228540
rect 553302 228528 553308 228540
rect 527600 228500 553308 228528
rect 527600 228488 527606 228500
rect 553302 228488 553308 228500
rect 553360 228488 553366 228540
rect 556798 228488 556804 228540
rect 556856 228528 556862 228540
rect 570598 228528 570604 228540
rect 556856 228500 570604 228528
rect 556856 228488 556862 228500
rect 570598 228488 570604 228500
rect 570656 228488 570662 228540
rect 402790 228352 402796 228404
rect 402848 228392 402854 228404
rect 411622 228392 411628 228404
rect 402848 228364 411628 228392
rect 402848 228352 402854 228364
rect 411622 228352 411628 228364
rect 411680 228352 411686 228404
rect 474458 228352 474464 228404
rect 474516 228392 474522 228404
rect 484486 228392 484492 228404
rect 474516 228364 484492 228392
rect 474516 228352 474522 228364
rect 484486 228352 484492 228364
rect 484544 228352 484550 228404
rect 490190 228352 490196 228404
rect 490248 228392 490254 228404
rect 505186 228392 505192 228404
rect 490248 228364 505192 228392
rect 490248 228352 490254 228364
rect 505186 228352 505192 228364
rect 505244 228352 505250 228404
rect 512086 228352 512092 228404
rect 512144 228392 512150 228404
rect 532970 228392 532976 228404
rect 512144 228364 532976 228392
rect 512144 228352 512150 228364
rect 532970 228352 532976 228364
rect 533028 228352 533034 228404
rect 537202 228352 537208 228404
rect 537260 228392 537266 228404
rect 565630 228392 565636 228404
rect 537260 228364 565636 228392
rect 537260 228352 537266 228364
rect 565630 228352 565636 228364
rect 565688 228352 565694 228404
rect 400140 228228 400260 228256
rect 400140 228132 400168 228228
rect 539410 228216 539416 228268
rect 539468 228256 539474 228268
rect 540790 228256 540796 228268
rect 539468 228228 540796 228256
rect 539468 228216 539474 228228
rect 540790 228216 540796 228228
rect 540848 228216 540854 228268
rect 119982 228080 119988 228132
rect 120040 228120 120046 228132
rect 181254 228120 181260 228132
rect 120040 228092 181260 228120
rect 120040 228080 120046 228092
rect 181254 228080 181260 228092
rect 181312 228080 181318 228132
rect 181438 228080 181444 228132
rect 181496 228120 181502 228132
rect 181496 228092 193076 228120
rect 181496 228080 181502 228092
rect 126698 227944 126704 227996
rect 126756 227984 126762 227996
rect 192846 227984 192852 227996
rect 126756 227956 192852 227984
rect 126756 227944 126762 227956
rect 192846 227944 192852 227956
rect 192904 227944 192910 227996
rect 193048 227984 193076 228092
rect 195238 228080 195244 228132
rect 195296 228120 195302 228132
rect 239030 228120 239036 228132
rect 195296 228092 239036 228120
rect 195296 228080 195302 228092
rect 239030 228080 239036 228092
rect 239088 228080 239094 228132
rect 246298 228080 246304 228132
rect 246356 228120 246362 228132
rect 253842 228120 253848 228132
rect 246356 228092 253848 228120
rect 246356 228080 246362 228092
rect 253842 228080 253848 228092
rect 253900 228080 253906 228132
rect 268930 228080 268936 228132
rect 268988 228120 268994 228132
rect 306006 228120 306012 228132
rect 268988 228092 306012 228120
rect 268988 228080 268994 228092
rect 306006 228080 306012 228092
rect 306064 228080 306070 228132
rect 400122 228080 400128 228132
rect 400180 228080 400186 228132
rect 415026 228012 415032 228064
rect 415084 228052 415090 228064
rect 421926 228052 421932 228064
rect 415084 228024 421932 228052
rect 415084 228012 415090 228024
rect 421926 228012 421932 228024
rect 421984 228012 421990 228064
rect 200298 227984 200304 227996
rect 193048 227956 200304 227984
rect 200298 227944 200304 227956
rect 200356 227944 200362 227996
rect 210418 227944 210424 227996
rect 210476 227984 210482 227996
rect 238386 227984 238392 227996
rect 210476 227956 238392 227984
rect 210476 227944 210482 227956
rect 238386 227944 238392 227956
rect 238444 227944 238450 227996
rect 416682 227876 416688 227928
rect 416740 227916 416746 227928
rect 420638 227916 420644 227928
rect 416740 227888 420644 227916
rect 416740 227876 416746 227888
rect 420638 227876 420644 227888
rect 420696 227876 420702 227928
rect 447042 227876 447048 227928
rect 447100 227916 447106 227928
rect 450538 227916 450544 227928
rect 447100 227888 450544 227916
rect 447100 227876 447106 227888
rect 450538 227876 450544 227888
rect 450596 227876 450602 227928
rect 88242 227808 88248 227860
rect 88300 227848 88306 227860
rect 95234 227848 95240 227860
rect 88300 227820 95240 227848
rect 88300 227808 88306 227820
rect 95234 227808 95240 227820
rect 95292 227808 95298 227860
rect 133506 227808 133512 227860
rect 133564 227848 133570 227860
rect 136634 227848 136640 227860
rect 133564 227820 136640 227848
rect 133564 227808 133570 227820
rect 136634 227808 136640 227820
rect 136692 227808 136698 227860
rect 136818 227808 136824 227860
rect 136876 227848 136882 227860
rect 141142 227848 141148 227860
rect 136876 227820 141148 227848
rect 136876 227808 136882 227820
rect 141142 227808 141148 227820
rect 141200 227808 141206 227860
rect 141510 227808 141516 227860
rect 141568 227848 141574 227860
rect 200482 227848 200488 227860
rect 141568 227820 200488 227848
rect 141568 227808 141574 227820
rect 200482 227808 200488 227820
rect 200540 227808 200546 227860
rect 200666 227808 200672 227860
rect 200724 227848 200730 227860
rect 210234 227848 210240 227860
rect 200724 227820 210240 227848
rect 200724 227808 200730 227820
rect 210234 227808 210240 227820
rect 210292 227808 210298 227860
rect 409046 227740 409052 227792
rect 409104 227780 409110 227792
rect 410334 227780 410340 227792
rect 409104 227752 410340 227780
rect 409104 227740 409110 227752
rect 410334 227740 410340 227752
rect 410392 227740 410398 227792
rect 411898 227740 411904 227792
rect 411956 227780 411962 227792
rect 413554 227780 413560 227792
rect 411956 227752 413560 227780
rect 411956 227740 411962 227752
rect 413554 227740 413560 227752
rect 413612 227740 413618 227792
rect 420638 227740 420644 227792
rect 420696 227780 420702 227792
rect 423858 227780 423864 227792
rect 420696 227752 423864 227780
rect 420696 227740 420702 227752
rect 423858 227740 423864 227752
rect 423916 227740 423922 227792
rect 471514 227740 471520 227792
rect 471572 227780 471578 227792
rect 479518 227780 479524 227792
rect 471572 227752 479524 227780
rect 471572 227740 471578 227752
rect 479518 227740 479524 227752
rect 479576 227740 479582 227792
rect 662046 227740 662052 227792
rect 662104 227780 662110 227792
rect 663886 227780 663892 227792
rect 662104 227752 663892 227780
rect 662104 227740 662110 227752
rect 663886 227740 663892 227752
rect 663944 227740 663950 227792
rect 42426 227672 42432 227724
rect 42484 227712 42490 227724
rect 43070 227712 43076 227724
rect 42484 227684 43076 227712
rect 42484 227672 42490 227684
rect 43070 227672 43076 227684
rect 43128 227672 43134 227724
rect 64782 227672 64788 227724
rect 64840 227712 64846 227724
rect 110322 227712 110328 227724
rect 64840 227684 110328 227712
rect 64840 227672 64846 227684
rect 110322 227672 110328 227684
rect 110380 227672 110386 227724
rect 110506 227672 110512 227724
rect 110564 227712 110570 227724
rect 182358 227712 182364 227724
rect 110564 227684 182364 227712
rect 110564 227672 110570 227684
rect 182358 227672 182364 227684
rect 182416 227672 182422 227724
rect 185394 227672 185400 227724
rect 185452 227712 185458 227724
rect 192662 227712 192668 227724
rect 185452 227684 192668 227712
rect 185452 227672 185458 227684
rect 192662 227672 192668 227684
rect 192720 227672 192726 227724
rect 214374 227712 214380 227724
rect 200086 227684 214380 227712
rect 60642 227536 60648 227588
rect 60700 227576 60706 227588
rect 102134 227576 102140 227588
rect 60700 227548 102140 227576
rect 60700 227536 60706 227548
rect 102134 227536 102140 227548
rect 102192 227536 102198 227588
rect 103422 227536 103428 227588
rect 103480 227576 103486 227588
rect 175366 227576 175372 227588
rect 103480 227548 175372 227576
rect 103480 227536 103486 227548
rect 175366 227536 175372 227548
rect 175424 227536 175430 227588
rect 181530 227536 181536 227588
rect 181588 227576 181594 227588
rect 181588 227548 185808 227576
rect 181588 227536 181594 227548
rect 175918 227508 175924 227520
rect 175660 227480 175924 227508
rect 96430 227400 96436 227452
rect 96488 227440 96494 227452
rect 170766 227440 170772 227452
rect 96488 227412 170772 227440
rect 96488 227400 96494 227412
rect 170766 227400 170772 227412
rect 170824 227400 170830 227452
rect 171088 227400 171094 227452
rect 171146 227440 171152 227452
rect 175660 227440 175688 227480
rect 175918 227468 175924 227480
rect 175976 227468 175982 227520
rect 185578 227440 185584 227452
rect 171146 227412 175688 227440
rect 176304 227412 185584 227440
rect 171146 227400 171152 227412
rect 176304 227372 176332 227412
rect 185578 227400 185584 227412
rect 185636 227400 185642 227452
rect 185780 227440 185808 227548
rect 186130 227536 186136 227588
rect 186188 227576 186194 227588
rect 200086 227576 200114 227684
rect 214374 227672 214380 227684
rect 214432 227672 214438 227724
rect 214742 227672 214748 227724
rect 214800 227712 214806 227724
rect 262214 227712 262220 227724
rect 214800 227684 262220 227712
rect 214800 227672 214806 227684
rect 262214 227672 262220 227684
rect 262272 227672 262278 227724
rect 277026 227672 277032 227724
rect 277084 227712 277090 227724
rect 311802 227712 311808 227724
rect 277084 227684 311808 227712
rect 277084 227672 277090 227684
rect 311802 227672 311808 227684
rect 311860 227672 311866 227724
rect 465902 227604 465908 227656
rect 465960 227644 465966 227656
rect 469858 227644 469864 227656
rect 465960 227616 469864 227644
rect 465960 227604 465966 227616
rect 469858 227604 469864 227616
rect 469916 227604 469922 227656
rect 186188 227548 200114 227576
rect 186188 227536 186194 227548
rect 200206 227536 200212 227588
rect 200264 227576 200270 227588
rect 251910 227576 251916 227588
rect 200264 227548 251916 227576
rect 200264 227536 200270 227548
rect 251910 227536 251916 227548
rect 251968 227536 251974 227588
rect 259270 227536 259276 227588
rect 259328 227576 259334 227588
rect 298278 227576 298284 227588
rect 259328 227548 298284 227576
rect 259328 227536 259334 227548
rect 298278 227536 298284 227548
rect 298336 227536 298342 227588
rect 301498 227536 301504 227588
rect 301556 227576 301562 227588
rect 308582 227576 308588 227588
rect 301556 227548 308588 227576
rect 301556 227536 301562 227548
rect 308582 227536 308588 227548
rect 308640 227536 308646 227588
rect 524598 227536 524604 227588
rect 524656 227576 524662 227588
rect 539962 227576 539968 227588
rect 524656 227548 539968 227576
rect 524656 227536 524662 227548
rect 539962 227536 539968 227548
rect 540020 227536 540026 227588
rect 219894 227440 219900 227452
rect 185780 227412 219900 227440
rect 219894 227400 219900 227412
rect 219952 227400 219958 227452
rect 220078 227400 220084 227452
rect 220136 227440 220142 227452
rect 241606 227440 241612 227452
rect 220136 227412 241612 227440
rect 220136 227400 220142 227412
rect 241606 227400 241612 227412
rect 241664 227400 241670 227452
rect 257798 227400 257804 227452
rect 257856 227440 257862 227452
rect 299566 227440 299572 227452
rect 257856 227412 299572 227440
rect 257856 227400 257862 227412
rect 299566 227400 299572 227412
rect 299624 227400 299630 227452
rect 304902 227400 304908 227452
rect 304960 227440 304966 227452
rect 333698 227440 333704 227452
rect 304960 227412 333704 227440
rect 304960 227400 304966 227412
rect 333698 227400 333704 227412
rect 333756 227400 333762 227452
rect 333882 227400 333888 227452
rect 333940 227440 333946 227452
rect 356238 227440 356244 227452
rect 333940 227412 356244 227440
rect 333940 227400 333946 227412
rect 356238 227400 356244 227412
rect 356296 227400 356302 227452
rect 357066 227400 357072 227452
rect 357124 227440 357130 227452
rect 374270 227440 374276 227452
rect 357124 227412 374276 227440
rect 357124 227400 357130 227412
rect 374270 227400 374276 227412
rect 374328 227400 374334 227452
rect 514018 227400 514024 227452
rect 514076 227440 514082 227452
rect 535730 227440 535736 227452
rect 514076 227412 535736 227440
rect 514076 227400 514082 227412
rect 535730 227400 535736 227412
rect 535788 227400 535794 227452
rect 538306 227400 538312 227452
rect 538364 227440 538370 227452
rect 556062 227440 556068 227452
rect 538364 227412 556068 227440
rect 538364 227400 538370 227412
rect 556062 227400 556068 227412
rect 556120 227400 556126 227452
rect 176120 227344 176332 227372
rect 89622 227264 89628 227316
rect 89680 227304 89686 227316
rect 161428 227304 161434 227316
rect 89680 227276 161434 227304
rect 89680 227264 89686 227276
rect 161428 227264 161434 227276
rect 161486 227264 161492 227316
rect 161566 227264 161572 227316
rect 161624 227304 161630 227316
rect 176120 227304 176148 227344
rect 161624 227276 176148 227304
rect 161624 227264 161630 227276
rect 176746 227264 176752 227316
rect 176804 227304 176810 227316
rect 228726 227304 228732 227316
rect 176804 227276 228732 227304
rect 176804 227264 176810 227276
rect 228726 227264 228732 227276
rect 228784 227264 228790 227316
rect 235810 227264 235816 227316
rect 235868 227304 235874 227316
rect 280246 227304 280252 227316
rect 235868 227276 280252 227304
rect 235868 227264 235874 227276
rect 280246 227264 280252 227276
rect 280304 227264 280310 227316
rect 306190 227264 306196 227316
rect 306248 227304 306254 227316
rect 336918 227304 336924 227316
rect 306248 227276 336924 227304
rect 306248 227264 306254 227276
rect 336918 227264 336924 227276
rect 336976 227264 336982 227316
rect 340690 227264 340696 227316
rect 340748 227304 340754 227316
rect 361390 227304 361396 227316
rect 340748 227276 361396 227304
rect 340748 227264 340754 227276
rect 361390 227264 361396 227276
rect 361448 227264 361454 227316
rect 382090 227264 382096 227316
rect 382148 227304 382154 227316
rect 392946 227304 392952 227316
rect 382148 227276 392952 227304
rect 382148 227264 382154 227276
rect 392946 227264 392952 227276
rect 393004 227264 393010 227316
rect 402606 227304 402612 227316
rect 393286 227276 402612 227304
rect 63034 227128 63040 227180
rect 63092 227168 63098 227180
rect 144822 227168 144828 227180
rect 63092 227140 144828 227168
rect 63092 227128 63098 227140
rect 144822 227128 144828 227140
rect 144880 227128 144886 227180
rect 150066 227128 150072 227180
rect 150124 227168 150130 227180
rect 213362 227168 213368 227180
rect 150124 227140 213368 227168
rect 150124 227128 150130 227140
rect 213362 227128 213368 227140
rect 213420 227128 213426 227180
rect 214374 227128 214380 227180
rect 214432 227168 214438 227180
rect 220078 227168 220084 227180
rect 214432 227140 220084 227168
rect 214432 227128 214438 227140
rect 220078 227128 220084 227140
rect 220136 227128 220142 227180
rect 220262 227128 220268 227180
rect 220320 227168 220326 227180
rect 223574 227168 223580 227180
rect 220320 227140 223580 227168
rect 220320 227128 220326 227140
rect 223574 227128 223580 227140
rect 223632 227128 223638 227180
rect 262858 227168 262864 227180
rect 224926 227140 262864 227168
rect 56502 226992 56508 227044
rect 56560 227032 56566 227044
rect 142430 227032 142436 227044
rect 56560 227004 142436 227032
rect 56560 226992 56566 227004
rect 142430 226992 142436 227004
rect 142488 226992 142494 227044
rect 143258 226992 143264 227044
rect 143316 227032 143322 227044
rect 208118 227032 208124 227044
rect 143316 227004 208124 227032
rect 143316 226992 143322 227004
rect 208118 226992 208124 227004
rect 208176 226992 208182 227044
rect 218422 227032 218428 227044
rect 209746 227004 218428 227032
rect 122742 226856 122748 226908
rect 122800 226896 122806 226908
rect 185394 226896 185400 226908
rect 122800 226868 185400 226896
rect 122800 226856 122806 226868
rect 185394 226856 185400 226868
rect 185452 226856 185458 226908
rect 185578 226856 185584 226908
rect 185636 226896 185642 226908
rect 209746 226896 209774 227004
rect 218422 226992 218428 227004
rect 218480 226992 218486 227044
rect 224926 227032 224954 227140
rect 262858 227128 262864 227140
rect 262916 227128 262922 227180
rect 263502 227128 263508 227180
rect 263560 227168 263566 227180
rect 277210 227168 277216 227180
rect 263560 227140 277216 227168
rect 263560 227128 263566 227140
rect 277210 227128 277216 227140
rect 277268 227128 277274 227180
rect 281350 227128 281356 227180
rect 281408 227168 281414 227180
rect 317598 227168 317604 227180
rect 281408 227140 317604 227168
rect 281408 227128 281414 227140
rect 317598 227128 317604 227140
rect 317656 227128 317662 227180
rect 322842 227128 322848 227180
rect 322900 227168 322906 227180
rect 349798 227168 349804 227180
rect 322900 227140 349804 227168
rect 322900 227128 322906 227140
rect 349798 227128 349804 227140
rect 349856 227128 349862 227180
rect 355870 227128 355876 227180
rect 355928 227168 355934 227180
rect 375558 227168 375564 227180
rect 355928 227140 375564 227168
rect 355928 227128 355934 227140
rect 375558 227128 375564 227140
rect 375616 227128 375622 227180
rect 376662 227128 376668 227180
rect 376720 227168 376726 227180
rect 389726 227168 389732 227180
rect 376720 227140 389732 227168
rect 376720 227128 376726 227140
rect 389726 227128 389732 227140
rect 389784 227128 389790 227180
rect 393130 227128 393136 227180
rect 393188 227168 393194 227180
rect 393286 227168 393314 227276
rect 402606 227264 402612 227276
rect 402664 227264 402670 227316
rect 494698 227264 494704 227316
rect 494756 227304 494762 227316
rect 494756 227276 504404 227304
rect 494756 227264 494762 227276
rect 393188 227140 393314 227168
rect 393188 227128 393194 227140
rect 402238 227128 402244 227180
rect 402296 227168 402302 227180
rect 408402 227168 408408 227180
rect 402296 227140 408408 227168
rect 402296 227128 402302 227140
rect 408402 227128 408408 227140
rect 408460 227128 408466 227180
rect 478598 227128 478604 227180
rect 478656 227168 478662 227180
rect 486786 227168 486792 227180
rect 478656 227140 486792 227168
rect 478656 227128 478662 227140
rect 486786 227128 486792 227140
rect 486844 227128 486850 227180
rect 489546 227128 489552 227180
rect 489604 227168 489610 227180
rect 504174 227168 504180 227180
rect 489604 227140 504180 227168
rect 489604 227128 489610 227140
rect 504174 227128 504180 227140
rect 504232 227128 504238 227180
rect 220096 227004 224954 227032
rect 185636 226868 209774 226896
rect 185636 226856 185642 226868
rect 213822 226856 213828 226908
rect 213880 226896 213886 226908
rect 220096 226896 220124 227004
rect 228910 226992 228916 227044
rect 228968 227032 228974 227044
rect 271230 227032 271236 227044
rect 228968 227004 271236 227032
rect 228968 226992 228974 227004
rect 271230 226992 271236 227004
rect 271288 226992 271294 227044
rect 271782 226992 271788 227044
rect 271840 227032 271846 227044
rect 301498 227032 301504 227044
rect 271840 227004 301504 227032
rect 271840 226992 271846 227004
rect 301498 226992 301504 227004
rect 301556 226992 301562 227044
rect 310422 226992 310428 227044
rect 310480 227032 310486 227044
rect 338206 227032 338212 227044
rect 310480 227004 338212 227032
rect 310480 226992 310486 227004
rect 338206 226992 338212 227004
rect 338264 226992 338270 227044
rect 338666 226992 338672 227044
rect 338724 227032 338730 227044
rect 360102 227032 360108 227044
rect 338724 227004 360108 227032
rect 338724 226992 338730 227004
rect 360102 226992 360108 227004
rect 360160 226992 360166 227044
rect 362770 226992 362776 227044
rect 362828 227032 362834 227044
rect 379422 227032 379428 227044
rect 362828 227004 379428 227032
rect 362828 226992 362834 227004
rect 379422 226992 379428 227004
rect 379480 226992 379486 227044
rect 391842 226992 391848 227044
rect 391900 227032 391906 227044
rect 403526 227032 403532 227044
rect 391900 227004 403532 227032
rect 391900 226992 391906 227004
rect 403526 226992 403532 227004
rect 403584 226992 403590 227044
rect 412542 226992 412548 227044
rect 412600 227032 412606 227044
rect 419350 227032 419356 227044
rect 412600 227004 419356 227032
rect 412600 226992 412606 227004
rect 419350 226992 419356 227004
rect 419408 226992 419414 227044
rect 486970 226992 486976 227044
rect 487028 227032 487034 227044
rect 500954 227032 500960 227044
rect 487028 227004 500960 227032
rect 487028 226992 487034 227004
rect 500954 226992 500960 227004
rect 501012 226992 501018 227044
rect 213880 226868 220124 226896
rect 213880 226856 213886 226868
rect 220262 226856 220268 226908
rect 220320 226896 220326 226908
rect 267366 226896 267372 226908
rect 220320 226868 267372 226896
rect 220320 226856 220326 226868
rect 267366 226856 267372 226868
rect 267424 226856 267430 226908
rect 293770 226856 293776 226908
rect 293828 226896 293834 226908
rect 324958 226896 324964 226908
rect 293828 226868 324964 226896
rect 293828 226856 293834 226868
rect 324958 226856 324964 226868
rect 325016 226856 325022 226908
rect 504376 226896 504404 227276
rect 510614 227264 510620 227316
rect 510672 227304 510678 227316
rect 524414 227304 524420 227316
rect 510672 227276 524420 227304
rect 510672 227264 510678 227276
rect 524414 227264 524420 227276
rect 524472 227264 524478 227316
rect 526254 227264 526260 227316
rect 526312 227304 526318 227316
rect 550910 227304 550916 227316
rect 526312 227276 550916 227304
rect 526312 227264 526318 227276
rect 550910 227264 550916 227276
rect 550968 227264 550974 227316
rect 506198 227128 506204 227180
rect 506256 227168 506262 227180
rect 525978 227168 525984 227180
rect 506256 227140 525984 227168
rect 506256 227128 506262 227140
rect 525978 227128 525984 227140
rect 526036 227128 526042 227180
rect 533338 227128 533344 227180
rect 533396 227168 533402 227180
rect 560938 227168 560944 227180
rect 533396 227140 560944 227168
rect 533396 227128 533402 227140
rect 560938 227128 560944 227140
rect 560996 227128 561002 227180
rect 505002 226992 505008 227044
rect 505060 227032 505066 227044
rect 523034 227032 523040 227044
rect 505060 227004 523040 227032
rect 505060 226992 505066 227004
rect 523034 226992 523040 227004
rect 523092 226992 523098 227044
rect 523678 226992 523684 227044
rect 523736 227032 523742 227044
rect 548334 227032 548340 227044
rect 523736 227004 548340 227032
rect 523736 226992 523742 227004
rect 548334 226992 548340 227004
rect 548392 226992 548398 227044
rect 555418 226992 555424 227044
rect 555476 227032 555482 227044
rect 633710 227032 633716 227044
rect 555476 227004 633716 227032
rect 555476 226992 555482 227004
rect 633710 226992 633716 227004
rect 633768 226992 633774 227044
rect 672810 227032 672816 227044
rect 669286 227004 672816 227032
rect 668578 226924 668584 226976
rect 668636 226964 668642 226976
rect 669286 226964 669314 227004
rect 672810 226992 672816 227004
rect 672868 226992 672874 227044
rect 668636 226936 669314 226964
rect 668636 226924 668642 226936
rect 510982 226896 510988 226908
rect 504376 226868 510988 226896
rect 510982 226856 510988 226868
rect 511040 226856 511046 226908
rect 676030 226788 676036 226840
rect 676088 226828 676094 226840
rect 678238 226828 678244 226840
rect 676088 226800 678244 226828
rect 676088 226788 676094 226800
rect 678238 226788 678244 226800
rect 678296 226788 678302 226840
rect 117222 226720 117228 226772
rect 117280 226760 117286 226772
rect 187510 226760 187516 226772
rect 117280 226732 187516 226760
rect 117280 226720 117286 226732
rect 187510 226720 187516 226732
rect 187568 226720 187574 226772
rect 189994 226720 190000 226772
rect 190052 226760 190058 226772
rect 233878 226760 233884 226772
rect 190052 226732 233884 226760
rect 190052 226720 190058 226732
rect 233878 226720 233884 226732
rect 233936 226720 233942 226772
rect 249610 226720 249616 226772
rect 249668 226760 249674 226772
rect 290550 226760 290556 226772
rect 249668 226732 290556 226760
rect 249668 226720 249674 226732
rect 290550 226720 290556 226732
rect 290608 226720 290614 226772
rect 243446 226652 243452 226704
rect 243504 226692 243510 226704
rect 248690 226692 248696 226704
rect 243504 226664 248696 226692
rect 243504 226652 243510 226664
rect 248690 226652 248696 226664
rect 248748 226652 248754 226704
rect 129550 226584 129556 226636
rect 129608 226624 129614 226636
rect 197354 226624 197360 226636
rect 129608 226596 197360 226624
rect 129608 226584 129614 226596
rect 197354 226584 197360 226596
rect 197412 226584 197418 226636
rect 203518 226584 203524 226636
rect 203576 226624 203582 226636
rect 203576 226596 215294 226624
rect 203576 226584 203582 226596
rect 136542 226448 136548 226500
rect 136600 226488 136606 226500
rect 141602 226488 141608 226500
rect 136600 226460 141608 226488
rect 136600 226448 136606 226460
rect 141602 226448 141608 226460
rect 141660 226448 141666 226500
rect 142246 226448 142252 226500
rect 142304 226488 142310 226500
rect 202966 226488 202972 226500
rect 142304 226460 202972 226488
rect 142304 226448 142310 226460
rect 202966 226448 202972 226460
rect 203024 226448 203030 226500
rect 212166 226448 212172 226500
rect 212224 226488 212230 226500
rect 214742 226488 214748 226500
rect 212224 226460 214748 226488
rect 212224 226448 212230 226460
rect 214742 226448 214748 226460
rect 214800 226448 214806 226500
rect 215266 226488 215294 226596
rect 219342 226584 219348 226636
rect 219400 226624 219406 226636
rect 220262 226624 220268 226636
rect 219400 226596 220268 226624
rect 219400 226584 219406 226596
rect 220262 226584 220268 226596
rect 220320 226584 220326 226636
rect 222930 226624 222936 226636
rect 220464 226596 222936 226624
rect 220464 226488 220492 226596
rect 222930 226584 222936 226596
rect 222988 226584 222994 226636
rect 231026 226584 231032 226636
rect 231084 226624 231090 226636
rect 243262 226624 243268 226636
rect 231084 226596 243268 226624
rect 231084 226584 231090 226596
rect 243262 226584 243268 226596
rect 243320 226584 243326 226636
rect 264238 226516 264244 226568
rect 264296 226556 264302 226568
rect 269298 226556 269304 226568
rect 264296 226528 269304 226556
rect 264296 226516 264302 226528
rect 269298 226516 269304 226528
rect 269356 226516 269362 226568
rect 673086 226556 673092 226568
rect 672842 226528 673092 226556
rect 673086 226516 673092 226528
rect 673144 226516 673150 226568
rect 215266 226460 220492 226488
rect 221826 226448 221832 226500
rect 221884 226488 221890 226500
rect 228910 226488 228916 226500
rect 221884 226460 228916 226488
rect 221884 226448 221890 226460
rect 228910 226448 228916 226460
rect 228968 226448 228974 226500
rect 351086 226448 351092 226500
rect 351144 226488 351150 226500
rect 353018 226488 353024 226500
rect 351144 226460 353024 226488
rect 351144 226448 351150 226460
rect 353018 226448 353024 226460
rect 353076 226448 353082 226500
rect 403986 226448 403992 226500
rect 404044 226488 404050 226500
rect 412266 226488 412272 226500
rect 404044 226460 412272 226488
rect 404044 226448 404050 226460
rect 412266 226448 412272 226460
rect 412324 226448 412330 226500
rect 474734 226448 474740 226500
rect 474792 226488 474798 226500
rect 482738 226488 482744 226500
rect 474792 226460 482744 226488
rect 474792 226448 474798 226460
rect 482738 226448 482744 226460
rect 482796 226448 482802 226500
rect 672724 226432 672776 226438
rect 141786 226380 141792 226432
rect 141844 226420 141850 226432
rect 142108 226420 142114 226432
rect 141844 226392 142114 226420
rect 141844 226380 141850 226392
rect 142108 226380 142114 226392
rect 142166 226380 142172 226432
rect 271138 226380 271144 226432
rect 271196 226420 271202 226432
rect 279602 226420 279608 226432
rect 271196 226392 279608 226420
rect 271196 226380 271202 226392
rect 279602 226380 279608 226392
rect 279660 226380 279666 226432
rect 672724 226374 672776 226380
rect 350258 226312 350264 226364
rect 350316 226352 350322 226364
rect 351730 226352 351736 226364
rect 350316 226324 351736 226352
rect 350316 226312 350322 226324
rect 351730 226312 351736 226324
rect 351788 226312 351794 226364
rect 388530 226312 388536 226364
rect 388588 226352 388594 226364
rect 391658 226352 391664 226364
rect 388588 226324 391664 226352
rect 388588 226312 388594 226324
rect 391658 226312 391664 226324
rect 391716 226312 391722 226364
rect 407758 226312 407764 226364
rect 407816 226352 407822 226364
rect 408678 226352 408684 226364
rect 407816 226324 408684 226352
rect 407816 226312 407822 226324
rect 408678 226312 408684 226324
rect 408736 226312 408742 226364
rect 481634 226312 481640 226364
rect 481692 226352 481698 226364
rect 487798 226352 487804 226364
rect 481692 226324 487804 226352
rect 481692 226312 481698 226324
rect 487798 226312 487804 226324
rect 487856 226312 487862 226364
rect 122558 226244 122564 226296
rect 122616 226284 122622 226296
rect 193950 226284 193956 226296
rect 122616 226256 193956 226284
rect 122616 226244 122622 226256
rect 193950 226244 193956 226256
rect 194008 226244 194014 226296
rect 194134 226244 194140 226296
rect 194192 226284 194198 226296
rect 244182 226284 244188 226296
rect 194192 226256 244188 226284
rect 194192 226244 194198 226256
rect 244182 226244 244188 226256
rect 244240 226244 244246 226296
rect 286318 226244 286324 226296
rect 286376 226284 286382 226296
rect 289906 226284 289912 226296
rect 286376 226256 289912 226284
rect 286376 226244 286382 226256
rect 289906 226244 289912 226256
rect 289964 226244 289970 226296
rect 291010 226244 291016 226296
rect 291068 226284 291074 226296
rect 322106 226284 322112 226296
rect 291068 226256 322112 226284
rect 291068 226244 291074 226256
rect 322106 226244 322112 226256
rect 322164 226244 322170 226296
rect 458634 226244 458640 226296
rect 458692 226284 458698 226296
rect 462958 226284 462964 226296
rect 458692 226256 462964 226284
rect 458692 226244 458698 226256
rect 462958 226244 462964 226256
rect 463016 226244 463022 226296
rect 672604 226160 672656 226166
rect 127618 226108 127624 226160
rect 127676 226148 127682 226160
rect 142108 226148 142114 226160
rect 127676 226120 142114 226148
rect 127676 226108 127682 226120
rect 142108 226108 142114 226120
rect 142166 226108 142172 226160
rect 142246 226108 142252 226160
rect 142304 226148 142310 226160
rect 203702 226148 203708 226160
rect 142304 226120 203708 226148
rect 142304 226108 142310 226120
rect 203702 226108 203708 226120
rect 203760 226108 203766 226160
rect 203886 226108 203892 226160
rect 203944 226148 203950 226160
rect 203944 226120 214604 226148
rect 203944 226108 203950 226120
rect 72418 225972 72424 226024
rect 72476 226012 72482 226024
rect 147582 226012 147588 226024
rect 72476 225984 147588 226012
rect 72476 225972 72482 225984
rect 147582 225972 147588 225984
rect 147640 225972 147646 226024
rect 147766 225972 147772 226024
rect 147824 226012 147830 226024
rect 149790 226012 149796 226024
rect 147824 225984 149796 226012
rect 147824 225972 147830 225984
rect 149790 225972 149796 225984
rect 149848 225972 149854 226024
rect 151906 225972 151912 226024
rect 151964 226012 151970 226024
rect 214374 226012 214380 226024
rect 151964 225984 214380 226012
rect 151964 225972 151970 225984
rect 214374 225972 214380 225984
rect 214432 225972 214438 226024
rect 214576 226012 214604 226120
rect 214742 226108 214748 226160
rect 214800 226148 214806 226160
rect 259638 226148 259644 226160
rect 214800 226120 259644 226148
rect 214800 226108 214806 226120
rect 259638 226108 259644 226120
rect 259696 226108 259702 226160
rect 261846 226108 261852 226160
rect 261904 226148 261910 226160
rect 300854 226148 300860 226160
rect 261904 226120 300860 226148
rect 261904 226108 261910 226120
rect 300854 226108 300860 226120
rect 300912 226108 300918 226160
rect 309042 226108 309048 226160
rect 309100 226148 309106 226160
rect 336274 226148 336280 226160
rect 309100 226120 336280 226148
rect 309100 226108 309106 226120
rect 336274 226108 336280 226120
rect 336332 226108 336338 226160
rect 528554 226108 528560 226160
rect 528612 226148 528618 226160
rect 542998 226148 543004 226160
rect 528612 226120 543004 226148
rect 528612 226108 528618 226120
rect 542998 226108 543004 226120
rect 543056 226108 543062 226160
rect 672604 226102 672656 226108
rect 220078 226012 220084 226024
rect 214576 225984 220084 226012
rect 220078 225972 220084 225984
rect 220136 225972 220142 226024
rect 220262 225972 220268 226024
rect 220320 226012 220326 226024
rect 266078 226012 266084 226024
rect 220320 225984 266084 226012
rect 220320 225972 220326 225984
rect 266078 225972 266084 225984
rect 266136 225972 266142 226024
rect 266998 225972 267004 226024
rect 267056 226012 267062 226024
rect 274450 226012 274456 226024
rect 267056 225984 274456 226012
rect 267056 225972 267062 225984
rect 274450 225972 274456 225984
rect 274508 225972 274514 226024
rect 278406 225972 278412 226024
rect 278464 226012 278470 226024
rect 313274 226012 313280 226024
rect 278464 225984 313280 226012
rect 278464 225972 278470 225984
rect 313274 225972 313280 225984
rect 313332 225972 313338 226024
rect 321370 225972 321376 226024
rect 321428 226012 321434 226024
rect 346578 226012 346584 226024
rect 321428 225984 346584 226012
rect 321428 225972 321434 225984
rect 346578 225972 346584 225984
rect 346636 225972 346642 226024
rect 352926 225972 352932 226024
rect 352984 226012 352990 226024
rect 371694 226012 371700 226024
rect 352984 225984 371700 226012
rect 352984 225972 352990 225984
rect 371694 225972 371700 225984
rect 371752 225972 371758 226024
rect 498102 225972 498108 226024
rect 498160 226012 498166 226024
rect 514294 226012 514300 226024
rect 498160 225984 514300 226012
rect 498160 225972 498166 225984
rect 514294 225972 514300 225984
rect 514352 225972 514358 226024
rect 516594 225972 516600 226024
rect 516652 226012 516658 226024
rect 538674 226012 538680 226024
rect 516652 225984 538680 226012
rect 516652 225972 516658 225984
rect 538674 225972 538680 225984
rect 538732 225972 538738 226024
rect 672494 225956 672546 225962
rect 672494 225898 672546 225904
rect 83458 225836 83464 225888
rect 83516 225876 83522 225888
rect 163038 225876 163044 225888
rect 83516 225848 163044 225876
rect 83516 225836 83522 225848
rect 163038 225836 163044 225848
rect 163096 225836 163102 225888
rect 193582 225836 193588 225888
rect 193640 225876 193646 225888
rect 194134 225876 194140 225888
rect 193640 225848 194140 225876
rect 193640 225836 193646 225848
rect 194134 225836 194140 225848
rect 194192 225836 194198 225888
rect 197998 225836 198004 225888
rect 198056 225876 198062 225888
rect 203886 225876 203892 225888
rect 198056 225848 203892 225876
rect 198056 225836 198062 225848
rect 203886 225836 203892 225848
rect 203944 225836 203950 225888
rect 204898 225836 204904 225888
rect 204956 225876 204962 225888
rect 231486 225876 231492 225888
rect 204956 225848 231492 225876
rect 204956 225836 204962 225848
rect 231486 225836 231492 225848
rect 231544 225836 231550 225888
rect 249334 225876 249340 225888
rect 233528 225848 249340 225876
rect 233528 225808 233556 225848
rect 249334 225836 249340 225848
rect 249392 225836 249398 225888
rect 252462 225836 252468 225888
rect 252520 225876 252526 225888
rect 293126 225876 293132 225888
rect 252520 225848 293132 225876
rect 252520 225836 252526 225848
rect 293126 225836 293132 225848
rect 293184 225836 293190 225888
rect 296438 225836 296444 225888
rect 296496 225876 296502 225888
rect 327902 225876 327908 225888
rect 296496 225848 327908 225876
rect 296496 225836 296502 225848
rect 327902 225836 327908 225848
rect 327960 225836 327966 225888
rect 329742 225836 329748 225888
rect 329800 225876 329806 225888
rect 353662 225876 353668 225888
rect 329800 225848 353668 225876
rect 329800 225836 329806 225848
rect 353662 225836 353668 225848
rect 353720 225836 353726 225888
rect 354582 225836 354588 225888
rect 354640 225876 354646 225888
rect 372338 225876 372344 225888
rect 354640 225848 372344 225876
rect 354640 225836 354646 225848
rect 372338 225836 372344 225848
rect 372396 225836 372402 225888
rect 373810 225836 373816 225888
rect 373868 225876 373874 225888
rect 377674 225876 377680 225888
rect 373868 225848 377680 225876
rect 373868 225836 373874 225848
rect 377674 225836 377680 225848
rect 377732 225836 377738 225888
rect 377858 225836 377864 225888
rect 377916 225876 377922 225888
rect 390370 225876 390376 225888
rect 377916 225848 390376 225876
rect 377916 225836 377922 225848
rect 390370 225836 390376 225848
rect 390428 225836 390434 225888
rect 394326 225836 394332 225888
rect 394384 225876 394390 225888
rect 403250 225876 403256 225888
rect 394384 225848 403256 225876
rect 394384 225836 394390 225848
rect 403250 225836 403256 225848
rect 403308 225836 403314 225888
rect 483750 225836 483756 225888
rect 483808 225876 483814 225888
rect 497274 225876 497280 225888
rect 483808 225848 497280 225876
rect 483808 225836 483814 225848
rect 497274 225836 497280 225848
rect 497332 225836 497338 225888
rect 501138 225836 501144 225888
rect 501196 225876 501202 225888
rect 519262 225876 519268 225888
rect 501196 225848 519268 225876
rect 501196 225836 501202 225848
rect 519262 225836 519268 225848
rect 519320 225836 519326 225888
rect 521746 225836 521752 225888
rect 521804 225876 521810 225888
rect 545758 225876 545764 225888
rect 521804 225848 545764 225876
rect 521804 225836 521810 225848
rect 545758 225836 545764 225848
rect 545816 225836 545822 225888
rect 558178 225836 558184 225888
rect 558236 225876 558242 225888
rect 571978 225876 571984 225888
rect 558236 225848 571984 225876
rect 558236 225836 558242 225848
rect 571978 225836 571984 225848
rect 572036 225836 572042 225888
rect 231964 225780 233556 225808
rect 76558 225700 76564 225752
rect 76616 225740 76622 225752
rect 151722 225740 151728 225752
rect 76616 225712 151728 225740
rect 76616 225700 76622 225712
rect 151722 225700 151728 225712
rect 151780 225700 151786 225752
rect 151906 225700 151912 225752
rect 151964 225740 151970 225752
rect 154298 225740 154304 225752
rect 151964 225712 154304 225740
rect 151964 225700 151970 225712
rect 154298 225700 154304 225712
rect 154356 225700 154362 225752
rect 184290 225740 184296 225752
rect 154500 225712 184296 225740
rect 66162 225564 66168 225616
rect 66220 225604 66226 225616
rect 142108 225604 142114 225616
rect 66220 225576 142114 225604
rect 66220 225564 66226 225576
rect 142108 225564 142114 225576
rect 142166 225564 142172 225616
rect 142246 225564 142252 225616
rect 142304 225604 142310 225616
rect 154500 225604 154528 225712
rect 184290 225700 184296 225712
rect 184348 225700 184354 225752
rect 184474 225700 184480 225752
rect 184532 225740 184538 225752
rect 212534 225740 212540 225752
rect 184532 225712 212540 225740
rect 184532 225700 184538 225712
rect 212534 225700 212540 225712
rect 212592 225700 212598 225752
rect 215202 225700 215208 225752
rect 215260 225740 215266 225752
rect 215260 225712 219940 225740
rect 215260 225700 215266 225712
rect 142304 225576 154528 225604
rect 142304 225564 142310 225576
rect 154666 225564 154672 225616
rect 154724 225604 154730 225616
rect 217134 225604 217140 225616
rect 154724 225576 217140 225604
rect 154724 225564 154730 225576
rect 217134 225564 217140 225576
rect 217192 225564 217198 225616
rect 219912 225604 219940 225712
rect 220078 225700 220084 225752
rect 220136 225740 220142 225752
rect 231964 225740 231992 225780
rect 672380 225752 672432 225758
rect 220136 225712 231992 225740
rect 220136 225700 220142 225712
rect 237282 225700 237288 225752
rect 237340 225740 237346 225752
rect 240318 225740 240324 225752
rect 237340 225712 240324 225740
rect 237340 225700 237346 225712
rect 240318 225700 240324 225712
rect 240376 225700 240382 225752
rect 255038 225700 255044 225752
rect 255096 225740 255102 225752
rect 296990 225740 296996 225752
rect 255096 225712 296996 225740
rect 255096 225700 255102 225712
rect 296990 225700 296996 225712
rect 297048 225700 297054 225752
rect 315666 225700 315672 225752
rect 315724 225740 315730 225752
rect 344646 225740 344652 225752
rect 315724 225712 344652 225740
rect 315724 225700 315730 225712
rect 344646 225700 344652 225712
rect 344704 225700 344710 225752
rect 347038 225700 347044 225752
rect 347096 225740 347102 225752
rect 367830 225740 367836 225752
rect 347096 225712 367836 225740
rect 347096 225700 347102 225712
rect 367830 225700 367836 225712
rect 367888 225700 367894 225752
rect 371786 225700 371792 225752
rect 371844 225740 371850 225752
rect 382734 225740 382740 225752
rect 371844 225712 382740 225740
rect 371844 225700 371850 225712
rect 382734 225700 382740 225712
rect 382792 225700 382798 225752
rect 382918 225700 382924 225752
rect 382976 225740 382982 225752
rect 396166 225740 396172 225752
rect 382976 225712 396172 225740
rect 382976 225700 382982 225712
rect 396166 225700 396172 225712
rect 396224 225700 396230 225752
rect 488902 225700 488908 225752
rect 488960 225740 488966 225752
rect 503622 225740 503628 225752
rect 488960 225712 503628 225740
rect 488960 225700 488966 225712
rect 503622 225700 503628 225712
rect 503680 225700 503686 225752
rect 508866 225700 508872 225752
rect 508924 225740 508930 225752
rect 529198 225740 529204 225752
rect 508924 225712 529204 225740
rect 508924 225700 508930 225712
rect 529198 225700 529204 225712
rect 529256 225700 529262 225752
rect 535914 225700 535920 225752
rect 535972 225740 535978 225752
rect 563974 225740 563980 225752
rect 535972 225712 563980 225740
rect 535972 225700 535978 225712
rect 563974 225700 563980 225712
rect 564032 225700 564038 225752
rect 672380 225694 672432 225700
rect 672264 225684 672316 225690
rect 672264 225626 672316 225632
rect 220262 225604 220268 225616
rect 219912 225576 220268 225604
rect 220262 225564 220268 225576
rect 220320 225564 220326 225616
rect 222010 225564 222016 225616
rect 222068 225604 222074 225616
rect 269942 225604 269948 225616
rect 222068 225576 269948 225604
rect 222068 225564 222074 225576
rect 269942 225564 269948 225576
rect 270000 225564 270006 225616
rect 270218 225564 270224 225616
rect 270276 225604 270282 225616
rect 282638 225604 282644 225616
rect 270276 225576 282644 225604
rect 270276 225564 270282 225576
rect 282638 225564 282644 225576
rect 282696 225564 282702 225616
rect 284110 225564 284116 225616
rect 284168 225604 284174 225616
rect 320174 225604 320180 225616
rect 284168 225576 320180 225604
rect 284168 225564 284174 225576
rect 320174 225564 320180 225576
rect 320232 225564 320238 225616
rect 332226 225564 332232 225616
rect 332284 225604 332290 225616
rect 357526 225604 357532 225616
rect 332284 225576 357532 225604
rect 332284 225564 332290 225576
rect 357526 225564 357532 225576
rect 357584 225564 357590 225616
rect 372522 225564 372528 225616
rect 372580 225604 372586 225616
rect 387426 225604 387432 225616
rect 372580 225576 387432 225604
rect 372580 225564 372586 225576
rect 387426 225564 387432 225576
rect 387484 225564 387490 225616
rect 390186 225564 390192 225616
rect 390244 225604 390250 225616
rect 401962 225604 401968 225616
rect 390244 225576 401968 225604
rect 390244 225564 390250 225576
rect 401962 225564 401968 225576
rect 402020 225564 402026 225616
rect 410978 225564 410984 225616
rect 411036 225604 411042 225616
rect 416130 225604 416136 225616
rect 411036 225576 416136 225604
rect 411036 225564 411042 225576
rect 416130 225564 416136 225576
rect 416188 225564 416194 225616
rect 467650 225564 467656 225616
rect 467708 225604 467714 225616
rect 476574 225604 476580 225616
rect 467708 225576 476580 225604
rect 467708 225564 467714 225576
rect 476574 225564 476580 225576
rect 476632 225564 476638 225616
rect 477310 225564 477316 225616
rect 477368 225604 477374 225616
rect 488810 225604 488816 225616
rect 477368 225576 488816 225604
rect 477368 225564 477374 225576
rect 488810 225564 488816 225576
rect 488868 225564 488874 225616
rect 494054 225564 494060 225616
rect 494112 225604 494118 225616
rect 509694 225604 509700 225616
rect 494112 225576 509700 225604
rect 494112 225564 494118 225576
rect 509694 225564 509700 225576
rect 509752 225564 509758 225616
rect 510154 225564 510160 225616
rect 510212 225604 510218 225616
rect 531038 225604 531044 225616
rect 510212 225576 531044 225604
rect 510212 225564 510218 225576
rect 531038 225564 531044 225576
rect 531096 225564 531102 225616
rect 531406 225564 531412 225616
rect 531464 225604 531470 225616
rect 558270 225604 558276 225616
rect 531464 225576 558276 225604
rect 531464 225564 531470 225576
rect 558270 225564 558276 225576
rect 558328 225564 558334 225616
rect 110138 225428 110144 225480
rect 110196 225468 110202 225480
rect 127618 225468 127624 225480
rect 110196 225440 127624 225468
rect 110196 225428 110202 225440
rect 127618 225428 127624 225440
rect 127676 225428 127682 225480
rect 196158 225468 196164 225480
rect 127820 225440 196164 225468
rect 125226 225292 125232 225344
rect 125284 225332 125290 225344
rect 127820 225332 127848 225440
rect 196158 225428 196164 225440
rect 196216 225428 196222 225480
rect 196342 225428 196348 225480
rect 196400 225468 196406 225480
rect 204898 225468 204904 225480
rect 196400 225440 204904 225468
rect 196400 225428 196406 225440
rect 204898 225428 204904 225440
rect 204956 225428 204962 225480
rect 208118 225428 208124 225480
rect 208176 225468 208182 225480
rect 257430 225468 257436 225480
rect 208176 225440 257436 225468
rect 208176 225428 208182 225440
rect 257430 225428 257436 225440
rect 257488 225428 257494 225480
rect 672156 225412 672208 225418
rect 463142 225360 463148 225412
rect 463200 225400 463206 225412
rect 467282 225400 467288 225412
rect 463200 225372 467288 225400
rect 463200 225360 463206 225372
rect 467282 225360 467288 225372
rect 467340 225360 467346 225412
rect 672156 225354 672208 225360
rect 125284 225304 127848 225332
rect 125284 225292 125290 225304
rect 129366 225292 129372 225344
rect 129424 225332 129430 225344
rect 199102 225332 199108 225344
rect 129424 225304 199108 225332
rect 129424 225292 129430 225304
rect 199102 225292 199108 225304
rect 199160 225292 199166 225344
rect 203702 225292 203708 225344
rect 203760 225332 203766 225344
rect 209406 225332 209412 225344
rect 203760 225304 209412 225332
rect 203760 225292 203766 225304
rect 209406 225292 209412 225304
rect 209464 225292 209470 225344
rect 209682 225292 209688 225344
rect 209740 225332 209746 225344
rect 214742 225332 214748 225344
rect 209740 225304 214748 225332
rect 209740 225292 209746 225304
rect 214742 225292 214748 225304
rect 214800 225292 214806 225344
rect 231486 225292 231492 225344
rect 231544 225332 231550 225344
rect 236454 225332 236460 225344
rect 231544 225304 236460 225332
rect 231544 225292 231550 225304
rect 236454 225292 236460 225304
rect 236512 225292 236518 225344
rect 241146 225292 241152 225344
rect 241204 225332 241210 225344
rect 286686 225332 286692 225344
rect 241204 225304 286692 225332
rect 241204 225292 241210 225304
rect 286686 225292 286692 225304
rect 286744 225292 286750 225344
rect 563026 225304 572714 225332
rect 135162 225156 135168 225208
rect 135220 225196 135226 225208
rect 204254 225196 204260 225208
rect 135220 225168 204260 225196
rect 135220 225156 135226 225168
rect 204254 225156 204260 225168
rect 204312 225156 204318 225208
rect 242710 225156 242716 225208
rect 242768 225196 242774 225208
rect 285398 225196 285404 225208
rect 242768 225168 285404 225196
rect 242768 225156 242774 225168
rect 285398 225156 285404 225168
rect 285456 225156 285462 225208
rect 132402 225020 132408 225072
rect 132460 225060 132466 225072
rect 201678 225060 201684 225072
rect 132460 225032 201684 225060
rect 132460 225020 132466 225032
rect 201678 225020 201684 225032
rect 201736 225020 201742 225072
rect 202230 225020 202236 225072
rect 202288 225060 202294 225072
rect 254486 225060 254492 225072
rect 202288 225032 254492 225060
rect 202288 225020 202294 225032
rect 254486 225020 254492 225032
rect 254544 225020 254550 225072
rect 297266 224952 297272 225004
rect 297324 224992 297330 225004
rect 305362 224992 305368 225004
rect 297324 224964 305368 224992
rect 297324 224952 297330 224964
rect 305362 224952 305368 224964
rect 305420 224952 305426 225004
rect 327718 224952 327724 225004
rect 327776 224992 327782 225004
rect 332042 224992 332048 225004
rect 327776 224964 332048 224992
rect 327776 224952 327782 224964
rect 332042 224952 332048 224964
rect 332100 224952 332106 225004
rect 369118 224952 369124 225004
rect 369176 224992 369182 225004
rect 373626 224992 373632 225004
rect 369176 224964 373632 224992
rect 369176 224952 369182 224964
rect 373626 224952 373632 224964
rect 373684 224952 373690 225004
rect 404170 224952 404176 225004
rect 404228 224992 404234 225004
rect 410610 224992 410616 225004
rect 404228 224964 410616 224992
rect 404228 224952 404234 224964
rect 410610 224952 410616 224964
rect 410668 224952 410674 225004
rect 416498 224952 416504 225004
rect 416556 224992 416562 225004
rect 422202 224992 422208 225004
rect 416556 224964 422208 224992
rect 416556 224952 416562 224964
rect 422202 224952 422208 224964
rect 422260 224952 422266 225004
rect 493594 224952 493600 225004
rect 493652 224992 493658 225004
rect 494698 224992 494704 225004
rect 493652 224964 494704 224992
rect 493652 224952 493658 224964
rect 494698 224952 494704 224964
rect 494756 224952 494762 225004
rect 495158 224952 495164 225004
rect 495216 224992 495222 225004
rect 563026 224992 563054 225304
rect 567010 225088 567016 225140
rect 567068 225128 567074 225140
rect 571426 225128 571432 225140
rect 567068 225100 571432 225128
rect 567068 225088 567074 225100
rect 571426 225088 571432 225100
rect 571484 225088 571490 225140
rect 495216 224964 563054 224992
rect 495216 224952 495222 224964
rect 563698 224952 563704 225004
rect 563756 224992 563762 225004
rect 572686 224992 572714 225304
rect 672034 225276 672086 225282
rect 672034 225218 672086 225224
rect 663766 225032 671968 225060
rect 630858 224992 630864 225004
rect 563756 224964 567148 224992
rect 572686 224964 630864 224992
rect 563756 224952 563762 224964
rect 96246 224884 96252 224936
rect 96304 224924 96310 224936
rect 173342 224924 173348 224936
rect 96304 224896 173348 224924
rect 96304 224884 96310 224896
rect 173342 224884 173348 224896
rect 173400 224884 173406 224936
rect 174906 224884 174912 224936
rect 174964 224924 174970 224936
rect 181346 224924 181352 224936
rect 174964 224896 181352 224924
rect 174964 224884 174970 224896
rect 181346 224884 181352 224896
rect 181404 224884 181410 224936
rect 181990 224884 181996 224936
rect 182048 224924 182054 224936
rect 182048 224896 185624 224924
rect 182048 224884 182054 224896
rect 102042 224748 102048 224800
rect 102100 224788 102106 224800
rect 178494 224788 178500 224800
rect 102100 224760 178500 224788
rect 102100 224748 102106 224760
rect 178494 224748 178500 224760
rect 178552 224748 178558 224800
rect 178770 224748 178776 224800
rect 178828 224788 178834 224800
rect 185394 224788 185400 224800
rect 178828 224760 185400 224788
rect 178828 224748 178834 224760
rect 185394 224748 185400 224760
rect 185452 224748 185458 224800
rect 185596 224788 185624 224896
rect 185762 224884 185768 224936
rect 185820 224924 185826 224936
rect 195238 224924 195244 224936
rect 185820 224896 195244 224924
rect 185820 224884 185826 224896
rect 195238 224884 195244 224896
rect 195296 224884 195302 224936
rect 195422 224884 195428 224936
rect 195480 224924 195486 224936
rect 242894 224924 242900 224936
rect 195480 224896 242900 224924
rect 195480 224884 195486 224896
rect 242894 224884 242900 224896
rect 242952 224884 242958 224936
rect 266170 224884 266176 224936
rect 266228 224924 266234 224936
rect 266228 224896 296714 224924
rect 266228 224884 266234 224896
rect 296686 224856 296714 224896
rect 460566 224884 460572 224936
rect 460624 224924 460630 224936
rect 463142 224924 463148 224936
rect 460624 224896 463148 224924
rect 460624 224884 460630 224896
rect 463142 224884 463148 224896
rect 463200 224884 463206 224936
rect 567120 224924 567148 224964
rect 630858 224952 630864 224964
rect 630916 224952 630922 225004
rect 658182 224952 658188 225004
rect 658240 224992 658246 225004
rect 663766 224992 663794 225032
rect 658240 224964 663794 224992
rect 658240 224952 658246 224964
rect 568942 224924 568948 224936
rect 567120 224896 568948 224924
rect 568942 224884 568948 224896
rect 569000 224884 569006 224936
rect 303430 224856 303436 224868
rect 296686 224828 303436 224856
rect 303430 224816 303436 224828
rect 303488 224816 303494 224868
rect 610986 224816 610992 224868
rect 611044 224856 611050 224868
rect 614942 224856 614948 224868
rect 611044 224828 614948 224856
rect 611044 224816 611050 224828
rect 614942 224816 614948 224828
rect 615000 224816 615006 224868
rect 204530 224788 204536 224800
rect 185596 224760 204536 224788
rect 204530 224748 204536 224760
rect 204588 224748 204594 224800
rect 204714 224748 204720 224800
rect 204772 224788 204778 224800
rect 204772 224760 224080 224788
rect 204772 224748 204778 224760
rect 79962 224612 79968 224664
rect 80020 224652 80026 224664
rect 160462 224652 160468 224664
rect 80020 224624 160468 224652
rect 80020 224612 80026 224624
rect 160462 224612 160468 224624
rect 160520 224612 160526 224664
rect 162762 224612 162768 224664
rect 162820 224652 162826 224664
rect 223850 224652 223856 224664
rect 162820 224624 223856 224652
rect 162820 224612 162826 224624
rect 223850 224612 223856 224624
rect 223908 224612 223914 224664
rect 224052 224652 224080 224760
rect 224218 224748 224224 224800
rect 224276 224788 224282 224800
rect 230014 224788 230020 224800
rect 224276 224760 230020 224788
rect 224276 224748 224282 224760
rect 230014 224748 230020 224760
rect 230072 224748 230078 224800
rect 232958 224748 232964 224800
rect 233016 224788 233022 224800
rect 237742 224788 237748 224800
rect 233016 224760 237748 224788
rect 233016 224748 233022 224760
rect 237742 224748 237748 224760
rect 237800 224748 237806 224800
rect 245286 224748 245292 224800
rect 245344 224788 245350 224800
rect 287974 224788 287980 224800
rect 245344 224760 287980 224788
rect 245344 224748 245350 224760
rect 287974 224748 287980 224760
rect 288032 224748 288038 224800
rect 311526 224748 311532 224800
rect 311584 224788 311590 224800
rect 338850 224788 338856 224800
rect 311584 224760 338856 224788
rect 311584 224748 311590 224760
rect 338850 224748 338856 224760
rect 338908 224748 338914 224800
rect 462498 224748 462504 224800
rect 462556 224788 462562 224800
rect 469306 224788 469312 224800
rect 462556 224760 469312 224788
rect 462556 224748 462562 224760
rect 469306 224748 469312 224760
rect 469364 224748 469370 224800
rect 506934 224748 506940 224800
rect 506992 224788 506998 224800
rect 526714 224788 526720 224800
rect 506992 224760 526720 224788
rect 506992 224748 506998 224760
rect 526714 224748 526720 224760
rect 526772 224748 526778 224800
rect 529934 224748 529940 224800
rect 529992 224788 529998 224800
rect 534534 224788 534540 224800
rect 529992 224760 534540 224788
rect 529992 224748 529998 224760
rect 534534 224748 534540 224760
rect 534592 224748 534598 224800
rect 557350 224788 557356 224800
rect 534736 224760 557356 224788
rect 366542 224720 366548 224732
rect 354646 224692 366548 224720
rect 224402 224652 224408 224664
rect 224052 224624 224408 224652
rect 224402 224612 224408 224624
rect 224460 224612 224466 224664
rect 224586 224612 224592 224664
rect 224644 224652 224650 224664
rect 270586 224652 270592 224664
rect 224644 224624 270592 224652
rect 224644 224612 224650 224624
rect 270586 224612 270592 224624
rect 270644 224612 270650 224664
rect 274266 224612 274272 224664
rect 274324 224652 274330 224664
rect 312446 224652 312452 224664
rect 274324 224624 312452 224652
rect 274324 224612 274330 224624
rect 312446 224612 312452 224624
rect 312504 224612 312510 224664
rect 319806 224612 319812 224664
rect 319864 224652 319870 224664
rect 345934 224652 345940 224664
rect 319864 224624 345940 224652
rect 319864 224612 319870 224624
rect 345934 224612 345940 224624
rect 345992 224612 345998 224664
rect 346210 224612 346216 224664
rect 346268 224652 346274 224664
rect 354646 224652 354674 224692
rect 366542 224680 366548 224692
rect 366600 224680 366606 224732
rect 346268 224624 354674 224652
rect 346268 224612 346274 224624
rect 505186 224612 505192 224664
rect 505244 224652 505250 224664
rect 534736 224652 534764 224760
rect 557350 224748 557356 224760
rect 557408 224748 557414 224800
rect 562134 224788 562140 224800
rect 557644 224760 562140 224788
rect 505244 224624 534764 224652
rect 505244 224612 505250 224624
rect 535270 224612 535276 224664
rect 535328 224652 535334 224664
rect 557644 224652 557672 224760
rect 562134 224748 562140 224760
rect 562192 224748 562198 224800
rect 562318 224748 562324 224800
rect 562376 224788 562382 224800
rect 567010 224788 567016 224800
rect 562376 224760 567016 224788
rect 562376 224748 562382 224760
rect 567010 224748 567016 224760
rect 567068 224748 567074 224800
rect 567838 224748 567844 224800
rect 567896 224788 567902 224800
rect 610802 224788 610808 224800
rect 567896 224760 610808 224788
rect 567896 224748 567902 224760
rect 610802 224748 610808 224760
rect 610860 224748 610866 224800
rect 671820 224732 671872 224738
rect 668486 224680 668492 224732
rect 668544 224720 668550 224732
rect 668544 224692 670740 224720
rect 668544 224680 668550 224692
rect 535328 224624 557672 224652
rect 535328 224612 535334 224624
rect 557810 224612 557816 224664
rect 557868 224652 557874 224664
rect 610434 224652 610440 224664
rect 557868 224624 610440 224652
rect 557868 224612 557874 224624
rect 610434 224612 610440 224624
rect 610492 224612 610498 224664
rect 610618 224612 610624 224664
rect 610676 224652 610682 224664
rect 616046 224652 616052 224664
rect 610676 224624 616052 224652
rect 610676 224612 610682 224624
rect 616046 224612 616052 224624
rect 616104 224612 616110 224664
rect 670712 224652 670740 224692
rect 671820 224674 671872 224680
rect 670712 224624 671738 224652
rect 85482 224476 85488 224528
rect 85540 224516 85546 224528
rect 165614 224516 165620 224528
rect 85540 224488 165620 224516
rect 85540 224476 85546 224488
rect 165614 224476 165620 224488
rect 165672 224476 165678 224528
rect 181346 224476 181352 224528
rect 181404 224516 181410 224528
rect 235166 224516 235172 224528
rect 181404 224488 235172 224516
rect 181404 224476 181410 224488
rect 235166 224476 235172 224488
rect 235224 224476 235230 224528
rect 251082 224476 251088 224528
rect 251140 224516 251146 224528
rect 294414 224516 294420 224528
rect 251140 224488 294420 224516
rect 251140 224476 251146 224488
rect 294414 224476 294420 224488
rect 294472 224476 294478 224528
rect 319990 224476 319996 224528
rect 320048 224516 320054 224528
rect 347222 224516 347228 224528
rect 320048 224488 347228 224516
rect 320048 224476 320054 224488
rect 347222 224476 347228 224488
rect 347280 224476 347286 224528
rect 363506 224476 363512 224528
rect 363564 224516 363570 224528
rect 368474 224516 368480 224528
rect 363564 224488 368480 224516
rect 363564 224476 363570 224488
rect 368474 224476 368480 224488
rect 368532 224476 368538 224528
rect 387702 224476 387708 224528
rect 387760 224516 387766 224528
rect 397822 224516 397828 224528
rect 387760 224488 397828 224516
rect 387760 224476 387766 224488
rect 397822 224476 397828 224488
rect 397880 224476 397886 224528
rect 456058 224476 456064 224528
rect 456116 224516 456122 224528
rect 459738 224516 459744 224528
rect 456116 224488 459744 224516
rect 456116 224476 456122 224488
rect 459738 224476 459744 224488
rect 459796 224476 459802 224528
rect 491294 224476 491300 224528
rect 491352 224516 491358 224528
rect 506106 224516 506112 224528
rect 491352 224488 506112 224516
rect 491352 224476 491358 224488
rect 506106 224476 506112 224488
rect 506164 224476 506170 224528
rect 515950 224476 515956 224528
rect 516008 224516 516014 224528
rect 530854 224516 530860 224528
rect 516008 224488 530860 224516
rect 516008 224476 516014 224488
rect 530854 224476 530860 224488
rect 530912 224476 530918 224528
rect 544102 224516 544108 224528
rect 532344 224488 544108 224516
rect 73706 224340 73712 224392
rect 73764 224380 73770 224392
rect 88978 224380 88984 224392
rect 73764 224352 88984 224380
rect 73764 224340 73770 224352
rect 88978 224340 88984 224352
rect 89036 224340 89042 224392
rect 89438 224340 89444 224392
rect 89496 224380 89502 224392
rect 167822 224380 167828 224392
rect 89496 224352 167828 224380
rect 89496 224340 89502 224352
rect 167822 224340 167828 224352
rect 167880 224340 167886 224392
rect 168282 224340 168288 224392
rect 168340 224380 168346 224392
rect 224218 224380 224224 224392
rect 168340 224352 224224 224380
rect 168340 224340 168346 224352
rect 224218 224340 224224 224352
rect 224276 224340 224282 224392
rect 224402 224340 224408 224392
rect 224460 224380 224466 224392
rect 232958 224380 232964 224392
rect 224460 224352 232964 224380
rect 224460 224340 224466 224352
rect 232958 224340 232964 224352
rect 233016 224340 233022 224392
rect 233142 224340 233148 224392
rect 233200 224380 233206 224392
rect 277670 224380 277676 224392
rect 233200 224352 277676 224380
rect 233200 224340 233206 224352
rect 277670 224340 277676 224352
rect 277728 224340 277734 224392
rect 299290 224340 299296 224392
rect 299348 224380 299354 224392
rect 331766 224380 331772 224392
rect 299348 224352 331772 224380
rect 299348 224340 299354 224352
rect 331766 224340 331772 224352
rect 331824 224340 331830 224392
rect 335170 224340 335176 224392
rect 335228 224380 335234 224392
rect 356882 224380 356888 224392
rect 335228 224352 356888 224380
rect 335228 224340 335234 224352
rect 356882 224340 356888 224352
rect 356940 224340 356946 224392
rect 361206 224340 361212 224392
rect 361264 224380 361270 224392
rect 377490 224380 377496 224392
rect 361264 224352 377496 224380
rect 361264 224340 361270 224352
rect 377490 224340 377496 224352
rect 377548 224340 377554 224392
rect 379238 224340 379244 224392
rect 379296 224380 379302 224392
rect 393590 224380 393596 224392
rect 379296 224352 393596 224380
rect 379296 224340 379302 224352
rect 393590 224340 393596 224352
rect 393648 224340 393654 224392
rect 480530 224340 480536 224392
rect 480588 224380 480594 224392
rect 492766 224380 492772 224392
rect 480588 224352 492772 224380
rect 480588 224340 480594 224352
rect 492766 224340 492772 224352
rect 492824 224340 492830 224392
rect 499206 224340 499212 224392
rect 499264 224380 499270 224392
rect 516778 224380 516784 224392
rect 499264 224352 516784 224380
rect 499264 224340 499270 224352
rect 516778 224340 516784 224352
rect 516836 224340 516842 224392
rect 520458 224340 520464 224392
rect 520516 224380 520522 224392
rect 532344 224380 532372 224488
rect 544102 224476 544108 224488
rect 544160 224476 544166 224528
rect 544286 224476 544292 224528
rect 544344 224516 544350 224528
rect 549990 224516 549996 224528
rect 544344 224488 549996 224516
rect 544344 224476 544350 224488
rect 549990 224476 549996 224488
rect 550048 224516 550054 224528
rect 550358 224516 550364 224528
rect 550048 224488 550364 224516
rect 550048 224476 550054 224488
rect 550358 224476 550364 224488
rect 550416 224476 550422 224528
rect 551186 224476 551192 224528
rect 551244 224516 551250 224528
rect 557166 224516 557172 224528
rect 551244 224488 557172 224516
rect 551244 224476 551250 224488
rect 557166 224476 557172 224488
rect 557224 224476 557230 224528
rect 625246 224516 625252 224528
rect 557506 224488 625252 224516
rect 550634 224380 550640 224392
rect 520516 224352 532372 224380
rect 532436 224352 550640 224380
rect 520516 224340 520522 224352
rect 426434 224272 426440 224324
rect 426492 224312 426498 224324
rect 426986 224312 426992 224324
rect 426492 224284 426992 224312
rect 426492 224272 426498 224284
rect 426986 224272 426992 224284
rect 427044 224272 427050 224324
rect 151630 224244 151636 224256
rect 84166 224216 151636 224244
rect 68922 224068 68928 224120
rect 68980 224108 68986 224120
rect 84166 224108 84194 224216
rect 151630 224204 151636 224216
rect 151688 224204 151694 224256
rect 151768 224204 151774 224256
rect 151826 224244 151832 224256
rect 155310 224244 155316 224256
rect 151826 224216 155316 224244
rect 151826 224204 151832 224216
rect 155310 224204 155316 224216
rect 155368 224204 155374 224256
rect 165522 224204 165528 224256
rect 165580 224244 165586 224256
rect 227438 224244 227444 224256
rect 165580 224216 227444 224244
rect 165580 224204 165586 224216
rect 227438 224204 227444 224216
rect 227496 224204 227502 224256
rect 231670 224204 231676 224256
rect 231728 224244 231734 224256
rect 278958 224244 278964 224256
rect 231728 224216 278964 224244
rect 231728 224204 231734 224216
rect 278958 224204 278964 224216
rect 279016 224204 279022 224256
rect 290826 224204 290832 224256
rect 290884 224244 290890 224256
rect 323670 224244 323676 224256
rect 290884 224216 323676 224244
rect 290884 224204 290890 224216
rect 323670 224204 323676 224216
rect 323728 224204 323734 224256
rect 323946 224204 323952 224256
rect 324004 224244 324010 224256
rect 334986 224244 334992 224256
rect 324004 224216 334992 224244
rect 324004 224204 324010 224216
rect 334986 224204 334992 224216
rect 335044 224204 335050 224256
rect 339402 224204 339408 224256
rect 339460 224244 339466 224256
rect 339460 224216 354674 224244
rect 339460 224204 339466 224216
rect 68980 224080 84194 224108
rect 68980 224068 68986 224080
rect 88978 224068 88984 224120
rect 89036 224108 89042 224120
rect 142108 224108 142114 224120
rect 89036 224080 142114 224108
rect 89036 224068 89042 224080
rect 142108 224068 142114 224080
rect 142166 224068 142172 224120
rect 142246 224068 142252 224120
rect 142304 224108 142310 224120
rect 194594 224108 194600 224120
rect 142304 224080 194600 224108
rect 142304 224068 142310 224080
rect 194594 224068 194600 224080
rect 194652 224068 194658 224120
rect 195238 224068 195244 224120
rect 195296 224108 195302 224120
rect 204714 224108 204720 224120
rect 195296 224080 204720 224108
rect 195296 224068 195302 224080
rect 204714 224068 204720 224080
rect 204772 224068 204778 224120
rect 204898 224068 204904 224120
rect 204956 224108 204962 224120
rect 250622 224108 250628 224120
rect 204956 224080 250628 224108
rect 204956 224068 204962 224080
rect 250622 224068 250628 224080
rect 250680 224068 250686 224120
rect 275094 224068 275100 224120
rect 275152 224108 275158 224120
rect 311158 224108 311164 224120
rect 275152 224080 311164 224108
rect 275152 224068 275158 224080
rect 311158 224068 311164 224080
rect 311216 224068 311222 224120
rect 354646 224108 354674 224216
rect 358078 224204 358084 224256
rect 358136 224244 358142 224256
rect 362954 224244 362960 224256
rect 358136 224216 362960 224244
rect 358136 224204 358142 224216
rect 362954 224204 362960 224216
rect 363012 224204 363018 224256
rect 366726 224204 366732 224256
rect 366784 224244 366790 224256
rect 381630 224244 381636 224256
rect 366784 224216 381636 224244
rect 366784 224204 366790 224216
rect 381630 224204 381636 224216
rect 381688 224204 381694 224256
rect 394510 224204 394516 224256
rect 394568 224244 394574 224256
rect 404538 224244 404544 224256
rect 394568 224216 404544 224244
rect 394568 224204 394574 224216
rect 404538 224204 404544 224216
rect 404596 224204 404602 224256
rect 405550 224204 405556 224256
rect 405608 224244 405614 224256
rect 414198 224244 414204 224256
rect 405608 224216 414204 224244
rect 405608 224204 405614 224216
rect 414198 224204 414204 224216
rect 414256 224204 414262 224256
rect 427906 224204 427912 224256
rect 427964 224244 427970 224256
rect 428734 224244 428740 224256
rect 427964 224216 428740 224244
rect 427964 224204 427970 224216
rect 428734 224204 428740 224216
rect 428792 224204 428798 224256
rect 470226 224204 470232 224256
rect 470284 224244 470290 224256
rect 480438 224244 480444 224256
rect 470284 224216 480444 224244
rect 470284 224204 470290 224216
rect 480438 224204 480444 224216
rect 480496 224204 480502 224256
rect 486602 224204 486608 224256
rect 486660 224244 486666 224256
rect 500402 224244 500408 224256
rect 486660 224216 500408 224244
rect 486660 224204 486666 224216
rect 500402 224204 500408 224216
rect 500460 224204 500466 224256
rect 504358 224204 504364 224256
rect 504416 224244 504422 224256
rect 523494 224244 523500 224256
rect 504416 224216 523500 224244
rect 504416 224204 504422 224216
rect 523494 224204 523500 224216
rect 523552 224204 523558 224256
rect 525610 224204 525616 224256
rect 525668 224244 525674 224256
rect 532436 224244 532464 224352
rect 550634 224340 550640 224352
rect 550692 224340 550698 224392
rect 550818 224340 550824 224392
rect 550876 224380 550882 224392
rect 557506 224380 557534 224488
rect 625246 224476 625252 224488
rect 625304 224476 625310 224528
rect 667750 224408 667756 224460
rect 667808 224448 667814 224460
rect 667808 224420 671622 224448
rect 667808 224408 667814 224420
rect 550876 224352 557534 224380
rect 550876 224340 550882 224352
rect 557810 224340 557816 224392
rect 557868 224380 557874 224392
rect 625430 224380 625436 224392
rect 557868 224352 625436 224380
rect 557868 224340 557874 224352
rect 625430 224340 625436 224352
rect 625488 224340 625494 224392
rect 525668 224216 532464 224244
rect 525668 224204 525674 224216
rect 532694 224204 532700 224256
rect 532752 224244 532758 224256
rect 619634 224244 619640 224256
rect 532752 224216 619640 224244
rect 532752 224204 532758 224216
rect 619634 224204 619640 224216
rect 619692 224204 619698 224256
rect 651282 224204 651288 224256
rect 651340 224244 651346 224256
rect 658182 224244 658188 224256
rect 651340 224216 658188 224244
rect 651340 224204 651346 224216
rect 658182 224204 658188 224216
rect 658240 224204 658246 224256
rect 671482 224120 671534 224126
rect 362310 224108 362316 224120
rect 354646 224080 362316 224108
rect 362310 224068 362316 224080
rect 362368 224068 362374 224120
rect 377398 224068 377404 224120
rect 377456 224108 377462 224120
rect 385862 224108 385868 224120
rect 377456 224080 385868 224108
rect 377456 224068 377462 224080
rect 385862 224068 385868 224080
rect 385920 224068 385926 224120
rect 519078 224068 519084 224120
rect 519136 224108 519142 224120
rect 530670 224108 530676 224120
rect 519136 224080 530676 224108
rect 519136 224068 519142 224080
rect 530670 224068 530676 224080
rect 530728 224068 530734 224120
rect 530854 224068 530860 224120
rect 530912 224108 530918 224120
rect 534350 224108 534356 224120
rect 530912 224080 534356 224108
rect 530912 224068 530918 224080
rect 534350 224068 534356 224080
rect 534408 224068 534414 224120
rect 534534 224068 534540 224120
rect 534592 224108 534598 224120
rect 543734 224108 543740 224120
rect 534592 224080 543740 224108
rect 534592 224068 534598 224080
rect 543734 224068 543740 224080
rect 543792 224068 543798 224120
rect 667014 224068 667020 224120
rect 667072 224108 667078 224120
rect 667072 224080 670832 224108
rect 667072 224068 667078 224080
rect 543918 224000 543924 224052
rect 543976 224040 543982 224052
rect 545022 224040 545028 224052
rect 543976 224012 545028 224040
rect 543976 224000 543982 224012
rect 545022 224000 545028 224012
rect 545080 224040 545086 224052
rect 623774 224040 623780 224052
rect 545080 224012 623780 224040
rect 545080 224000 545086 224012
rect 623774 224000 623780 224012
rect 623832 224000 623838 224052
rect 670804 224040 670832 224080
rect 671482 224062 671534 224068
rect 670804 224012 671398 224040
rect 105998 223932 106004 223984
rect 106056 223972 106062 223984
rect 181070 223972 181076 223984
rect 106056 223944 181076 223972
rect 106056 223932 106062 223944
rect 181070 223932 181076 223944
rect 181128 223932 181134 223984
rect 201218 223932 201224 223984
rect 201276 223972 201282 223984
rect 255774 223972 255780 223984
rect 201276 223944 255780 223972
rect 201276 223932 201282 223944
rect 255774 223932 255780 223944
rect 255832 223932 255838 223984
rect 286686 223932 286692 223984
rect 286744 223972 286750 223984
rect 319530 223972 319536 223984
rect 286744 223944 319536 223972
rect 286744 223932 286750 223944
rect 319530 223932 319536 223944
rect 319588 223932 319594 223984
rect 667750 223932 667756 223984
rect 667808 223972 667814 223984
rect 667808 223944 670740 223972
rect 667808 223932 667814 223944
rect 279418 223864 279424 223916
rect 279476 223904 279482 223916
rect 284754 223904 284760 223916
rect 279476 223876 284760 223904
rect 279476 223864 279482 223876
rect 284754 223864 284760 223876
rect 284812 223864 284818 223916
rect 509694 223864 509700 223916
rect 509752 223904 509758 223916
rect 510154 223904 510160 223916
rect 509752 223876 510160 223904
rect 509752 223864 509758 223876
rect 510154 223864 510160 223876
rect 510212 223904 510218 223916
rect 610618 223904 610624 223916
rect 510212 223876 610624 223904
rect 510212 223864 510218 223876
rect 610618 223864 610624 223876
rect 610676 223864 610682 223916
rect 610802 223864 610808 223916
rect 610860 223904 610866 223916
rect 622670 223904 622676 223916
rect 610860 223876 622676 223904
rect 610860 223864 610866 223876
rect 622670 223864 622676 223876
rect 622728 223864 622734 223916
rect 108666 223796 108672 223848
rect 108724 223836 108730 223848
rect 183830 223836 183836 223848
rect 108724 223808 183836 223836
rect 108724 223796 108730 223808
rect 183830 223796 183836 223808
rect 183888 223796 183894 223848
rect 184842 223796 184848 223848
rect 184900 223836 184906 223848
rect 184900 223808 186314 223836
rect 184900 223796 184906 223808
rect 112806 223660 112812 223712
rect 112864 223700 112870 223712
rect 185946 223700 185952 223712
rect 112864 223672 185952 223700
rect 112864 223660 112870 223672
rect 185946 223660 185952 223672
rect 186004 223660 186010 223712
rect 186286 223700 186314 223808
rect 186958 223796 186964 223848
rect 187016 223836 187022 223848
rect 217778 223836 217784 223848
rect 187016 223808 217784 223836
rect 187016 223796 187022 223808
rect 217778 223796 217784 223808
rect 217836 223796 217842 223848
rect 228726 223796 228732 223848
rect 228784 223836 228790 223848
rect 274910 223836 274916 223848
rect 228784 223808 274916 223836
rect 228784 223796 228790 223808
rect 274910 223796 274916 223808
rect 274968 223796 274974 223848
rect 670712 223836 670740 223944
rect 670712 223808 671278 223836
rect 524414 223728 524420 223780
rect 524472 223768 524478 223780
rect 525058 223768 525064 223780
rect 524472 223740 525064 223768
rect 524472 223728 524478 223740
rect 525058 223728 525064 223740
rect 525116 223768 525122 223780
rect 532694 223768 532700 223780
rect 525116 223740 532700 223768
rect 525116 223728 525122 223740
rect 532694 223728 532700 223740
rect 532752 223728 532758 223780
rect 534994 223768 535000 223780
rect 534046 223740 535000 223768
rect 195422 223700 195428 223712
rect 186286 223672 195428 223700
rect 195422 223660 195428 223672
rect 195480 223660 195486 223712
rect 195882 223660 195888 223712
rect 195940 223700 195946 223712
rect 204898 223700 204904 223712
rect 195940 223672 204904 223700
rect 195940 223660 195946 223672
rect 204898 223660 204904 223672
rect 204956 223660 204962 223712
rect 238018 223660 238024 223712
rect 238076 223700 238082 223712
rect 266722 223700 266728 223712
rect 238076 223672 266728 223700
rect 238076 223660 238082 223672
rect 266722 223660 266728 223672
rect 266780 223660 266786 223712
rect 319622 223660 319628 223712
rect 319680 223700 319686 223712
rect 319990 223700 319996 223712
rect 319680 223672 319996 223700
rect 319680 223660 319686 223672
rect 319990 223660 319996 223672
rect 320048 223660 320054 223712
rect 530670 223592 530676 223644
rect 530728 223632 530734 223644
rect 534046 223632 534074 223740
rect 534994 223728 535000 223740
rect 535052 223768 535058 223780
rect 621566 223768 621572 223780
rect 535052 223740 621572 223768
rect 535052 223728 535058 223740
rect 621566 223728 621572 223740
rect 621624 223728 621630 223780
rect 530728 223604 534074 223632
rect 530728 223592 530734 223604
rect 534350 223592 534356 223644
rect 534408 223632 534414 223644
rect 538306 223632 538312 223644
rect 534408 223604 538312 223632
rect 534408 223592 534414 223604
rect 538306 223592 538312 223604
rect 538364 223592 538370 223644
rect 539962 223592 539968 223644
rect 540020 223632 540026 223644
rect 567838 223632 567844 223644
rect 540020 223604 567844 223632
rect 540020 223592 540026 223604
rect 567838 223592 567844 223604
rect 567896 223592 567902 223644
rect 568298 223592 568304 223644
rect 568356 223632 568362 223644
rect 628742 223632 628748 223644
rect 568356 223604 628748 223632
rect 568356 223592 568362 223604
rect 628742 223592 628748 223604
rect 628800 223592 628806 223644
rect 670418 223592 670424 223644
rect 670476 223632 670482 223644
rect 670476 223604 671186 223632
rect 670476 223592 670482 223604
rect 78582 223524 78588 223576
rect 78640 223564 78646 223576
rect 154022 223564 154028 223576
rect 78640 223536 154028 223564
rect 78640 223524 78646 223536
rect 154022 223524 154028 223536
rect 154080 223524 154086 223576
rect 154206 223524 154212 223576
rect 154264 223564 154270 223576
rect 161934 223564 161940 223576
rect 154264 223536 161940 223564
rect 154264 223524 154270 223536
rect 161934 223524 161940 223536
rect 161992 223524 161998 223576
rect 162118 223524 162124 223576
rect 162176 223564 162182 223576
rect 186590 223564 186596 223576
rect 162176 223536 186596 223564
rect 162176 223524 162182 223536
rect 186590 223524 186596 223536
rect 186648 223524 186654 223576
rect 187326 223524 187332 223576
rect 187384 223564 187390 223576
rect 242250 223564 242256 223576
rect 187384 223536 242256 223564
rect 187384 223524 187390 223536
rect 242250 223524 242256 223536
rect 242308 223524 242314 223576
rect 250898 223524 250904 223576
rect 250956 223564 250962 223576
rect 291194 223564 291200 223576
rect 250956 223536 291200 223564
rect 250956 223524 250962 223536
rect 291194 223524 291200 223536
rect 291252 223524 291258 223576
rect 297910 223524 297916 223576
rect 297968 223564 297974 223576
rect 303246 223564 303252 223576
rect 297968 223536 303252 223564
rect 297968 223524 297974 223536
rect 303246 223524 303252 223536
rect 303304 223524 303310 223576
rect 307662 223524 307668 223576
rect 307720 223564 307726 223576
rect 335630 223564 335636 223576
rect 307720 223536 335636 223564
rect 307720 223524 307726 223536
rect 335630 223524 335636 223536
rect 335688 223524 335694 223576
rect 406746 223524 406752 223576
rect 406804 223564 406810 223576
rect 414842 223564 414848 223576
rect 406804 223536 414848 223564
rect 406804 223524 406810 223536
rect 414842 223524 414848 223536
rect 414900 223524 414906 223576
rect 454862 223524 454868 223576
rect 454920 223564 454926 223576
rect 460474 223564 460480 223576
rect 454920 223536 460480 223564
rect 454920 223524 454926 223536
rect 460474 223524 460480 223536
rect 460532 223524 460538 223576
rect 473446 223524 473452 223576
rect 473504 223564 473510 223576
rect 475562 223564 475568 223576
rect 473504 223536 475568 223564
rect 473504 223524 473510 223536
rect 475562 223524 475568 223536
rect 475620 223524 475626 223576
rect 342070 223496 342076 223508
rect 335832 223468 342076 223496
rect 75822 223388 75828 223440
rect 75880 223428 75886 223440
rect 154942 223428 154948 223440
rect 75880 223400 154948 223428
rect 75880 223388 75886 223400
rect 154942 223388 154948 223400
rect 155000 223388 155006 223440
rect 155494 223388 155500 223440
rect 155552 223428 155558 223440
rect 159174 223428 159180 223440
rect 155552 223400 159180 223428
rect 155552 223388 155558 223400
rect 159174 223388 159180 223400
rect 159232 223388 159238 223440
rect 159358 223388 159364 223440
rect 159416 223428 159422 223440
rect 181806 223428 181812 223440
rect 159416 223400 181812 223428
rect 159416 223388 159422 223400
rect 181806 223388 181812 223400
rect 181864 223388 181870 223440
rect 184014 223388 184020 223440
rect 184072 223428 184078 223440
rect 239674 223428 239680 223440
rect 184072 223400 239680 223428
rect 184072 223388 184078 223400
rect 239674 223388 239680 223400
rect 239732 223388 239738 223440
rect 244090 223388 244096 223440
rect 244148 223428 244154 223440
rect 286042 223428 286048 223440
rect 244148 223400 286048 223428
rect 244148 223388 244154 223400
rect 286042 223388 286048 223400
rect 286100 223388 286106 223440
rect 304718 223388 304724 223440
rect 304776 223428 304782 223440
rect 308122 223428 308128 223440
rect 304776 223400 308128 223428
rect 304776 223388 304782 223400
rect 308122 223388 308128 223400
rect 308180 223388 308186 223440
rect 312906 223388 312912 223440
rect 312964 223428 312970 223440
rect 312964 223400 335354 223428
rect 312964 223388 312970 223400
rect 335326 223360 335354 223400
rect 335832 223360 335860 223468
rect 342070 223456 342076 223468
rect 342128 223456 342134 223508
rect 666646 223456 666652 223508
rect 666704 223496 666710 223508
rect 666704 223468 671048 223496
rect 666704 223456 666710 223468
rect 342806 223388 342812 223440
rect 342864 223428 342870 223440
rect 347866 223428 347872 223440
rect 342864 223400 347872 223428
rect 342864 223388 342870 223400
rect 347866 223388 347872 223400
rect 347924 223388 347930 223440
rect 517514 223388 517520 223440
rect 517572 223428 517578 223440
rect 531498 223428 531504 223440
rect 517572 223400 531504 223428
rect 517572 223388 517578 223400
rect 531498 223388 531504 223400
rect 531556 223388 531562 223440
rect 534718 223388 534724 223440
rect 534776 223428 534782 223440
rect 547414 223428 547420 223440
rect 534776 223400 547420 223428
rect 534776 223388 534782 223400
rect 547414 223388 547420 223400
rect 547472 223388 547478 223440
rect 561950 223388 561956 223440
rect 562008 223428 562014 223440
rect 568758 223428 568764 223440
rect 562008 223400 568764 223428
rect 562008 223388 562014 223400
rect 568758 223388 568764 223400
rect 568816 223388 568822 223440
rect 335326 223332 335860 223360
rect 335998 223320 336004 223372
rect 336056 223360 336062 223372
rect 342254 223360 342260 223372
rect 336056 223332 342260 223360
rect 336056 223320 336062 223332
rect 342254 223320 342260 223332
rect 342312 223320 342318 223372
rect 66898 223252 66904 223304
rect 66956 223292 66962 223304
rect 146662 223292 146668 223304
rect 66956 223264 146668 223292
rect 66956 223252 66962 223264
rect 146662 223252 146668 223264
rect 146720 223252 146726 223304
rect 147306 223252 147312 223304
rect 147364 223292 147370 223304
rect 176654 223292 176660 223304
rect 147364 223264 176660 223292
rect 147364 223252 147370 223264
rect 176654 223252 176660 223264
rect 176712 223252 176718 223304
rect 188890 223252 188896 223304
rect 188948 223292 188954 223304
rect 245102 223292 245108 223304
rect 188948 223264 245108 223292
rect 188948 223252 188954 223264
rect 245102 223252 245108 223264
rect 245160 223252 245166 223304
rect 246850 223252 246856 223304
rect 246908 223292 246914 223304
rect 288618 223292 288624 223304
rect 246908 223264 288624 223292
rect 246908 223252 246914 223264
rect 288618 223252 288624 223264
rect 288676 223252 288682 223304
rect 289722 223252 289728 223304
rect 289780 223292 289786 223304
rect 297726 223292 297732 223304
rect 289780 223264 297732 223292
rect 289780 223252 289786 223264
rect 297726 223252 297732 223264
rect 297784 223252 297790 223304
rect 299106 223252 299112 223304
rect 299164 223292 299170 223304
rect 328546 223292 328552 223304
rect 299164 223264 328552 223292
rect 299164 223252 299170 223264
rect 328546 223252 328552 223264
rect 328604 223252 328610 223304
rect 347222 223252 347228 223304
rect 347280 223292 347286 223304
rect 357894 223292 357900 223304
rect 347280 223264 357900 223292
rect 347280 223252 347286 223264
rect 357894 223252 357900 223264
rect 357952 223252 357958 223304
rect 483106 223252 483112 223304
rect 483164 223292 483170 223304
rect 496078 223292 496084 223304
rect 483164 223264 496084 223292
rect 483164 223252 483170 223264
rect 496078 223252 496084 223264
rect 496136 223252 496142 223304
rect 503346 223252 503352 223304
rect 503404 223292 503410 223304
rect 503404 223264 514064 223292
rect 503404 223252 503410 223264
rect 69566 223116 69572 223168
rect 69624 223156 69630 223168
rect 149514 223156 149520 223168
rect 69624 223128 149520 223156
rect 69624 223116 69630 223128
rect 149514 223116 149520 223128
rect 149572 223116 149578 223168
rect 152090 223156 152096 223168
rect 151786 223128 152096 223156
rect 71406 222980 71412 223032
rect 71464 223020 71470 223032
rect 151786 223020 151814 223128
rect 152090 223116 152096 223128
rect 152148 223116 152154 223168
rect 154390 223116 154396 223168
rect 154448 223156 154454 223168
rect 216214 223156 216220 223168
rect 154448 223128 216220 223156
rect 154448 223116 154454 223128
rect 216214 223116 216220 223128
rect 216272 223116 216278 223168
rect 241330 223116 241336 223168
rect 241388 223156 241394 223168
rect 283466 223156 283472 223168
rect 241388 223128 283472 223156
rect 241388 223116 241394 223128
rect 283466 223116 283472 223128
rect 283524 223116 283530 223168
rect 288250 223116 288256 223168
rect 288308 223156 288314 223168
rect 321094 223156 321100 223168
rect 288308 223128 321100 223156
rect 288308 223116 288314 223128
rect 321094 223116 321100 223128
rect 321152 223116 321158 223168
rect 344646 223116 344652 223168
rect 344704 223156 344710 223168
rect 364610 223156 364616 223168
rect 344704 223128 364616 223156
rect 344704 223116 344710 223128
rect 364610 223116 364616 223128
rect 364668 223116 364674 223168
rect 365530 223116 365536 223168
rect 365588 223156 365594 223168
rect 379606 223156 379612 223168
rect 365588 223128 379612 223156
rect 365588 223116 365594 223128
rect 379606 223116 379612 223128
rect 379664 223116 379670 223168
rect 380066 223116 380072 223168
rect 380124 223156 380130 223168
rect 386506 223156 386512 223168
rect 380124 223128 386512 223156
rect 380124 223116 380130 223128
rect 386506 223116 386512 223128
rect 386564 223116 386570 223168
rect 488626 223116 488632 223168
rect 488684 223156 488690 223168
rect 503162 223156 503168 223168
rect 488684 223128 503168 223156
rect 488684 223116 488690 223128
rect 503162 223116 503168 223128
rect 503220 223116 503226 223168
rect 508222 223116 508228 223168
rect 508280 223156 508286 223168
rect 514036 223156 514064 223264
rect 514662 223252 514668 223304
rect 514720 223292 514726 223304
rect 536282 223292 536288 223304
rect 514720 223264 536288 223292
rect 514720 223252 514726 223264
rect 536282 223252 536288 223264
rect 536340 223252 536346 223304
rect 554038 223252 554044 223304
rect 554096 223292 554102 223304
rect 562502 223292 562508 223304
rect 554096 223264 562508 223292
rect 554096 223252 554102 223264
rect 562502 223252 562508 223264
rect 562560 223252 562566 223304
rect 566826 223252 566832 223304
rect 566884 223292 566890 223304
rect 568298 223292 568304 223304
rect 566884 223264 568304 223292
rect 566884 223252 566890 223264
rect 568298 223252 568304 223264
rect 568356 223252 568362 223304
rect 586974 223252 586980 223304
rect 587032 223292 587038 223304
rect 593966 223292 593972 223304
rect 587032 223264 593972 223292
rect 587032 223252 587038 223264
rect 593966 223252 593972 223264
rect 594024 223252 594030 223304
rect 521746 223156 521752 223168
rect 508280 223128 509234 223156
rect 514036 223128 521752 223156
rect 508280 223116 508286 223128
rect 71464 222992 151814 223020
rect 71464 222980 71470 222992
rect 153654 222980 153660 223032
rect 153712 223020 153718 223032
rect 155494 223020 155500 223032
rect 153712 222992 155500 223020
rect 153712 222980 153718 222992
rect 155494 222980 155500 222992
rect 155552 222980 155558 223032
rect 155678 222980 155684 223032
rect 155736 223020 155742 223032
rect 219526 223020 219532 223032
rect 155736 222992 219532 223020
rect 155736 222980 155742 222992
rect 219526 222980 219532 222992
rect 219584 222980 219590 223032
rect 230198 222980 230204 223032
rect 230256 223020 230262 223032
rect 275462 223020 275468 223032
rect 230256 222992 275468 223020
rect 230256 222980 230262 222992
rect 275462 222980 275468 222992
rect 275520 222980 275526 223032
rect 278590 222980 278596 223032
rect 278648 223020 278654 223032
rect 315022 223020 315028 223032
rect 278648 222992 315028 223020
rect 278648 222980 278654 222992
rect 315022 222980 315028 222992
rect 315080 222980 315086 223032
rect 316678 222980 316684 223032
rect 316736 223020 316742 223032
rect 327258 223020 327264 223032
rect 316736 222992 327264 223020
rect 316736 222980 316742 222992
rect 327258 222980 327264 222992
rect 327316 222980 327322 223032
rect 328086 222980 328092 223032
rect 328144 223020 328150 223032
rect 351454 223020 351460 223032
rect 328144 222992 351460 223020
rect 328144 222980 328150 222992
rect 351454 222980 351460 222992
rect 351512 222980 351518 223032
rect 353938 222980 353944 223032
rect 353996 223020 354002 223032
rect 365898 223020 365904 223032
rect 353996 222992 365904 223020
rect 353996 222980 354002 222992
rect 365898 222980 365904 222992
rect 365956 222980 365962 223032
rect 366910 222980 366916 223032
rect 366968 223020 366974 223032
rect 383838 223020 383844 223032
rect 366968 222992 383844 223020
rect 366968 222980 366974 222992
rect 383838 222980 383844 222992
rect 383896 222980 383902 223032
rect 384206 222980 384212 223032
rect 384264 223020 384270 223032
rect 393958 223020 393964 223032
rect 384264 222992 393964 223020
rect 384264 222980 384270 222992
rect 393958 222980 393964 222992
rect 394016 222980 394022 223032
rect 493042 222980 493048 223032
rect 493100 223020 493106 223032
rect 508498 223020 508504 223032
rect 493100 222992 508504 223020
rect 493100 222980 493106 222992
rect 508498 222980 508504 222992
rect 508556 222980 508562 223032
rect 509206 223020 509234 223128
rect 521746 223116 521752 223128
rect 521804 223116 521810 223168
rect 532050 223116 532056 223168
rect 532108 223156 532114 223168
rect 559006 223156 559012 223168
rect 532108 223128 559012 223156
rect 532108 223116 532114 223128
rect 559006 223116 559012 223128
rect 559064 223116 559070 223168
rect 559834 223116 559840 223168
rect 559892 223156 559898 223168
rect 567654 223156 567660 223168
rect 559892 223128 567660 223156
rect 559892 223116 559898 223128
rect 567654 223116 567660 223128
rect 567712 223116 567718 223168
rect 620646 223156 620652 223168
rect 567856 223128 592034 223156
rect 527818 223020 527824 223032
rect 509206 222992 527824 223020
rect 527818 222980 527824 222992
rect 527876 222980 527882 223032
rect 529474 222980 529480 223032
rect 529532 223020 529538 223032
rect 555694 223020 555700 223032
rect 529532 222992 555700 223020
rect 529532 222980 529538 222992
rect 555694 222980 555700 222992
rect 555752 222980 555758 223032
rect 559374 222980 559380 223032
rect 559432 223020 559438 223032
rect 567856 223020 567884 223128
rect 559432 222992 567884 223020
rect 559432 222980 559438 222992
rect 568298 222980 568304 223032
rect 568356 223020 568362 223032
rect 587158 223020 587164 223032
rect 568356 222992 587164 223020
rect 568356 222980 568362 222992
rect 587158 222980 587164 222992
rect 587216 222980 587222 223032
rect 592006 223020 592034 223128
rect 605806 223128 620652 223156
rect 605806 223020 605834 223128
rect 620646 223116 620652 223128
rect 620704 223116 620710 223168
rect 667014 223116 667020 223168
rect 667072 223156 667078 223168
rect 667072 223128 670956 223156
rect 667072 223116 667078 223128
rect 592006 222992 605834 223020
rect 617334 222980 617340 223032
rect 617392 223020 617398 223032
rect 625614 223020 625620 223032
rect 617392 222992 625620 223020
rect 617392 222980 617398 222992
rect 625614 222980 625620 222992
rect 625672 222980 625678 223032
rect 62758 222844 62764 222896
rect 62816 222884 62822 222896
rect 141970 222884 141976 222896
rect 62816 222856 141976 222884
rect 62816 222844 62822 222856
rect 141970 222844 141976 222856
rect 142028 222844 142034 222896
rect 142154 222844 142160 222896
rect 142212 222884 142218 222896
rect 143994 222884 144000 222896
rect 142212 222856 144000 222884
rect 142212 222844 142218 222856
rect 143994 222844 144000 222856
rect 144052 222844 144058 222896
rect 146018 222844 146024 222896
rect 146076 222884 146082 222896
rect 211982 222884 211988 222896
rect 146076 222856 211988 222884
rect 146076 222844 146082 222856
rect 211982 222844 211988 222856
rect 212040 222844 212046 222896
rect 215938 222844 215944 222896
rect 215996 222884 216002 222896
rect 233326 222884 233332 222896
rect 215996 222856 233332 222884
rect 215996 222844 216002 222856
rect 233326 222844 233332 222856
rect 233384 222844 233390 222896
rect 234522 222844 234528 222896
rect 234580 222884 234586 222896
rect 281534 222884 281540 222896
rect 234580 222856 281540 222884
rect 234580 222844 234586 222856
rect 281534 222844 281540 222856
rect 281592 222844 281598 222896
rect 282454 222844 282460 222896
rect 282512 222884 282518 222896
rect 316310 222884 316316 222896
rect 282512 222856 316316 222884
rect 282512 222844 282518 222856
rect 316310 222844 316316 222856
rect 316368 222844 316374 222896
rect 324130 222844 324136 222896
rect 324188 222884 324194 222896
rect 348510 222884 348516 222896
rect 324188 222856 348516 222884
rect 324188 222844 324194 222856
rect 348510 222844 348516 222856
rect 348568 222844 348574 222896
rect 349062 222844 349068 222896
rect 349120 222884 349126 222896
rect 367186 222884 367192 222896
rect 349120 222856 367192 222884
rect 349120 222844 349126 222856
rect 367186 222844 367192 222856
rect 367244 222844 367250 222896
rect 368382 222844 368388 222896
rect 368440 222884 368446 222896
rect 382366 222884 382372 222896
rect 368440 222856 382372 222884
rect 368440 222844 368446 222856
rect 382366 222844 382372 222856
rect 382424 222844 382430 222896
rect 383470 222844 383476 222896
rect 383528 222884 383534 222896
rect 394878 222884 394884 222896
rect 383528 222856 394884 222884
rect 383528 222844 383534 222856
rect 394878 222844 394884 222856
rect 394936 222844 394942 222896
rect 395798 222844 395804 222896
rect 395856 222884 395862 222896
rect 406470 222884 406476 222896
rect 395856 222856 406476 222884
rect 395856 222844 395862 222856
rect 406470 222844 406476 222856
rect 406528 222844 406534 222896
rect 420822 222844 420828 222896
rect 420880 222884 420886 222896
rect 425146 222884 425152 222896
rect 420880 222856 425152 222884
rect 420880 222844 420886 222856
rect 425146 222844 425152 222856
rect 425204 222844 425210 222896
rect 459922 222844 459928 222896
rect 459980 222884 459986 222896
rect 467098 222884 467104 222896
rect 459980 222856 467104 222884
rect 459980 222844 459986 222856
rect 467098 222844 467104 222856
rect 467156 222844 467162 222896
rect 467466 222844 467472 222896
rect 467524 222884 467530 222896
rect 473722 222884 473728 222896
rect 467524 222856 473728 222884
rect 467524 222844 467530 222856
rect 473722 222844 473728 222856
rect 473780 222844 473786 222896
rect 479886 222844 479892 222896
rect 479944 222884 479950 222896
rect 491938 222884 491944 222896
rect 479944 222856 491944 222884
rect 479944 222844 479950 222856
rect 491938 222844 491944 222856
rect 491996 222844 492002 222896
rect 500770 222844 500776 222896
rect 500828 222884 500834 222896
rect 517514 222884 517520 222896
rect 500828 222856 517520 222884
rect 500828 222844 500834 222856
rect 517514 222844 517520 222856
rect 517572 222844 517578 222896
rect 519814 222844 519820 222896
rect 519872 222884 519878 222896
rect 542354 222884 542360 222896
rect 519872 222856 542360 222884
rect 519872 222844 519878 222856
rect 542354 222844 542360 222856
rect 542412 222844 542418 222896
rect 543826 222844 543832 222896
rect 543884 222884 543890 222896
rect 552474 222884 552480 222896
rect 543884 222856 552480 222884
rect 543884 222844 543890 222856
rect 552474 222844 552480 222856
rect 552532 222884 552538 222896
rect 562318 222884 562324 222896
rect 552532 222856 562324 222884
rect 552532 222844 552538 222856
rect 562318 222844 562324 222856
rect 562376 222844 562382 222896
rect 562502 222844 562508 222896
rect 562560 222884 562566 222896
rect 632698 222884 632704 222896
rect 562560 222856 632704 222884
rect 562560 222844 562566 222856
rect 632698 222844 632704 222856
rect 632756 222844 632762 222896
rect 81342 222708 81348 222760
rect 81400 222748 81406 222760
rect 153654 222748 153660 222760
rect 81400 222720 153660 222748
rect 81400 222708 81406 222720
rect 153654 222708 153660 222720
rect 153712 222708 153718 222760
rect 154022 222708 154028 222760
rect 154080 222748 154086 222760
rect 156966 222748 156972 222760
rect 154080 222720 156972 222748
rect 154080 222708 154086 222720
rect 156966 222708 156972 222720
rect 157024 222708 157030 222760
rect 166258 222708 166264 222760
rect 166316 222748 166322 222760
rect 192018 222748 192024 222760
rect 166316 222720 192024 222748
rect 166316 222708 166322 222720
rect 192018 222708 192024 222720
rect 192076 222708 192082 222760
rect 194502 222708 194508 222760
rect 194560 222748 194566 222760
rect 247402 222748 247408 222760
rect 194560 222720 247408 222748
rect 194560 222708 194566 222720
rect 247402 222708 247408 222720
rect 247460 222708 247466 222760
rect 264790 222708 264796 222760
rect 264848 222748 264854 222760
rect 304350 222748 304356 222760
rect 264848 222720 304356 222748
rect 264848 222708 264854 222720
rect 304350 222708 304356 222720
rect 304408 222708 304414 222760
rect 482738 222708 482744 222760
rect 482796 222748 482802 222760
rect 586974 222748 586980 222760
rect 482796 222720 586980 222748
rect 482796 222708 482802 222720
rect 586974 222708 586980 222720
rect 587032 222708 587038 222760
rect 587158 222708 587164 222760
rect 587216 222748 587222 222760
rect 587216 222720 620324 222748
rect 587216 222708 587222 222720
rect 99282 222572 99288 222624
rect 99340 222612 99346 222624
rect 175734 222612 175740 222624
rect 99340 222584 175740 222612
rect 99340 222572 99346 222584
rect 175734 222572 175740 222584
rect 175792 222572 175798 222624
rect 197170 222572 197176 222624
rect 197228 222612 197234 222624
rect 249978 222612 249984 222624
rect 197228 222584 249984 222612
rect 197228 222572 197234 222584
rect 249978 222572 249984 222584
rect 250036 222572 250042 222624
rect 557534 222572 557540 222624
rect 557592 222612 557598 222624
rect 559834 222612 559840 222624
rect 557592 222584 559840 222612
rect 557592 222572 557598 222584
rect 559834 222572 559840 222584
rect 559892 222572 559898 222624
rect 562318 222572 562324 222624
rect 562376 222612 562382 222624
rect 617334 222612 617340 222624
rect 562376 222584 617340 222612
rect 562376 222572 562382 222584
rect 617334 222572 617340 222584
rect 617392 222572 617398 222624
rect 620296 222612 620324 222720
rect 620462 222708 620468 222760
rect 620520 222748 620526 222760
rect 627086 222748 627092 222760
rect 620520 222720 627092 222748
rect 620520 222708 620526 222720
rect 627086 222708 627092 222720
rect 627144 222708 627150 222760
rect 629846 222612 629852 222624
rect 620296 222584 629852 222612
rect 629846 222572 629852 222584
rect 629904 222572 629910 222624
rect 175918 222504 175924 222556
rect 175976 222544 175982 222556
rect 175976 222516 190454 222544
rect 175976 222504 175982 222516
rect 87966 222436 87972 222488
rect 88024 222476 88030 222488
rect 164970 222476 164976 222488
rect 88024 222448 164976 222476
rect 88024 222436 88030 222448
rect 164970 222436 164976 222448
rect 165028 222436 165034 222488
rect 190426 222476 190454 222516
rect 207474 222476 207480 222488
rect 190426 222448 207480 222476
rect 207474 222436 207480 222448
rect 207532 222436 207538 222488
rect 207658 222436 207664 222488
rect 207716 222476 207722 222488
rect 258350 222476 258356 222488
rect 207716 222448 258356 222476
rect 207716 222436 207722 222448
rect 258350 222436 258356 222448
rect 258408 222436 258414 222488
rect 489914 222436 489920 222488
rect 489972 222476 489978 222488
rect 491110 222476 491116 222488
rect 489972 222448 491116 222476
rect 489972 222436 489978 222448
rect 491110 222436 491116 222448
rect 491168 222476 491174 222488
rect 491168 222448 499574 222476
rect 491168 222436 491174 222448
rect 172146 222368 172152 222420
rect 172204 222408 172210 222420
rect 172204 222380 186314 222408
rect 172204 222368 172210 222380
rect 85298 222300 85304 222352
rect 85356 222340 85362 222352
rect 154206 222340 154212 222352
rect 85356 222312 154212 222340
rect 85356 222300 85362 222312
rect 154206 222300 154212 222312
rect 154264 222300 154270 222352
rect 186286 222340 186314 222380
rect 199746 222340 199752 222352
rect 186286 222312 199752 222340
rect 199746 222300 199752 222312
rect 199804 222300 199810 222352
rect 211798 222300 211804 222352
rect 211856 222340 211862 222352
rect 228082 222340 228088 222352
rect 211856 222312 228088 222340
rect 211856 222300 211862 222312
rect 228082 222300 228088 222312
rect 228140 222300 228146 222352
rect 287882 222300 287888 222352
rect 287940 222340 287946 222352
rect 295058 222340 295064 222352
rect 287940 222312 295064 222340
rect 287940 222300 287946 222312
rect 295058 222300 295064 222312
rect 295116 222300 295122 222352
rect 484486 222300 484492 222352
rect 484544 222340 484550 222352
rect 499546 222340 499574 222448
rect 504358 222436 504364 222488
rect 504416 222476 504422 222488
rect 523678 222476 523684 222488
rect 504416 222448 523684 222476
rect 504416 222436 504422 222448
rect 523678 222436 523684 222448
rect 523736 222436 523742 222488
rect 529842 222436 529848 222488
rect 529900 222476 529906 222488
rect 619910 222476 619916 222488
rect 529900 222448 619916 222476
rect 529900 222436 529906 222448
rect 619910 222436 619916 222448
rect 619968 222436 619974 222488
rect 568298 222340 568304 222352
rect 484544 222312 485774 222340
rect 499546 222312 568304 222340
rect 484544 222300 484550 222312
rect 156616 222244 179276 222272
rect 118418 222164 118424 222216
rect 118476 222204 118482 222216
rect 141970 222204 141976 222216
rect 118476 222176 141976 222204
rect 118476 222164 118482 222176
rect 141970 222164 141976 222176
rect 142028 222164 142034 222216
rect 142154 222164 142160 222216
rect 142212 222204 142218 222216
rect 156616 222204 156644 222244
rect 142212 222176 156644 222204
rect 179248 222204 179276 222244
rect 191006 222204 191012 222216
rect 179248 222176 191012 222204
rect 142212 222164 142218 222176
rect 191006 222164 191012 222176
rect 191064 222164 191070 222216
rect 485746 222204 485774 222312
rect 568298 222300 568304 222312
rect 568356 222300 568362 222352
rect 568758 222300 568764 222352
rect 568816 222340 568822 222352
rect 627914 222340 627920 222352
rect 568816 222312 627920 222340
rect 568816 222300 568822 222312
rect 627914 222300 627920 222312
rect 627972 222300 627978 222352
rect 504358 222204 504364 222216
rect 485746 222176 504364 222204
rect 504358 222164 504364 222176
rect 504416 222164 504422 222216
rect 523678 222164 523684 222216
rect 523736 222204 523742 222216
rect 559374 222204 559380 222216
rect 523736 222176 559380 222204
rect 523736 222164 523742 222176
rect 559374 222164 559380 222176
rect 559432 222164 559438 222216
rect 567654 222164 567660 222216
rect 567712 222204 567718 222216
rect 620462 222204 620468 222216
rect 567712 222176 620468 222204
rect 567712 222164 567718 222176
rect 620462 222164 620468 222176
rect 620520 222164 620526 222216
rect 620646 222164 620652 222216
rect 620704 222204 620710 222216
rect 631502 222204 631508 222216
rect 620704 222176 631508 222204
rect 620704 222164 620710 222176
rect 631502 222164 631508 222176
rect 631560 222164 631566 222216
rect 160830 222096 160836 222148
rect 160888 222136 160894 222148
rect 166074 222136 166080 222148
rect 160888 222108 166080 222136
rect 160888 222096 160894 222108
rect 166074 222096 166080 222108
rect 166132 222096 166138 222148
rect 172698 222136 172704 222148
rect 166276 222108 172704 222136
rect 97902 221960 97908 222012
rect 97960 222000 97966 222012
rect 166276 222000 166304 222108
rect 172698 222096 172704 222108
rect 172756 222096 172762 222148
rect 174078 222096 174084 222148
rect 174136 222136 174142 222148
rect 174136 222108 179184 222136
rect 174136 222096 174142 222108
rect 179156 222068 179184 222108
rect 191466 222096 191472 222148
rect 191524 222136 191530 222148
rect 247586 222136 247592 222148
rect 191524 222108 247592 222136
rect 191524 222096 191530 222108
rect 247586 222096 247592 222108
rect 247644 222096 247650 222148
rect 258074 222096 258080 222148
rect 258132 222136 258138 222148
rect 263686 222136 263692 222148
rect 258132 222108 263692 222136
rect 258132 222096 258138 222108
rect 263686 222096 263692 222108
rect 263744 222096 263750 222148
rect 270034 222096 270040 222148
rect 270092 222136 270098 222148
rect 306374 222136 306380 222148
rect 270092 222108 306380 222136
rect 270092 222096 270098 222108
rect 306374 222096 306380 222108
rect 306432 222096 306438 222148
rect 310698 222096 310704 222148
rect 310756 222136 310762 222148
rect 312630 222136 312636 222148
rect 310756 222108 312636 222136
rect 310756 222096 310762 222108
rect 312630 222096 312636 222108
rect 312688 222096 312694 222148
rect 331398 222096 331404 222148
rect 331456 222136 331462 222148
rect 353754 222136 353760 222148
rect 331456 222108 353760 222136
rect 331456 222096 331462 222108
rect 353754 222096 353760 222108
rect 353812 222096 353818 222148
rect 424962 222096 424968 222148
rect 425020 222136 425026 222148
rect 429286 222136 429292 222148
rect 425020 222108 429292 222136
rect 425020 222096 425026 222108
rect 429286 222096 429292 222108
rect 429344 222096 429350 222148
rect 452562 222096 452568 222148
rect 452620 222136 452626 222148
rect 455598 222136 455604 222148
rect 452620 222108 455604 222136
rect 452620 222096 452626 222108
rect 455598 222096 455604 222108
rect 455656 222096 455662 222148
rect 462130 222096 462136 222148
rect 462188 222136 462194 222148
rect 468754 222136 468760 222148
rect 462188 222108 468760 222136
rect 462188 222096 462194 222108
rect 468754 222096 468760 222108
rect 468812 222096 468818 222148
rect 471882 222096 471888 222148
rect 471940 222136 471946 222148
rect 477862 222136 477868 222148
rect 471940 222108 477868 222136
rect 471940 222096 471946 222108
rect 477862 222096 477868 222108
rect 477920 222096 477926 222148
rect 559558 222096 559564 222148
rect 559616 222136 559622 222148
rect 564802 222136 564808 222148
rect 559616 222108 564808 222136
rect 559616 222096 559622 222108
rect 564802 222096 564808 222108
rect 564860 222096 564866 222148
rect 179156 222040 186314 222068
rect 97960 221972 166304 222000
rect 97960 221960 97966 221972
rect 166994 221960 167000 222012
rect 167052 222000 167058 222012
rect 169754 222000 169760 222012
rect 167052 221972 169760 222000
rect 167052 221960 167058 221972
rect 169754 221960 169760 221972
rect 169812 221960 169818 222012
rect 171778 221960 171784 222012
rect 171836 222000 171842 222012
rect 178954 222000 178960 222012
rect 171836 221972 178960 222000
rect 171836 221960 171842 221972
rect 178954 221960 178960 221972
rect 179012 221960 179018 222012
rect 186286 222000 186314 222040
rect 495158 222028 495164 222080
rect 495216 222068 495222 222080
rect 497734 222068 497740 222080
rect 495216 222040 497740 222068
rect 495216 222028 495222 222040
rect 497734 222028 497740 222040
rect 497792 222028 497798 222080
rect 515490 222028 515496 222080
rect 515548 222068 515554 222080
rect 529842 222068 529848 222080
rect 515548 222040 529848 222068
rect 515548 222028 515554 222040
rect 529842 222028 529848 222040
rect 529900 222028 529906 222080
rect 533982 222028 533988 222080
rect 534040 222068 534046 222080
rect 559374 222068 559380 222080
rect 534040 222040 559380 222068
rect 534040 222028 534046 222040
rect 559374 222028 559380 222040
rect 559432 222028 559438 222080
rect 592034 222028 592040 222080
rect 592092 222068 592098 222080
rect 596634 222068 596640 222080
rect 592092 222040 596640 222068
rect 592092 222028 592098 222040
rect 596634 222028 596640 222040
rect 596692 222028 596698 222080
rect 596818 222028 596824 222080
rect 596876 222068 596882 222080
rect 605006 222068 605012 222080
rect 596876 222040 605012 222068
rect 596876 222028 596882 222040
rect 605006 222028 605012 222040
rect 605064 222028 605070 222080
rect 231854 222000 231860 222012
rect 186286 221972 231860 222000
rect 231854 221960 231860 221972
rect 231912 221960 231918 222012
rect 233694 221960 233700 222012
rect 233752 222000 233758 222012
rect 277946 222000 277952 222012
rect 233752 221972 277952 222000
rect 233752 221960 233758 221972
rect 277946 221960 277952 221972
rect 278004 221960 278010 222012
rect 280062 221960 280068 222012
rect 280120 222000 280126 222012
rect 314010 222000 314016 222012
rect 280120 221972 314016 222000
rect 280120 221960 280126 221972
rect 314010 221960 314016 221972
rect 314068 221960 314074 222012
rect 318242 221960 318248 222012
rect 318300 222000 318306 222012
rect 343818 222000 343824 222012
rect 318300 221972 343824 222000
rect 318300 221960 318306 221972
rect 343818 221960 343824 221972
rect 343876 221960 343882 222012
rect 367646 221960 367652 222012
rect 367704 222000 367710 222012
rect 380250 222000 380256 222012
rect 367704 221972 380256 222000
rect 367704 221960 367710 221972
rect 380250 221960 380256 221972
rect 380308 221960 380314 222012
rect 536098 221892 536104 221944
rect 536156 221932 536162 221944
rect 543688 221932 543694 221944
rect 536156 221904 543694 221932
rect 536156 221892 536162 221904
rect 543688 221892 543694 221904
rect 543746 221892 543752 221944
rect 557166 221892 557172 221944
rect 557224 221932 557230 221944
rect 608594 221932 608600 221944
rect 557224 221904 608600 221932
rect 557224 221892 557230 221904
rect 608594 221892 608600 221904
rect 608652 221892 608658 221944
rect 104526 221824 104532 221876
rect 104584 221864 104590 221876
rect 176286 221864 176292 221876
rect 104584 221836 176292 221864
rect 104584 221824 104590 221836
rect 176286 221824 176292 221836
rect 176344 221824 176350 221876
rect 182634 221864 182640 221876
rect 176626 221836 182640 221864
rect 80514 221688 80520 221740
rect 80572 221728 80578 221740
rect 86218 221728 86224 221740
rect 80572 221700 86224 221728
rect 80572 221688 80578 221700
rect 86218 221688 86224 221700
rect 86276 221688 86282 221740
rect 94682 221688 94688 221740
rect 94740 221728 94746 221740
rect 161428 221728 161434 221740
rect 94740 221700 161434 221728
rect 94740 221688 94746 221700
rect 161428 221688 161434 221700
rect 161486 221688 161492 221740
rect 161566 221688 161572 221740
rect 161624 221728 161630 221740
rect 167178 221728 167184 221740
rect 161624 221700 167184 221728
rect 161624 221688 161630 221700
rect 167178 221688 167184 221700
rect 167236 221688 167242 221740
rect 167454 221688 167460 221740
rect 167512 221728 167518 221740
rect 171410 221728 171416 221740
rect 167512 221700 171416 221728
rect 167512 221688 167518 221700
rect 171410 221688 171416 221700
rect 171468 221688 171474 221740
rect 171594 221688 171600 221740
rect 171652 221728 171658 221740
rect 176626 221728 176654 221836
rect 182634 221824 182640 221836
rect 182692 221824 182698 221876
rect 182818 221824 182824 221876
rect 182876 221864 182882 221876
rect 240134 221864 240140 221876
rect 182876 221836 240140 221864
rect 182876 221824 182882 221836
rect 240134 221824 240140 221836
rect 240192 221824 240198 221876
rect 263318 221824 263324 221876
rect 263376 221864 263382 221876
rect 301222 221864 301228 221876
rect 263376 221836 301228 221864
rect 263376 221824 263382 221836
rect 301222 221824 301228 221836
rect 301280 221824 301286 221876
rect 301406 221824 301412 221876
rect 301464 221864 301470 221876
rect 310882 221864 310888 221876
rect 301464 221836 310888 221864
rect 301464 221824 301470 221836
rect 310882 221824 310888 221836
rect 310940 221824 310946 221876
rect 313182 221824 313188 221876
rect 313240 221864 313246 221876
rect 340414 221864 340420 221876
rect 313240 221836 340420 221864
rect 313240 221824 313246 221836
rect 340414 221824 340420 221836
rect 340472 221824 340478 221876
rect 351270 221824 351276 221876
rect 351328 221864 351334 221876
rect 369302 221864 369308 221876
rect 351328 221836 369308 221864
rect 351328 221824 351334 221836
rect 369302 221824 369308 221836
rect 369360 221824 369366 221876
rect 509878 221824 509884 221876
rect 509936 221864 509942 221876
rect 522666 221864 522672 221876
rect 509936 221836 522672 221864
rect 509936 221824 509942 221836
rect 522666 221824 522672 221836
rect 522724 221824 522730 221876
rect 546586 221864 546592 221876
rect 544166 221836 546592 221864
rect 544166 221796 544194 221836
rect 546586 221824 546592 221836
rect 546644 221824 546650 221876
rect 547138 221824 547144 221876
rect 547196 221864 547202 221876
rect 556798 221864 556804 221876
rect 547196 221836 556804 221864
rect 547196 221824 547202 221836
rect 556798 221824 556804 221836
rect 556856 221824 556862 221876
rect 543844 221768 544194 221796
rect 171652 221700 176654 221728
rect 171652 221688 171658 221700
rect 178954 221688 178960 221740
rect 179012 221728 179018 221740
rect 232222 221728 232228 221740
rect 179012 221700 232228 221728
rect 179012 221688 179018 221700
rect 232222 221688 232228 221700
rect 232280 221688 232286 221740
rect 239214 221688 239220 221740
rect 239272 221728 239278 221740
rect 283650 221728 283656 221740
rect 239272 221700 283656 221728
rect 239272 221688 239278 221700
rect 283650 221688 283656 221700
rect 283708 221688 283714 221740
rect 303246 221688 303252 221740
rect 303304 221728 303310 221740
rect 332778 221728 332784 221740
rect 303304 221700 332784 221728
rect 303304 221688 303310 221700
rect 332778 221688 332784 221700
rect 332836 221688 332842 221740
rect 357158 221688 357164 221740
rect 357216 221728 357222 221740
rect 374638 221728 374644 221740
rect 357216 221700 374644 221728
rect 357216 221688 357222 221700
rect 374638 221688 374644 221700
rect 374696 221688 374702 221740
rect 391014 221688 391020 221740
rect 391072 221728 391078 221740
rect 400306 221728 400312 221740
rect 391072 221700 400312 221728
rect 391072 221688 391078 221700
rect 400306 221688 400312 221700
rect 400364 221688 400370 221740
rect 475838 221688 475844 221740
rect 475896 221728 475902 221740
rect 486142 221728 486148 221740
rect 475896 221700 486148 221728
rect 475896 221688 475902 221700
rect 486142 221688 486148 221700
rect 486200 221688 486206 221740
rect 496262 221688 496268 221740
rect 496320 221728 496326 221740
rect 513558 221728 513564 221740
rect 496320 221700 513564 221728
rect 496320 221688 496326 221700
rect 513558 221688 513564 221700
rect 513616 221688 513622 221740
rect 522850 221688 522856 221740
rect 522908 221728 522914 221740
rect 543844 221728 543872 221768
rect 522908 221700 543872 221728
rect 522908 221688 522914 221700
rect 549254 221688 549260 221740
rect 549312 221728 549318 221740
rect 606662 221728 606668 221740
rect 549312 221700 606668 221728
rect 549312 221688 549318 221700
rect 606662 221688 606668 221700
rect 606720 221688 606726 221740
rect 59354 221552 59360 221604
rect 59412 221592 59418 221604
rect 138290 221592 138296 221604
rect 59412 221564 138296 221592
rect 59412 221552 59418 221564
rect 138290 221552 138296 221564
rect 138348 221552 138354 221604
rect 138474 221552 138480 221604
rect 138532 221592 138538 221604
rect 140774 221592 140780 221604
rect 138532 221564 140780 221592
rect 138532 221552 138538 221564
rect 140774 221552 140780 221564
rect 140832 221552 140838 221604
rect 140958 221552 140964 221604
rect 141016 221592 141022 221604
rect 205910 221592 205916 221604
rect 141016 221564 205916 221592
rect 141016 221552 141022 221564
rect 205910 221552 205916 221564
rect 205968 221552 205974 221604
rect 208394 221552 208400 221604
rect 208452 221592 208458 221604
rect 260834 221592 260840 221604
rect 208452 221564 260840 221592
rect 208452 221552 208458 221564
rect 260834 221552 260840 221564
rect 260892 221552 260898 221604
rect 261018 221552 261024 221604
rect 261076 221592 261082 221604
rect 301774 221592 301780 221604
rect 261076 221564 301780 221592
rect 261076 221552 261082 221564
rect 301774 221552 301780 221564
rect 301832 221552 301838 221604
rect 308858 221552 308864 221604
rect 308916 221592 308922 221604
rect 339678 221592 339684 221604
rect 308916 221564 339684 221592
rect 308916 221552 308922 221564
rect 339678 221552 339684 221564
rect 339736 221552 339742 221604
rect 341334 221552 341340 221604
rect 341392 221592 341398 221604
rect 361758 221592 361764 221604
rect 341392 221564 361764 221592
rect 341392 221552 341398 221564
rect 361758 221552 361764 221564
rect 361816 221552 361822 221604
rect 369486 221552 369492 221604
rect 369544 221592 369550 221604
rect 384022 221592 384028 221604
rect 369544 221564 384028 221592
rect 369544 221552 369550 221564
rect 384022 221552 384028 221564
rect 384080 221552 384086 221604
rect 384390 221552 384396 221604
rect 384448 221592 384454 221604
rect 395154 221592 395160 221604
rect 384448 221564 395160 221592
rect 384448 221552 384454 221564
rect 395154 221552 395160 221564
rect 395212 221552 395218 221604
rect 400766 221552 400772 221604
rect 400824 221592 400830 221604
rect 405734 221592 405740 221604
rect 400824 221564 405740 221592
rect 400824 221552 400830 221564
rect 405734 221552 405740 221564
rect 405792 221552 405798 221604
rect 480806 221552 480812 221604
rect 480864 221592 480870 221604
rect 492950 221592 492956 221604
rect 480864 221564 492956 221592
rect 480864 221552 480870 221564
rect 492950 221552 492956 221564
rect 493008 221552 493014 221604
rect 497458 221552 497464 221604
rect 497516 221592 497522 221604
rect 515122 221592 515128 221604
rect 497516 221564 515128 221592
rect 497516 221552 497522 221564
rect 515122 221552 515128 221564
rect 515180 221552 515186 221604
rect 524230 221552 524236 221604
rect 524288 221592 524294 221604
rect 524288 221564 533476 221592
rect 524288 221552 524294 221564
rect 73890 221416 73896 221468
rect 73948 221456 73954 221468
rect 82078 221456 82084 221468
rect 73948 221428 82084 221456
rect 73948 221416 73954 221428
rect 82078 221416 82084 221428
rect 82136 221416 82142 221468
rect 86310 221416 86316 221468
rect 86368 221456 86374 221468
rect 86368 221428 161612 221456
rect 86368 221416 86374 221428
rect 91278 221280 91284 221332
rect 91336 221320 91342 221332
rect 91336 221292 118004 221320
rect 91336 221280 91342 221292
rect 117976 221184 118004 221292
rect 118142 221280 118148 221332
rect 118200 221320 118206 221332
rect 127434 221320 127440 221332
rect 118200 221292 127440 221320
rect 118200 221280 118206 221292
rect 127434 221280 127440 221292
rect 127492 221280 127498 221332
rect 161428 221320 161434 221332
rect 127636 221292 161434 221320
rect 127636 221184 127664 221292
rect 161428 221280 161434 221292
rect 161486 221280 161492 221332
rect 161584 221320 161612 221428
rect 161750 221416 161756 221468
rect 161808 221456 161814 221468
rect 161808 221428 171824 221456
rect 161808 221416 161814 221428
rect 164418 221320 164424 221332
rect 161584 221292 164424 221320
rect 164418 221280 164424 221292
rect 164476 221280 164482 221332
rect 171594 221320 171600 221332
rect 164712 221292 171600 221320
rect 164712 221184 164740 221292
rect 171594 221280 171600 221292
rect 171652 221280 171658 221332
rect 171796 221320 171824 221428
rect 171962 221416 171968 221468
rect 172020 221456 172026 221468
rect 226518 221456 226524 221468
rect 172020 221428 226524 221456
rect 172020 221416 172026 221428
rect 226518 221416 226524 221428
rect 226576 221416 226582 221468
rect 227898 221416 227904 221468
rect 227956 221456 227962 221468
rect 276106 221456 276112 221468
rect 227956 221428 276112 221456
rect 227956 221416 227962 221428
rect 276106 221416 276112 221428
rect 276164 221416 276170 221468
rect 292482 221416 292488 221468
rect 292540 221456 292546 221468
rect 326246 221456 326252 221468
rect 292540 221428 326252 221456
rect 292540 221416 292546 221428
rect 326246 221416 326252 221428
rect 326304 221416 326310 221468
rect 342162 221416 342168 221468
rect 342220 221456 342226 221468
rect 364794 221456 364800 221468
rect 342220 221428 364800 221456
rect 342220 221416 342226 221428
rect 364794 221416 364800 221428
rect 364852 221416 364858 221468
rect 375282 221416 375288 221468
rect 375340 221456 375346 221468
rect 390738 221456 390744 221468
rect 375340 221428 390744 221456
rect 375340 221416 375346 221428
rect 390738 221416 390744 221428
rect 390796 221416 390802 221468
rect 396810 221416 396816 221468
rect 396868 221456 396874 221468
rect 407298 221456 407304 221468
rect 396868 221428 407304 221456
rect 396868 221416 396874 221428
rect 407298 221416 407304 221428
rect 407356 221416 407362 221468
rect 408402 221416 408408 221468
rect 408460 221456 408466 221468
rect 416866 221456 416872 221468
rect 408460 221428 416872 221456
rect 408460 221416 408466 221428
rect 416866 221416 416872 221428
rect 416924 221416 416930 221468
rect 468938 221416 468944 221468
rect 468996 221456 469002 221468
rect 476206 221456 476212 221468
rect 468996 221428 476212 221456
rect 468996 221416 469002 221428
rect 476206 221416 476212 221428
rect 476264 221416 476270 221468
rect 483750 221416 483756 221468
rect 483808 221456 483814 221468
rect 533246 221456 533252 221468
rect 483808 221428 533252 221456
rect 483808 221416 483814 221428
rect 533246 221416 533252 221428
rect 533304 221416 533310 221468
rect 533448 221456 533476 221564
rect 533614 221552 533620 221604
rect 533672 221592 533678 221604
rect 601970 221592 601976 221604
rect 533672 221564 601976 221592
rect 533672 221552 533678 221564
rect 601970 221552 601976 221564
rect 602028 221552 602034 221604
rect 533448 221428 536696 221456
rect 536668 221388 536696 221428
rect 543706 221428 548748 221456
rect 536668 221360 536788 221388
rect 193306 221320 193312 221332
rect 171796 221292 193312 221320
rect 193306 221280 193312 221292
rect 193364 221280 193370 221332
rect 204162 221280 204168 221332
rect 204220 221320 204226 221332
rect 252738 221320 252744 221332
rect 204220 221292 252744 221320
rect 204220 221280 204226 221292
rect 252738 221280 252744 221292
rect 252796 221280 252802 221332
rect 266814 221280 266820 221332
rect 266872 221320 266878 221332
rect 303798 221320 303804 221332
rect 266872 221292 303804 221320
rect 266872 221280 266878 221292
rect 303798 221280 303804 221292
rect 303856 221280 303862 221332
rect 523494 221280 523500 221332
rect 523552 221320 523558 221332
rect 533154 221320 533160 221332
rect 523552 221292 533160 221320
rect 523552 221280 523558 221292
rect 533154 221280 533160 221292
rect 533212 221280 533218 221332
rect 536760 221252 536788 221360
rect 538674 221348 538680 221400
rect 538732 221388 538738 221400
rect 543706 221388 543734 221428
rect 538732 221360 543734 221388
rect 538732 221348 538738 221360
rect 543642 221252 543648 221264
rect 536760 221224 543648 221252
rect 543642 221212 543648 221224
rect 543700 221212 543706 221264
rect 543826 221212 543832 221264
rect 543884 221252 543890 221264
rect 548518 221252 548524 221264
rect 543884 221224 548524 221252
rect 543884 221212 543890 221224
rect 548518 221212 548524 221224
rect 548576 221212 548582 221264
rect 548720 221252 548748 221428
rect 597002 221416 597008 221468
rect 597060 221456 597066 221468
rect 633434 221456 633440 221468
rect 597060 221428 633440 221456
rect 597060 221416 597066 221428
rect 633434 221416 633440 221428
rect 633492 221416 633498 221468
rect 548886 221348 548892 221400
rect 548944 221388 548950 221400
rect 596818 221388 596824 221400
rect 548944 221360 596824 221388
rect 548944 221348 548950 221360
rect 596818 221348 596824 221360
rect 596876 221348 596882 221400
rect 669774 221348 669780 221400
rect 669832 221348 669838 221400
rect 604638 221252 604644 221264
rect 548720 221224 604644 221252
rect 604638 221212 604644 221224
rect 604696 221212 604702 221264
rect 117976 221156 127664 221184
rect 127728 221156 164740 221184
rect 111150 221008 111156 221060
rect 111208 221048 111214 221060
rect 118142 221048 118148 221060
rect 111208 221020 118148 221048
rect 111208 221008 111214 221020
rect 118142 221008 118148 221020
rect 118200 221008 118206 221060
rect 124398 221008 124404 221060
rect 124456 221048 124462 221060
rect 127250 221048 127256 221060
rect 124456 221020 127256 221048
rect 124456 221008 124462 221020
rect 127250 221008 127256 221020
rect 127308 221008 127314 221060
rect 127434 221008 127440 221060
rect 127492 221048 127498 221060
rect 127728 221048 127756 221156
rect 166074 221144 166080 221196
rect 166132 221184 166138 221196
rect 221274 221184 221280 221196
rect 166132 221156 221280 221184
rect 166132 221144 166138 221156
rect 221274 221144 221280 221156
rect 221332 221144 221338 221196
rect 222746 221144 222752 221196
rect 222804 221184 222810 221196
rect 268286 221184 268292 221196
rect 222804 221156 268292 221184
rect 222804 221144 222810 221156
rect 268286 221144 268292 221156
rect 268344 221144 268350 221196
rect 669792 221128 669820 221348
rect 521102 221076 521108 221128
rect 521160 221116 521166 221128
rect 591942 221116 591948 221128
rect 521160 221088 591948 221116
rect 521160 221076 521166 221088
rect 591942 221076 591948 221088
rect 592000 221076 592006 221128
rect 592126 221076 592132 221128
rect 592184 221116 592190 221128
rect 600406 221116 600412 221128
rect 592184 221088 600412 221116
rect 592184 221076 592190 221088
rect 600406 221076 600412 221088
rect 600464 221076 600470 221128
rect 669774 221076 669780 221128
rect 669832 221076 669838 221128
rect 127492 221020 127756 221048
rect 127492 221008 127498 221020
rect 127894 221008 127900 221060
rect 127952 221048 127958 221060
rect 127952 221020 145788 221048
rect 127952 221008 127958 221020
rect 145760 220980 145788 221020
rect 146386 221008 146392 221060
rect 146444 221048 146450 221060
rect 206462 221048 206468 221060
rect 146444 221020 206468 221048
rect 146444 221008 146450 221020
rect 206462 221008 206468 221020
rect 206520 221008 206526 221060
rect 219802 221008 219808 221060
rect 219860 221048 219866 221060
rect 263042 221048 263048 221060
rect 219860 221020 263048 221048
rect 219860 221008 219866 221020
rect 263042 221008 263048 221020
rect 263100 221008 263106 221060
rect 145760 220952 145880 220980
rect 82998 220872 83004 220924
rect 83056 220912 83062 220924
rect 142108 220912 142114 220924
rect 83056 220884 142114 220912
rect 83056 220872 83062 220884
rect 142108 220872 142114 220884
rect 142166 220872 142172 220924
rect 142246 220872 142252 220924
rect 142304 220912 142310 220924
rect 145558 220912 145564 220924
rect 142304 220884 145564 220912
rect 142304 220872 142310 220884
rect 145558 220872 145564 220884
rect 145616 220872 145622 220924
rect 145852 220912 145880 220952
rect 525978 220940 525984 220992
rect 526036 220980 526042 220992
rect 601786 220980 601792 220992
rect 526036 220952 601792 220980
rect 526036 220940 526042 220952
rect 601786 220940 601792 220952
rect 601844 220940 601850 220992
rect 161428 220912 161434 220924
rect 145852 220884 161434 220912
rect 161428 220872 161434 220884
rect 161486 220872 161492 220924
rect 161566 220872 161572 220924
rect 161624 220912 161630 220924
rect 222286 220912 222292 220924
rect 161624 220884 222292 220912
rect 161624 220872 161630 220884
rect 222286 220872 222292 220884
rect 222344 220872 222350 220924
rect 282638 220872 282644 220924
rect 282696 220912 282702 220924
rect 287698 220912 287704 220924
rect 282696 220884 287704 220912
rect 282696 220872 282702 220884
rect 287698 220872 287704 220884
rect 287756 220872 287762 220924
rect 456702 220872 456708 220924
rect 456760 220912 456766 220924
rect 456760 220884 460934 220912
rect 456760 220872 456766 220884
rect 253842 220804 253848 220856
rect 253900 220844 253906 220856
rect 258626 220844 258632 220856
rect 253900 220816 258632 220844
rect 253900 220804 253906 220816
rect 258626 220804 258632 220816
rect 258684 220804 258690 220856
rect 418338 220804 418344 220856
rect 418396 220844 418402 220856
rect 424042 220844 424048 220856
rect 418396 220816 424048 220844
rect 418396 220804 418402 220816
rect 424042 220804 424048 220816
rect 424100 220804 424106 220856
rect 460906 220844 460934 220884
rect 466086 220872 466092 220924
rect 466144 220912 466150 220924
rect 471422 220912 471428 220924
rect 466144 220884 471428 220912
rect 466144 220872 466150 220884
rect 471422 220872 471428 220884
rect 471480 220872 471486 220924
rect 669406 220872 669412 220924
rect 669464 220872 669470 220924
rect 462130 220844 462136 220856
rect 460906 220816 462136 220844
rect 462130 220804 462136 220816
rect 462188 220804 462194 220856
rect 517514 220804 517520 220856
rect 517572 220844 517578 220856
rect 518526 220844 518532 220856
rect 517572 220816 518532 220844
rect 517572 220804 517578 220816
rect 518526 220804 518532 220816
rect 518584 220844 518590 220856
rect 592034 220844 592040 220856
rect 518584 220816 592040 220844
rect 518584 220804 518590 220816
rect 592034 220804 592040 220816
rect 592092 220804 592098 220856
rect 596910 220804 596916 220856
rect 596968 220844 596974 220856
rect 600682 220844 600688 220856
rect 596968 220816 600688 220844
rect 596968 220804 596974 220816
rect 600682 220804 600688 220816
rect 600740 220804 600746 220856
rect 669424 220788 669452 220872
rect 114278 220736 114284 220788
rect 114336 220776 114342 220788
rect 145834 220776 145840 220788
rect 114336 220748 145840 220776
rect 114336 220736 114342 220748
rect 145834 220736 145840 220748
rect 145892 220736 145898 220788
rect 146938 220736 146944 220788
rect 146996 220776 147002 220788
rect 177206 220776 177212 220788
rect 146996 220748 177212 220776
rect 146996 220736 147002 220748
rect 177206 220736 177212 220748
rect 177264 220736 177270 220788
rect 177390 220736 177396 220788
rect 177448 220776 177454 220788
rect 181254 220776 181260 220788
rect 177448 220748 181260 220776
rect 177448 220736 177454 220748
rect 181254 220736 181260 220748
rect 181312 220736 181318 220788
rect 181438 220736 181444 220788
rect 181496 220776 181502 220788
rect 190362 220776 190368 220788
rect 181496 220748 190368 220776
rect 181496 220736 181502 220748
rect 190362 220736 190368 220748
rect 190420 220736 190426 220788
rect 190546 220736 190552 220788
rect 190604 220776 190610 220788
rect 236638 220776 236644 220788
rect 190604 220748 236644 220776
rect 190604 220736 190610 220748
rect 236638 220736 236644 220748
rect 236696 220736 236702 220788
rect 242618 220736 242624 220788
rect 242676 220776 242682 220788
rect 246482 220776 246488 220788
rect 242676 220748 246488 220776
rect 242676 220736 242682 220748
rect 246482 220736 246488 220748
rect 246540 220736 246546 220788
rect 260190 220736 260196 220788
rect 260248 220776 260254 220788
rect 298554 220776 298560 220788
rect 260248 220748 298560 220776
rect 260248 220736 260254 220748
rect 298554 220736 298560 220748
rect 298612 220736 298618 220788
rect 302418 220736 302424 220788
rect 302476 220776 302482 220788
rect 334066 220776 334072 220788
rect 302476 220748 334072 220776
rect 302476 220736 302482 220748
rect 334066 220736 334072 220748
rect 334124 220736 334130 220788
rect 385218 220736 385224 220788
rect 385276 220776 385282 220788
rect 388714 220776 388720 220788
rect 385276 220748 388720 220776
rect 385276 220736 385282 220748
rect 388714 220736 388720 220748
rect 388772 220736 388778 220788
rect 414198 220736 414204 220788
rect 414256 220776 414262 220788
rect 418154 220776 418160 220788
rect 414256 220748 418160 220776
rect 414256 220736 414262 220748
rect 418154 220736 418160 220748
rect 418212 220736 418218 220788
rect 455322 220736 455328 220788
rect 455380 220776 455386 220788
rect 458818 220776 458824 220788
rect 455380 220748 458824 220776
rect 455380 220736 455386 220748
rect 458818 220736 458824 220748
rect 458876 220736 458882 220788
rect 465718 220736 465724 220788
rect 465776 220776 465782 220788
rect 469582 220776 469588 220788
rect 465776 220748 469588 220776
rect 465776 220736 465782 220748
rect 469582 220736 469588 220748
rect 469640 220736 469646 220788
rect 473998 220736 474004 220788
rect 474056 220776 474062 220788
rect 475378 220776 475384 220788
rect 474056 220748 475384 220776
rect 474056 220736 474062 220748
rect 475378 220736 475384 220748
rect 475436 220736 475442 220788
rect 476758 220736 476764 220788
rect 476816 220776 476822 220788
rect 478690 220776 478696 220788
rect 476816 220748 478696 220776
rect 476816 220736 476822 220748
rect 478690 220736 478696 220748
rect 478748 220736 478754 220788
rect 511810 220736 511816 220788
rect 511868 220776 511874 220788
rect 596726 220776 596732 220788
rect 511868 220748 512040 220776
rect 511868 220736 511874 220748
rect 512012 220708 512040 220748
rect 592236 220748 596732 220776
rect 512012 220680 518894 220708
rect 101214 220600 101220 220652
rect 101272 220640 101278 220652
rect 175090 220640 175096 220652
rect 101272 220612 175096 220640
rect 101272 220600 101278 220612
rect 175090 220600 175096 220612
rect 175148 220600 175154 220652
rect 175274 220600 175280 220652
rect 175332 220640 175338 220652
rect 224218 220640 224224 220652
rect 175332 220612 224224 220640
rect 175332 220600 175338 220612
rect 224218 220600 224224 220612
rect 224276 220600 224282 220652
rect 253566 220600 253572 220652
rect 253624 220640 253630 220652
rect 293310 220640 293316 220652
rect 253624 220612 293316 220640
rect 253624 220600 253630 220612
rect 293310 220600 293316 220612
rect 293368 220600 293374 220652
rect 294966 220600 294972 220652
rect 295024 220640 295030 220652
rect 325878 220640 325884 220652
rect 295024 220612 325884 220640
rect 295024 220600 295030 220612
rect 325878 220600 325884 220612
rect 325936 220600 325942 220652
rect 357894 220600 357900 220652
rect 357952 220640 357958 220652
rect 374454 220640 374460 220652
rect 357952 220612 374460 220640
rect 357952 220600 357958 220612
rect 374454 220600 374460 220612
rect 374512 220600 374518 220652
rect 500218 220600 500224 220652
rect 500276 220640 500282 220652
rect 511810 220640 511816 220652
rect 500276 220612 511816 220640
rect 500276 220600 500282 220612
rect 511810 220600 511816 220612
rect 511868 220600 511874 220652
rect 332686 220532 332692 220584
rect 332744 220572 332750 220584
rect 337194 220572 337200 220584
rect 332744 220544 337200 220572
rect 332744 220532 332750 220544
rect 337194 220532 337200 220544
rect 337252 220532 337258 220584
rect 69750 220464 69756 220516
rect 69808 220504 69814 220516
rect 136910 220504 136916 220516
rect 69808 220476 136916 220504
rect 69808 220464 69814 220476
rect 136910 220464 136916 220476
rect 136968 220464 136974 220516
rect 137094 220464 137100 220516
rect 137152 220504 137158 220516
rect 146938 220504 146944 220516
rect 137152 220476 146944 220504
rect 137152 220464 137158 220476
rect 146938 220464 146944 220476
rect 146996 220464 147002 220516
rect 147122 220464 147128 220516
rect 147180 220504 147186 220516
rect 208578 220504 208584 220516
rect 147180 220476 208584 220504
rect 147180 220464 147186 220476
rect 208578 220464 208584 220476
rect 208636 220464 208642 220516
rect 210510 220464 210516 220516
rect 210568 220504 210574 220516
rect 259914 220504 259920 220516
rect 210568 220476 259920 220504
rect 210568 220464 210574 220476
rect 259914 220464 259920 220476
rect 259972 220464 259978 220516
rect 267642 220464 267648 220516
rect 267700 220504 267706 220516
rect 306834 220504 306840 220516
rect 267700 220476 306840 220504
rect 267700 220464 267706 220476
rect 306834 220464 306840 220476
rect 306892 220464 306898 220516
rect 338022 220464 338028 220516
rect 338080 220504 338086 220516
rect 358998 220504 359004 220516
rect 338080 220476 359004 220504
rect 338080 220464 338086 220476
rect 358998 220464 359004 220476
rect 359056 220464 359062 220516
rect 469122 220464 469128 220516
rect 469180 220504 469186 220516
rect 474550 220504 474556 220516
rect 469180 220476 474556 220504
rect 469180 220464 469186 220476
rect 474550 220464 474556 220476
rect 474608 220464 474614 220516
rect 488442 220464 488448 220516
rect 488500 220504 488506 220516
rect 501874 220504 501880 220516
rect 488500 220476 501880 220504
rect 488500 220464 488506 220476
rect 501874 220464 501880 220476
rect 501932 220464 501938 220516
rect 518866 220504 518894 220680
rect 543642 220668 543648 220720
rect 543700 220708 543706 220720
rect 549070 220708 549076 220720
rect 543700 220680 549076 220708
rect 543700 220668 543706 220680
rect 549070 220668 549076 220680
rect 549128 220668 549134 220720
rect 520918 220600 520924 220652
rect 520976 220640 520982 220652
rect 537478 220640 537484 220652
rect 520976 220612 537484 220640
rect 520976 220600 520982 220612
rect 537478 220600 537484 220612
rect 537536 220600 537542 220652
rect 551002 220600 551008 220652
rect 551060 220640 551066 220652
rect 554222 220640 554228 220652
rect 551060 220612 554228 220640
rect 551060 220600 551066 220612
rect 554222 220600 554228 220612
rect 554280 220600 554286 220652
rect 555694 220600 555700 220652
rect 555752 220640 555758 220652
rect 562870 220640 562876 220652
rect 555752 220612 562876 220640
rect 555752 220600 555758 220612
rect 562870 220600 562876 220612
rect 562928 220600 562934 220652
rect 563054 220600 563060 220652
rect 563112 220640 563118 220652
rect 587342 220640 587348 220652
rect 563112 220612 587348 220640
rect 563112 220600 563118 220612
rect 587342 220600 587348 220612
rect 587400 220600 587406 220652
rect 587526 220600 587532 220652
rect 587584 220640 587590 220652
rect 592236 220640 592264 220748
rect 596726 220736 596732 220748
rect 596784 220736 596790 220788
rect 669406 220736 669412 220788
rect 669464 220736 669470 220788
rect 669866 220736 669872 220788
rect 669924 220776 669930 220788
rect 670234 220776 670240 220788
rect 669924 220748 670240 220776
rect 669924 220736 669930 220748
rect 670234 220736 670240 220748
rect 670292 220736 670298 220788
rect 587584 220612 592264 220640
rect 587584 220600 587590 220612
rect 538306 220532 538312 220584
rect 538364 220572 538370 220584
rect 543826 220572 543832 220584
rect 538364 220544 543832 220572
rect 538364 220532 538370 220544
rect 543826 220532 543832 220544
rect 543884 220532 543890 220584
rect 531682 220504 531688 220516
rect 518866 220476 531688 220504
rect 531682 220464 531688 220476
rect 531740 220464 531746 220516
rect 556522 220504 556528 220516
rect 546650 220476 556528 220504
rect 73062 220328 73068 220380
rect 73120 220368 73126 220380
rect 145650 220368 145656 220380
rect 73120 220340 145656 220368
rect 73120 220328 73126 220340
rect 145650 220328 145656 220340
rect 145708 220328 145714 220380
rect 145834 220328 145840 220380
rect 145892 220368 145898 220380
rect 153470 220368 153476 220380
rect 145892 220340 153476 220368
rect 145892 220328 145898 220340
rect 153470 220328 153476 220340
rect 153528 220328 153534 220380
rect 154390 220328 154396 220380
rect 154448 220368 154454 220380
rect 214098 220368 214104 220380
rect 154448 220340 214104 220368
rect 154448 220328 154454 220340
rect 214098 220328 214104 220340
rect 214156 220328 214162 220380
rect 214282 220328 214288 220380
rect 214340 220368 214346 220380
rect 214340 220340 224264 220368
rect 214340 220328 214346 220340
rect 79686 220192 79692 220244
rect 79744 220232 79750 220244
rect 158898 220232 158904 220244
rect 79744 220204 158904 220232
rect 79744 220192 79750 220204
rect 158898 220192 158904 220204
rect 158956 220192 158962 220244
rect 164142 220192 164148 220244
rect 164200 220232 164206 220244
rect 223666 220232 223672 220244
rect 164200 220204 223672 220232
rect 164200 220192 164206 220204
rect 223666 220192 223672 220204
rect 223724 220192 223730 220244
rect 224236 220232 224264 220340
rect 224402 220328 224408 220380
rect 224460 220368 224466 220380
rect 267918 220368 267924 220380
rect 224460 220340 267924 220368
rect 224460 220328 224466 220340
rect 267918 220328 267924 220340
rect 267976 220328 267982 220380
rect 273438 220328 273444 220380
rect 273496 220368 273502 220380
rect 309226 220368 309232 220380
rect 273496 220340 309232 220368
rect 273496 220328 273502 220340
rect 309226 220328 309232 220340
rect 309284 220328 309290 220380
rect 314838 220328 314844 220380
rect 314896 220368 314902 220380
rect 341058 220368 341064 220380
rect 314896 220340 341064 220368
rect 314896 220328 314902 220340
rect 341058 220328 341064 220340
rect 341116 220328 341122 220380
rect 342990 220328 342996 220380
rect 343048 220368 343054 220380
rect 363322 220368 363328 220380
rect 343048 220340 363328 220368
rect 343048 220328 343054 220340
rect 363322 220328 363328 220340
rect 363380 220328 363386 220380
rect 472986 220328 472992 220380
rect 473044 220368 473050 220380
rect 481174 220368 481180 220380
rect 473044 220340 481180 220368
rect 473044 220328 473050 220340
rect 481174 220328 481180 220340
rect 481232 220328 481238 220380
rect 496446 220328 496452 220380
rect 496504 220368 496510 220380
rect 509326 220368 509332 220380
rect 496504 220340 509332 220368
rect 496504 220328 496510 220340
rect 509326 220328 509332 220340
rect 509384 220328 509390 220380
rect 516962 220328 516968 220380
rect 517020 220368 517026 220380
rect 527542 220368 527548 220380
rect 517020 220340 527548 220368
rect 517020 220328 517026 220340
rect 527542 220328 527548 220340
rect 527600 220328 527606 220380
rect 531222 220328 531228 220380
rect 531280 220368 531286 220380
rect 546650 220368 546678 220476
rect 556522 220464 556528 220476
rect 556580 220464 556586 220516
rect 562134 220504 562140 220516
rect 557506 220476 562140 220504
rect 554038 220368 554044 220380
rect 531280 220340 546678 220368
rect 548536 220340 554044 220368
rect 531280 220328 531286 220340
rect 234154 220232 234160 220244
rect 224236 220204 234160 220232
rect 234154 220192 234160 220204
rect 234212 220192 234218 220244
rect 237006 220192 237012 220244
rect 237064 220232 237070 220244
rect 280430 220232 280436 220244
rect 237064 220204 280436 220232
rect 237064 220192 237070 220204
rect 280430 220192 280436 220204
rect 280488 220192 280494 220244
rect 283374 220192 283380 220244
rect 283432 220232 283438 220244
rect 316494 220232 316500 220244
rect 283432 220204 316500 220232
rect 283432 220192 283438 220204
rect 316494 220192 316500 220204
rect 316552 220192 316558 220244
rect 321646 220192 321652 220244
rect 321704 220232 321710 220244
rect 324498 220232 324504 220244
rect 321704 220204 324504 220232
rect 321704 220192 321710 220204
rect 324498 220192 324504 220204
rect 324556 220192 324562 220244
rect 342622 220232 342628 220244
rect 324700 220204 342628 220232
rect 76374 220056 76380 220108
rect 76432 220096 76438 220108
rect 156138 220096 156144 220108
rect 76432 220068 156144 220096
rect 76432 220056 76438 220068
rect 156138 220056 156144 220068
rect 156196 220056 156202 220108
rect 157518 220056 157524 220108
rect 157576 220096 157582 220108
rect 214098 220096 214104 220108
rect 157576 220068 214104 220096
rect 157576 220056 157582 220068
rect 214098 220056 214104 220068
rect 214156 220056 214162 220108
rect 244274 220096 244280 220108
rect 214484 220068 244280 220096
rect 107838 219920 107844 219972
rect 107896 219960 107902 219972
rect 114278 219960 114284 219972
rect 107896 219932 114284 219960
rect 107896 219920 107902 219932
rect 114278 219920 114284 219932
rect 114336 219920 114342 219972
rect 114462 219920 114468 219972
rect 114520 219960 114526 219972
rect 114520 219932 126744 219960
rect 114520 219920 114526 219932
rect 121086 219784 121092 219836
rect 121144 219824 121150 219836
rect 126716 219824 126744 219932
rect 127618 219920 127624 219972
rect 127676 219960 127682 219972
rect 181438 219960 181444 219972
rect 127676 219932 181444 219960
rect 127676 219920 127682 219932
rect 181438 219920 181444 219932
rect 181496 219920 181502 219972
rect 181622 219920 181628 219972
rect 181680 219960 181686 219972
rect 214282 219960 214288 219972
rect 181680 219932 214288 219960
rect 181680 219920 181686 219932
rect 214282 219920 214288 219932
rect 214340 219920 214346 219972
rect 137094 219824 137100 219836
rect 121144 219796 122834 219824
rect 126716 219796 137100 219824
rect 121144 219784 121150 219796
rect 122806 219688 122834 219796
rect 137094 219784 137100 219796
rect 137152 219784 137158 219836
rect 197630 219824 197636 219836
rect 137296 219796 197636 219824
rect 127618 219688 127624 219700
rect 122806 219660 127624 219688
rect 127618 219648 127624 219660
rect 127676 219648 127682 219700
rect 131022 219648 131028 219700
rect 131080 219688 131086 219700
rect 137296 219688 137324 219796
rect 197630 219784 197636 219796
rect 197688 219784 197694 219836
rect 197814 219784 197820 219836
rect 197872 219824 197878 219836
rect 214484 219824 214512 220068
rect 244274 220056 244280 220068
rect 244332 220056 244338 220108
rect 244458 220056 244464 220108
rect 244516 220096 244522 220108
rect 288526 220096 288532 220108
rect 244516 220068 288532 220096
rect 244516 220056 244522 220068
rect 288526 220056 288532 220068
rect 288584 220056 288590 220108
rect 288710 220056 288716 220108
rect 288768 220096 288774 220108
rect 288768 220068 316034 220096
rect 288768 220056 288774 220068
rect 254762 219960 254768 219972
rect 197872 219796 214512 219824
rect 214576 219932 254768 219960
rect 197872 219784 197878 219796
rect 144638 219688 144644 219700
rect 131080 219660 137324 219688
rect 137388 219660 144644 219688
rect 131080 219648 131086 219660
rect 136910 219512 136916 219564
rect 136968 219552 136974 219564
rect 137388 219552 137416 219660
rect 144638 219648 144644 219660
rect 144696 219648 144702 219700
rect 144822 219648 144828 219700
rect 144880 219688 144886 219700
rect 146754 219688 146760 219700
rect 144880 219660 146760 219688
rect 144880 219648 144886 219660
rect 146754 219648 146760 219660
rect 146812 219648 146818 219700
rect 203150 219688 203156 219700
rect 146956 219660 203156 219688
rect 136968 219524 137416 219552
rect 136968 219512 136974 219524
rect 137646 219512 137652 219564
rect 137704 219552 137710 219564
rect 146956 219552 146984 219660
rect 203150 219648 203156 219660
rect 203208 219648 203214 219700
rect 203886 219648 203892 219700
rect 203944 219688 203950 219700
rect 214576 219688 214604 219932
rect 254762 219920 254768 219932
rect 254820 219920 254826 219972
rect 316006 219960 316034 220068
rect 316494 220056 316500 220108
rect 316552 220096 316558 220108
rect 324700 220096 324728 220204
rect 342622 220192 342628 220204
rect 342680 220192 342686 220244
rect 348786 220192 348792 220244
rect 348844 220232 348850 220244
rect 369946 220232 369952 220244
rect 348844 220204 369952 220232
rect 348844 220192 348850 220204
rect 369946 220192 369952 220204
rect 370004 220192 370010 220244
rect 370498 220192 370504 220244
rect 370556 220232 370562 220244
rect 381078 220232 381084 220244
rect 370556 220204 381084 220232
rect 370556 220192 370562 220204
rect 381078 220192 381084 220204
rect 381136 220192 381142 220244
rect 388714 220192 388720 220244
rect 388772 220232 388778 220244
rect 400950 220232 400956 220244
rect 388772 220204 400956 220232
rect 388772 220192 388778 220204
rect 400950 220192 400956 220204
rect 401008 220192 401014 220244
rect 432230 220192 432236 220244
rect 432288 220232 432294 220244
rect 434806 220232 434812 220244
rect 432288 220204 434812 220232
rect 432288 220192 432294 220204
rect 434806 220192 434812 220204
rect 434864 220192 434870 220244
rect 459462 220192 459468 220244
rect 459520 220232 459526 220244
rect 465442 220232 465448 220244
rect 459520 220204 465448 220232
rect 459520 220192 459526 220204
rect 465442 220192 465448 220204
rect 465500 220192 465506 220244
rect 473170 220192 473176 220244
rect 473228 220232 473234 220244
rect 482002 220232 482008 220244
rect 473228 220204 482008 220232
rect 473228 220192 473234 220204
rect 482002 220192 482008 220204
rect 482060 220192 482066 220244
rect 482922 220192 482928 220244
rect 482980 220232 482986 220244
rect 495250 220232 495256 220244
rect 482980 220204 495256 220232
rect 482980 220192 482986 220204
rect 495250 220192 495256 220204
rect 495308 220192 495314 220244
rect 501322 220192 501328 220244
rect 501380 220232 501386 220244
rect 520182 220232 520188 220244
rect 501380 220204 520188 220232
rect 501380 220192 501386 220204
rect 520182 220192 520188 220204
rect 520240 220192 520246 220244
rect 528370 220192 528376 220244
rect 528428 220232 528434 220244
rect 548536 220232 548564 220340
rect 554038 220328 554044 220340
rect 554096 220328 554102 220380
rect 554222 220328 554228 220380
rect 554280 220368 554286 220380
rect 557506 220368 557534 220476
rect 562134 220464 562140 220476
rect 562192 220464 562198 220516
rect 562428 220476 567516 220504
rect 554280 220340 557534 220368
rect 554280 220328 554286 220340
rect 558270 220328 558276 220380
rect 558328 220368 558334 220380
rect 561766 220368 561772 220380
rect 558328 220340 561772 220368
rect 558328 220328 558334 220340
rect 561766 220328 561772 220340
rect 561824 220328 561830 220380
rect 562428 220300 562456 220476
rect 566826 220328 566832 220380
rect 566884 220368 566890 220380
rect 567286 220368 567292 220380
rect 566884 220340 567292 220368
rect 566884 220328 566890 220340
rect 567286 220328 567292 220340
rect 567344 220328 567350 220380
rect 567488 220368 567516 220476
rect 568574 220464 568580 220516
rect 568632 220504 568638 220516
rect 569770 220504 569776 220516
rect 568632 220476 569776 220504
rect 568632 220464 568638 220476
rect 569770 220464 569776 220476
rect 569828 220464 569834 220516
rect 572668 220464 572674 220516
rect 572726 220504 572732 220516
rect 610526 220504 610532 220516
rect 572726 220476 610532 220504
rect 572726 220464 572732 220476
rect 610526 220464 610532 220476
rect 610584 220464 610590 220516
rect 572346 220368 572352 220380
rect 567488 220340 572352 220368
rect 572346 220328 572352 220340
rect 572404 220328 572410 220380
rect 574738 220328 574744 220380
rect 574796 220368 574802 220380
rect 611446 220368 611452 220380
rect 574796 220340 611452 220368
rect 574796 220328 574802 220340
rect 611446 220328 611452 220340
rect 611504 220328 611510 220380
rect 562382 220272 562456 220300
rect 528428 220204 548564 220232
rect 528428 220192 528434 220204
rect 548702 220192 548708 220244
rect 548760 220232 548766 220244
rect 562382 220232 562410 220272
rect 548760 220204 562410 220232
rect 548760 220192 548766 220204
rect 562870 220192 562876 220244
rect 562928 220232 562934 220244
rect 608962 220232 608968 220244
rect 562928 220204 608968 220232
rect 562928 220192 562934 220204
rect 608962 220192 608968 220204
rect 609020 220192 609026 220244
rect 316552 220068 324728 220096
rect 316552 220056 316558 220068
rect 325602 220056 325608 220108
rect 325660 220096 325666 220108
rect 352098 220096 352104 220108
rect 325660 220068 352104 220096
rect 325660 220056 325666 220068
rect 352098 220056 352104 220068
rect 352156 220056 352162 220108
rect 358814 220056 358820 220108
rect 358872 220096 358878 220108
rect 378318 220096 378324 220108
rect 358872 220068 378324 220096
rect 358872 220056 358878 220068
rect 378318 220056 378324 220068
rect 378376 220056 378382 220108
rect 379422 220056 379428 220108
rect 379480 220096 379486 220108
rect 392118 220096 392124 220108
rect 379480 220068 392124 220096
rect 379480 220056 379486 220068
rect 392118 220056 392124 220068
rect 392176 220056 392182 220108
rect 395982 220056 395988 220108
rect 396040 220096 396046 220108
rect 404722 220096 404728 220108
rect 396040 220068 404728 220096
rect 396040 220056 396046 220068
rect 404722 220056 404728 220068
rect 404780 220056 404786 220108
rect 421650 220056 421656 220108
rect 421708 220096 421714 220108
rect 426802 220096 426808 220108
rect 421708 220068 426808 220096
rect 421708 220056 421714 220068
rect 426802 220056 426808 220068
rect 426860 220056 426866 220108
rect 478322 220056 478328 220108
rect 478380 220096 478386 220108
rect 489454 220096 489460 220108
rect 478380 220068 489460 220096
rect 478380 220056 478386 220068
rect 489454 220056 489460 220068
rect 489512 220056 489518 220108
rect 492490 220056 492496 220108
rect 492548 220096 492554 220108
rect 506842 220096 506848 220108
rect 492548 220068 506848 220096
rect 492548 220056 492554 220068
rect 506842 220056 506848 220068
rect 506900 220056 506906 220108
rect 513098 220056 513104 220108
rect 513156 220096 513162 220108
rect 534166 220096 534172 220108
rect 513156 220068 534172 220096
rect 513156 220056 513162 220068
rect 534166 220056 534172 220068
rect 534224 220056 534230 220108
rect 538122 220056 538128 220108
rect 538180 220096 538186 220108
rect 561766 220096 561772 220108
rect 538180 220068 561772 220096
rect 538180 220056 538186 220068
rect 561766 220056 561772 220068
rect 561824 220056 561830 220108
rect 587342 220056 587348 220108
rect 587400 220096 587406 220108
rect 608778 220096 608784 220108
rect 587400 220068 608784 220096
rect 587400 220056 587406 220068
rect 608778 220056 608784 220068
rect 608836 220056 608842 220108
rect 562134 219988 562140 220040
rect 562192 220028 562198 220040
rect 562192 220000 587204 220028
rect 562192 219988 562198 220000
rect 322382 219960 322388 219972
rect 316006 219932 322388 219960
rect 322382 219920 322388 219932
rect 322440 219920 322446 219972
rect 587176 219960 587204 220000
rect 587176 219932 592034 219960
rect 503622 219852 503628 219904
rect 503680 219892 503686 219904
rect 586974 219892 586980 219904
rect 503680 219864 586980 219892
rect 503680 219852 503686 219864
rect 586974 219852 586980 219864
rect 587032 219852 587038 219904
rect 592006 219892 592034 219932
rect 607306 219892 607312 219904
rect 592006 219864 607312 219892
rect 607306 219852 607312 219864
rect 607364 219852 607370 219904
rect 217134 219784 217140 219836
rect 217192 219824 217198 219836
rect 265158 219824 265164 219836
rect 217192 219796 265164 219824
rect 217192 219784 217198 219796
rect 265158 219784 265164 219796
rect 265216 219784 265222 219836
rect 548702 219756 548708 219768
rect 528526 219728 548708 219756
rect 203944 219660 214604 219688
rect 203944 219648 203950 219660
rect 220446 219648 220452 219700
rect 220504 219688 220510 219700
rect 224402 219688 224408 219700
rect 220504 219660 224408 219688
rect 220504 219648 220510 219660
rect 224402 219648 224408 219660
rect 224460 219648 224466 219700
rect 227070 219648 227076 219700
rect 227128 219688 227134 219700
rect 272702 219688 272708 219700
rect 227128 219660 272708 219688
rect 227128 219648 227134 219660
rect 272702 219648 272708 219660
rect 272760 219648 272766 219700
rect 464982 219580 464988 219632
rect 465040 219620 465046 219632
rect 472066 219620 472072 219632
rect 465040 219592 472072 219620
rect 465040 219580 465046 219592
rect 472066 219580 472072 219592
rect 472124 219580 472130 219632
rect 527542 219580 527548 219632
rect 527600 219620 527606 219632
rect 528526 219620 528554 219728
rect 548702 219716 548708 219728
rect 548760 219716 548766 219768
rect 548886 219716 548892 219768
rect 548944 219756 548950 219768
rect 595622 219756 595628 219768
rect 548944 219728 595628 219756
rect 548944 219716 548950 219728
rect 595622 219716 595628 219728
rect 595680 219716 595686 219768
rect 606018 219756 606024 219768
rect 595824 219728 606024 219756
rect 527600 219592 528554 219620
rect 527600 219580 527606 219592
rect 540790 219580 540796 219632
rect 540848 219620 540854 219632
rect 595824 219620 595852 219728
rect 606018 219716 606024 219728
rect 606076 219716 606082 219768
rect 620094 219620 620100 219632
rect 540848 219592 595852 219620
rect 595916 219592 620100 219620
rect 540848 219580 540854 219592
rect 137704 219524 146984 219552
rect 137704 219512 137710 219524
rect 147582 219512 147588 219564
rect 147640 219552 147646 219564
rect 211338 219552 211344 219564
rect 147640 219524 211344 219552
rect 147640 219512 147646 219524
rect 211338 219512 211344 219524
rect 211396 219512 211402 219564
rect 214098 219512 214104 219564
rect 214156 219552 214162 219564
rect 218698 219552 218704 219564
rect 214156 219524 218704 219552
rect 214156 219512 214162 219524
rect 218698 219512 218704 219524
rect 218756 219512 218762 219564
rect 224218 219512 224224 219564
rect 224276 219552 224282 219564
rect 229278 219552 229284 219564
rect 224276 219524 229284 219552
rect 224276 219512 224282 219524
rect 229278 219512 229284 219524
rect 229336 219512 229342 219564
rect 432046 219552 432052 219564
rect 431926 219524 432052 219552
rect 405918 219444 405924 219496
rect 405976 219484 405982 219496
rect 412726 219484 412732 219496
rect 405976 219456 412732 219484
rect 405976 219444 405982 219456
rect 412726 219444 412732 219456
rect 412784 219444 412790 219496
rect 421006 219484 421012 219496
rect 418172 219456 421012 219484
rect 70578 219376 70584 219428
rect 70636 219416 70642 219428
rect 117590 219416 117596 219428
rect 70636 219388 117596 219416
rect 70636 219376 70642 219388
rect 117590 219376 117596 219388
rect 117648 219376 117654 219428
rect 117774 219376 117780 219428
rect 117832 219416 117838 219428
rect 118694 219416 118700 219428
rect 117832 219388 118700 219416
rect 117832 219376 117838 219388
rect 118694 219376 118700 219388
rect 118752 219376 118758 219428
rect 131850 219376 131856 219428
rect 131908 219416 131914 219428
rect 132402 219416 132408 219428
rect 131908 219388 132408 219416
rect 131908 219376 131914 219388
rect 132402 219376 132408 219388
rect 132460 219376 132466 219428
rect 132586 219376 132592 219428
rect 132644 219416 132650 219428
rect 168926 219416 168932 219428
rect 132644 219388 168932 219416
rect 132644 219376 132650 219388
rect 168926 219376 168932 219388
rect 168984 219376 168990 219428
rect 169110 219376 169116 219428
rect 169168 219416 169174 219428
rect 169570 219416 169576 219428
rect 169168 219388 169576 219416
rect 169168 219376 169174 219388
rect 169570 219376 169576 219388
rect 169628 219376 169634 219428
rect 169754 219376 169760 219428
rect 169812 219416 169818 219428
rect 172146 219416 172152 219428
rect 169812 219388 172152 219416
rect 169812 219376 169818 219388
rect 172146 219376 172152 219388
rect 172204 219376 172210 219428
rect 172422 219376 172428 219428
rect 172480 219416 172486 219428
rect 173158 219416 173164 219428
rect 172480 219388 173164 219416
rect 172480 219376 172486 219388
rect 173158 219376 173164 219388
rect 173216 219376 173222 219428
rect 178218 219376 178224 219428
rect 178276 219416 178282 219428
rect 178770 219416 178776 219428
rect 178276 219388 178776 219416
rect 178276 219376 178282 219388
rect 178770 219376 178776 219388
rect 178828 219376 178834 219428
rect 181622 219376 181628 219428
rect 181680 219416 181686 219428
rect 182082 219416 182088 219428
rect 181680 219388 182088 219416
rect 181680 219376 181686 219388
rect 182082 219376 182088 219388
rect 182140 219376 182146 219428
rect 182266 219376 182272 219428
rect 182324 219416 182330 219428
rect 184474 219416 184480 219428
rect 182324 219388 184480 219416
rect 182324 219376 182330 219388
rect 184474 219376 184480 219388
rect 184532 219376 184538 219428
rect 185670 219376 185676 219428
rect 185728 219416 185734 219428
rect 186130 219416 186136 219428
rect 185728 219388 186136 219416
rect 185728 219376 185734 219388
rect 186130 219376 186136 219388
rect 186188 219376 186194 219428
rect 186268 219376 186274 219428
rect 186326 219416 186332 219428
rect 215938 219416 215944 219428
rect 186326 219388 215944 219416
rect 186326 219376 186332 219388
rect 215938 219376 215944 219388
rect 215996 219376 216002 219428
rect 219618 219376 219624 219428
rect 219676 219416 219682 219428
rect 261202 219416 261208 219428
rect 219676 219388 261208 219416
rect 219676 219376 219682 219388
rect 261202 219376 261208 219388
rect 261260 219376 261266 219428
rect 262674 219376 262680 219428
rect 262732 219416 262738 219428
rect 263594 219416 263600 219428
rect 262732 219388 263600 219416
rect 262732 219376 262738 219388
rect 263594 219376 263600 219388
rect 263652 219376 263658 219428
rect 272334 219376 272340 219428
rect 272392 219416 272398 219428
rect 301406 219416 301412 219428
rect 272392 219388 301412 219416
rect 272392 219376 272398 219388
rect 301406 219376 301412 219388
rect 301464 219376 301470 219428
rect 308214 219376 308220 219428
rect 308272 219416 308278 219428
rect 309134 219416 309140 219428
rect 308272 219388 309140 219416
rect 308272 219376 308278 219388
rect 309134 219376 309140 219388
rect 309192 219376 309198 219428
rect 314010 219376 314016 219428
rect 314068 219416 314074 219428
rect 330294 219416 330300 219428
rect 314068 219388 330300 219416
rect 314068 219376 314074 219388
rect 330294 219376 330300 219388
rect 330352 219376 330358 219428
rect 333698 219376 333704 219428
rect 333756 219416 333762 219428
rect 347222 219416 347228 219428
rect 333756 219388 347228 219416
rect 333756 219376 333762 219388
rect 347222 219376 347228 219388
rect 347280 219376 347286 219428
rect 349614 219376 349620 219428
rect 349672 219416 349678 219428
rect 350534 219416 350540 219428
rect 349672 219388 350540 219416
rect 349672 219376 349678 219388
rect 350534 219376 350540 219388
rect 350592 219376 350598 219428
rect 352098 219376 352104 219428
rect 352156 219416 352162 219428
rect 355318 219416 355324 219428
rect 352156 219388 355324 219416
rect 352156 219376 352162 219388
rect 355318 219376 355324 219388
rect 355376 219376 355382 219428
rect 362034 219376 362040 219428
rect 362092 219416 362098 219428
rect 367646 219416 367652 219428
rect 362092 219388 367652 219416
rect 362092 219376 362098 219388
rect 367646 219376 367652 219388
rect 367704 219376 367710 219428
rect 380250 219376 380256 219428
rect 380308 219416 380314 219428
rect 384206 219416 384212 219428
rect 380308 219388 384212 219416
rect 380308 219376 380314 219388
rect 384206 219376 384212 219388
rect 384264 219376 384270 219428
rect 399294 219376 399300 219428
rect 399352 219416 399358 219428
rect 400214 219416 400220 219428
rect 399352 219388 400220 219416
rect 399352 219376 399358 219388
rect 400214 219376 400220 219388
rect 400272 219376 400278 219428
rect 415854 219376 415860 219428
rect 415912 219416 415918 219428
rect 416774 219416 416780 219428
rect 415912 219388 416780 219416
rect 415912 219376 415918 219388
rect 416774 219376 416780 219388
rect 416832 219376 416838 219428
rect 417510 219376 417516 219428
rect 417568 219416 417574 219428
rect 418172 219416 418200 219456
rect 421006 219444 421012 219456
rect 421064 219444 421070 219496
rect 431926 219484 431954 219524
rect 432046 219512 432052 219524
rect 432104 219512 432110 219564
rect 501138 219512 501144 219564
rect 501196 219552 501202 219564
rect 501196 219524 509234 219552
rect 501196 219512 501202 219524
rect 429212 219456 431954 219484
rect 509206 219484 509234 219524
rect 582374 219484 582380 219496
rect 509206 219456 582380 219484
rect 417568 219388 418200 219416
rect 417568 219376 417574 219388
rect 428274 219376 428280 219428
rect 428332 219416 428338 219428
rect 429212 219416 429240 219456
rect 582374 219444 582380 219456
rect 582432 219444 582438 219496
rect 595916 219484 595944 219592
rect 620094 219580 620100 219592
rect 620152 219580 620158 219632
rect 607490 219484 607496 219496
rect 582760 219456 595944 219484
rect 596008 219456 607496 219484
rect 428332 219388 429240 219416
rect 428332 219376 428338 219388
rect 562042 219348 562048 219360
rect 560266 219320 562048 219348
rect 93762 219240 93768 219292
rect 93820 219280 93826 219292
rect 94406 219280 94412 219292
rect 93820 219252 94412 219280
rect 93820 219240 93826 219252
rect 94406 219240 94412 219252
rect 94464 219240 94470 219292
rect 117958 219240 117964 219292
rect 118016 219280 118022 219292
rect 159358 219280 159364 219292
rect 118016 219252 159364 219280
rect 118016 219240 118022 219252
rect 159358 219240 159364 219252
rect 159416 219240 159422 219292
rect 162486 219240 162492 219292
rect 162544 219280 162550 219292
rect 171594 219280 171600 219292
rect 162544 219252 171600 219280
rect 162544 219240 162550 219252
rect 171594 219240 171600 219252
rect 171652 219240 171658 219292
rect 180058 219280 180064 219292
rect 171796 219252 180064 219280
rect 64598 219104 64604 219156
rect 64656 219144 64662 219156
rect 66898 219144 66904 219156
rect 64656 219116 66904 219144
rect 64656 219104 64662 219116
rect 66898 219104 66904 219116
rect 66956 219104 66962 219156
rect 83826 219104 83832 219156
rect 83884 219144 83890 219156
rect 157978 219144 157984 219156
rect 83884 219116 157984 219144
rect 83884 219104 83890 219116
rect 157978 219104 157984 219116
rect 158036 219104 158042 219156
rect 165798 219104 165804 219156
rect 165856 219144 165862 219156
rect 171796 219144 171824 219252
rect 180058 219240 180064 219252
rect 180116 219240 180122 219292
rect 181438 219240 181444 219292
rect 181496 219280 181502 219292
rect 189994 219280 190000 219292
rect 181496 219252 190000 219280
rect 181496 219240 181502 219252
rect 189994 219240 190000 219252
rect 190052 219240 190058 219292
rect 190638 219240 190644 219292
rect 190696 219280 190702 219292
rect 194870 219280 194876 219292
rect 190696 219252 194876 219280
rect 190696 219240 190702 219252
rect 194870 219240 194876 219252
rect 194928 219240 194934 219292
rect 195054 219240 195060 219292
rect 195112 219280 195118 219292
rect 224034 219280 224040 219292
rect 195112 219252 224040 219280
rect 195112 219240 195118 219252
rect 224034 219240 224040 219252
rect 224092 219240 224098 219292
rect 237834 219240 237840 219292
rect 237892 219280 237898 219292
rect 239214 219280 239220 219292
rect 237892 219252 239220 219280
rect 237892 219240 237898 219252
rect 239214 219240 239220 219252
rect 239272 219240 239278 219292
rect 239490 219240 239496 219292
rect 239548 219280 239554 219292
rect 272886 219280 272892 219292
rect 239548 219252 272892 219280
rect 239548 219240 239554 219252
rect 272886 219240 272892 219252
rect 272944 219240 272950 219292
rect 285858 219240 285864 219292
rect 285916 219280 285922 219292
rect 313826 219280 313832 219292
rect 285916 219252 313832 219280
rect 285916 219240 285922 219252
rect 313826 219240 313832 219252
rect 313884 219240 313890 219292
rect 419166 219240 419172 219292
rect 419224 219280 419230 219292
rect 422662 219280 422668 219292
rect 419224 219252 422668 219280
rect 419224 219240 419230 219252
rect 422662 219240 422668 219252
rect 422720 219240 422726 219292
rect 536190 219240 536196 219292
rect 536248 219280 536254 219292
rect 536650 219280 536656 219292
rect 536248 219252 536656 219280
rect 536248 219240 536254 219252
rect 536650 219240 536656 219252
rect 536708 219240 536714 219292
rect 548886 219280 548892 219292
rect 543706 219252 548892 219280
rect 165856 219116 171824 219144
rect 165856 219104 165862 219116
rect 171962 219104 171968 219156
rect 172020 219144 172026 219156
rect 175918 219144 175924 219156
rect 172020 219116 175924 219144
rect 172020 219104 172026 219116
rect 175918 219104 175924 219116
rect 175976 219104 175982 219156
rect 207842 219144 207848 219156
rect 176626 219116 207848 219144
rect 62298 218968 62304 219020
rect 62356 219008 62362 219020
rect 72418 219008 72424 219020
rect 62356 218980 72424 219008
rect 62356 218968 62362 218980
rect 72418 218968 72424 218980
rect 72476 218968 72482 219020
rect 77202 218968 77208 219020
rect 77260 219008 77266 219020
rect 150618 219008 150624 219020
rect 77260 218980 150624 219008
rect 77260 218968 77266 218980
rect 150618 218968 150624 218980
rect 150676 218968 150682 219020
rect 152366 218968 152372 219020
rect 152424 219008 152430 219020
rect 153838 219008 153844 219020
rect 152424 218980 153844 219008
rect 152424 218968 152430 218980
rect 153838 218968 153844 218980
rect 153896 218968 153902 219020
rect 154022 218968 154028 219020
rect 154080 219008 154086 219020
rect 160186 219008 160192 219020
rect 154080 218980 160192 219008
rect 154080 218968 154086 218980
rect 160186 218968 160192 218980
rect 160244 218968 160250 219020
rect 161474 218968 161480 219020
rect 161532 219008 161538 219020
rect 166258 219008 166264 219020
rect 161532 218980 166264 219008
rect 161532 218968 161538 218980
rect 166258 218968 166264 218980
rect 166316 218968 166322 219020
rect 169754 218968 169760 219020
rect 169812 219008 169818 219020
rect 176626 219008 176654 219116
rect 207842 219104 207848 219116
rect 207900 219104 207906 219156
rect 208854 219104 208860 219156
rect 208912 219144 208918 219156
rect 209682 219144 209688 219156
rect 208912 219116 209688 219144
rect 208912 219104 208918 219116
rect 209682 219104 209688 219116
rect 209740 219104 209746 219156
rect 211338 219104 211344 219156
rect 211396 219144 211402 219156
rect 217318 219144 217324 219156
rect 211396 219116 217324 219144
rect 211396 219104 211402 219116
rect 217318 219104 217324 219116
rect 217376 219104 217382 219156
rect 218790 219104 218796 219156
rect 218848 219144 218854 219156
rect 219342 219144 219348 219156
rect 218848 219116 219348 219144
rect 218848 219104 218854 219116
rect 219342 219104 219348 219116
rect 219400 219104 219406 219156
rect 224218 219104 224224 219156
rect 224276 219144 224282 219156
rect 253382 219144 253388 219156
rect 224276 219116 253388 219144
rect 224276 219104 224282 219116
rect 253382 219104 253388 219116
rect 253440 219104 253446 219156
rect 261202 219104 261208 219156
rect 261260 219144 261266 219156
rect 264238 219144 264244 219156
rect 261260 219116 264244 219144
rect 261260 219104 261266 219116
rect 264238 219104 264244 219116
rect 264296 219104 264302 219156
rect 264422 219104 264428 219156
rect 264480 219144 264486 219156
rect 266998 219144 267004 219156
rect 264480 219116 267004 219144
rect 264480 219104 264486 219116
rect 266998 219104 267004 219116
rect 267056 219104 267062 219156
rect 272702 219104 272708 219156
rect 272760 219144 272766 219156
rect 272760 219116 287054 219144
rect 272760 219104 272766 219116
rect 169812 218980 176654 219008
rect 169812 218968 169818 218980
rect 179046 218968 179052 219020
rect 179104 219008 179110 219020
rect 196250 219008 196256 219020
rect 179104 218980 196256 219008
rect 179104 218968 179110 218980
rect 196250 218968 196256 218980
rect 196308 218968 196314 219020
rect 200206 218968 200212 219020
rect 200264 219008 200270 219020
rect 204162 219008 204168 219020
rect 200264 218980 204168 219008
rect 200264 218968 200270 218980
rect 204162 218968 204168 218980
rect 204220 218968 204226 219020
rect 204714 218968 204720 219020
rect 204772 219008 204778 219020
rect 246298 219008 246304 219020
rect 204772 218980 246304 219008
rect 204772 218968 204778 218980
rect 246298 218968 246304 218980
rect 246356 218968 246362 219020
rect 252738 218968 252744 219020
rect 252796 219008 252802 219020
rect 282178 219008 282184 219020
rect 252796 218980 282184 219008
rect 252796 218968 252802 218980
rect 282178 218968 282184 218980
rect 282236 218968 282242 219020
rect 287026 219008 287054 219116
rect 295794 219104 295800 219156
rect 295852 219144 295858 219156
rect 296714 219144 296720 219156
rect 295852 219116 296720 219144
rect 295852 219104 295858 219116
rect 296714 219104 296720 219116
rect 296772 219104 296778 219156
rect 320634 219104 320640 219156
rect 320692 219144 320698 219156
rect 342806 219144 342812 219156
rect 320692 219116 342812 219144
rect 320692 219104 320698 219116
rect 342806 219104 342812 219116
rect 342864 219104 342870 219156
rect 343818 219104 343824 219156
rect 343876 219144 343882 219156
rect 353938 219144 353944 219156
rect 343876 219116 353944 219144
rect 343876 219104 343882 219116
rect 353938 219104 353944 219116
rect 353996 219104 354002 219156
rect 363690 219104 363696 219156
rect 363748 219144 363754 219156
rect 370498 219144 370504 219156
rect 363748 219116 370504 219144
rect 363748 219104 363754 219116
rect 370498 219104 370504 219116
rect 370556 219104 370562 219156
rect 542538 219104 542544 219156
rect 542596 219144 542602 219156
rect 542998 219144 543004 219156
rect 542596 219116 543004 219144
rect 542596 219104 542602 219116
rect 542998 219104 543004 219116
rect 543056 219144 543062 219156
rect 543706 219144 543734 219252
rect 548886 219240 548892 219252
rect 548944 219240 548950 219292
rect 557350 219240 557356 219292
rect 557408 219280 557414 219292
rect 560266 219280 560294 219320
rect 562042 219308 562048 219320
rect 562100 219308 562106 219360
rect 572530 219348 572536 219360
rect 563164 219320 572536 219348
rect 557408 219252 560294 219280
rect 557408 219240 557414 219252
rect 561306 219144 561312 219156
rect 543056 219116 543734 219144
rect 547248 219116 561312 219144
rect 543056 219104 543062 219116
rect 297266 219008 297272 219020
rect 287026 218980 297272 219008
rect 297266 218968 297272 218980
rect 297324 218968 297330 219020
rect 307386 218968 307392 219020
rect 307444 219008 307450 219020
rect 307444 218980 329236 219008
rect 307444 218968 307450 218980
rect 59814 218832 59820 218884
rect 59872 218872 59878 218884
rect 139946 218872 139952 218884
rect 59872 218844 139952 218872
rect 59872 218832 59878 218844
rect 139946 218832 139952 218844
rect 140004 218832 140010 218884
rect 142246 218832 142252 218884
rect 142304 218872 142310 218884
rect 146938 218872 146944 218884
rect 142304 218844 146944 218872
rect 142304 218832 142310 218844
rect 146938 218832 146944 218844
rect 146996 218832 147002 218884
rect 150894 218832 150900 218884
rect 150952 218872 150958 218884
rect 154390 218872 154396 218884
rect 150952 218844 154396 218872
rect 150952 218832 150958 218844
rect 154390 218832 154396 218844
rect 154448 218832 154454 218884
rect 159818 218832 159824 218884
rect 159876 218872 159882 218884
rect 203518 218872 203524 218884
rect 159876 218844 203524 218872
rect 159876 218832 159882 218844
rect 203518 218832 203524 218844
rect 203576 218832 203582 218884
rect 206462 218832 206468 218884
rect 206520 218872 206526 218884
rect 253842 218872 253848 218884
rect 206520 218844 253848 218872
rect 206520 218832 206526 218844
rect 253842 218832 253848 218844
rect 253900 218832 253906 218884
rect 259086 218832 259092 218884
rect 259144 218872 259150 218884
rect 259144 218844 287054 218872
rect 259144 218832 259150 218844
rect 58986 218696 58992 218748
rect 59044 218736 59050 218748
rect 145098 218736 145104 218748
rect 59044 218708 145104 218736
rect 59044 218696 59050 218708
rect 145098 218696 145104 218708
rect 145156 218696 145162 218748
rect 146754 218696 146760 218748
rect 146812 218736 146818 218748
rect 180518 218736 180524 218748
rect 146812 218708 180524 218736
rect 146812 218696 146818 218708
rect 180518 218696 180524 218708
rect 180576 218696 180582 218748
rect 180702 218696 180708 218748
rect 180760 218736 180766 218748
rect 185946 218736 185952 218748
rect 180760 218708 185952 218736
rect 180760 218696 180766 218708
rect 185946 218696 185952 218708
rect 186004 218696 186010 218748
rect 186498 218696 186504 218748
rect 186556 218736 186562 218748
rect 195054 218736 195060 218748
rect 186556 218708 195060 218736
rect 186556 218696 186562 218708
rect 195054 218696 195060 218708
rect 195112 218696 195118 218748
rect 195606 218696 195612 218748
rect 195664 218736 195670 218748
rect 197998 218736 198004 218748
rect 195664 218708 198004 218736
rect 195664 218696 195670 218708
rect 197998 218696 198004 218708
rect 198056 218696 198062 218748
rect 198274 218696 198280 218748
rect 198332 218736 198338 218748
rect 243446 218736 243452 218748
rect 198332 218708 243452 218736
rect 198332 218696 198338 218708
rect 243446 218696 243452 218708
rect 243504 218696 243510 218748
rect 253198 218696 253204 218748
rect 253256 218736 253262 218748
rect 286318 218736 286324 218748
rect 253256 218708 286324 218736
rect 253256 218696 253262 218708
rect 286318 218696 286324 218708
rect 286376 218696 286382 218748
rect 287026 218736 287054 218844
rect 291654 218832 291660 218884
rect 291712 218872 291718 218884
rect 291712 218844 296714 218872
rect 291712 218832 291718 218844
rect 291838 218736 291844 218748
rect 287026 218708 291844 218736
rect 291838 218696 291844 218708
rect 291896 218696 291902 218748
rect 296686 218736 296714 218844
rect 300486 218832 300492 218884
rect 300544 218872 300550 218884
rect 327718 218872 327724 218884
rect 300544 218844 327724 218872
rect 300544 218832 300550 218844
rect 327718 218832 327724 218844
rect 327776 218832 327782 218884
rect 329208 218872 329236 218980
rect 330294 218968 330300 219020
rect 330352 219008 330358 219020
rect 335998 219008 336004 219020
rect 330352 218980 336004 219008
rect 330352 218968 330358 218980
rect 335998 218968 336004 218980
rect 336056 218968 336062 219020
rect 337194 218968 337200 219020
rect 337252 219008 337258 219020
rect 345658 219008 345664 219020
rect 337252 218980 345664 219008
rect 337252 218968 337258 218980
rect 345658 218968 345664 218980
rect 345716 218968 345722 219020
rect 347222 218968 347228 219020
rect 347280 219008 347286 219020
rect 363506 219008 363512 219020
rect 347280 218980 363512 219008
rect 347280 218968 347286 218980
rect 363506 218968 363512 218980
rect 363564 218968 363570 219020
rect 368658 218968 368664 219020
rect 368716 219008 368722 219020
rect 377398 219008 377404 219020
rect 368716 218980 377404 219008
rect 368716 218968 368722 218980
rect 377398 218968 377404 218980
rect 377456 218968 377462 219020
rect 377600 218980 383654 219008
rect 332686 218872 332692 218884
rect 329208 218844 332692 218872
rect 332686 218832 332692 218844
rect 332744 218832 332750 218884
rect 340506 218832 340512 218884
rect 340564 218872 340570 218884
rect 358078 218872 358084 218884
rect 340564 218844 358084 218872
rect 340564 218832 340570 218844
rect 358078 218832 358084 218844
rect 358136 218832 358142 218884
rect 376938 218832 376944 218884
rect 376996 218872 377002 218884
rect 377600 218872 377628 218980
rect 376996 218844 377628 218872
rect 376996 218832 377002 218844
rect 382734 218832 382740 218884
rect 382792 218872 382798 218884
rect 383470 218872 383476 218884
rect 382792 218844 383476 218872
rect 382792 218832 382798 218844
rect 383470 218832 383476 218844
rect 383528 218832 383534 218884
rect 383626 218872 383654 218980
rect 386874 218968 386880 219020
rect 386932 219008 386938 219020
rect 398098 219008 398104 219020
rect 386932 218980 398104 219008
rect 386932 218968 386938 218980
rect 398098 218968 398104 218980
rect 398156 218968 398162 219020
rect 388530 218872 388536 218884
rect 383626 218844 388536 218872
rect 388530 218832 388536 218844
rect 388588 218832 388594 218884
rect 402606 218832 402612 218884
rect 402664 218872 402670 218884
rect 409046 218872 409052 218884
rect 402664 218844 409052 218872
rect 402664 218832 402670 218844
rect 409046 218832 409052 218844
rect 409104 218832 409110 218884
rect 411714 218832 411720 218884
rect 411772 218872 411778 218884
rect 412542 218872 412548 218884
rect 411772 218844 412548 218872
rect 411772 218832 411778 218844
rect 412542 218832 412548 218844
rect 412600 218832 412606 218884
rect 512730 218832 512736 218884
rect 512788 218872 512794 218884
rect 547248 218872 547276 219116
rect 561306 219104 561312 219116
rect 561364 219104 561370 219156
rect 563164 219144 563192 219320
rect 572530 219308 572536 219320
rect 572588 219308 572594 219360
rect 576826 219320 582374 219348
rect 572668 219240 572674 219292
rect 572726 219280 572732 219292
rect 576826 219280 576854 219320
rect 572726 219252 576854 219280
rect 582346 219280 582374 219320
rect 582760 219280 582788 219456
rect 595622 219308 595628 219360
rect 595680 219348 595686 219360
rect 596008 219348 596036 219456
rect 607490 219444 607496 219456
rect 607548 219444 607554 219496
rect 595680 219320 596036 219348
rect 595680 219308 595686 219320
rect 582346 219252 582788 219280
rect 572726 219240 572732 219252
rect 586974 219172 586980 219224
rect 587032 219212 587038 219224
rect 597554 219212 597560 219224
rect 587032 219184 597560 219212
rect 587032 219172 587038 219184
rect 597554 219172 597560 219184
rect 597612 219172 597618 219224
rect 574554 219144 574560 219156
rect 562336 219116 563192 219144
rect 563348 219116 574560 219144
rect 548702 218968 548708 219020
rect 548760 219008 548766 219020
rect 562336 219008 562364 219116
rect 563348 219020 563376 219116
rect 574554 219104 574560 219116
rect 574612 219104 574618 219156
rect 563146 219008 563152 219020
rect 548760 218980 562364 219008
rect 562428 218980 563152 219008
rect 548760 218968 548766 218980
rect 512788 218844 528554 218872
rect 512788 218832 512794 218844
rect 321646 218736 321652 218748
rect 296686 218708 321652 218736
rect 321646 218696 321652 218708
rect 321704 218696 321710 218748
rect 327258 218696 327264 218748
rect 327316 218736 327322 218748
rect 351086 218736 351092 218748
rect 327316 218708 351092 218736
rect 327316 218696 327322 218708
rect 351086 218696 351092 218708
rect 351144 218696 351150 218748
rect 353754 218696 353760 218748
rect 353812 218736 353818 218748
rect 369118 218736 369124 218748
rect 353812 218708 369124 218736
rect 353812 218696 353818 218708
rect 369118 218696 369124 218708
rect 369176 218696 369182 218748
rect 370314 218696 370320 218748
rect 370372 218736 370378 218748
rect 380066 218736 380072 218748
rect 370372 218708 380072 218736
rect 370372 218696 370378 218708
rect 380066 218696 380072 218708
rect 380124 218696 380130 218748
rect 383562 218696 383568 218748
rect 383620 218736 383626 218748
rect 396258 218736 396264 218748
rect 383620 218708 396264 218736
rect 383620 218696 383626 218708
rect 396258 218696 396264 218708
rect 396316 218696 396322 218748
rect 412542 218696 412548 218748
rect 412600 218736 412606 218748
rect 417142 218736 417148 218748
rect 412600 218708 417148 218736
rect 412600 218696 412606 218708
rect 417142 218696 417148 218708
rect 417200 218696 417206 218748
rect 482738 218696 482744 218748
rect 482796 218736 482802 218748
rect 485314 218736 485320 218748
rect 482796 218708 485320 218736
rect 482796 218696 482802 218708
rect 485314 218696 485320 218708
rect 485372 218696 485378 218748
rect 500402 218696 500408 218748
rect 500460 218736 500466 218748
rect 508038 218736 508044 218748
rect 500460 218708 508044 218736
rect 500460 218696 500466 218708
rect 508038 218696 508044 218708
rect 508096 218696 508102 218748
rect 517698 218696 517704 218748
rect 517756 218736 517762 218748
rect 518158 218736 518164 218748
rect 517756 218708 518164 218736
rect 517756 218696 517762 218708
rect 518158 218696 518164 218708
rect 518216 218736 518222 218748
rect 519998 218736 520004 218748
rect 518216 218708 520004 218736
rect 518216 218696 518222 218708
rect 519998 218696 520004 218708
rect 520056 218696 520062 218748
rect 528526 218736 528554 218844
rect 534046 218844 547276 218872
rect 534046 218736 534074 218844
rect 547414 218832 547420 218884
rect 547472 218872 547478 218884
rect 562428 218872 562456 218980
rect 563146 218968 563152 218980
rect 563204 218968 563210 219020
rect 563330 218968 563336 219020
rect 563388 218968 563394 219020
rect 563514 218968 563520 219020
rect 563572 219008 563578 219020
rect 572346 219008 572352 219020
rect 563572 218980 572352 219008
rect 563572 218968 563578 218980
rect 572346 218968 572352 218980
rect 572404 218968 572410 219020
rect 572668 218968 572674 219020
rect 572726 219008 572732 219020
rect 603074 219008 603080 219020
rect 572726 218980 603080 219008
rect 572726 218968 572732 218980
rect 603074 218968 603080 218980
rect 603132 218968 603138 219020
rect 547472 218844 562456 218872
rect 547472 218832 547478 218844
rect 562594 218832 562600 218884
rect 562652 218872 562658 218884
rect 562962 218872 562968 218884
rect 562652 218844 562968 218872
rect 562652 218832 562658 218844
rect 562962 218832 562968 218844
rect 563020 218832 563026 218884
rect 563330 218832 563336 218884
rect 563388 218872 563394 218884
rect 614114 218872 614120 218884
rect 563388 218844 614120 218872
rect 563388 218832 563394 218844
rect 614114 218832 614120 218844
rect 614172 218832 614178 218884
rect 528526 218708 534074 218736
rect 537478 218696 537484 218748
rect 537536 218736 537542 218748
rect 598106 218736 598112 218748
rect 537536 218708 562824 218736
rect 537536 218696 537542 218708
rect 562796 218668 562824 218708
rect 563164 218708 598112 218736
rect 562796 218640 562916 218668
rect 107010 218560 107016 218612
rect 107068 218600 107074 218612
rect 117958 218600 117964 218612
rect 107068 218572 117964 218600
rect 107068 218560 107074 218572
rect 117958 218560 117964 218572
rect 118016 218560 118022 218612
rect 118142 218560 118148 218612
rect 118200 218600 118206 218612
rect 162118 218600 162124 218612
rect 118200 218572 162124 218600
rect 118200 218560 118206 218572
rect 162118 218560 162124 218572
rect 162176 218560 162182 218612
rect 166626 218560 166632 218612
rect 166684 218600 166690 218612
rect 169754 218600 169760 218612
rect 166684 218572 169760 218600
rect 166684 218560 166690 218572
rect 169754 218560 169760 218572
rect 169812 218560 169818 218612
rect 169938 218560 169944 218612
rect 169996 218600 170002 218612
rect 170950 218600 170956 218612
rect 169996 218572 170956 218600
rect 169996 218560 170002 218572
rect 170950 218560 170956 218572
rect 171008 218560 171014 218612
rect 171594 218560 171600 218612
rect 171652 218600 171658 218612
rect 181070 218600 181076 218612
rect 171652 218572 181076 218600
rect 171652 218560 171658 218572
rect 181070 218560 181076 218572
rect 181128 218560 181134 218612
rect 182358 218560 182364 218612
rect 182416 218600 182422 218612
rect 189718 218600 189724 218612
rect 182416 218572 189724 218600
rect 182416 218560 182422 218572
rect 189718 218560 189724 218572
rect 189776 218560 189782 218612
rect 192846 218560 192852 218612
rect 192904 218600 192910 218612
rect 192904 218572 195468 218600
rect 192904 218560 192910 218572
rect 142246 218464 142252 218476
rect 103486 218436 142252 218464
rect 100386 218288 100392 218340
rect 100444 218328 100450 218340
rect 103486 218328 103514 218436
rect 142246 218424 142252 218436
rect 142304 218424 142310 218476
rect 142430 218424 142436 218476
rect 142488 218464 142494 218476
rect 150434 218464 150440 218476
rect 142488 218436 150440 218464
rect 142488 218424 142494 218436
rect 150434 218424 150440 218436
rect 150492 218424 150498 218476
rect 150618 218424 150624 218476
rect 150676 218464 150682 218476
rect 152366 218464 152372 218476
rect 150676 218436 152372 218464
rect 150676 218424 150682 218436
rect 152366 218424 152372 218436
rect 152424 218424 152430 218476
rect 152550 218424 152556 218476
rect 152608 218464 152614 218476
rect 153102 218464 153108 218476
rect 152608 218436 153108 218464
rect 152608 218424 152614 218436
rect 153102 218424 153108 218436
rect 153160 218424 153166 218476
rect 153378 218424 153384 218476
rect 153436 218464 153442 218476
rect 154022 218464 154028 218476
rect 153436 218436 154028 218464
rect 153436 218424 153442 218436
rect 154022 218424 154028 218436
rect 154080 218424 154086 218476
rect 155034 218424 155040 218476
rect 155092 218464 155098 218476
rect 155678 218464 155684 218476
rect 155092 218436 155684 218464
rect 155092 218424 155098 218436
rect 155678 218424 155684 218436
rect 155736 218424 155742 218476
rect 156690 218424 156696 218476
rect 156748 218464 156754 218476
rect 157242 218464 157248 218476
rect 156748 218436 157248 218464
rect 156748 218424 156754 218436
rect 157242 218424 157248 218436
rect 157300 218424 157306 218476
rect 159174 218424 159180 218476
rect 159232 218464 159238 218476
rect 160002 218464 160008 218476
rect 159232 218436 160008 218464
rect 159232 218424 159238 218436
rect 160002 218424 160008 218436
rect 160060 218424 160066 218476
rect 160186 218424 160192 218476
rect 160244 218464 160250 218476
rect 186958 218464 186964 218476
rect 160244 218436 186964 218464
rect 160244 218424 160250 218436
rect 186958 218424 186964 218436
rect 187016 218424 187022 218476
rect 189810 218424 189816 218476
rect 189868 218464 189874 218476
rect 195238 218464 195244 218476
rect 189868 218436 195244 218464
rect 189868 218424 189874 218436
rect 195238 218424 195244 218436
rect 195296 218424 195302 218476
rect 195440 218464 195468 218572
rect 198090 218560 198096 218612
rect 198148 218600 198154 218612
rect 200206 218600 200212 218612
rect 198148 218572 200212 218600
rect 198148 218560 198154 218572
rect 200206 218560 200212 218572
rect 200264 218560 200270 218612
rect 200390 218560 200396 218612
rect 200448 218600 200454 218612
rect 210326 218600 210332 218612
rect 200448 218572 210332 218600
rect 200448 218560 200454 218572
rect 210326 218560 210332 218572
rect 210384 218560 210390 218612
rect 212994 218560 213000 218612
rect 213052 218600 213058 218612
rect 224218 218600 224224 218612
rect 213052 218572 224224 218600
rect 213052 218560 213058 218572
rect 224218 218560 224224 218572
rect 224276 218560 224282 218612
rect 225966 218560 225972 218612
rect 226024 218600 226030 218612
rect 264422 218600 264428 218612
rect 226024 218572 264428 218600
rect 226024 218560 226030 218572
rect 264422 218560 264428 218572
rect 264480 218560 264486 218612
rect 265986 218560 265992 218612
rect 266044 218600 266050 218612
rect 272702 218600 272708 218612
rect 266044 218572 272708 218600
rect 266044 218560 266050 218572
rect 272702 218560 272708 218572
rect 272760 218560 272766 218612
rect 272886 218560 272892 218612
rect 272944 218600 272950 218612
rect 279418 218600 279424 218612
rect 272944 218572 279424 218600
rect 272944 218560 272950 218572
rect 279418 218560 279424 218572
rect 279476 218560 279482 218612
rect 305546 218600 305552 218612
rect 280080 218572 305552 218600
rect 198274 218464 198280 218476
rect 195440 218436 198280 218464
rect 198274 218424 198280 218436
rect 198332 218424 198338 218476
rect 199746 218424 199752 218476
rect 199804 218464 199810 218476
rect 204714 218464 204720 218476
rect 199804 218436 204720 218464
rect 199804 218424 199810 218436
rect 204714 218424 204720 218436
rect 204772 218424 204778 218476
rect 204916 218436 214604 218464
rect 100444 218300 103514 218328
rect 100444 218288 100450 218300
rect 113634 218288 113640 218340
rect 113692 218328 113698 218340
rect 118142 218328 118148 218340
rect 113692 218300 118148 218328
rect 113692 218288 113698 218300
rect 118142 218288 118148 218300
rect 118200 218288 118206 218340
rect 120258 218288 120264 218340
rect 120316 218328 120322 218340
rect 161474 218328 161480 218340
rect 120316 218300 161480 218328
rect 120316 218288 120322 218300
rect 161474 218288 161480 218300
rect 161532 218288 161538 218340
rect 161658 218288 161664 218340
rect 161716 218328 161722 218340
rect 162762 218328 162768 218340
rect 161716 218300 162768 218328
rect 161716 218288 161722 218300
rect 162762 218288 162768 218300
rect 162820 218288 162826 218340
rect 163314 218288 163320 218340
rect 163372 218328 163378 218340
rect 163958 218328 163964 218340
rect 163372 218300 163964 218328
rect 163372 218288 163378 218300
rect 163958 218288 163964 218300
rect 164016 218288 164022 218340
rect 164970 218288 164976 218340
rect 165028 218328 165034 218340
rect 165522 218328 165528 218340
rect 165028 218300 165528 218328
rect 165028 218288 165034 218300
rect 165522 218288 165528 218300
rect 165580 218288 165586 218340
rect 170766 218288 170772 218340
rect 170824 218328 170830 218340
rect 175274 218328 175280 218340
rect 170824 218300 175280 218328
rect 170824 218288 170830 218300
rect 175274 218288 175280 218300
rect 175332 218288 175338 218340
rect 175734 218288 175740 218340
rect 175792 218328 175798 218340
rect 181438 218328 181444 218340
rect 175792 218300 181444 218328
rect 175792 218288 175798 218300
rect 181438 218288 181444 218300
rect 181496 218288 181502 218340
rect 192018 218288 192024 218340
rect 192076 218328 192082 218340
rect 193582 218328 193588 218340
rect 192076 218300 193588 218328
rect 192076 218288 192082 218300
rect 193582 218288 193588 218300
rect 193640 218288 193646 218340
rect 196434 218288 196440 218340
rect 196492 218328 196498 218340
rect 204916 218328 204944 218436
rect 196492 218300 204944 218328
rect 196492 218288 196498 218300
rect 209682 218288 209688 218340
rect 209740 218328 209746 218340
rect 213178 218328 213184 218340
rect 209740 218300 213184 218328
rect 209740 218288 209746 218300
rect 213178 218288 213184 218300
rect 213236 218288 213242 218340
rect 214576 218328 214604 218436
rect 216306 218424 216312 218476
rect 216364 218464 216370 218476
rect 216364 218436 216904 218464
rect 216364 218424 216370 218436
rect 216876 218328 216904 218436
rect 217318 218424 217324 218476
rect 217376 218464 217382 218476
rect 219802 218464 219808 218476
rect 217376 218436 219808 218464
rect 217376 218424 217382 218436
rect 219802 218424 219808 218436
rect 219860 218424 219866 218476
rect 224034 218424 224040 218476
rect 224092 218464 224098 218476
rect 231026 218464 231032 218476
rect 224092 218436 231032 218464
rect 224092 218424 224098 218436
rect 231026 218424 231032 218436
rect 231084 218424 231090 218476
rect 238018 218464 238024 218476
rect 232700 218436 238024 218464
rect 232700 218328 232728 218436
rect 238018 218424 238024 218436
rect 238076 218424 238082 218476
rect 271138 218464 271144 218476
rect 238726 218436 271144 218464
rect 214576 218300 216628 218328
rect 216876 218300 232728 218328
rect 55674 218152 55680 218204
rect 55732 218192 55738 218204
rect 56502 218192 56508 218204
rect 55732 218164 56508 218192
rect 55732 218152 55738 218164
rect 56502 218152 56508 218164
rect 56560 218152 56566 218204
rect 57422 218152 57428 218204
rect 57480 218192 57486 218204
rect 61378 218192 61384 218204
rect 57480 218164 61384 218192
rect 57480 218152 57486 218164
rect 61378 218152 61384 218164
rect 61436 218152 61442 218204
rect 66438 218152 66444 218204
rect 66496 218192 66502 218204
rect 67542 218192 67548 218204
rect 66496 218164 67548 218192
rect 66496 218152 66502 218164
rect 67542 218152 67548 218164
rect 67600 218152 67606 218204
rect 68094 218152 68100 218204
rect 68152 218192 68158 218204
rect 69566 218192 69572 218204
rect 68152 218164 69572 218192
rect 68152 218152 68158 218164
rect 69566 218152 69572 218164
rect 69624 218152 69630 218204
rect 75546 218152 75552 218204
rect 75604 218192 75610 218204
rect 76558 218192 76564 218204
rect 75604 218164 76564 218192
rect 75604 218152 75610 218164
rect 76558 218152 76564 218164
rect 76616 218152 76622 218204
rect 97074 218152 97080 218204
rect 97132 218192 97138 218204
rect 97132 218164 100892 218192
rect 97132 218152 97138 218164
rect 56502 218016 56508 218068
rect 56560 218056 56566 218068
rect 57238 218056 57244 218068
rect 56560 218028 57244 218056
rect 56560 218016 56566 218028
rect 57238 218016 57244 218028
rect 57296 218016 57302 218068
rect 58158 218016 58164 218068
rect 58216 218056 58222 218068
rect 59354 218056 59360 218068
rect 58216 218028 59360 218056
rect 58216 218016 58222 218028
rect 59354 218016 59360 218028
rect 59412 218016 59418 218068
rect 61470 218016 61476 218068
rect 61528 218056 61534 218068
rect 62758 218056 62764 218068
rect 61528 218028 62764 218056
rect 61528 218016 61534 218028
rect 62758 218016 62764 218028
rect 62816 218016 62822 218068
rect 63954 218016 63960 218068
rect 64012 218056 64018 218068
rect 64782 218056 64788 218068
rect 64012 218028 64788 218056
rect 64012 218016 64018 218028
rect 64782 218016 64788 218028
rect 64840 218016 64846 218068
rect 65610 218016 65616 218068
rect 65668 218056 65674 218068
rect 66162 218056 66168 218068
rect 65668 218028 66168 218056
rect 65668 218016 65674 218028
rect 66162 218016 66168 218028
rect 66220 218016 66226 218068
rect 67266 218016 67272 218068
rect 67324 218056 67330 218068
rect 68278 218056 68284 218068
rect 67324 218028 68284 218056
rect 67324 218016 67330 218028
rect 68278 218016 68284 218028
rect 68336 218016 68342 218068
rect 72234 218016 72240 218068
rect 72292 218056 72298 218068
rect 73706 218056 73712 218068
rect 72292 218028 73712 218056
rect 72292 218016 72298 218028
rect 73706 218016 73712 218028
rect 73764 218016 73770 218068
rect 74718 218016 74724 218068
rect 74776 218056 74782 218068
rect 75822 218056 75828 218068
rect 74776 218028 75828 218056
rect 74776 218016 74782 218028
rect 75822 218016 75828 218028
rect 75880 218016 75886 218068
rect 78030 218016 78036 218068
rect 78088 218056 78094 218068
rect 78582 218056 78588 218068
rect 78088 218028 78588 218056
rect 78088 218016 78094 218028
rect 78582 218016 78588 218028
rect 78640 218016 78646 218068
rect 78858 218016 78864 218068
rect 78916 218056 78922 218068
rect 79962 218056 79968 218068
rect 78916 218028 79968 218056
rect 78916 218016 78922 218028
rect 79962 218016 79968 218028
rect 80020 218016 80026 218068
rect 82170 218016 82176 218068
rect 82228 218056 82234 218068
rect 83458 218056 83464 218068
rect 82228 218028 83464 218056
rect 82228 218016 82234 218028
rect 83458 218016 83464 218028
rect 83516 218016 83522 218068
rect 84654 218016 84660 218068
rect 84712 218056 84718 218068
rect 85298 218056 85304 218068
rect 84712 218028 85304 218056
rect 84712 218016 84718 218028
rect 85298 218016 85304 218028
rect 85356 218016 85362 218068
rect 87138 218016 87144 218068
rect 87196 218056 87202 218068
rect 88242 218056 88248 218068
rect 87196 218028 88248 218056
rect 87196 218016 87202 218028
rect 88242 218016 88248 218028
rect 88300 218016 88306 218068
rect 88794 218016 88800 218068
rect 88852 218056 88858 218068
rect 89438 218056 89444 218068
rect 88852 218028 89444 218056
rect 88852 218016 88858 218028
rect 89438 218016 89444 218028
rect 89496 218016 89502 218068
rect 92934 218016 92940 218068
rect 92992 218056 92998 218068
rect 93578 218056 93584 218068
rect 92992 218028 93584 218056
rect 92992 218016 92998 218028
rect 93578 218016 93584 218028
rect 93636 218016 93642 218068
rect 95418 218016 95424 218068
rect 95476 218056 95482 218068
rect 96246 218056 96252 218068
rect 95476 218028 96252 218056
rect 95476 218016 95482 218028
rect 96246 218016 96252 218028
rect 96304 218016 96310 218068
rect 98730 218016 98736 218068
rect 98788 218056 98794 218068
rect 99282 218056 99288 218068
rect 98788 218028 99288 218056
rect 98788 218016 98794 218028
rect 99282 218016 99288 218028
rect 99340 218016 99346 218068
rect 99558 218016 99564 218068
rect 99616 218056 99622 218068
rect 100662 218056 100668 218068
rect 99616 218028 100668 218056
rect 99616 218016 99622 218028
rect 100662 218016 100668 218028
rect 100720 218016 100726 218068
rect 100864 217988 100892 218164
rect 117590 218152 117596 218204
rect 117648 218192 117654 218204
rect 123386 218192 123392 218204
rect 117648 218164 123392 218192
rect 117648 218152 117654 218164
rect 123386 218152 123392 218164
rect 123444 218152 123450 218204
rect 123570 218152 123576 218204
rect 123628 218192 123634 218204
rect 123628 218164 136772 218192
rect 123628 218152 123634 218164
rect 102870 218084 102876 218136
rect 102928 218124 102934 218136
rect 103422 218124 103428 218136
rect 102928 218096 103428 218124
rect 102928 218084 102934 218096
rect 103422 218084 103428 218096
rect 103480 218084 103486 218136
rect 103698 218016 103704 218068
rect 103756 218056 103762 218068
rect 104802 218056 104808 218068
rect 103756 218028 104808 218056
rect 103756 218016 103762 218028
rect 104802 218016 104808 218028
rect 104860 218016 104866 218068
rect 105354 218016 105360 218068
rect 105412 218056 105418 218068
rect 105998 218056 106004 218068
rect 105412 218028 106004 218056
rect 105412 218016 105418 218028
rect 105998 218016 106004 218028
rect 106056 218016 106062 218068
rect 109494 218016 109500 218068
rect 109552 218056 109558 218068
rect 110414 218056 110420 218068
rect 109552 218028 110420 218056
rect 109552 218016 109558 218028
rect 110414 218016 110420 218028
rect 110472 218016 110478 218068
rect 111978 218016 111984 218068
rect 112036 218056 112042 218068
rect 112806 218056 112812 218068
rect 112036 218028 112812 218056
rect 112036 218016 112042 218028
rect 112806 218016 112812 218028
rect 112864 218016 112870 218068
rect 116118 218016 116124 218068
rect 116176 218056 116182 218068
rect 117222 218056 117228 218068
rect 116176 218028 117228 218056
rect 116176 218016 116182 218028
rect 117222 218016 117228 218028
rect 117280 218016 117286 218068
rect 119430 218016 119436 218068
rect 119488 218056 119494 218068
rect 119982 218056 119988 218068
rect 119488 218028 119988 218056
rect 119488 218016 119494 218028
rect 119982 218016 119988 218028
rect 120040 218016 120046 218068
rect 121914 218016 121920 218068
rect 121972 218056 121978 218068
rect 122558 218056 122564 218068
rect 121972 218028 122564 218056
rect 121972 218016 121978 218028
rect 122558 218016 122564 218028
rect 122616 218016 122622 218068
rect 126054 218016 126060 218068
rect 126112 218056 126118 218068
rect 126698 218056 126704 218068
rect 126112 218028 126704 218056
rect 126112 218016 126118 218028
rect 126698 218016 126704 218028
rect 126756 218016 126762 218068
rect 127710 218016 127716 218068
rect 127768 218056 127774 218068
rect 128262 218056 128268 218068
rect 127768 218028 128268 218056
rect 127768 218016 127774 218028
rect 128262 218016 128268 218028
rect 128320 218016 128326 218068
rect 128538 218016 128544 218068
rect 128596 218056 128602 218068
rect 129366 218056 129372 218068
rect 128596 218028 129372 218056
rect 128596 218016 128602 218028
rect 129366 218016 129372 218028
rect 129424 218016 129430 218068
rect 130194 218016 130200 218068
rect 130252 218056 130258 218068
rect 132494 218056 132500 218068
rect 130252 218028 132500 218056
rect 130252 218016 130258 218028
rect 132494 218016 132500 218028
rect 132552 218016 132558 218068
rect 132678 218016 132684 218068
rect 132736 218056 132742 218068
rect 133506 218056 133512 218068
rect 132736 218028 133512 218056
rect 132736 218016 132742 218028
rect 133506 218016 133512 218028
rect 133564 218016 133570 218068
rect 135990 218016 135996 218068
rect 136048 218056 136054 218068
rect 136542 218056 136548 218068
rect 136048 218028 136548 218056
rect 136048 218016 136054 218028
rect 136542 218016 136548 218028
rect 136600 218016 136606 218068
rect 136744 218056 136772 218164
rect 136910 218152 136916 218204
rect 136968 218192 136974 218204
rect 136968 218164 150296 218192
rect 136968 218152 136974 218164
rect 137278 218056 137284 218068
rect 136744 218028 137284 218056
rect 137278 218016 137284 218028
rect 137336 218016 137342 218068
rect 140130 218016 140136 218068
rect 140188 218056 140194 218068
rect 142430 218056 142436 218068
rect 140188 218028 142436 218056
rect 140188 218016 140194 218028
rect 142430 218016 142436 218028
rect 142488 218016 142494 218068
rect 142614 218016 142620 218068
rect 142672 218056 142678 218068
rect 143258 218056 143264 218068
rect 142672 218028 143264 218056
rect 142672 218016 142678 218028
rect 143258 218016 143264 218028
rect 143316 218016 143322 218068
rect 144270 218016 144276 218068
rect 144328 218056 144334 218068
rect 144822 218056 144828 218068
rect 144328 218028 144828 218056
rect 144328 218016 144334 218028
rect 144822 218016 144828 218028
rect 144880 218016 144886 218068
rect 145098 218016 145104 218068
rect 145156 218056 145162 218068
rect 145926 218056 145932 218068
rect 145156 218028 145932 218056
rect 145156 218016 145162 218028
rect 145926 218016 145932 218028
rect 145984 218016 145990 218068
rect 148410 218016 148416 218068
rect 148468 218056 148474 218068
rect 148870 218056 148876 218068
rect 148468 218028 148876 218056
rect 148468 218016 148474 218028
rect 148870 218016 148876 218028
rect 148928 218016 148934 218068
rect 149238 218016 149244 218068
rect 149296 218056 149302 218068
rect 150066 218056 150072 218068
rect 149296 218028 150072 218056
rect 149296 218016 149302 218028
rect 150066 218016 150072 218028
rect 150124 218016 150130 218068
rect 150268 218056 150296 218164
rect 150434 218152 150440 218204
rect 150492 218192 150498 218204
rect 171410 218192 171416 218204
rect 150492 218164 171416 218192
rect 150492 218152 150498 218164
rect 171410 218152 171416 218164
rect 171468 218152 171474 218204
rect 179322 218192 179328 218204
rect 171796 218164 179328 218192
rect 171796 218124 171824 218164
rect 179322 218152 179328 218164
rect 179380 218152 179386 218204
rect 179874 218152 179880 218204
rect 179932 218192 179938 218204
rect 200390 218192 200396 218204
rect 179932 218164 200396 218192
rect 179932 218152 179938 218164
rect 200390 218152 200396 218164
rect 200448 218152 200454 218204
rect 200574 218152 200580 218204
rect 200632 218192 200638 218204
rect 201494 218192 201500 218204
rect 200632 218164 201500 218192
rect 200632 218152 200638 218164
rect 201494 218152 201500 218164
rect 201552 218152 201558 218204
rect 204714 218152 204720 218204
rect 204772 218192 204778 218204
rect 207658 218192 207664 218204
rect 204772 218164 207664 218192
rect 204772 218152 204778 218164
rect 207658 218152 207664 218164
rect 207716 218152 207722 218204
rect 207842 218152 207848 218204
rect 207900 218192 207906 218204
rect 211798 218192 211804 218204
rect 207900 218164 211804 218192
rect 207900 218152 207906 218164
rect 211798 218152 211804 218164
rect 211856 218152 211862 218204
rect 171704 218096 171824 218124
rect 216600 218124 216628 218300
rect 232866 218288 232872 218340
rect 232924 218328 232930 218340
rect 238726 218328 238754 218436
rect 271138 218424 271144 218436
rect 271196 218424 271202 218476
rect 279234 218424 279240 218476
rect 279292 218464 279298 218476
rect 280080 218464 280108 218572
rect 305546 218560 305552 218572
rect 305604 218560 305610 218612
rect 398466 218560 398472 218612
rect 398524 218600 398530 218612
rect 407758 218600 407764 218612
rect 398524 218572 407764 218600
rect 398524 218560 398530 218572
rect 407758 218560 407764 218572
rect 407816 218560 407822 218612
rect 429930 218560 429936 218612
rect 429988 218600 429994 218612
rect 432690 218600 432696 218612
rect 429988 218572 432696 218600
rect 429988 218560 429994 218572
rect 432690 218560 432696 218572
rect 432748 218560 432754 218612
rect 469858 218560 469864 218612
rect 469916 218600 469922 218612
rect 471238 218600 471244 218612
rect 469916 218572 471244 218600
rect 469916 218560 469922 218572
rect 471238 218560 471244 218572
rect 471296 218560 471302 218612
rect 475562 218560 475568 218612
rect 475620 218600 475626 218612
rect 482830 218600 482836 218612
rect 475620 218572 482836 218600
rect 475620 218560 475626 218572
rect 482830 218560 482836 218572
rect 482888 218560 482894 218612
rect 507670 218560 507676 218612
rect 507728 218600 507734 218612
rect 548702 218600 548708 218612
rect 507728 218572 548708 218600
rect 507728 218560 507734 218572
rect 548702 218560 548708 218572
rect 548760 218560 548766 218612
rect 548886 218560 548892 218612
rect 548944 218600 548950 218612
rect 562594 218600 562600 218612
rect 548944 218572 562600 218600
rect 548944 218560 548950 218572
rect 562594 218560 562600 218572
rect 562652 218560 562658 218612
rect 562888 218600 562916 218640
rect 563164 218600 563192 218708
rect 598106 218696 598112 218708
rect 598164 218696 598170 218748
rect 562888 218572 563192 218600
rect 564158 218560 564164 218612
rect 564216 218600 564222 218612
rect 572530 218600 572536 218612
rect 564216 218572 572536 218600
rect 564216 218560 564222 218572
rect 572530 218560 572536 218572
rect 572588 218560 572594 218612
rect 572668 218560 572674 218612
rect 572726 218600 572732 218612
rect 610710 218600 610716 218612
rect 572726 218572 610716 218600
rect 572726 218560 572732 218572
rect 610710 218560 610716 218572
rect 610768 218560 610774 218612
rect 279292 218436 280108 218464
rect 279292 218424 279298 218436
rect 282178 218424 282184 218476
rect 282236 218464 282242 218476
rect 287882 218464 287888 218476
rect 282236 218436 287888 218464
rect 282236 218424 282242 218436
rect 287882 218424 287888 218436
rect 287940 218424 287946 218476
rect 294138 218424 294144 218476
rect 294196 218464 294202 218476
rect 316678 218464 316684 218476
rect 294196 218436 316684 218464
rect 294196 218424 294202 218436
rect 316678 218424 316684 218436
rect 316736 218424 316742 218476
rect 502794 218424 502800 218476
rect 502852 218464 502858 218476
rect 503162 218464 503168 218476
rect 502852 218436 503168 218464
rect 502852 218424 502858 218436
rect 503162 218424 503168 218436
rect 503220 218464 503226 218476
rect 507854 218464 507860 218476
rect 503220 218436 507860 218464
rect 503220 218424 503226 218436
rect 507854 218424 507860 218436
rect 507912 218424 507918 218476
rect 508038 218424 508044 218476
rect 508096 218464 508102 218476
rect 604454 218464 604460 218476
rect 508096 218436 604460 218464
rect 508096 218424 508102 218436
rect 604454 218424 604460 218436
rect 604512 218424 604518 218476
rect 458174 218356 458180 218408
rect 458232 218396 458238 218408
rect 458232 218368 460934 218396
rect 458232 218356 458238 218368
rect 232924 218300 238754 218328
rect 232924 218288 232930 218300
rect 246114 218288 246120 218340
rect 246172 218328 246178 218340
rect 253198 218328 253204 218340
rect 246172 218300 253204 218328
rect 246172 218288 246178 218300
rect 253198 218288 253204 218300
rect 253256 218288 253262 218340
rect 253382 218288 253388 218340
rect 253440 218328 253446 218340
rect 258074 218328 258080 218340
rect 253440 218300 258080 218328
rect 253440 218288 253446 218300
rect 258074 218288 258080 218300
rect 258132 218288 258138 218340
rect 426618 218288 426624 218340
rect 426676 218328 426682 218340
rect 429562 218328 429568 218340
rect 426676 218300 429568 218328
rect 426676 218288 426682 218300
rect 429562 218288 429568 218300
rect 429620 218288 429626 218340
rect 434898 218288 434904 218340
rect 434956 218328 434962 218340
rect 436646 218328 436652 218340
rect 434956 218300 436652 218328
rect 434956 218288 434962 218300
rect 436646 218288 436652 218300
rect 436704 218288 436710 218340
rect 450722 218288 450728 218340
rect 450780 218328 450786 218340
rect 453850 218328 453856 218340
rect 450780 218300 453856 218328
rect 450780 218288 450786 218300
rect 453850 218288 453856 218300
rect 453908 218288 453914 218340
rect 460906 218328 460934 218368
rect 461302 218328 461308 218340
rect 460906 218300 461308 218328
rect 461302 218288 461308 218300
rect 461360 218288 461366 218340
rect 497458 218288 497464 218340
rect 497516 218328 497522 218340
rect 595990 218328 595996 218340
rect 497516 218300 595996 218328
rect 497516 218288 497522 218300
rect 595990 218288 595996 218300
rect 596048 218288 596054 218340
rect 217962 218152 217968 218204
rect 218020 218192 218026 218204
rect 222746 218192 222752 218204
rect 218020 218164 222752 218192
rect 218020 218152 218026 218164
rect 222746 218152 222752 218164
rect 222804 218152 222810 218204
rect 222930 218152 222936 218204
rect 222988 218192 222994 218204
rect 225598 218192 225604 218204
rect 222988 218164 225604 218192
rect 222988 218152 222994 218164
rect 225598 218152 225604 218164
rect 225656 218152 225662 218204
rect 241974 218152 241980 218204
rect 242032 218192 242038 218204
rect 242894 218192 242900 218204
rect 242032 218164 242900 218192
rect 242032 218152 242038 218164
rect 242894 218152 242900 218164
rect 242952 218152 242958 218204
rect 249426 218152 249432 218204
rect 249484 218192 249490 218204
rect 251726 218192 251732 218204
rect 249484 218164 251732 218192
rect 249484 218152 249490 218164
rect 251726 218152 251732 218164
rect 251784 218152 251790 218204
rect 328914 218152 328920 218204
rect 328972 218192 328978 218204
rect 330478 218192 330484 218204
rect 328972 218164 330484 218192
rect 328972 218152 328978 218164
rect 330478 218152 330484 218164
rect 330536 218152 330542 218204
rect 365346 218152 365352 218204
rect 365404 218192 365410 218204
rect 371786 218192 371792 218204
rect 365404 218164 371792 218192
rect 365404 218152 365410 218164
rect 371786 218152 371792 218164
rect 371844 218152 371850 218204
rect 374454 218152 374460 218204
rect 374512 218192 374518 218204
rect 376018 218192 376024 218204
rect 374512 218164 376024 218192
rect 374512 218152 374518 218164
rect 376018 218152 376024 218164
rect 376076 218152 376082 218204
rect 381906 218152 381912 218204
rect 381964 218192 381970 218204
rect 382918 218192 382924 218204
rect 381964 218164 382924 218192
rect 381964 218152 381970 218164
rect 382918 218152 382924 218164
rect 382976 218152 382982 218204
rect 401778 218152 401784 218204
rect 401836 218192 401842 218204
rect 402790 218192 402796 218204
rect 401836 218164 402796 218192
rect 401836 218152 401842 218164
rect 402790 218152 402796 218164
rect 402848 218152 402854 218204
rect 407574 218152 407580 218204
rect 407632 218192 407638 218204
rect 411898 218192 411904 218204
rect 407632 218164 411904 218192
rect 407632 218152 407638 218164
rect 411898 218152 411904 218164
rect 411956 218152 411962 218204
rect 422478 218152 422484 218204
rect 422536 218192 422542 218204
rect 425422 218192 425428 218204
rect 422536 218164 425428 218192
rect 422536 218152 422542 218164
rect 425422 218152 425428 218164
rect 425480 218152 425486 218204
rect 425790 218152 425796 218204
rect 425848 218192 425854 218204
rect 428458 218192 428464 218204
rect 425848 218164 428464 218192
rect 425848 218152 425854 218164
rect 428458 218152 428464 218164
rect 428516 218152 428522 218204
rect 433242 218152 433248 218204
rect 433300 218192 433306 218204
rect 435266 218192 435272 218204
rect 433300 218164 435272 218192
rect 433300 218152 433306 218164
rect 435266 218152 435272 218164
rect 435324 218152 435330 218204
rect 461946 218152 461952 218204
rect 462004 218192 462010 218204
rect 466270 218192 466276 218204
rect 462004 218164 466276 218192
rect 462004 218152 462010 218164
rect 466270 218152 466276 218164
rect 466328 218152 466334 218204
rect 491938 218152 491944 218204
rect 491996 218192 492002 218204
rect 502242 218192 502248 218204
rect 491996 218164 502248 218192
rect 491996 218152 492002 218164
rect 502242 218152 502248 218164
rect 502300 218152 502306 218204
rect 507118 218152 507124 218204
rect 507176 218192 507182 218204
rect 507670 218192 507676 218204
rect 507176 218164 507676 218192
rect 507176 218152 507182 218164
rect 507670 218152 507676 218164
rect 507728 218152 507734 218204
rect 507854 218152 507860 218204
rect 507912 218192 507918 218204
rect 563054 218192 563060 218204
rect 507912 218164 563060 218192
rect 507912 218152 507918 218164
rect 563054 218152 563060 218164
rect 563112 218152 563118 218204
rect 572668 218152 572674 218204
rect 572726 218192 572732 218204
rect 572726 218164 614068 218192
rect 572726 218152 572732 218164
rect 216600 218096 216720 218124
rect 171704 218056 171732 218096
rect 150268 218028 171732 218056
rect 173250 218016 173256 218068
rect 173308 218056 173314 218068
rect 186222 218056 186228 218068
rect 173308 218028 186228 218056
rect 173308 218016 173314 218028
rect 186222 218016 186228 218028
rect 186280 218016 186286 218068
rect 188154 218016 188160 218068
rect 188212 218056 188218 218068
rect 188890 218056 188896 218068
rect 188212 218028 188896 218056
rect 188212 218016 188218 218028
rect 188890 218016 188896 218028
rect 188948 218016 188954 218068
rect 192018 218056 192024 218068
rect 189092 218028 192024 218056
rect 100864 217960 103514 217988
rect 103486 217920 103514 217960
rect 174262 217920 174268 217932
rect 103486 217892 174268 217920
rect 174262 217880 174268 217892
rect 174320 217880 174326 217932
rect 188890 217880 188896 217932
rect 188948 217920 188954 217932
rect 189092 217920 189120 218028
rect 192018 218016 192024 218028
rect 192076 218016 192082 218068
rect 192294 218016 192300 218068
rect 192352 218056 192358 218068
rect 193030 218056 193036 218068
rect 192352 218028 193036 218056
rect 192352 218016 192358 218028
rect 193030 218016 193036 218028
rect 193088 218016 193094 218068
rect 193950 218016 193956 218068
rect 194008 218056 194014 218068
rect 194502 218056 194508 218068
rect 194008 218028 194508 218056
rect 194008 218016 194014 218028
rect 194502 218016 194508 218028
rect 194560 218016 194566 218068
rect 194778 218016 194784 218068
rect 194836 218056 194842 218068
rect 195882 218056 195888 218068
rect 194836 218028 195888 218056
rect 194836 218016 194842 218028
rect 195882 218016 195888 218028
rect 195940 218016 195946 218068
rect 198918 218016 198924 218068
rect 198976 218056 198982 218068
rect 200022 218056 200028 218068
rect 198976 218028 200028 218056
rect 198976 218016 198982 218028
rect 200022 218016 200028 218028
rect 200080 218016 200086 218068
rect 203058 218016 203064 218068
rect 203116 218056 203122 218068
rect 206278 218056 206284 218068
rect 203116 218028 206284 218056
rect 203116 218016 203122 218028
rect 206278 218016 206284 218028
rect 206336 218016 206342 218068
rect 207198 218016 207204 218068
rect 207256 218056 207262 218068
rect 208118 218056 208124 218068
rect 207256 218028 208124 218056
rect 207256 218016 207262 218028
rect 208118 218016 208124 218028
rect 208176 218016 208182 218068
rect 214650 218016 214656 218068
rect 214708 218056 214714 218068
rect 215202 218056 215208 218068
rect 214708 218028 215208 218056
rect 214708 218016 214714 218028
rect 215202 218016 215208 218028
rect 215260 218016 215266 218068
rect 215478 218016 215484 218068
rect 215536 218056 215542 218068
rect 216122 218056 216128 218068
rect 215536 218028 216128 218056
rect 215536 218016 215542 218028
rect 216122 218016 216128 218028
rect 216180 218016 216186 218068
rect 216692 218056 216720 218096
rect 563210 218096 572576 218124
rect 220078 218056 220084 218068
rect 216692 218028 220084 218056
rect 220078 218016 220084 218028
rect 220136 218016 220142 218068
rect 221274 218016 221280 218068
rect 221332 218056 221338 218068
rect 221826 218056 221832 218068
rect 221332 218028 221832 218056
rect 221332 218016 221338 218028
rect 221826 218016 221832 218028
rect 221884 218016 221890 218068
rect 223758 218016 223764 218068
rect 223816 218056 223822 218068
rect 224586 218056 224592 218068
rect 223816 218028 224592 218056
rect 223816 218016 223822 218028
rect 224586 218016 224592 218028
rect 224644 218016 224650 218068
rect 225414 218016 225420 218068
rect 225472 218056 225478 218068
rect 226150 218056 226156 218068
rect 225472 218028 226156 218056
rect 225472 218016 225478 218028
rect 226150 218016 226156 218028
rect 226208 218016 226214 218068
rect 229554 218016 229560 218068
rect 229612 218056 229618 218068
rect 230474 218056 230480 218068
rect 229612 218028 230480 218056
rect 229612 218016 229618 218028
rect 230474 218016 230480 218028
rect 230532 218016 230538 218068
rect 231210 218016 231216 218068
rect 231268 218056 231274 218068
rect 231670 218056 231676 218068
rect 231268 218028 231676 218056
rect 231268 218016 231274 218028
rect 231670 218016 231676 218028
rect 231728 218016 231734 218068
rect 232038 218016 232044 218068
rect 232096 218056 232102 218068
rect 233142 218056 233148 218068
rect 232096 218028 233148 218056
rect 232096 218016 232102 218028
rect 233142 218016 233148 218028
rect 233200 218016 233206 218068
rect 235350 218016 235356 218068
rect 235408 218056 235414 218068
rect 235810 218056 235816 218068
rect 235408 218028 235816 218056
rect 235408 218016 235414 218028
rect 235810 218016 235816 218028
rect 235868 218016 235874 218068
rect 236178 218016 236184 218068
rect 236236 218056 236242 218068
rect 237282 218056 237288 218068
rect 236236 218028 237288 218056
rect 236236 218016 236242 218028
rect 237282 218016 237288 218028
rect 237340 218016 237346 218068
rect 240318 218016 240324 218068
rect 240376 218056 240382 218068
rect 241330 218056 241336 218068
rect 240376 218028 241336 218056
rect 240376 218016 240382 218028
rect 241330 218016 241336 218028
rect 241388 218016 241394 218068
rect 243630 218016 243636 218068
rect 243688 218056 243694 218068
rect 244090 218056 244096 218068
rect 243688 218028 244096 218056
rect 243688 218016 243694 218028
rect 244090 218016 244096 218028
rect 244148 218016 244154 218068
rect 247770 218016 247776 218068
rect 247828 218056 247834 218068
rect 248230 218056 248236 218068
rect 247828 218028 248236 218056
rect 247828 218016 247834 218028
rect 248230 218016 248236 218028
rect 248288 218016 248294 218068
rect 248598 218016 248604 218068
rect 248656 218056 248662 218068
rect 249610 218056 249616 218068
rect 248656 218028 249616 218056
rect 248656 218016 248662 218028
rect 249610 218016 249616 218028
rect 249668 218016 249674 218068
rect 250254 218016 250260 218068
rect 250312 218056 250318 218068
rect 250898 218056 250904 218068
rect 250312 218028 250904 218056
rect 250312 218016 250318 218028
rect 250898 218016 250904 218028
rect 250956 218016 250962 218068
rect 251910 218016 251916 218068
rect 251968 218056 251974 218068
rect 252462 218056 252468 218068
rect 251968 218028 252468 218056
rect 251968 218016 251974 218028
rect 252462 218016 252468 218028
rect 252520 218016 252526 218068
rect 254394 218016 254400 218068
rect 254452 218056 254458 218068
rect 255038 218056 255044 218068
rect 254452 218028 255044 218056
rect 254452 218016 254458 218028
rect 255038 218016 255044 218028
rect 255096 218016 255102 218068
rect 256050 218016 256056 218068
rect 256108 218056 256114 218068
rect 256510 218056 256516 218068
rect 256108 218028 256516 218056
rect 256108 218016 256114 218028
rect 256510 218016 256516 218028
rect 256568 218016 256574 218068
rect 256878 218016 256884 218068
rect 256936 218056 256942 218068
rect 257522 218056 257528 218068
rect 256936 218028 257528 218056
rect 256936 218016 256942 218028
rect 257522 218016 257528 218028
rect 257580 218016 257586 218068
rect 258534 218016 258540 218068
rect 258592 218056 258598 218068
rect 259270 218056 259276 218068
rect 258592 218028 259276 218056
rect 258592 218016 258598 218028
rect 259270 218016 259276 218028
rect 259328 218016 259334 218068
rect 264330 218016 264336 218068
rect 264388 218056 264394 218068
rect 264790 218056 264796 218068
rect 264388 218028 264796 218056
rect 264388 218016 264394 218028
rect 264790 218016 264796 218028
rect 264848 218016 264854 218068
rect 265158 218016 265164 218068
rect 265216 218056 265222 218068
rect 266170 218056 266176 218068
rect 265216 218028 266176 218056
rect 265216 218016 265222 218028
rect 266170 218016 266176 218028
rect 266228 218016 266234 218068
rect 268470 218016 268476 218068
rect 268528 218056 268534 218068
rect 268930 218056 268936 218068
rect 268528 218028 268936 218056
rect 268528 218016 268534 218028
rect 268930 218016 268936 218028
rect 268988 218016 268994 218068
rect 269298 218016 269304 218068
rect 269356 218056 269362 218068
rect 270218 218056 270224 218068
rect 269356 218028 270224 218056
rect 269356 218016 269362 218028
rect 270218 218016 270224 218028
rect 270276 218016 270282 218068
rect 270954 218016 270960 218068
rect 271012 218056 271018 218068
rect 272518 218056 272524 218068
rect 271012 218028 272524 218056
rect 271012 218016 271018 218028
rect 272518 218016 272524 218028
rect 272576 218016 272582 218068
rect 276750 218016 276756 218068
rect 276808 218056 276814 218068
rect 277210 218056 277216 218068
rect 276808 218028 277216 218056
rect 276808 218016 276814 218028
rect 277210 218016 277216 218028
rect 277268 218016 277274 218068
rect 277578 218016 277584 218068
rect 277636 218056 277642 218068
rect 278590 218056 278596 218068
rect 277636 218028 278596 218056
rect 277636 218016 277642 218028
rect 278590 218016 278596 218028
rect 278648 218016 278654 218068
rect 280890 218016 280896 218068
rect 280948 218056 280954 218068
rect 281442 218056 281448 218068
rect 280948 218028 281448 218056
rect 280948 218016 280954 218028
rect 281442 218016 281448 218028
rect 281500 218016 281506 218068
rect 281718 218016 281724 218068
rect 281776 218056 281782 218068
rect 282454 218056 282460 218068
rect 281776 218028 282460 218056
rect 281776 218016 281782 218028
rect 282454 218016 282460 218028
rect 282512 218016 282518 218068
rect 285030 218016 285036 218068
rect 285088 218056 285094 218068
rect 285490 218056 285496 218068
rect 285088 218028 285496 218056
rect 285088 218016 285094 218028
rect 285490 218016 285496 218028
rect 285548 218016 285554 218068
rect 287514 218016 287520 218068
rect 287572 218056 287578 218068
rect 288710 218056 288716 218068
rect 287572 218028 288716 218056
rect 287572 218016 287578 218028
rect 288710 218016 288716 218028
rect 288768 218016 288774 218068
rect 289170 218016 289176 218068
rect 289228 218056 289234 218068
rect 289722 218056 289728 218068
rect 289228 218028 289728 218056
rect 289228 218016 289234 218028
rect 289722 218016 289728 218028
rect 289780 218016 289786 218068
rect 289998 218016 290004 218068
rect 290056 218056 290062 218068
rect 291102 218056 291108 218068
rect 290056 218028 291108 218056
rect 290056 218016 290062 218028
rect 291102 218016 291108 218028
rect 291160 218016 291166 218068
rect 293310 218016 293316 218068
rect 293368 218056 293374 218068
rect 293770 218056 293776 218068
rect 293368 218028 293776 218056
rect 293368 218016 293374 218028
rect 293770 218016 293776 218028
rect 293828 218016 293834 218068
rect 297450 218016 297456 218068
rect 297508 218056 297514 218068
rect 297910 218056 297916 218068
rect 297508 218028 297916 218056
rect 297508 218016 297514 218028
rect 297910 218016 297916 218028
rect 297968 218016 297974 218068
rect 298278 218016 298284 218068
rect 298336 218056 298342 218068
rect 299106 218056 299112 218068
rect 298336 218028 299112 218056
rect 298336 218016 298342 218028
rect 299106 218016 299112 218028
rect 299164 218016 299170 218068
rect 299934 218016 299940 218068
rect 299992 218056 299998 218068
rect 300670 218056 300676 218068
rect 299992 218028 300676 218056
rect 299992 218016 299998 218028
rect 300670 218016 300676 218028
rect 300728 218016 300734 218068
rect 301590 218016 301596 218068
rect 301648 218056 301654 218068
rect 302142 218056 302148 218068
rect 301648 218028 302148 218056
rect 301648 218016 301654 218028
rect 302142 218016 302148 218028
rect 302200 218016 302206 218068
rect 304074 218016 304080 218068
rect 304132 218056 304138 218068
rect 304718 218056 304724 218068
rect 304132 218028 304724 218056
rect 304132 218016 304138 218028
rect 304718 218016 304724 218028
rect 304776 218016 304782 218068
rect 305730 218016 305736 218068
rect 305788 218056 305794 218068
rect 306190 218056 306196 218068
rect 305788 218028 306196 218056
rect 305788 218016 305794 218028
rect 306190 218016 306196 218028
rect 306248 218016 306254 218068
rect 306558 218016 306564 218068
rect 306616 218056 306622 218068
rect 307662 218056 307668 218068
rect 306616 218028 307668 218056
rect 306616 218016 306622 218028
rect 307662 218016 307668 218028
rect 307720 218016 307726 218068
rect 309870 218016 309876 218068
rect 309928 218056 309934 218068
rect 310422 218056 310428 218068
rect 309928 218028 310428 218056
rect 309928 218016 309934 218028
rect 310422 218016 310428 218028
rect 310480 218016 310486 218068
rect 312354 218016 312360 218068
rect 312412 218056 312418 218068
rect 312906 218056 312912 218068
rect 312412 218028 312912 218056
rect 312412 218016 312418 218028
rect 312906 218016 312912 218028
rect 312964 218016 312970 218068
rect 317322 218016 317328 218068
rect 317380 218056 317386 218068
rect 317966 218056 317972 218068
rect 317380 218028 317972 218056
rect 317380 218016 317386 218028
rect 317966 218016 317972 218028
rect 318024 218016 318030 218068
rect 318978 218016 318984 218068
rect 319036 218056 319042 218068
rect 319622 218056 319628 218068
rect 319036 218028 319628 218056
rect 319036 218016 319042 218028
rect 319622 218016 319628 218028
rect 319680 218016 319686 218068
rect 322290 218016 322296 218068
rect 322348 218056 322354 218068
rect 322842 218056 322848 218068
rect 322348 218028 322848 218056
rect 322348 218016 322354 218028
rect 322842 218016 322848 218028
rect 322900 218016 322906 218068
rect 323118 218016 323124 218068
rect 323176 218056 323182 218068
rect 324130 218056 324136 218068
rect 323176 218028 324136 218056
rect 323176 218016 323182 218028
rect 324130 218016 324136 218028
rect 324188 218016 324194 218068
rect 324774 218016 324780 218068
rect 324832 218056 324838 218068
rect 325418 218056 325424 218068
rect 324832 218028 325424 218056
rect 324832 218016 324838 218028
rect 325418 218016 325424 218028
rect 325476 218016 325482 218068
rect 326430 218016 326436 218068
rect 326488 218056 326494 218068
rect 326890 218056 326896 218068
rect 326488 218028 326896 218056
rect 326488 218016 326494 218028
rect 326890 218016 326896 218028
rect 326948 218016 326954 218068
rect 330570 218016 330576 218068
rect 330628 218056 330634 218068
rect 331030 218056 331036 218068
rect 330628 218028 331036 218056
rect 330628 218016 330634 218028
rect 331030 218016 331036 218028
rect 331088 218016 331094 218068
rect 333054 218016 333060 218068
rect 333112 218056 333118 218068
rect 333882 218056 333888 218068
rect 333112 218028 333888 218056
rect 333112 218016 333118 218028
rect 333882 218016 333888 218028
rect 333940 218016 333946 218068
rect 334710 218016 334716 218068
rect 334768 218056 334774 218068
rect 335170 218056 335176 218068
rect 334768 218028 335176 218056
rect 334768 218016 334774 218028
rect 335170 218016 335176 218028
rect 335228 218016 335234 218068
rect 335538 218016 335544 218068
rect 335596 218056 335602 218068
rect 338666 218056 338672 218068
rect 335596 218028 338672 218056
rect 335596 218016 335602 218028
rect 338666 218016 338672 218028
rect 338724 218016 338730 218068
rect 338850 218016 338856 218068
rect 338908 218056 338914 218068
rect 339402 218056 339408 218068
rect 338908 218028 339408 218056
rect 338908 218016 338914 218028
rect 339402 218016 339408 218028
rect 339460 218016 339466 218068
rect 339678 218016 339684 218068
rect 339736 218056 339742 218068
rect 340690 218056 340696 218068
rect 339736 218028 340696 218056
rect 339736 218016 339742 218028
rect 340690 218016 340696 218028
rect 340748 218016 340754 218068
rect 345474 218016 345480 218068
rect 345532 218056 345538 218068
rect 347038 218056 347044 218068
rect 345532 218028 347044 218056
rect 345532 218016 345538 218028
rect 347038 218016 347044 218028
rect 347096 218016 347102 218068
rect 347958 218016 347964 218068
rect 348016 218056 348022 218068
rect 349062 218056 349068 218068
rect 348016 218028 349068 218056
rect 348016 218016 348022 218028
rect 349062 218016 349068 218028
rect 349120 218016 349126 218068
rect 355410 218016 355416 218068
rect 355468 218056 355474 218068
rect 355870 218056 355876 218068
rect 355468 218028 355876 218056
rect 355468 218016 355474 218028
rect 355870 218016 355876 218028
rect 355928 218016 355934 218068
rect 356238 218016 356244 218068
rect 356296 218056 356302 218068
rect 356974 218056 356980 218068
rect 356296 218028 356980 218056
rect 356296 218016 356302 218028
rect 356974 218016 356980 218028
rect 357032 218016 357038 218068
rect 359550 218016 359556 218068
rect 359608 218056 359614 218068
rect 360102 218056 360108 218068
rect 359608 218028 360108 218056
rect 359608 218016 359614 218028
rect 360102 218016 360108 218028
rect 360160 218016 360166 218068
rect 360378 218016 360384 218068
rect 360436 218056 360442 218068
rect 361022 218056 361028 218068
rect 360436 218028 361028 218056
rect 360436 218016 360442 218028
rect 361022 218016 361028 218028
rect 361080 218016 361086 218068
rect 364518 218016 364524 218068
rect 364576 218056 364582 218068
rect 365530 218056 365536 218068
rect 364576 218028 365536 218056
rect 364576 218016 364582 218028
rect 365530 218016 365536 218028
rect 365588 218016 365594 218068
rect 366174 218016 366180 218068
rect 366232 218056 366238 218068
rect 366726 218056 366732 218068
rect 366232 218028 366732 218056
rect 366232 218016 366238 218028
rect 366726 218016 366732 218028
rect 366784 218016 366790 218068
rect 367830 218016 367836 218068
rect 367888 218056 367894 218068
rect 368382 218056 368388 218068
rect 367888 218028 368388 218056
rect 367888 218016 367894 218028
rect 368382 218016 368388 218028
rect 368440 218016 368446 218068
rect 371970 218016 371976 218068
rect 372028 218056 372034 218068
rect 372522 218056 372528 218068
rect 372028 218028 372528 218056
rect 372028 218016 372034 218028
rect 372522 218016 372528 218028
rect 372580 218016 372586 218068
rect 372798 218016 372804 218068
rect 372856 218056 372862 218068
rect 373442 218056 373448 218068
rect 372856 218028 373448 218056
rect 372856 218016 372862 218028
rect 373442 218016 373448 218028
rect 373500 218016 373506 218068
rect 376110 218016 376116 218068
rect 376168 218056 376174 218068
rect 376662 218056 376668 218068
rect 376168 218028 376668 218056
rect 376168 218016 376174 218028
rect 376662 218016 376668 218028
rect 376720 218016 376726 218068
rect 378594 218016 378600 218068
rect 378652 218056 378658 218068
rect 379238 218056 379244 218068
rect 378652 218028 379244 218056
rect 378652 218016 378658 218028
rect 379238 218016 379244 218028
rect 379296 218016 379302 218068
rect 381078 218016 381084 218068
rect 381136 218056 381142 218068
rect 382090 218056 382096 218068
rect 381136 218028 382096 218056
rect 381136 218016 381142 218028
rect 382090 218016 382096 218028
rect 382148 218016 382154 218068
rect 389358 218016 389364 218068
rect 389416 218056 389422 218068
rect 390002 218056 390008 218068
rect 389416 218028 390008 218056
rect 389416 218016 389422 218028
rect 390002 218016 390008 218028
rect 390060 218016 390066 218068
rect 392670 218016 392676 218068
rect 392728 218056 392734 218068
rect 393130 218056 393136 218068
rect 392728 218028 393136 218056
rect 392728 218016 392734 218028
rect 393130 218016 393136 218028
rect 393188 218016 393194 218068
rect 393498 218016 393504 218068
rect 393556 218056 393562 218068
rect 394510 218056 394516 218068
rect 393556 218028 394516 218056
rect 393556 218016 393562 218028
rect 394510 218016 394516 218028
rect 394568 218016 394574 218068
rect 395154 218016 395160 218068
rect 395212 218056 395218 218068
rect 395798 218056 395804 218068
rect 395212 218028 395804 218056
rect 395212 218016 395218 218028
rect 395798 218016 395804 218028
rect 395856 218016 395862 218068
rect 397638 218016 397644 218068
rect 397696 218056 397702 218068
rect 400766 218056 400772 218068
rect 397696 218028 400772 218056
rect 397696 218016 397702 218028
rect 400766 218016 400772 218028
rect 400824 218016 400830 218068
rect 400950 218016 400956 218068
rect 401008 218056 401014 218068
rect 402238 218056 402244 218068
rect 401008 218028 402244 218056
rect 401008 218016 401014 218028
rect 402238 218016 402244 218028
rect 402296 218016 402302 218068
rect 403434 218016 403440 218068
rect 403492 218056 403498 218068
rect 403986 218056 403992 218068
rect 403492 218028 403992 218056
rect 403492 218016 403498 218028
rect 403986 218016 403992 218028
rect 404044 218016 404050 218068
rect 405090 218016 405096 218068
rect 405148 218056 405154 218068
rect 405550 218056 405556 218068
rect 405148 218028 405556 218056
rect 405148 218016 405154 218028
rect 405550 218016 405556 218028
rect 405608 218016 405614 218068
rect 409230 218016 409236 218068
rect 409288 218056 409294 218068
rect 409782 218056 409788 218068
rect 409288 218028 409788 218056
rect 409288 218016 409294 218028
rect 409782 218016 409788 218028
rect 409840 218016 409846 218068
rect 410058 218016 410064 218068
rect 410116 218056 410122 218068
rect 410702 218056 410708 218068
rect 410116 218028 410708 218056
rect 410116 218016 410122 218028
rect 410702 218016 410708 218028
rect 410760 218016 410766 218068
rect 413370 218016 413376 218068
rect 413428 218056 413434 218068
rect 413830 218056 413836 218068
rect 413428 218028 413836 218056
rect 413428 218016 413434 218028
rect 413830 218016 413836 218028
rect 413888 218016 413894 218068
rect 419994 218016 420000 218068
rect 420052 218056 420058 218068
rect 420914 218056 420920 218068
rect 420052 218028 420920 218056
rect 420052 218016 420058 218028
rect 420914 218016 420920 218028
rect 420972 218016 420978 218068
rect 424134 218016 424140 218068
rect 424192 218056 424198 218068
rect 426986 218056 426992 218068
rect 424192 218028 426992 218056
rect 424192 218016 424198 218028
rect 426986 218016 426992 218028
rect 427044 218016 427050 218068
rect 427446 218016 427452 218068
rect 427504 218056 427510 218068
rect 427906 218056 427912 218068
rect 427504 218028 427912 218056
rect 427504 218016 427510 218028
rect 427906 218016 427912 218028
rect 427964 218016 427970 218068
rect 429102 218016 429108 218068
rect 429160 218056 429166 218068
rect 430574 218056 430580 218068
rect 429160 218028 430580 218056
rect 429160 218016 429166 218028
rect 430574 218016 430580 218028
rect 430632 218016 430638 218068
rect 432414 218016 432420 218068
rect 432472 218056 432478 218068
rect 433702 218056 433708 218068
rect 432472 218028 433708 218056
rect 432472 218016 432478 218028
rect 433702 218016 433708 218028
rect 433760 218016 433766 218068
rect 435726 218016 435732 218068
rect 435784 218056 435790 218068
rect 436278 218056 436284 218068
rect 435784 218028 436284 218056
rect 435784 218016 435790 218028
rect 436278 218016 436284 218028
rect 436336 218016 436342 218068
rect 436554 218016 436560 218068
rect 436612 218056 436618 218068
rect 437474 218056 437480 218068
rect 436612 218028 437480 218056
rect 436612 218016 436618 218028
rect 437474 218016 437480 218028
rect 437532 218016 437538 218068
rect 438210 218016 438216 218068
rect 438268 218056 438274 218068
rect 438854 218056 438860 218068
rect 438268 218028 438860 218056
rect 438268 218016 438274 218028
rect 438854 218016 438860 218028
rect 438912 218016 438918 218068
rect 439866 218016 439872 218068
rect 439924 218056 439930 218068
rect 440326 218056 440332 218068
rect 439924 218028 440332 218056
rect 439924 218016 439930 218028
rect 440326 218016 440332 218028
rect 440384 218016 440390 218068
rect 453298 218016 453304 218068
rect 453356 218056 453362 218068
rect 455414 218056 455420 218068
rect 453356 218028 455420 218056
rect 453356 218016 453362 218028
rect 455414 218016 455420 218028
rect 455472 218016 455478 218068
rect 455598 218016 455604 218068
rect 455656 218056 455662 218068
rect 457162 218056 457168 218068
rect 455656 218028 457168 218056
rect 455656 218016 455662 218028
rect 457162 218016 457168 218028
rect 457220 218016 457226 218068
rect 463142 218016 463148 218068
rect 463200 218056 463206 218068
rect 464614 218056 464620 218068
rect 463200 218028 464620 218056
rect 463200 218016 463206 218028
rect 464614 218016 464620 218028
rect 464672 218016 464678 218068
rect 467282 218016 467288 218068
rect 467340 218056 467346 218068
rect 467926 218056 467932 218068
rect 467340 218028 467932 218056
rect 467340 218016 467346 218028
rect 467926 218016 467932 218028
rect 467984 218016 467990 218068
rect 471422 218016 471428 218068
rect 471480 218056 471486 218068
rect 472894 218056 472900 218068
rect 471480 218028 472900 218056
rect 471480 218016 471486 218028
rect 472894 218016 472900 218028
rect 472952 218016 472958 218068
rect 490374 218016 490380 218068
rect 490432 218056 490438 218068
rect 490432 218028 496860 218056
rect 490432 218016 490438 218028
rect 188948 217892 189120 217920
rect 496832 217920 496860 218028
rect 496998 218016 497004 218068
rect 497056 218056 497062 218068
rect 497458 218056 497464 218068
rect 497056 218028 497464 218056
rect 497056 218016 497062 218028
rect 497458 218016 497464 218028
rect 497516 218016 497522 218068
rect 563210 218056 563238 218096
rect 497660 218028 563238 218056
rect 572548 218056 572576 218096
rect 572548 218028 605834 218056
rect 497660 217920 497688 218028
rect 563330 217948 563336 218000
rect 563388 217988 563394 218000
rect 572346 217988 572352 218000
rect 563388 217960 572352 217988
rect 563388 217948 563394 217960
rect 572346 217948 572352 217960
rect 572404 217948 572410 218000
rect 605806 217988 605834 218028
rect 612274 217988 612280 218000
rect 605806 217960 612280 217988
rect 612274 217948 612280 217960
rect 612332 217948 612338 218000
rect 614040 217988 614068 218164
rect 644934 218016 644940 218068
rect 644992 218056 644998 218068
rect 653582 218056 653588 218068
rect 644992 218028 653588 218056
rect 644992 218016 644998 218028
rect 653582 218016 653588 218028
rect 653640 218016 653646 218068
rect 614482 217988 614488 218000
rect 614040 217960 614488 217988
rect 614482 217948 614488 217960
rect 614540 217948 614546 218000
rect 496832 217892 497688 217920
rect 188948 217880 188954 217892
rect 523034 217812 523040 217864
rect 523092 217852 523098 217864
rect 524230 217852 524236 217864
rect 523092 217824 524236 217852
rect 523092 217812 523098 217824
rect 524230 217812 524236 217824
rect 524288 217812 524294 217864
rect 603994 217852 604000 217864
rect 534046 217824 604000 217852
rect 533430 217676 533436 217728
rect 533488 217716 533494 217728
rect 534046 217716 534074 217824
rect 603994 217812 604000 217824
rect 604052 217812 604058 217864
rect 603442 217716 603448 217728
rect 533488 217688 534074 217716
rect 538048 217688 603448 217716
rect 533488 217676 533494 217688
rect 116946 217540 116952 217592
rect 117004 217580 117010 217592
rect 189166 217580 189172 217592
rect 117004 217552 189172 217580
rect 117004 217540 117010 217552
rect 189166 217540 189172 217552
rect 189224 217540 189230 217592
rect 530946 217540 530952 217592
rect 531004 217580 531010 217592
rect 538048 217580 538076 217688
rect 603442 217676 603448 217688
rect 603500 217676 603506 217728
rect 604454 217676 604460 217728
rect 604512 217716 604518 217728
rect 614298 217716 614304 217728
rect 604512 217688 614304 217716
rect 604512 217676 604518 217688
rect 614298 217676 614304 217688
rect 614356 217676 614362 217728
rect 531004 217552 538076 217580
rect 531004 217540 531010 217552
rect 542354 217540 542360 217592
rect 542412 217580 542418 217592
rect 543274 217580 543280 217592
rect 542412 217552 543280 217580
rect 542412 217540 542418 217552
rect 543274 217540 543280 217552
rect 543332 217580 543338 217592
rect 606202 217580 606208 217592
rect 543332 217552 606208 217580
rect 543332 217540 543338 217552
rect 606202 217540 606208 217552
rect 606260 217540 606266 217592
rect 614114 217540 614120 217592
rect 614172 217580 614178 217592
rect 626626 217580 626632 217592
rect 614172 217552 626632 217580
rect 614172 217540 614178 217552
rect 626626 217540 626632 217552
rect 626684 217540 626690 217592
rect 115290 217404 115296 217456
rect 115348 217444 115354 217456
rect 187970 217444 187976 217456
rect 115348 217416 187976 217444
rect 115348 217404 115354 217416
rect 187970 217404 187976 217416
rect 188028 217404 188034 217456
rect 527818 217404 527824 217456
rect 527876 217444 527882 217456
rect 528462 217444 528468 217456
rect 527876 217416 528468 217444
rect 527876 217404 527882 217416
rect 528462 217404 528468 217416
rect 528520 217444 528526 217456
rect 596910 217444 596916 217456
rect 528520 217416 596916 217444
rect 528520 217404 528526 217416
rect 596910 217404 596916 217416
rect 596968 217404 596974 217456
rect 603074 217404 603080 217456
rect 603132 217444 603138 217456
rect 628282 217444 628288 217456
rect 603132 217416 628288 217444
rect 603132 217404 603138 217416
rect 628282 217404 628288 217416
rect 628340 217404 628346 217456
rect 168558 217308 168564 217320
rect 93826 217280 168564 217308
rect 90404 217200 90410 217252
rect 90462 217240 90468 217252
rect 93826 217240 93854 217280
rect 168558 217268 168564 217280
rect 168616 217268 168622 217320
rect 506106 217268 506112 217320
rect 506164 217308 506170 217320
rect 506164 217280 563238 217308
rect 506164 217268 506170 217280
rect 90462 217212 93854 217240
rect 90462 217200 90468 217212
rect 436094 217200 436100 217252
rect 436152 217240 436158 217252
rect 437336 217240 437342 217252
rect 436152 217212 437342 217240
rect 436152 217200 436158 217212
rect 437336 217200 437342 217212
rect 437394 217200 437400 217252
rect 447134 217200 447140 217252
rect 447192 217240 447198 217252
rect 448100 217240 448106 217252
rect 447192 217212 448106 217240
rect 447192 217200 447198 217212
rect 448100 217200 448106 217212
rect 448158 217200 448164 217252
rect 469306 217200 469312 217252
rect 469364 217240 469370 217252
rect 470456 217240 470462 217252
rect 469364 217212 470462 217240
rect 469364 217200 469370 217212
rect 470456 217200 470462 217212
rect 470514 217200 470520 217252
rect 498194 217200 498200 217252
rect 498252 217240 498258 217252
rect 499436 217240 499442 217252
rect 498252 217212 499442 217240
rect 498252 217200 498258 217212
rect 499436 217200 499442 217212
rect 499494 217200 499500 217252
rect 508544 217132 508550 217184
rect 508602 217172 508608 217184
rect 563054 217172 563060 217184
rect 508602 217144 563060 217172
rect 508602 217132 508608 217144
rect 563054 217132 563060 217144
rect 563112 217132 563118 217184
rect 563210 217172 563238 217280
rect 563330 217268 563336 217320
rect 563388 217308 563394 217320
rect 571978 217308 571984 217320
rect 563388 217280 571984 217308
rect 563388 217268 563394 217280
rect 571978 217268 571984 217280
rect 572036 217268 572042 217320
rect 597922 217308 597928 217320
rect 572548 217280 597928 217308
rect 572548 217240 572576 217280
rect 597922 217268 597928 217280
rect 597980 217268 597986 217320
rect 598106 217268 598112 217320
rect 598164 217308 598170 217320
rect 622394 217308 622400 217320
rect 598164 217280 622400 217308
rect 598164 217268 598170 217280
rect 622394 217268 622400 217280
rect 622452 217268 622458 217320
rect 572180 217212 572576 217240
rect 572180 217172 572208 217212
rect 563210 217144 572208 217172
rect 572668 217132 572674 217184
rect 572726 217172 572732 217184
rect 596542 217172 596548 217184
rect 572726 217144 596548 217172
rect 572726 217132 572732 217144
rect 596542 217132 596548 217144
rect 596600 217132 596606 217184
rect 596910 217132 596916 217184
rect 596968 217172 596974 217184
rect 603074 217172 603080 217184
rect 596968 217144 603080 217172
rect 596968 217132 596974 217144
rect 603074 217132 603080 217144
rect 603132 217132 603138 217184
rect 498608 217064 498614 217116
rect 498666 217104 498672 217116
rect 498666 217076 499574 217104
rect 498666 217064 498672 217076
rect 499546 217036 499574 217076
rect 499546 217008 574048 217036
rect 574020 216900 574048 217008
rect 574186 216996 574192 217048
rect 574244 217036 574250 217048
rect 610066 217036 610072 217048
rect 574244 217008 610072 217036
rect 574244 216996 574250 217008
rect 610066 216996 610072 217008
rect 610124 216996 610130 217048
rect 596358 216900 596364 216912
rect 574020 216872 596364 216900
rect 596358 216860 596364 216872
rect 596416 216860 596422 216912
rect 596542 216860 596548 216912
rect 596600 216900 596606 216912
rect 598474 216900 598480 216912
rect 596600 216872 598480 216900
rect 596600 216860 596606 216872
rect 598474 216860 598480 216872
rect 598532 216860 598538 216912
rect 613378 216900 613384 216912
rect 605806 216872 613384 216900
rect 595990 216724 595996 216776
rect 596048 216764 596054 216776
rect 605806 216764 605834 216872
rect 613378 216860 613384 216872
rect 613436 216860 613442 216912
rect 596048 216736 605834 216764
rect 596048 216724 596054 216736
rect 610710 216724 610716 216776
rect 610768 216764 610774 216776
rect 615678 216764 615684 216776
rect 610768 216736 615684 216764
rect 610768 216724 610774 216736
rect 615678 216724 615684 216736
rect 615736 216724 615742 216776
rect 646314 216044 646320 216096
rect 646372 216084 646378 216096
rect 654778 216084 654784 216096
rect 646372 216056 654784 216084
rect 646372 216044 646378 216056
rect 654778 216044 654784 216056
rect 654836 216044 654842 216096
rect 649626 215908 649632 215960
rect 649684 215948 649690 215960
rect 659102 215948 659108 215960
rect 649684 215920 659108 215948
rect 649684 215908 649690 215920
rect 659102 215908 659108 215920
rect 659160 215908 659166 215960
rect 675846 215364 675852 215416
rect 675904 215404 675910 215416
rect 676950 215404 676956 215416
rect 675904 215376 676956 215404
rect 675904 215364 675910 215376
rect 676950 215364 676956 215376
rect 677008 215364 677014 215416
rect 574738 214820 574744 214872
rect 574796 214860 574802 214872
rect 616874 214860 616880 214872
rect 574796 214832 616880 214860
rect 574796 214820 574802 214832
rect 616874 214820 616880 214832
rect 616932 214820 616938 214872
rect 574370 214684 574376 214736
rect 574428 214724 574434 214736
rect 623314 214724 623320 214736
rect 574428 214696 623320 214724
rect 574428 214684 574434 214696
rect 623314 214684 623320 214696
rect 623372 214684 623378 214736
rect 574554 214548 574560 214600
rect 574612 214588 574618 214600
rect 574612 214560 605834 214588
rect 574612 214548 574618 214560
rect 601786 214412 601792 214464
rect 601844 214452 601850 214464
rect 602338 214452 602344 214464
rect 601844 214424 602344 214452
rect 601844 214412 601850 214424
rect 602338 214412 602344 214424
rect 602396 214412 602402 214464
rect 605806 214452 605834 214560
rect 607306 214548 607312 214600
rect 607364 214588 607370 214600
rect 607858 214588 607864 214600
rect 607364 214560 607864 214588
rect 607364 214548 607370 214560
rect 607858 214548 607864 214560
rect 607916 214548 607922 214600
rect 608778 214548 608784 214600
rect 608836 214588 608842 214600
rect 609514 214588 609520 214600
rect 608836 214560 609520 214588
rect 608836 214548 608842 214560
rect 609514 214548 609520 214560
rect 609572 214548 609578 214600
rect 618254 214548 618260 214600
rect 618312 214588 618318 214600
rect 618898 214588 618904 214600
rect 618312 214560 618904 214588
rect 618312 214548 618318 214560
rect 618898 214548 618904 214560
rect 618956 214548 618962 214600
rect 619910 214548 619916 214600
rect 619968 214588 619974 214600
rect 620554 214588 620560 214600
rect 619968 214560 620560 214588
rect 619968 214548 619974 214560
rect 620554 214548 620560 214560
rect 620612 214548 620618 214600
rect 623958 214548 623964 214600
rect 624016 214588 624022 214600
rect 624016 214560 625154 214588
rect 624016 214548 624022 214560
rect 624418 214452 624424 214464
rect 605806 214424 624424 214452
rect 624418 214412 624424 214424
rect 624476 214412 624482 214464
rect 625126 214452 625154 214560
rect 625430 214548 625436 214600
rect 625488 214588 625494 214600
rect 626074 214588 626080 214600
rect 625488 214560 626080 214588
rect 625488 214548 625494 214560
rect 626074 214548 626080 214560
rect 626132 214548 626138 214600
rect 630030 214548 630036 214600
rect 630088 214588 630094 214600
rect 632882 214588 632888 214600
rect 630088 214560 632888 214588
rect 630088 214548 630094 214560
rect 632882 214548 632888 214560
rect 632940 214548 632946 214600
rect 648246 214548 648252 214600
rect 648304 214588 648310 214600
rect 664438 214588 664444 214600
rect 648304 214560 664444 214588
rect 648304 214548 648310 214560
rect 664438 214548 664444 214560
rect 664496 214548 664502 214600
rect 664806 214548 664812 214600
rect 664864 214588 664870 214600
rect 666002 214588 666008 214600
rect 664864 214560 666008 214588
rect 664864 214548 664870 214560
rect 666002 214548 666008 214560
rect 666060 214548 666066 214600
rect 629386 214452 629392 214464
rect 625126 214424 629392 214452
rect 629386 214412 629392 214424
rect 629444 214412 629450 214464
rect 35802 213936 35808 213988
rect 35860 213976 35866 213988
rect 41690 213976 41696 213988
rect 35860 213948 41696 213976
rect 35860 213936 35866 213948
rect 41690 213936 41696 213948
rect 41748 213936 41754 213988
rect 646038 213868 646044 213920
rect 646096 213908 646102 213920
rect 646498 213908 646504 213920
rect 646096 213880 646504 213908
rect 646096 213868 646102 213880
rect 646498 213868 646504 213880
rect 646556 213868 646562 213920
rect 653214 213868 653220 213920
rect 653272 213908 653278 213920
rect 656158 213908 656164 213920
rect 653272 213880 656164 213908
rect 653272 213868 653278 213880
rect 656158 213868 656164 213880
rect 656216 213868 656222 213920
rect 645486 213732 645492 213784
rect 645544 213772 645550 213784
rect 649810 213772 649816 213784
rect 645544 213744 649816 213772
rect 645544 213732 645550 213744
rect 649810 213732 649816 213744
rect 649868 213732 649874 213784
rect 654134 213732 654140 213784
rect 654192 213772 654198 213784
rect 654778 213772 654784 213784
rect 654192 213744 654784 213772
rect 654192 213732 654198 213744
rect 654778 213732 654784 213744
rect 654836 213732 654842 213784
rect 663150 213732 663156 213784
rect 663208 213772 663214 213784
rect 665818 213772 665824 213784
rect 663208 213744 665824 213772
rect 663208 213732 663214 213744
rect 665818 213732 665824 213744
rect 665876 213732 665882 213784
rect 654594 213256 654600 213308
rect 654652 213296 654658 213308
rect 657538 213296 657544 213308
rect 654652 213268 657544 213296
rect 654652 213256 654658 213268
rect 657538 213256 657544 213268
rect 657596 213256 657602 213308
rect 673730 213256 673736 213308
rect 673788 213256 673794 213308
rect 575474 213188 575480 213240
rect 575532 213228 575538 213240
rect 594794 213228 594800 213240
rect 575532 213200 594800 213228
rect 575532 213188 575538 213200
rect 594794 213188 594800 213200
rect 594852 213188 594858 213240
rect 643830 213188 643836 213240
rect 643888 213228 643894 213240
rect 653398 213228 653404 213240
rect 643888 213200 653404 213228
rect 643888 213188 643894 213200
rect 653398 213188 653404 213200
rect 653456 213188 653462 213240
rect 673546 213228 673552 213240
rect 673380 213200 673552 213228
rect 600682 213120 600688 213172
rect 600740 213160 600746 213172
rect 601234 213160 601240 213172
rect 600740 213132 601240 213160
rect 600740 213120 600746 213132
rect 601234 213120 601240 213132
rect 601292 213120 601298 213172
rect 632698 212984 632704 213036
rect 632756 213024 632762 213036
rect 634354 213024 634360 213036
rect 632756 212996 634360 213024
rect 632756 212984 632762 212996
rect 634354 212984 634360 212996
rect 634412 212984 634418 213036
rect 664254 212984 664260 213036
rect 664312 213024 664318 213036
rect 665082 213024 665088 213036
rect 664312 212996 665088 213024
rect 664312 212984 664318 212996
rect 665082 212984 665088 212996
rect 665140 212984 665146 213036
rect 673380 212956 673408 213200
rect 673546 213188 673552 213200
rect 673604 213188 673610 213240
rect 673546 213052 673552 213104
rect 673604 213092 673610 213104
rect 673748 213092 673776 213256
rect 673604 213064 673776 213092
rect 673604 213052 673610 213064
rect 673730 212956 673736 212968
rect 673380 212928 673736 212956
rect 673730 212916 673736 212928
rect 673788 212916 673794 212968
rect 658182 212848 658188 212900
rect 658240 212888 658246 212900
rect 658918 212888 658924 212900
rect 658240 212860 658924 212888
rect 658240 212848 658246 212860
rect 658918 212848 658924 212860
rect 658976 212848 658982 212900
rect 650454 212712 650460 212764
rect 650512 212752 650518 212764
rect 651282 212752 651288 212764
rect 650512 212724 651288 212752
rect 650512 212712 650518 212724
rect 651282 212712 651288 212724
rect 651340 212712 651346 212764
rect 35802 212644 35808 212696
rect 35860 212684 35866 212696
rect 39574 212684 39580 212696
rect 35860 212656 39580 212684
rect 35860 212644 35866 212656
rect 39574 212644 39580 212656
rect 39632 212644 39638 212696
rect 591298 212644 591304 212696
rect 591356 212684 591362 212696
rect 639874 212684 639880 212696
rect 591356 212656 639880 212684
rect 591356 212644 591362 212656
rect 639874 212644 639880 212656
rect 639932 212644 639938 212696
rect 659562 212644 659568 212696
rect 659620 212684 659626 212696
rect 662414 212684 662420 212696
rect 659620 212656 662420 212684
rect 659620 212644 659626 212656
rect 662414 212644 662420 212656
rect 662472 212644 662478 212696
rect 592678 212508 592684 212560
rect 592736 212548 592742 212560
rect 641714 212548 641720 212560
rect 592736 212520 641720 212548
rect 592736 212508 592742 212520
rect 641714 212508 641720 212520
rect 641772 212508 641778 212560
rect 656526 212508 656532 212560
rect 656584 212548 656590 212560
rect 657906 212548 657912 212560
rect 656584 212520 657912 212548
rect 656584 212508 656590 212520
rect 657906 212508 657912 212520
rect 657964 212508 657970 212560
rect 578510 211148 578516 211200
rect 578568 211188 578574 211200
rect 580902 211188 580908 211200
rect 578568 211160 580908 211188
rect 578568 211148 578574 211160
rect 580902 211148 580908 211160
rect 580960 211148 580966 211200
rect 600406 210400 600412 210452
rect 600464 210440 600470 210452
rect 601004 210440 601010 210452
rect 600464 210412 601010 210440
rect 600464 210400 600470 210412
rect 601004 210400 601010 210412
rect 601062 210400 601068 210452
rect 35802 209924 35808 209976
rect 35860 209964 35866 209976
rect 40126 209964 40132 209976
rect 35860 209936 40132 209964
rect 35860 209924 35866 209936
rect 40126 209924 40132 209936
rect 40184 209924 40190 209976
rect 579522 209788 579528 209840
rect 579580 209828 579586 209840
rect 582282 209828 582288 209840
rect 579580 209800 582288 209828
rect 579580 209788 579586 209800
rect 582282 209788 582288 209800
rect 582340 209788 582346 209840
rect 632146 209556 632152 209568
rect 625126 209528 632152 209556
rect 35618 208632 35624 208684
rect 35676 208672 35682 208684
rect 39758 208672 39764 208684
rect 35676 208644 39764 208672
rect 35676 208632 35682 208644
rect 39758 208632 39764 208644
rect 39816 208632 39822 208684
rect 581638 208564 581644 208616
rect 581696 208604 581702 208616
rect 625126 208604 625154 209528
rect 632146 209516 632152 209528
rect 632204 209516 632210 209568
rect 652018 209516 652024 209568
rect 652076 209556 652082 209568
rect 652076 209528 654134 209556
rect 652076 209516 652082 209528
rect 654106 209080 654134 209528
rect 667014 209080 667020 209092
rect 654106 209052 667020 209080
rect 667014 209040 667020 209052
rect 667072 209040 667078 209092
rect 581696 208576 625154 208604
rect 581696 208564 581702 208576
rect 35802 208360 35808 208412
rect 35860 208400 35866 208412
rect 40034 208400 40040 208412
rect 35860 208372 40040 208400
rect 35860 208360 35866 208372
rect 40034 208360 40040 208372
rect 40092 208360 40098 208412
rect 578878 208292 578884 208344
rect 578936 208332 578942 208344
rect 589458 208332 589464 208344
rect 578936 208304 589464 208332
rect 578936 208292 578942 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 35802 207136 35808 207188
rect 35860 207176 35866 207188
rect 40126 207176 40132 207188
rect 35860 207148 40132 207176
rect 35860 207136 35866 207148
rect 40126 207136 40132 207148
rect 40184 207136 40190 207188
rect 580902 206864 580908 206916
rect 580960 206904 580966 206916
rect 589458 206904 589464 206916
rect 580960 206876 589464 206904
rect 580960 206864 580966 206876
rect 589458 206864 589464 206876
rect 589516 206864 589522 206916
rect 35802 205776 35808 205828
rect 35860 205816 35866 205828
rect 40218 205816 40224 205828
rect 35860 205788 40224 205816
rect 35860 205776 35866 205788
rect 40218 205776 40224 205788
rect 40276 205776 40282 205828
rect 579522 205776 579528 205828
rect 579580 205816 579586 205828
rect 580994 205816 581000 205828
rect 579580 205788 581000 205816
rect 579580 205776 579586 205788
rect 580994 205776 581000 205788
rect 581052 205776 581058 205828
rect 582282 205504 582288 205556
rect 582340 205544 582346 205556
rect 589458 205544 589464 205556
rect 582340 205516 589464 205544
rect 582340 205504 582346 205516
rect 589458 205504 589464 205516
rect 589516 205504 589522 205556
rect 35802 204416 35808 204468
rect 35860 204456 35866 204468
rect 41506 204456 41512 204468
rect 35860 204428 41512 204456
rect 35860 204416 35866 204428
rect 41506 204416 41512 204428
rect 41564 204416 41570 204468
rect 35618 204280 35624 204332
rect 35676 204320 35682 204332
rect 41690 204320 41696 204332
rect 35676 204292 41696 204320
rect 35676 204280 35682 204292
rect 41690 204280 41696 204292
rect 41748 204280 41754 204332
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 35802 202852 35808 202904
rect 35860 202892 35866 202904
rect 37918 202892 37924 202904
rect 35860 202864 37924 202892
rect 35860 202852 35866 202864
rect 37918 202852 37924 202864
rect 37976 202852 37982 202904
rect 578326 202852 578332 202904
rect 578384 202892 578390 202904
rect 580258 202892 580264 202904
rect 578384 202864 580264 202892
rect 578384 202852 578390 202864
rect 580258 202852 580264 202864
rect 580316 202852 580322 202904
rect 580994 202784 581000 202836
rect 581052 202824 581058 202836
rect 589458 202824 589464 202836
rect 581052 202796 589464 202824
rect 581052 202784 581058 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 578786 200132 578792 200184
rect 578844 200172 578850 200184
rect 590378 200172 590384 200184
rect 578844 200144 590384 200172
rect 578844 200132 578850 200144
rect 590378 200132 590384 200144
rect 590436 200132 590442 200184
rect 580258 199996 580264 200048
rect 580316 200036 580322 200048
rect 589458 200036 589464 200048
rect 580316 200008 589464 200036
rect 580316 199996 580322 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 579522 198704 579528 198756
rect 579580 198744 579586 198756
rect 589458 198744 589464 198756
rect 579580 198716 589464 198744
rect 579580 198704 579586 198716
rect 589458 198704 589464 198716
rect 589516 198704 589522 198756
rect 578510 195984 578516 196036
rect 578568 196024 578574 196036
rect 589274 196024 589280 196036
rect 578568 195996 589280 196024
rect 578568 195984 578574 195996
rect 589274 195984 589280 195996
rect 589332 195984 589338 196036
rect 579522 194556 579528 194608
rect 579580 194596 579586 194608
rect 589458 194596 589464 194608
rect 579580 194568 589464 194596
rect 579580 194556 579586 194568
rect 589458 194556 589464 194568
rect 589516 194556 589522 194608
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 589458 191876 589464 191888
rect 579580 191848 589464 191876
rect 579580 191836 579586 191848
rect 589458 191836 589464 191848
rect 589516 191836 589522 191888
rect 579522 190476 579528 190528
rect 579580 190516 579586 190528
rect 590562 190516 590568 190528
rect 579580 190488 590568 190516
rect 579580 190476 579586 190488
rect 590562 190476 590568 190488
rect 590620 190476 590626 190528
rect 579522 187688 579528 187740
rect 579580 187728 579586 187740
rect 589458 187728 589464 187740
rect 579580 187700 589464 187728
rect 579580 187688 579586 187700
rect 589458 187688 589464 187700
rect 589516 187688 589522 187740
rect 42426 187416 42432 187468
rect 42484 187456 42490 187468
rect 43254 187456 43260 187468
rect 42484 187428 43260 187456
rect 42484 187416 42490 187428
rect 43254 187416 43260 187428
rect 43312 187416 43318 187468
rect 579522 186260 579528 186312
rect 579580 186300 579586 186312
rect 589642 186300 589648 186312
rect 579580 186272 589648 186300
rect 579580 186260 579586 186272
rect 589642 186260 589648 186272
rect 589700 186260 589706 186312
rect 579522 184832 579528 184884
rect 579580 184872 579586 184884
rect 589458 184872 589464 184884
rect 579580 184844 589464 184872
rect 579580 184832 579586 184844
rect 589458 184832 589464 184844
rect 589516 184832 589522 184884
rect 669222 184832 669228 184884
rect 669280 184872 669286 184884
rect 670694 184872 670700 184884
rect 669280 184844 670700 184872
rect 669280 184832 669286 184844
rect 670694 184832 670700 184844
rect 670752 184832 670758 184884
rect 42150 183472 42156 183524
rect 42208 183512 42214 183524
rect 42978 183512 42984 183524
rect 42208 183484 42984 183512
rect 42208 183472 42214 183484
rect 42978 183472 42984 183484
rect 43036 183472 43042 183524
rect 579522 182112 579528 182164
rect 579580 182152 579586 182164
rect 589458 182152 589464 182164
rect 579580 182124 589464 182152
rect 579580 182112 579586 182124
rect 589458 182112 589464 182124
rect 589516 182112 589522 182164
rect 578786 180752 578792 180804
rect 578844 180792 578850 180804
rect 590562 180792 590568 180804
rect 578844 180764 590568 180792
rect 578844 180752 578850 180764
rect 590562 180752 590568 180764
rect 590620 180752 590626 180804
rect 578786 178032 578792 178084
rect 578844 178072 578850 178084
rect 589458 178072 589464 178084
rect 578844 178044 589464 178072
rect 578844 178032 578850 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 668210 177964 668216 178016
rect 668268 178004 668274 178016
rect 670786 178004 670792 178016
rect 668268 177976 670792 178004
rect 668268 177964 668274 177976
rect 670786 177964 670792 177976
rect 670844 177964 670850 178016
rect 579522 177896 579528 177948
rect 579580 177936 579586 177948
rect 589642 177936 589648 177948
rect 579580 177908 589648 177936
rect 579580 177896 579586 177908
rect 589642 177896 589648 177908
rect 589700 177896 589706 177948
rect 589458 175352 589464 175364
rect 586486 175324 589464 175352
rect 579982 175244 579988 175296
rect 580040 175284 580046 175296
rect 586486 175284 586514 175324
rect 589458 175312 589464 175324
rect 589516 175312 589522 175364
rect 580040 175256 586514 175284
rect 580040 175244 580046 175256
rect 667934 174700 667940 174752
rect 667992 174740 667998 174752
rect 669590 174740 669596 174752
rect 667992 174712 669596 174740
rect 667992 174700 667998 174712
rect 669590 174700 669596 174712
rect 669648 174700 669654 174752
rect 578418 174496 578424 174548
rect 578476 174536 578482 174548
rect 589642 174536 589648 174548
rect 578476 174508 589648 174536
rect 578476 174496 578482 174508
rect 589642 174496 589648 174508
rect 589700 174496 589706 174548
rect 578234 172864 578240 172916
rect 578292 172904 578298 172916
rect 579982 172904 579988 172916
rect 578292 172876 579988 172904
rect 578292 172864 578298 172876
rect 579982 172864 579988 172876
rect 580040 172864 580046 172916
rect 580902 172524 580908 172576
rect 580960 172564 580966 172576
rect 589458 172564 589464 172576
rect 580960 172536 589464 172564
rect 580960 172524 580966 172536
rect 589458 172524 589464 172536
rect 589516 172524 589522 172576
rect 580258 171096 580264 171148
rect 580316 171136 580322 171148
rect 589458 171136 589464 171148
rect 580316 171108 589464 171136
rect 580316 171096 580322 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 578694 169736 578700 169788
rect 578752 169776 578758 169788
rect 580902 169776 580908 169788
rect 578752 169748 580908 169776
rect 578752 169736 578758 169748
rect 580902 169736 580908 169748
rect 580960 169736 580966 169788
rect 667934 169668 667940 169720
rect 667992 169708 667998 169720
rect 669774 169708 669780 169720
rect 667992 169680 669780 169708
rect 667992 169668 667998 169680
rect 669774 169668 669780 169680
rect 669832 169668 669838 169720
rect 582374 168376 582380 168428
rect 582432 168416 582438 168428
rect 589458 168416 589464 168428
rect 582432 168388 589464 168416
rect 582432 168376 582438 168388
rect 589458 168376 589464 168388
rect 589516 168376 589522 168428
rect 578234 167288 578240 167340
rect 578292 167328 578298 167340
rect 580258 167328 580264 167340
rect 578292 167300 580264 167328
rect 578292 167288 578298 167300
rect 580258 167288 580264 167300
rect 580316 167288 580322 167340
rect 579982 167016 579988 167068
rect 580040 167056 580046 167068
rect 589458 167056 589464 167068
rect 580040 167028 589464 167056
rect 580040 167016 580046 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 579522 166268 579528 166320
rect 579580 166308 579586 166320
rect 589642 166308 589648 166320
rect 579580 166280 589648 166308
rect 579580 166268 579586 166280
rect 589642 166268 589648 166280
rect 589700 166268 589706 166320
rect 579338 165180 579344 165232
rect 579396 165220 579402 165232
rect 582374 165220 582380 165232
rect 579396 165192 582380 165220
rect 579396 165180 579402 165192
rect 582374 165180 582380 165192
rect 582432 165180 582438 165232
rect 668026 164908 668032 164960
rect 668084 164948 668090 164960
rect 670326 164948 670332 164960
rect 668084 164920 670332 164948
rect 668084 164908 668090 164920
rect 670326 164908 670332 164920
rect 670384 164908 670390 164960
rect 582466 164228 582472 164280
rect 582524 164268 582530 164280
rect 589458 164268 589464 164280
rect 582524 164240 589464 164268
rect 582524 164228 582530 164240
rect 589458 164228 589464 164240
rect 589516 164228 589522 164280
rect 578234 163616 578240 163668
rect 578292 163656 578298 163668
rect 579982 163656 579988 163668
rect 578292 163628 579988 163656
rect 578292 163616 578298 163628
rect 579982 163616 579988 163628
rect 580040 163616 580046 163668
rect 675846 163208 675852 163260
rect 675904 163248 675910 163260
rect 679618 163248 679624 163260
rect 675904 163220 679624 163248
rect 675904 163208 675910 163220
rect 679618 163208 679624 163220
rect 679676 163208 679682 163260
rect 580902 162868 580908 162920
rect 580960 162908 580966 162920
rect 589458 162908 589464 162920
rect 580960 162880 589464 162908
rect 580960 162868 580966 162880
rect 589458 162868 589464 162880
rect 589516 162868 589522 162920
rect 676030 162732 676036 162784
rect 676088 162772 676094 162784
rect 680998 162772 681004 162784
rect 676088 162744 681004 162772
rect 676088 162732 676094 162744
rect 680998 162732 681004 162744
rect 681056 162732 681062 162784
rect 578418 162664 578424 162716
rect 578476 162704 578482 162716
rect 582466 162704 582472 162716
rect 578476 162676 582472 162704
rect 578476 162664 578482 162676
rect 582466 162664 582472 162676
rect 582524 162664 582530 162716
rect 580534 161440 580540 161492
rect 580592 161480 580598 161492
rect 589458 161480 589464 161492
rect 580592 161452 589464 161480
rect 580592 161440 580598 161452
rect 589458 161440 589464 161452
rect 589516 161440 589522 161492
rect 580718 160080 580724 160132
rect 580776 160120 580782 160132
rect 589458 160120 589464 160132
rect 580776 160092 589464 160120
rect 580776 160080 580782 160092
rect 589458 160080 589464 160092
rect 589516 160080 589522 160132
rect 668210 160012 668216 160064
rect 668268 160052 668274 160064
rect 670786 160052 670792 160064
rect 668268 160024 670792 160052
rect 668268 160012 668274 160024
rect 670786 160012 670792 160024
rect 670844 160012 670850 160064
rect 578878 158720 578884 158772
rect 578936 158760 578942 158772
rect 580902 158760 580908 158772
rect 578936 158732 580908 158760
rect 578936 158720 578942 158732
rect 580902 158720 580908 158732
rect 580960 158720 580966 158772
rect 585778 158720 585784 158772
rect 585836 158760 585842 158772
rect 589458 158760 589464 158772
rect 585836 158732 589464 158760
rect 585836 158720 585842 158732
rect 589458 158720 589464 158732
rect 589516 158720 589522 158772
rect 587158 157360 587164 157412
rect 587216 157400 587222 157412
rect 589274 157400 589280 157412
rect 587216 157372 589280 157400
rect 587216 157360 587222 157372
rect 589274 157360 589280 157372
rect 589332 157360 589338 157412
rect 668210 155116 668216 155168
rect 668268 155156 668274 155168
rect 670786 155156 670792 155168
rect 668268 155128 670792 155156
rect 668268 155116 668274 155128
rect 670786 155116 670792 155128
rect 670844 155116 670850 155168
rect 578326 154776 578332 154828
rect 578384 154816 578390 154828
rect 580534 154816 580540 154828
rect 578384 154788 580540 154816
rect 578384 154776 578390 154788
rect 580534 154776 580540 154788
rect 580592 154776 580598 154828
rect 584398 154572 584404 154624
rect 584456 154612 584462 154624
rect 589458 154612 589464 154624
rect 584456 154584 589464 154612
rect 584456 154572 584462 154584
rect 589458 154572 589464 154584
rect 589516 154572 589522 154624
rect 583018 153212 583024 153264
rect 583076 153252 583082 153264
rect 589458 153252 589464 153264
rect 583076 153224 589464 153252
rect 583076 153212 583082 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 578234 152736 578240 152788
rect 578292 152776 578298 152788
rect 580718 152776 580724 152788
rect 578292 152748 580724 152776
rect 578292 152736 578298 152748
rect 580718 152736 580724 152748
rect 580776 152736 580782 152788
rect 580258 151784 580264 151836
rect 580316 151824 580322 151836
rect 589458 151824 589464 151836
rect 580316 151796 589464 151824
rect 580316 151784 580322 151796
rect 589458 151784 589464 151796
rect 589516 151784 589522 151836
rect 578878 150560 578884 150612
rect 578936 150600 578942 150612
rect 585778 150600 585784 150612
rect 578936 150572 585784 150600
rect 578936 150560 578942 150572
rect 585778 150560 585784 150572
rect 585836 150560 585842 150612
rect 585134 149064 585140 149116
rect 585192 149104 585198 149116
rect 589458 149104 589464 149116
rect 585192 149076 589464 149104
rect 585192 149064 585198 149076
rect 589458 149064 589464 149076
rect 589516 149064 589522 149116
rect 579522 148316 579528 148368
rect 579580 148356 579586 148368
rect 587158 148356 587164 148368
rect 579580 148328 587164 148356
rect 579580 148316 579586 148328
rect 587158 148316 587164 148328
rect 587216 148316 587222 148368
rect 578878 146276 578884 146328
rect 578936 146316 578942 146328
rect 585134 146316 585140 146328
rect 578936 146288 585140 146316
rect 578936 146276 578942 146288
rect 585134 146276 585140 146288
rect 585192 146276 585198 146328
rect 668762 146004 668768 146056
rect 668820 146044 668826 146056
rect 670786 146044 670792 146056
rect 668820 146016 670792 146044
rect 668820 146004 668826 146016
rect 670786 146004 670792 146016
rect 670844 146004 670850 146056
rect 584766 144916 584772 144968
rect 584824 144956 584830 144968
rect 589458 144956 589464 144968
rect 584824 144928 589464 144956
rect 584824 144916 584830 144928
rect 589458 144916 589464 144928
rect 589516 144916 589522 144968
rect 579246 144644 579252 144696
rect 579304 144684 579310 144696
rect 584398 144684 584404 144696
rect 579304 144656 584404 144684
rect 579304 144644 579310 144656
rect 584398 144644 584404 144656
rect 584456 144644 584462 144696
rect 585962 143556 585968 143608
rect 586020 143596 586026 143608
rect 589458 143596 589464 143608
rect 586020 143568 589464 143596
rect 586020 143556 586026 143568
rect 589458 143556 589464 143568
rect 589516 143556 589522 143608
rect 579522 143420 579528 143472
rect 579580 143460 579586 143472
rect 583018 143460 583024 143472
rect 579580 143432 583024 143460
rect 579580 143420 579586 143432
rect 583018 143420 583024 143432
rect 583076 143420 583082 143472
rect 587158 142400 587164 142452
rect 587216 142440 587222 142452
rect 589826 142440 589832 142452
rect 587216 142412 589832 142440
rect 587216 142400 587222 142412
rect 589826 142400 589832 142412
rect 589884 142400 589890 142452
rect 580442 140768 580448 140820
rect 580500 140808 580506 140820
rect 589458 140808 589464 140820
rect 580500 140780 589464 140808
rect 580500 140768 580506 140780
rect 589458 140768 589464 140780
rect 589516 140768 589522 140820
rect 578602 140700 578608 140752
rect 578660 140740 578666 140752
rect 580258 140740 580264 140752
rect 578660 140712 580264 140740
rect 578660 140700 578666 140712
rect 580258 140700 580264 140712
rect 580316 140700 580322 140752
rect 583018 139408 583024 139460
rect 583076 139448 583082 139460
rect 589458 139448 589464 139460
rect 583076 139420 589464 139448
rect 583076 139408 583082 139420
rect 589458 139408 589464 139420
rect 589516 139408 589522 139460
rect 578602 139272 578608 139324
rect 578660 139312 578666 139324
rect 589918 139312 589924 139324
rect 578660 139284 589924 139312
rect 578660 139272 578666 139284
rect 589918 139272 589924 139284
rect 589976 139272 589982 139324
rect 579522 138660 579528 138712
rect 579580 138700 579586 138712
rect 588538 138700 588544 138712
rect 579580 138672 588544 138700
rect 579580 138660 579586 138672
rect 588538 138660 588544 138672
rect 588596 138660 588602 138712
rect 579062 137300 579068 137352
rect 579120 137340 579126 137352
rect 584766 137340 584772 137352
rect 579120 137312 584772 137340
rect 579120 137300 579126 137312
rect 584766 137300 584772 137312
rect 584824 137300 584830 137352
rect 584582 136620 584588 136672
rect 584640 136660 584646 136672
rect 589458 136660 589464 136672
rect 584640 136632 589464 136660
rect 584640 136620 584646 136632
rect 589458 136620 589464 136632
rect 589516 136620 589522 136672
rect 580258 134512 580264 134564
rect 580316 134552 580322 134564
rect 589458 134552 589464 134564
rect 580316 134524 589464 134552
rect 580316 134512 580322 134524
rect 589458 134512 589464 134524
rect 589516 134512 589522 134564
rect 667934 133764 667940 133816
rect 667992 133804 667998 133816
rect 669958 133804 669964 133816
rect 667992 133776 669964 133804
rect 667992 133764 667998 133776
rect 669958 133764 669964 133776
rect 670016 133764 670022 133816
rect 585778 132472 585784 132524
rect 585836 132512 585842 132524
rect 589458 132512 589464 132524
rect 585836 132484 589464 132512
rect 585836 132472 585842 132484
rect 589458 132472 589464 132484
rect 589516 132472 589522 132524
rect 581822 131248 581828 131300
rect 581880 131288 581886 131300
rect 589458 131288 589464 131300
rect 581880 131260 589464 131288
rect 581880 131248 581886 131260
rect 589458 131248 589464 131260
rect 589516 131248 589522 131300
rect 578878 131112 578884 131164
rect 578936 131152 578942 131164
rect 585962 131152 585968 131164
rect 578936 131124 585968 131152
rect 578936 131112 578942 131124
rect 585962 131112 585968 131124
rect 586020 131112 586026 131164
rect 668670 130636 668676 130688
rect 668728 130676 668734 130688
rect 670786 130676 670792 130688
rect 668728 130648 670792 130676
rect 668728 130636 668734 130648
rect 670786 130636 670792 130648
rect 670844 130636 670850 130688
rect 667934 129548 667940 129600
rect 667992 129588 667998 129600
rect 670142 129588 670148 129600
rect 667992 129560 670148 129588
rect 667992 129548 667998 129560
rect 670142 129548 670148 129560
rect 670200 129548 670206 129600
rect 583202 129140 583208 129192
rect 583260 129180 583266 129192
rect 590378 129180 590384 129192
rect 583260 129152 590384 129180
rect 583260 129140 583266 129152
rect 590378 129140 590384 129152
rect 590436 129140 590442 129192
rect 579522 129004 579528 129056
rect 579580 129044 579586 129056
rect 587158 129044 587164 129056
rect 579580 129016 587164 129044
rect 579580 129004 579586 129016
rect 587158 129004 587164 129016
rect 587216 129004 587222 129056
rect 579062 126964 579068 127016
rect 579120 127004 579126 127016
rect 589458 127004 589464 127016
rect 579120 126976 589464 127004
rect 579120 126964 579126 126976
rect 589458 126964 589464 126976
rect 589516 126964 589522 127016
rect 578326 125604 578332 125656
rect 578384 125644 578390 125656
rect 580442 125644 580448 125656
rect 578384 125616 580448 125644
rect 578384 125604 578390 125616
rect 580442 125604 580448 125616
rect 580500 125604 580506 125656
rect 580442 124176 580448 124228
rect 580500 124216 580506 124228
rect 589458 124216 589464 124228
rect 580500 124188 589464 124216
rect 580500 124176 580506 124188
rect 589458 124176 589464 124188
rect 589516 124176 589522 124228
rect 578418 123564 578424 123616
rect 578476 123604 578482 123616
rect 583018 123604 583024 123616
rect 578476 123576 583024 123604
rect 578476 123564 578482 123576
rect 583018 123564 583024 123576
rect 583076 123564 583082 123616
rect 584398 122816 584404 122868
rect 584456 122856 584462 122868
rect 589458 122856 589464 122868
rect 584456 122828 589464 122856
rect 584456 122816 584462 122828
rect 589458 122816 589464 122828
rect 589516 122816 589522 122868
rect 578878 122136 578884 122188
rect 578936 122176 578942 122188
rect 584582 122176 584588 122188
rect 578936 122148 584588 122176
rect 578936 122136 578942 122148
rect 584582 122136 584588 122148
rect 584640 122136 584646 122188
rect 580626 122000 580632 122052
rect 580684 122040 580690 122052
rect 589918 122040 589924 122052
rect 580684 122012 589924 122040
rect 580684 122000 580690 122012
rect 589918 122000 589924 122012
rect 589976 122000 589982 122052
rect 675846 120028 675852 120080
rect 675904 120068 675910 120080
rect 676398 120068 676404 120080
rect 675904 120040 676404 120068
rect 675904 120028 675910 120040
rect 676398 120028 676404 120040
rect 676456 120028 676462 120080
rect 587342 118668 587348 118720
rect 587400 118708 587406 118720
rect 590010 118708 590016 118720
rect 587400 118680 590016 118708
rect 587400 118668 587406 118680
rect 590010 118668 590016 118680
rect 590068 118668 590074 118720
rect 578510 118396 578516 118448
rect 578568 118436 578574 118448
rect 580258 118436 580264 118448
rect 578568 118408 580264 118436
rect 578568 118396 578574 118408
rect 580258 118396 580264 118408
rect 580316 118396 580322 118448
rect 579522 116900 579528 116952
rect 579580 116940 579586 116952
rect 583202 116940 583208 116952
rect 579580 116912 583208 116940
rect 579580 116900 579586 116912
rect 583202 116900 583208 116912
rect 583260 116900 583266 116952
rect 586146 115948 586152 116000
rect 586204 115988 586210 116000
rect 589458 115988 589464 116000
rect 586204 115960 589464 115988
rect 586204 115948 586210 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 583202 115200 583208 115252
rect 583260 115240 583266 115252
rect 589642 115240 589648 115252
rect 583260 115212 589648 115240
rect 583260 115200 583266 115212
rect 589642 115200 589648 115212
rect 589700 115200 589706 115252
rect 579246 114452 579252 114504
rect 579304 114492 579310 114504
rect 581638 114492 581644 114504
rect 579304 114464 581644 114492
rect 579304 114452 579310 114464
rect 581638 114452 581644 114464
rect 581696 114452 581702 114504
rect 583018 113160 583024 113212
rect 583076 113200 583082 113212
rect 589458 113200 589464 113212
rect 583076 113172 589464 113200
rect 583076 113160 583082 113172
rect 589458 113160 589464 113172
rect 589516 113160 589522 113212
rect 668118 112888 668124 112940
rect 668176 112928 668182 112940
rect 670142 112928 670148 112940
rect 668176 112900 670148 112928
rect 668176 112888 668182 112900
rect 670142 112888 670148 112900
rect 670200 112888 670206 112940
rect 579522 112820 579528 112872
rect 579580 112860 579586 112872
rect 585778 112860 585784 112872
rect 579580 112832 585784 112860
rect 579580 112820 579586 112832
rect 585778 112820 585784 112832
rect 585836 112820 585842 112872
rect 585962 112412 585968 112464
rect 586020 112452 586026 112464
rect 590102 112452 590108 112464
rect 586020 112424 590108 112452
rect 586020 112412 586026 112424
rect 590102 112412 590108 112424
rect 590160 112412 590166 112464
rect 581638 110440 581644 110492
rect 581696 110480 581702 110492
rect 589458 110480 589464 110492
rect 581696 110452 589464 110480
rect 581696 110440 581702 110452
rect 589458 110440 589464 110452
rect 589516 110440 589522 110492
rect 579338 110100 579344 110152
rect 579396 110140 579402 110152
rect 581822 110140 581828 110152
rect 579396 110112 581828 110140
rect 579396 110100 579402 110112
rect 581822 110100 581828 110112
rect 581880 110100 581886 110152
rect 584582 109012 584588 109064
rect 584640 109052 584646 109064
rect 589274 109052 589280 109064
rect 584640 109024 589280 109052
rect 584640 109012 584646 109024
rect 589274 109012 589280 109024
rect 589332 109012 589338 109064
rect 578326 108672 578332 108724
rect 578384 108712 578390 108724
rect 580626 108712 580632 108724
rect 578384 108684 580632 108712
rect 578384 108672 578390 108684
rect 580626 108672 580632 108684
rect 580684 108672 580690 108724
rect 668394 107992 668400 108044
rect 668452 108032 668458 108044
rect 670786 108032 670792 108044
rect 668452 108004 670792 108032
rect 668452 107992 668458 108004
rect 670786 107992 670792 108004
rect 670844 107992 670850 108044
rect 589458 107692 589464 107704
rect 579632 107664 589464 107692
rect 578878 107584 578884 107636
rect 578936 107624 578942 107636
rect 579632 107624 579660 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 578936 107596 579660 107624
rect 578936 107584 578942 107596
rect 587158 106292 587164 106344
rect 587216 106332 587222 106344
rect 589826 106332 589832 106344
rect 587216 106304 589832 106332
rect 587216 106292 587222 106304
rect 589826 106292 589832 106304
rect 589884 106292 589890 106344
rect 580258 104864 580264 104916
rect 580316 104904 580322 104916
rect 589458 104904 589464 104916
rect 580316 104876 589464 104904
rect 580316 104864 580322 104876
rect 589458 104864 589464 104876
rect 589516 104864 589522 104916
rect 667934 104524 667940 104576
rect 667992 104564 667998 104576
rect 669958 104564 669964 104576
rect 667992 104536 669964 104564
rect 667992 104524 667998 104536
rect 669958 104524 669964 104536
rect 670016 104524 670022 104576
rect 579522 103436 579528 103488
rect 579580 103476 579586 103488
rect 588538 103476 588544 103488
rect 579580 103448 588544 103476
rect 579580 103436 579586 103448
rect 588538 103436 588544 103448
rect 588596 103436 588602 103488
rect 579522 101804 579528 101856
rect 579580 101844 579586 101856
rect 584398 101844 584404 101856
rect 579580 101816 584404 101844
rect 579580 101804 579586 101816
rect 584398 101804 584404 101816
rect 584456 101804 584462 101856
rect 584398 100104 584404 100156
rect 584456 100144 584462 100156
rect 589458 100144 589464 100156
rect 584456 100116 589464 100144
rect 584456 100104 584462 100116
rect 589458 100104 589464 100116
rect 589516 100104 589522 100156
rect 579062 99356 579068 99408
rect 579120 99396 579126 99408
rect 586146 99396 586152 99408
rect 579120 99368 586152 99396
rect 579120 99356 579126 99368
rect 586146 99356 586152 99368
rect 586204 99356 586210 99408
rect 622302 99288 622308 99340
rect 622360 99328 622366 99340
rect 630766 99328 630772 99340
rect 622360 99300 630772 99328
rect 622360 99288 622366 99300
rect 630766 99288 630772 99300
rect 630824 99288 630830 99340
rect 578602 99220 578608 99272
rect 578660 99260 578666 99272
rect 580442 99260 580448 99272
rect 578660 99232 580448 99260
rect 578660 99220 578666 99232
rect 580442 99220 580448 99232
rect 580500 99220 580506 99272
rect 623682 99152 623688 99204
rect 623740 99192 623746 99204
rect 633434 99192 633440 99204
rect 623740 99164 633440 99192
rect 623740 99152 623746 99164
rect 633434 99152 633440 99164
rect 633492 99152 633498 99204
rect 577498 99084 577504 99136
rect 577556 99124 577562 99136
rect 595254 99124 595260 99136
rect 577556 99096 595260 99124
rect 577556 99084 577562 99096
rect 595254 99084 595260 99096
rect 595312 99084 595318 99136
rect 625062 99016 625068 99068
rect 625120 99056 625126 99068
rect 636286 99056 636292 99068
rect 625120 99028 636292 99056
rect 625120 99016 625126 99028
rect 636286 99016 636292 99028
rect 636344 99016 636350 99068
rect 628282 98880 628288 98932
rect 628340 98920 628346 98932
rect 642174 98920 642180 98932
rect 628340 98892 642180 98920
rect 628340 98880 628346 98892
rect 642174 98880 642180 98892
rect 642232 98880 642238 98932
rect 629018 98744 629024 98796
rect 629076 98784 629082 98796
rect 643646 98784 643652 98796
rect 629076 98756 643652 98784
rect 629076 98744 629082 98756
rect 643646 98744 643652 98756
rect 643704 98744 643710 98796
rect 647142 98608 647148 98660
rect 647200 98648 647206 98660
rect 661954 98648 661960 98660
rect 647200 98620 661960 98648
rect 647200 98608 647206 98620
rect 661954 98608 661960 98620
rect 662012 98608 662018 98660
rect 630490 98472 630496 98524
rect 630548 98512 630554 98524
rect 646590 98512 646596 98524
rect 630548 98484 646596 98512
rect 630548 98472 630554 98484
rect 646590 98472 646596 98484
rect 646648 98472 646654 98524
rect 631042 98200 631048 98252
rect 631100 98240 631106 98252
rect 631100 98212 634814 98240
rect 631100 98200 631106 98212
rect 634786 98172 634814 98212
rect 640702 98172 640708 98184
rect 634786 98144 640708 98172
rect 640702 98132 640708 98144
rect 640760 98132 640766 98184
rect 631980 98076 632192 98104
rect 578326 97928 578332 97980
rect 578384 97968 578390 97980
rect 587342 97968 587348 97980
rect 578384 97940 587348 97968
rect 578384 97928 578390 97940
rect 587342 97928 587348 97940
rect 587400 97928 587406 97980
rect 620186 97928 620192 97980
rect 620244 97968 620250 97980
rect 626258 97968 626264 97980
rect 620244 97940 626264 97968
rect 620244 97928 620250 97940
rect 626258 97928 626264 97940
rect 626316 97928 626322 97980
rect 629754 97928 629760 97980
rect 629812 97968 629818 97980
rect 631980 97968 632008 98076
rect 632164 98036 632192 98076
rect 645302 98036 645308 98048
rect 632164 98008 645308 98036
rect 645302 97996 645308 98008
rect 645360 97996 645366 98048
rect 629812 97940 632008 97968
rect 629812 97928 629818 97940
rect 659194 97928 659200 97980
rect 659252 97968 659258 97980
rect 663886 97968 663892 97980
rect 659252 97940 663892 97968
rect 659252 97928 659258 97940
rect 663886 97928 663892 97940
rect 663944 97928 663950 97980
rect 618714 97792 618720 97844
rect 618772 97832 618778 97844
rect 625798 97832 625804 97844
rect 618772 97804 625804 97832
rect 618772 97792 618778 97804
rect 625798 97792 625804 97804
rect 625856 97792 625862 97844
rect 627546 97792 627552 97844
rect 627604 97832 627610 97844
rect 631042 97832 631048 97844
rect 627604 97804 631048 97832
rect 627604 97792 627610 97804
rect 631042 97792 631048 97804
rect 631100 97792 631106 97844
rect 634170 97792 634176 97844
rect 634228 97832 634234 97844
rect 650546 97832 650552 97844
rect 634228 97804 650552 97832
rect 634228 97792 634234 97804
rect 650546 97792 650552 97804
rect 650604 97792 650610 97844
rect 655422 97792 655428 97844
rect 655480 97832 655486 97844
rect 655480 97804 659792 97832
rect 655480 97792 655486 97804
rect 634722 97656 634728 97708
rect 634780 97696 634786 97708
rect 650178 97696 650184 97708
rect 634780 97668 650184 97696
rect 634780 97656 634786 97668
rect 650178 97656 650184 97668
rect 650236 97656 650242 97708
rect 651834 97656 651840 97708
rect 651892 97696 651898 97708
rect 659562 97696 659568 97708
rect 651892 97668 659568 97696
rect 651892 97656 651898 97668
rect 659562 97656 659568 97668
rect 659620 97656 659626 97708
rect 659764 97696 659792 97804
rect 659930 97792 659936 97844
rect 659988 97832 659994 97844
rect 665174 97832 665180 97844
rect 659988 97804 665180 97832
rect 659988 97792 659994 97804
rect 665174 97792 665180 97804
rect 665232 97792 665238 97844
rect 662506 97696 662512 97708
rect 659764 97668 662512 97696
rect 662506 97656 662512 97668
rect 662564 97656 662570 97708
rect 621658 97520 621664 97572
rect 621716 97560 621722 97572
rect 629294 97560 629300 97572
rect 621716 97532 629300 97560
rect 621716 97520 621722 97532
rect 629294 97520 629300 97532
rect 629352 97520 629358 97572
rect 631962 97520 631968 97572
rect 632020 97560 632026 97572
rect 647510 97560 647516 97572
rect 632020 97532 647516 97560
rect 632020 97520 632026 97532
rect 647510 97520 647516 97532
rect 647568 97520 647574 97572
rect 650362 97452 650368 97504
rect 650420 97492 650426 97504
rect 658274 97492 658280 97504
rect 650420 97464 658280 97492
rect 650420 97452 650426 97464
rect 658274 97452 658280 97464
rect 658332 97452 658338 97504
rect 612642 97384 612648 97436
rect 612700 97424 612706 97436
rect 618898 97424 618904 97436
rect 612700 97396 618904 97424
rect 612700 97384 612706 97396
rect 618898 97384 618904 97396
rect 618956 97384 618962 97436
rect 623130 97384 623136 97436
rect 623188 97424 623194 97436
rect 632054 97424 632060 97436
rect 623188 97396 632060 97424
rect 623188 97384 623194 97396
rect 632054 97384 632060 97396
rect 632112 97384 632118 97436
rect 633250 97384 633256 97436
rect 633308 97424 633314 97436
rect 648614 97424 648620 97436
rect 633308 97396 648620 97424
rect 633308 97384 633314 97396
rect 648614 97384 648620 97396
rect 648672 97384 648678 97436
rect 658090 97316 658096 97368
rect 658148 97356 658154 97368
rect 663058 97356 663064 97368
rect 658148 97328 663064 97356
rect 658148 97316 658154 97328
rect 663058 97316 663064 97328
rect 663116 97316 663122 97368
rect 605466 97248 605472 97300
rect 605524 97288 605530 97300
rect 611906 97288 611912 97300
rect 605524 97260 611912 97288
rect 605524 97248 605530 97260
rect 611906 97248 611912 97260
rect 611964 97248 611970 97300
rect 626074 97248 626080 97300
rect 626132 97288 626138 97300
rect 637758 97288 637764 97300
rect 626132 97260 637764 97288
rect 626132 97248 626138 97260
rect 637758 97248 637764 97260
rect 637816 97248 637822 97300
rect 644290 97248 644296 97300
rect 644348 97288 644354 97300
rect 644348 97260 656710 97288
rect 644348 97248 644354 97260
rect 626810 97112 626816 97164
rect 626868 97152 626874 97164
rect 639230 97152 639236 97164
rect 626868 97124 639236 97152
rect 626868 97112 626874 97124
rect 639230 97112 639236 97124
rect 639288 97112 639294 97164
rect 643002 97112 643008 97164
rect 643060 97152 643066 97164
rect 643060 97124 656572 97152
rect 643060 97112 643066 97124
rect 624602 96976 624608 97028
rect 624660 97016 624666 97028
rect 634998 97016 635004 97028
rect 624660 96988 635004 97016
rect 624660 96976 624666 96988
rect 634998 96976 635004 96988
rect 635056 96976 635062 97028
rect 635550 96976 635556 97028
rect 635608 97016 635614 97028
rect 647694 97016 647700 97028
rect 635608 96988 647700 97016
rect 635608 96976 635614 96988
rect 647694 96976 647700 96988
rect 647752 96976 647758 97028
rect 598934 96908 598940 96960
rect 598992 96948 598998 96960
rect 599670 96948 599676 96960
rect 598992 96920 599676 96948
rect 598992 96908 598998 96920
rect 599670 96908 599676 96920
rect 599728 96908 599734 96960
rect 606202 96908 606208 96960
rect 606260 96948 606266 96960
rect 607122 96948 607128 96960
rect 606260 96920 607128 96948
rect 606260 96908 606266 96920
rect 607122 96908 607128 96920
rect 607180 96908 607186 96960
rect 615770 96908 615776 96960
rect 615828 96948 615834 96960
rect 616782 96948 616788 96960
rect 615828 96920 616788 96948
rect 615828 96908 615834 96920
rect 616782 96908 616788 96920
rect 616840 96908 616846 96960
rect 612090 96840 612096 96892
rect 612148 96880 612154 96892
rect 612642 96880 612648 96892
rect 612148 96852 612648 96880
rect 612148 96840 612154 96852
rect 612642 96840 612648 96852
rect 612700 96840 612706 96892
rect 617242 96840 617248 96892
rect 617300 96880 617306 96892
rect 618162 96880 618168 96892
rect 617300 96852 618168 96880
rect 617300 96840 617306 96852
rect 618162 96840 618168 96852
rect 618220 96840 618226 96892
rect 632698 96840 632704 96892
rect 632756 96880 632762 96892
rect 648246 96880 648252 96892
rect 632756 96852 648252 96880
rect 632756 96840 632762 96852
rect 648246 96840 648252 96852
rect 648304 96840 648310 96892
rect 653950 96840 653956 96892
rect 654008 96880 654014 96892
rect 654594 96880 654600 96892
rect 654008 96852 654600 96880
rect 654008 96840 654014 96852
rect 654594 96840 654600 96852
rect 654652 96840 654658 96892
rect 654778 96840 654784 96892
rect 654836 96880 654842 96892
rect 655422 96880 655428 96892
rect 654836 96852 655428 96880
rect 654836 96840 654842 96852
rect 655422 96840 655428 96852
rect 655480 96840 655486 96892
rect 656544 96812 656572 97124
rect 656682 97084 656710 97260
rect 656802 97180 656808 97232
rect 656860 97220 656866 97232
rect 661402 97220 661408 97232
rect 656860 97192 661408 97220
rect 656860 97180 656866 97192
rect 661402 97180 661408 97192
rect 661460 97180 661466 97232
rect 658826 97084 658832 97096
rect 656682 97056 658832 97084
rect 658826 97044 658832 97056
rect 658884 97044 658890 97096
rect 656710 96908 656716 96960
rect 656768 96948 656774 96960
rect 660114 96948 660120 96960
rect 656768 96920 660120 96948
rect 656768 96908 656774 96920
rect 660114 96908 660120 96920
rect 660172 96908 660178 96960
rect 660114 96812 660120 96824
rect 656544 96784 660120 96812
rect 660114 96772 660120 96784
rect 660172 96772 660178 96824
rect 610618 96704 610624 96756
rect 610676 96744 610682 96756
rect 611262 96744 611268 96756
rect 610676 96716 611268 96744
rect 610676 96704 610682 96716
rect 611262 96704 611268 96716
rect 611320 96704 611326 96756
rect 647878 96744 647884 96756
rect 645596 96716 647884 96744
rect 640518 96568 640524 96620
rect 640576 96608 640582 96620
rect 645596 96608 645624 96716
rect 647878 96704 647884 96716
rect 647936 96704 647942 96756
rect 640576 96580 645624 96608
rect 640576 96568 640582 96580
rect 645762 96568 645768 96620
rect 645820 96608 645826 96620
rect 656342 96608 656348 96620
rect 645820 96580 656348 96608
rect 645820 96568 645826 96580
rect 656342 96568 656348 96580
rect 656400 96568 656406 96620
rect 639046 96432 639052 96484
rect 639104 96472 639110 96484
rect 645118 96472 645124 96484
rect 639104 96444 645124 96472
rect 639104 96432 639110 96444
rect 645118 96432 645124 96444
rect 645176 96432 645182 96484
rect 646406 96432 646412 96484
rect 646464 96472 646470 96484
rect 652018 96472 652024 96484
rect 646464 96444 652024 96472
rect 646464 96432 646470 96444
rect 652018 96432 652024 96444
rect 652076 96432 652082 96484
rect 652570 96432 652576 96484
rect 652628 96472 652634 96484
rect 665542 96472 665548 96484
rect 652628 96444 665548 96472
rect 652628 96432 652634 96444
rect 665542 96432 665548 96444
rect 665600 96432 665606 96484
rect 631226 96296 631232 96348
rect 631284 96336 631290 96348
rect 647142 96336 647148 96348
rect 631284 96308 647148 96336
rect 631284 96296 631290 96308
rect 647142 96296 647148 96308
rect 647200 96296 647206 96348
rect 648890 96296 648896 96348
rect 648948 96336 648954 96348
rect 664162 96336 664168 96348
rect 648948 96308 664168 96336
rect 648948 96296 648954 96308
rect 664162 96296 664168 96308
rect 664220 96296 664226 96348
rect 637574 96160 637580 96212
rect 637632 96200 637638 96212
rect 660666 96200 660672 96212
rect 637632 96172 660672 96200
rect 637632 96160 637638 96172
rect 660666 96160 660672 96172
rect 660724 96160 660730 96212
rect 611078 96024 611084 96076
rect 611136 96064 611142 96076
rect 622118 96064 622124 96076
rect 611136 96036 622124 96064
rect 611136 96024 611142 96036
rect 622118 96024 622124 96036
rect 622176 96024 622182 96076
rect 649902 96024 649908 96076
rect 649960 96064 649966 96076
rect 663702 96064 663708 96076
rect 649960 96036 663708 96064
rect 649960 96024 649966 96036
rect 663702 96024 663708 96036
rect 663760 96024 663766 96076
rect 644934 95956 644940 96008
rect 644992 95996 644998 96008
rect 649074 95996 649080 96008
rect 644992 95968 649080 95996
rect 644992 95956 644998 95968
rect 649074 95956 649080 95968
rect 649132 95956 649138 96008
rect 607674 95888 607680 95940
rect 607732 95928 607738 95940
rect 624970 95928 624976 95940
rect 607732 95900 624976 95928
rect 607732 95888 607738 95900
rect 624970 95888 624976 95900
rect 625028 95888 625034 95940
rect 665358 95928 665364 95940
rect 656866 95900 665364 95928
rect 643462 95820 643468 95872
rect 643520 95860 643526 95872
rect 649258 95860 649264 95872
rect 643520 95832 649264 95860
rect 643520 95820 643526 95832
rect 649258 95820 649264 95832
rect 649316 95820 649322 95872
rect 656866 95860 656894 95900
rect 665358 95888 665364 95900
rect 665416 95888 665422 95940
rect 649460 95832 656894 95860
rect 638586 95684 638592 95736
rect 638644 95724 638650 95736
rect 647326 95724 647332 95736
rect 638644 95696 647332 95724
rect 638644 95684 638650 95696
rect 647326 95684 647332 95696
rect 647384 95684 647390 95736
rect 647878 95684 647884 95736
rect 647936 95724 647942 95736
rect 649460 95724 649488 95832
rect 647936 95696 649488 95724
rect 647936 95684 647942 95696
rect 653306 95616 653312 95668
rect 653364 95656 653370 95668
rect 664346 95656 664352 95668
rect 653364 95628 664352 95656
rect 653364 95616 653370 95628
rect 664346 95616 664352 95628
rect 664404 95616 664410 95668
rect 640058 95548 640064 95600
rect 640116 95588 640122 95600
rect 647878 95588 647884 95600
rect 640116 95560 647884 95588
rect 640116 95548 640122 95560
rect 647878 95548 647884 95560
rect 647936 95548 647942 95600
rect 641530 95412 641536 95464
rect 641588 95412 641594 95464
rect 645118 95412 645124 95464
rect 645176 95452 645182 95464
rect 651834 95452 651840 95464
rect 645176 95424 651840 95452
rect 645176 95412 645182 95424
rect 651834 95412 651840 95424
rect 651892 95412 651898 95464
rect 641548 95316 641576 95412
rect 649902 95316 649908 95328
rect 641548 95288 649908 95316
rect 649902 95276 649908 95288
rect 649960 95276 649966 95328
rect 620922 95140 620928 95192
rect 620980 95180 620986 95192
rect 626442 95180 626448 95192
rect 620980 95152 626448 95180
rect 620980 95140 620986 95152
rect 626442 95140 626448 95152
rect 626500 95140 626506 95192
rect 647694 95140 647700 95192
rect 647752 95180 647758 95192
rect 648798 95180 648804 95192
rect 647752 95152 648804 95180
rect 647752 95140 647758 95152
rect 648798 95140 648804 95152
rect 648856 95140 648862 95192
rect 579522 95004 579528 95056
rect 579580 95044 579586 95056
rect 583202 95044 583208 95056
rect 579580 95016 583208 95044
rect 579580 95004 579586 95016
rect 583202 95004 583208 95016
rect 583260 95004 583266 95056
rect 616506 95004 616512 95056
rect 616564 95044 616570 95056
rect 623038 95044 623044 95056
rect 616564 95016 623044 95044
rect 616564 95004 616570 95016
rect 623038 95004 623044 95016
rect 623096 95004 623102 95056
rect 609146 94460 609152 94512
rect 609204 94500 609210 94512
rect 620278 94500 620284 94512
rect 609204 94472 620284 94500
rect 609204 94460 609210 94472
rect 620278 94460 620284 94472
rect 620336 94460 620342 94512
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626442 93820 626448 93832
rect 619600 93792 626448 93820
rect 619600 93780 619606 93792
rect 626442 93780 626448 93792
rect 626500 93780 626506 93832
rect 651282 93508 651288 93560
rect 651340 93548 651346 93560
rect 655422 93548 655428 93560
rect 651340 93520 655428 93548
rect 651340 93508 651346 93520
rect 655422 93508 655428 93520
rect 655480 93508 655486 93560
rect 578510 93440 578516 93492
rect 578568 93480 578574 93492
rect 585962 93480 585968 93492
rect 578568 93452 585968 93480
rect 578568 93440 578574 93452
rect 585962 93440 585968 93452
rect 586020 93440 586026 93492
rect 649074 93236 649080 93288
rect 649132 93276 649138 93288
rect 656158 93276 656164 93288
rect 649132 93248 656164 93276
rect 649132 93236 649138 93248
rect 656158 93236 656164 93248
rect 656216 93236 656222 93288
rect 611262 93100 611268 93152
rect 611320 93140 611326 93152
rect 619266 93140 619272 93152
rect 611320 93112 619272 93140
rect 611320 93100 611326 93112
rect 619266 93100 619272 93112
rect 619324 93100 619330 93152
rect 606938 92828 606944 92880
rect 606996 92868 607002 92880
rect 610066 92868 610072 92880
rect 606996 92840 610072 92868
rect 606996 92828 607002 92840
rect 610066 92828 610072 92840
rect 610124 92828 610130 92880
rect 648614 92488 648620 92540
rect 648672 92528 648678 92540
rect 649994 92528 650000 92540
rect 648672 92500 650000 92528
rect 648672 92488 648678 92500
rect 649994 92488 650000 92500
rect 650052 92488 650058 92540
rect 617978 92420 617984 92472
rect 618036 92460 618042 92472
rect 626442 92460 626448 92472
rect 618036 92432 626448 92460
rect 618036 92420 618042 92432
rect 626442 92420 626448 92432
rect 626500 92420 626506 92472
rect 647326 92352 647332 92404
rect 647384 92392 647390 92404
rect 654318 92392 654324 92404
rect 647384 92364 654324 92392
rect 647384 92352 647390 92364
rect 654318 92352 654324 92364
rect 654376 92352 654382 92404
rect 579338 91060 579344 91112
rect 579396 91100 579402 91112
rect 584582 91100 584588 91112
rect 579396 91072 584588 91100
rect 579396 91060 579402 91072
rect 584582 91060 584588 91072
rect 584640 91060 584646 91112
rect 618162 90992 618168 91044
rect 618220 91032 618226 91044
rect 626442 91032 626448 91044
rect 618220 91004 626448 91032
rect 618220 90992 618226 91004
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 651834 90652 651840 90704
rect 651892 90692 651898 90704
rect 655422 90692 655428 90704
rect 651892 90664 655428 90692
rect 651892 90652 651898 90664
rect 655422 90652 655428 90664
rect 655480 90652 655486 90704
rect 623038 89632 623044 89684
rect 623096 89672 623102 89684
rect 623096 89644 625154 89672
rect 623096 89632 623102 89644
rect 625126 89604 625154 89644
rect 626442 89604 626448 89616
rect 625126 89576 626448 89604
rect 626442 89564 626448 89576
rect 626500 89564 626506 89616
rect 585134 88952 585140 89004
rect 585192 88992 585198 89004
rect 589918 88992 589924 89004
rect 585192 88964 589924 88992
rect 585192 88952 585198 88964
rect 589918 88952 589924 88964
rect 589976 88952 589982 89004
rect 649718 88748 649724 88800
rect 649776 88788 649782 88800
rect 658550 88788 658556 88800
rect 649776 88760 658556 88788
rect 649776 88748 649782 88760
rect 658550 88748 658556 88760
rect 658608 88748 658614 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 663886 88788 663892 88800
rect 662380 88760 663892 88788
rect 662380 88748 662386 88760
rect 663886 88748 663892 88760
rect 663944 88748 663950 88800
rect 656342 88612 656348 88664
rect 656400 88652 656406 88664
rect 657446 88652 657452 88664
rect 656400 88624 657452 88652
rect 656400 88612 656406 88624
rect 657446 88612 657452 88624
rect 657504 88612 657510 88664
rect 610066 88272 610072 88324
rect 610124 88312 610130 88324
rect 626442 88312 626448 88324
rect 610124 88284 626448 88312
rect 610124 88272 610130 88284
rect 626442 88272 626448 88284
rect 626500 88272 626506 88324
rect 655238 88272 655244 88324
rect 655296 88312 655302 88324
rect 658458 88312 658464 88324
rect 655296 88284 658464 88312
rect 655296 88272 655302 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 622118 88136 622124 88188
rect 622176 88176 622182 88188
rect 626258 88176 626264 88188
rect 622176 88148 626264 88176
rect 622176 88136 622182 88148
rect 626258 88136 626264 88148
rect 626316 88136 626322 88188
rect 579522 88068 579528 88120
rect 579580 88108 579586 88120
rect 585134 88108 585140 88120
rect 579580 88080 585140 88108
rect 579580 88068 579586 88080
rect 585134 88068 585140 88080
rect 585192 88068 585198 88120
rect 648430 86980 648436 87032
rect 648488 87020 648494 87032
rect 662506 87020 662512 87032
rect 648488 86992 662512 87020
rect 648488 86980 648494 86992
rect 662506 86980 662512 86992
rect 662564 86980 662570 87032
rect 656710 86844 656716 86896
rect 656768 86884 656774 86896
rect 659562 86884 659568 86896
rect 656768 86856 659568 86884
rect 656768 86844 656774 86856
rect 659562 86844 659568 86856
rect 659620 86844 659626 86896
rect 649258 86708 649264 86760
rect 649316 86748 649322 86760
rect 661402 86748 661408 86760
rect 649316 86720 661408 86748
rect 649316 86708 649322 86720
rect 661402 86708 661408 86720
rect 661460 86708 661466 86760
rect 647878 86572 647884 86624
rect 647936 86612 647942 86624
rect 660114 86612 660120 86624
rect 647936 86584 660120 86612
rect 647936 86572 647942 86584
rect 660114 86572 660120 86584
rect 660172 86572 660178 86624
rect 656158 86436 656164 86488
rect 656216 86476 656222 86488
rect 660666 86476 660672 86488
rect 656216 86448 660672 86476
rect 656216 86436 656222 86448
rect 660666 86436 660672 86448
rect 660724 86436 660730 86488
rect 619266 86300 619272 86352
rect 619324 86340 619330 86352
rect 626442 86340 626448 86352
rect 619324 86312 626448 86340
rect 619324 86300 619330 86312
rect 626442 86300 626448 86312
rect 626500 86300 626506 86352
rect 652018 86300 652024 86352
rect 652076 86340 652082 86352
rect 657170 86340 657176 86352
rect 652076 86312 657176 86340
rect 652076 86300 652082 86312
rect 657170 86300 657176 86312
rect 657228 86300 657234 86352
rect 620278 85484 620284 85536
rect 620336 85524 620342 85536
rect 626442 85524 626448 85536
rect 620336 85496 626448 85524
rect 620336 85484 620342 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 609882 85348 609888 85400
rect 609940 85388 609946 85400
rect 609940 85360 625154 85388
rect 609940 85348 609946 85360
rect 625126 85320 625154 85360
rect 625338 85320 625344 85332
rect 625126 85292 625344 85320
rect 625338 85280 625344 85292
rect 625396 85280 625402 85332
rect 579154 84124 579160 84176
rect 579212 84164 579218 84176
rect 581638 84164 581644 84176
rect 579212 84136 581644 84164
rect 579212 84124 579218 84136
rect 581638 84124 581644 84136
rect 581696 84124 581702 84176
rect 608502 84124 608508 84176
rect 608560 84164 608566 84176
rect 625798 84164 625804 84176
rect 608560 84136 625804 84164
rect 608560 84124 608566 84136
rect 625798 84124 625804 84136
rect 625856 84124 625862 84176
rect 579062 82356 579068 82408
rect 579120 82396 579126 82408
rect 583018 82396 583024 82408
rect 579120 82368 583024 82396
rect 579120 82356 579126 82368
rect 583018 82356 583024 82368
rect 583076 82356 583082 82408
rect 579522 82084 579528 82136
rect 579580 82124 579586 82136
rect 587158 82124 587164 82136
rect 579580 82096 587164 82124
rect 579580 82084 579586 82096
rect 587158 82084 587164 82096
rect 587216 82084 587222 82136
rect 628742 80928 628748 80980
rect 628800 80968 628806 80980
rect 642450 80968 642456 80980
rect 628800 80940 642456 80968
rect 628800 80928 628806 80940
rect 642450 80928 642456 80940
rect 642508 80928 642514 80980
rect 612642 80792 612648 80844
rect 612700 80832 612706 80844
rect 647418 80832 647424 80844
rect 612700 80804 647424 80832
rect 612700 80792 612706 80804
rect 647418 80792 647424 80804
rect 647476 80792 647482 80844
rect 595438 80656 595444 80708
rect 595496 80696 595502 80708
rect 636746 80696 636752 80708
rect 595496 80668 636752 80696
rect 595496 80656 595502 80668
rect 636746 80656 636752 80668
rect 636804 80656 636810 80708
rect 629202 79976 629208 80028
rect 629260 80016 629266 80028
rect 633434 80016 633440 80028
rect 629260 79988 633440 80016
rect 629260 79976 629266 79988
rect 633434 79976 633440 79988
rect 633492 79976 633498 80028
rect 613746 79432 613752 79484
rect 613804 79472 613810 79484
rect 645946 79472 645952 79484
rect 613804 79444 645952 79472
rect 613804 79432 613810 79444
rect 645946 79432 645952 79444
rect 646004 79432 646010 79484
rect 579062 79296 579068 79348
rect 579120 79336 579126 79348
rect 588722 79336 588728 79348
rect 579120 79308 588728 79336
rect 579120 79296 579126 79308
rect 588722 79296 588728 79308
rect 588780 79296 588786 79348
rect 613930 79296 613936 79348
rect 613988 79336 613994 79348
rect 646498 79336 646504 79348
rect 613988 79308 646504 79336
rect 613988 79296 613994 79308
rect 646498 79296 646504 79308
rect 646556 79296 646562 79348
rect 633434 78072 633440 78124
rect 633492 78112 633498 78124
rect 645302 78112 645308 78124
rect 633492 78084 645308 78112
rect 633492 78072 633498 78084
rect 645302 78072 645308 78084
rect 645360 78072 645366 78124
rect 631042 77936 631048 77988
rect 631100 77976 631106 77988
rect 643094 77976 643100 77988
rect 631100 77948 643100 77976
rect 631100 77936 631106 77948
rect 643094 77936 643100 77948
rect 643152 77936 643158 77988
rect 628466 77732 628472 77784
rect 628524 77772 628530 77784
rect 632790 77772 632796 77784
rect 628524 77744 632796 77772
rect 628524 77732 628530 77744
rect 632790 77732 632796 77744
rect 632848 77732 632854 77784
rect 625798 77256 625804 77308
rect 625856 77296 625862 77308
rect 631042 77296 631048 77308
rect 625856 77268 631048 77296
rect 625856 77256 625862 77268
rect 631042 77256 631048 77268
rect 631100 77256 631106 77308
rect 616782 76644 616788 76696
rect 616840 76684 616846 76696
rect 646314 76684 646320 76696
rect 616840 76656 646320 76684
rect 616840 76644 616846 76656
rect 646314 76644 646320 76656
rect 646372 76644 646378 76696
rect 611998 76508 612004 76560
rect 612056 76548 612062 76560
rect 662414 76548 662420 76560
rect 612056 76520 662420 76548
rect 612056 76508 612062 76520
rect 662414 76508 662420 76520
rect 662472 76508 662478 76560
rect 578234 75828 578240 75880
rect 578292 75868 578298 75880
rect 580258 75868 580264 75880
rect 578292 75840 580264 75868
rect 578292 75828 578298 75840
rect 580258 75828 580264 75840
rect 580316 75828 580322 75880
rect 618898 75420 618904 75472
rect 618956 75460 618962 75472
rect 648614 75460 648620 75472
rect 618956 75432 648620 75460
rect 618956 75420 618962 75432
rect 648614 75420 648620 75432
rect 648672 75420 648678 75472
rect 615402 75284 615408 75336
rect 615460 75324 615466 75336
rect 646866 75324 646872 75336
rect 615460 75296 646872 75324
rect 615460 75284 615466 75296
rect 646866 75284 646872 75296
rect 646924 75284 646930 75336
rect 607122 75148 607128 75200
rect 607180 75188 607186 75200
rect 646130 75188 646136 75200
rect 607180 75160 646136 75188
rect 607180 75148 607186 75160
rect 646130 75148 646136 75160
rect 646188 75148 646194 75200
rect 578878 72428 578884 72480
rect 578936 72468 578942 72480
rect 601694 72468 601700 72480
rect 578936 72440 601700 72468
rect 578936 72428 578942 72440
rect 601694 72428 601700 72440
rect 601752 72428 601758 72480
rect 579062 71340 579068 71392
rect 579120 71380 579126 71392
rect 584398 71380 584404 71392
rect 579120 71352 584404 71380
rect 579120 71340 579126 71352
rect 584398 71340 584404 71352
rect 584456 71340 584462 71392
rect 580258 68280 580264 68332
rect 580316 68320 580322 68332
rect 604454 68320 604460 68332
rect 580316 68292 604460 68320
rect 580316 68280 580322 68292
rect 604454 68280 604460 68292
rect 604512 68280 604518 68332
rect 577498 59984 577504 60036
rect 577556 60024 577562 60036
rect 603074 60024 603080 60036
rect 577556 59996 603080 60024
rect 577556 59984 577562 59996
rect 603074 59984 603080 59996
rect 603132 59984 603138 60036
rect 576118 58624 576124 58676
rect 576176 58664 576182 58676
rect 601878 58664 601884 58676
rect 576176 58636 601884 58664
rect 576176 58624 576182 58636
rect 601878 58624 601884 58636
rect 601936 58624 601942 58676
rect 574922 57196 574928 57248
rect 574980 57236 574986 57248
rect 600498 57236 600504 57248
rect 574980 57208 600504 57236
rect 574980 57196 574986 57208
rect 600498 57196 600504 57208
rect 600556 57196 600562 57248
rect 574554 55972 574560 56024
rect 574612 56012 574618 56024
rect 598934 56012 598940 56024
rect 574612 55984 598940 56012
rect 574612 55972 574618 55984
rect 598934 55972 598940 55984
rect 598992 55972 598998 56024
rect 574738 55836 574744 55888
rect 574796 55876 574802 55888
rect 600314 55876 600320 55888
rect 574796 55848 600320 55876
rect 574796 55836 574802 55848
rect 600314 55836 600320 55848
rect 600372 55836 600378 55888
rect 463298 55372 471974 55400
rect 463298 53644 463326 55372
rect 464172 55236 470732 55264
rect 464172 53768 464200 55236
rect 470704 55060 470732 55236
rect 471946 55196 471974 55372
rect 596450 55196 596456 55208
rect 471946 55168 596456 55196
rect 596450 55156 596456 55168
rect 596508 55156 596514 55208
rect 597646 55060 597652 55072
rect 470704 55032 597652 55060
rect 597646 55020 597652 55032
rect 597704 55020 597710 55072
rect 597922 54924 597928 54936
rect 464632 54896 597928 54924
rect 464632 53904 464660 54896
rect 597922 54884 597928 54896
rect 597980 54884 597986 54936
rect 599118 54788 599124 54800
rect 464080 53740 464200 53768
rect 464264 53876 464660 53904
rect 464816 54760 599124 54788
rect 464080 53644 464108 53740
rect 464264 53644 464292 53876
rect 463234 53592 463240 53644
rect 463292 53604 463326 53644
rect 463292 53592 463298 53604
rect 464062 53592 464068 53644
rect 464120 53592 464126 53644
rect 464246 53592 464252 53644
rect 464304 53592 464310 53644
rect 459462 53456 459468 53508
rect 459520 53496 459526 53508
rect 464816 53496 464844 54760
rect 599118 54748 599124 54760
rect 599176 54748 599182 54800
rect 624418 54652 624424 54664
rect 465368 54624 470364 54652
rect 465368 53768 465396 54624
rect 470336 54584 470364 54624
rect 470796 54624 624424 54652
rect 470796 54584 470824 54624
rect 624418 54612 624424 54624
rect 624476 54612 624482 54664
rect 470336 54556 470824 54584
rect 625798 54516 625804 54528
rect 470888 54488 625804 54516
rect 470888 54448 470916 54488
rect 625798 54476 625804 54488
rect 625856 54476 625862 54528
rect 465276 53740 465396 53768
rect 465460 54420 470916 54448
rect 465276 53644 465304 53740
rect 465460 53644 465488 54420
rect 596174 54380 596180 54392
rect 470980 54352 596180 54380
rect 470980 54312 471008 54352
rect 596174 54340 596180 54352
rect 596232 54340 596238 54392
rect 465828 54284 471008 54312
rect 465258 53592 465264 53644
rect 465316 53592 465322 53644
rect 465442 53592 465448 53644
rect 465500 53592 465506 53644
rect 459520 53468 464844 53496
rect 459520 53456 459526 53468
rect 464982 53456 464988 53508
rect 465040 53496 465046 53508
rect 465828 53496 465856 54284
rect 581638 54244 581644 54256
rect 471164 54216 581644 54244
rect 471164 54176 471192 54216
rect 581638 54204 581644 54216
rect 581696 54204 581702 54256
rect 471072 54148 471192 54176
rect 471072 54040 471100 54148
rect 574738 54108 574744 54120
rect 467024 54012 471100 54040
rect 471348 54080 574744 54108
rect 467024 53768 467052 54012
rect 471348 53836 471376 54080
rect 574738 54068 574744 54080
rect 574796 54068 574802 54120
rect 574554 53972 574560 53984
rect 466380 53740 467052 53768
rect 467116 53808 471376 53836
rect 471946 53944 574560 53972
rect 466380 53644 466408 53740
rect 467116 53644 467144 53808
rect 466362 53592 466368 53644
rect 466420 53592 466426 53644
rect 467098 53592 467104 53644
rect 467156 53592 467162 53644
rect 471054 53592 471060 53644
rect 471112 53632 471118 53644
rect 471946 53632 471974 53944
rect 574554 53932 574560 53944
rect 574612 53932 574618 53984
rect 574922 53836 574928 53848
rect 471112 53604 471974 53632
rect 473326 53808 574928 53836
rect 471112 53592 471118 53604
rect 465040 53468 465856 53496
rect 465040 53456 465046 53468
rect 463050 53320 463056 53372
rect 463108 53360 463114 53372
rect 473326 53360 473354 53808
rect 574922 53796 574928 53808
rect 574980 53796 574986 53848
rect 463108 53332 473354 53360
rect 463108 53320 463114 53332
rect 50522 53184 50528 53236
rect 50580 53224 50586 53236
rect 130378 53224 130384 53236
rect 50580 53196 130384 53224
rect 50580 53184 50586 53196
rect 130378 53184 130384 53196
rect 130436 53184 130442 53236
rect 463234 53184 463240 53236
rect 463292 53224 463298 53236
rect 463786 53224 463792 53236
rect 463292 53196 463792 53224
rect 463292 53184 463298 53196
rect 463786 53184 463792 53196
rect 463844 53184 463850 53236
rect 312354 53116 312360 53168
rect 312412 53156 312418 53168
rect 313734 53156 313740 53168
rect 312412 53128 313740 53156
rect 312412 53116 312418 53128
rect 313734 53116 313740 53128
rect 313792 53116 313798 53168
rect 316310 53116 316316 53168
rect 316368 53156 316374 53168
rect 317690 53156 317696 53168
rect 316368 53128 317696 53156
rect 316368 53116 316374 53128
rect 317690 53116 317696 53128
rect 317748 53116 317754 53168
rect 48958 53048 48964 53100
rect 49016 53088 49022 53100
rect 130562 53088 130568 53100
rect 49016 53060 130568 53088
rect 49016 53048 49022 53060
rect 130562 53048 130568 53060
rect 130620 53048 130626 53100
rect 463602 53048 463608 53100
rect 463660 53088 463666 53100
rect 464246 53088 464252 53100
rect 463660 53060 464252 53088
rect 463660 53048 463666 53060
rect 464246 53048 464252 53060
rect 464304 53048 464310 53100
rect 465442 53048 465448 53100
rect 465500 53088 465506 53100
rect 466362 53088 466368 53100
rect 465500 53060 466368 53088
rect 465500 53048 465506 53060
rect 466362 53048 466368 53060
rect 466420 53048 466426 53100
rect 461302 52912 461308 52964
rect 461360 52952 461366 52964
rect 471054 52952 471060 52964
rect 461360 52924 471060 52952
rect 461360 52912 461366 52924
rect 471054 52912 471060 52924
rect 471112 52912 471118 52964
rect 461900 52776 461906 52828
rect 461958 52816 461964 52828
rect 467098 52816 467104 52828
rect 461958 52788 467104 52816
rect 461958 52776 461964 52788
rect 467098 52776 467104 52788
rect 467156 52776 467162 52828
rect 47578 51960 47584 52012
rect 47636 52000 47642 52012
rect 130746 52000 130752 52012
rect 47636 51972 130752 52000
rect 47636 51960 47642 51972
rect 130746 51960 130752 51972
rect 130804 51960 130810 52012
rect 50338 51824 50344 51876
rect 50396 51864 50402 51876
rect 128998 51864 129004 51876
rect 50396 51836 129004 51864
rect 50396 51824 50402 51836
rect 128998 51824 129004 51836
rect 129056 51824 129062 51876
rect 129642 51824 129648 51876
rect 129700 51864 129706 51876
rect 591298 51864 591304 51876
rect 129700 51836 591304 51864
rect 129700 51824 129706 51836
rect 591298 51824 591304 51836
rect 591356 51824 591362 51876
rect 128814 51688 128820 51740
rect 128872 51728 128878 51740
rect 592678 51728 592684 51740
rect 128872 51700 592684 51728
rect 128872 51688 128878 51700
rect 592678 51688 592684 51700
rect 592736 51688 592742 51740
rect 318334 50464 318340 50516
rect 318392 50504 318398 50516
rect 458174 50504 458180 50516
rect 318392 50476 458180 50504
rect 318392 50464 318398 50476
rect 458174 50464 458180 50476
rect 458232 50464 458238 50516
rect 46198 50328 46204 50380
rect 46256 50368 46262 50380
rect 131022 50368 131028 50380
rect 46256 50340 131028 50368
rect 46256 50328 46262 50340
rect 131022 50328 131028 50340
rect 131080 50328 131086 50380
rect 314010 50328 314016 50380
rect 314068 50368 314074 50380
rect 458358 50368 458364 50380
rect 314068 50340 458364 50368
rect 314068 50328 314074 50340
rect 458358 50328 458364 50340
rect 458416 50328 458422 50380
rect 522942 50328 522948 50380
rect 523000 50368 523006 50380
rect 544010 50368 544016 50380
rect 523000 50340 544016 50368
rect 523000 50328 523006 50340
rect 544010 50328 544016 50340
rect 544068 50328 544074 50380
rect 49142 49104 49148 49156
rect 49200 49144 49206 49156
rect 129274 49144 129280 49156
rect 49200 49116 129280 49144
rect 49200 49104 49206 49116
rect 129274 49104 129280 49116
rect 129332 49104 129338 49156
rect 45462 48968 45468 49020
rect 45520 49008 45526 49020
rect 129458 49008 129464 49020
rect 45520 48980 129464 49008
rect 45520 48968 45526 48980
rect 129458 48968 129464 48980
rect 129516 48968 129522 49020
rect 130562 46044 130568 46096
rect 130620 46084 130626 46096
rect 132310 46084 132316 46096
rect 130620 46056 132316 46084
rect 130620 46044 130626 46056
rect 132310 46044 132316 46056
rect 132368 46044 132374 46096
rect 130746 45500 130752 45552
rect 130804 45540 130810 45552
rect 132586 45540 132592 45552
rect 130804 45512 132592 45540
rect 130804 45500 130810 45512
rect 132586 45500 132592 45512
rect 132644 45500 132650 45552
rect 129458 45364 129464 45416
rect 129516 45404 129522 45416
rect 129516 45376 131390 45404
rect 129516 45364 129522 45376
rect 131362 45090 131390 45376
rect 129642 45024 129648 45076
rect 129700 45064 129706 45076
rect 129700 45036 131068 45064
rect 129700 45024 129706 45036
rect 131040 45020 131068 45036
rect 131040 44992 131330 45020
rect 129274 44888 129280 44940
rect 129332 44928 129338 44940
rect 131224 44928 131606 44936
rect 129332 44908 131606 44928
rect 129332 44900 131252 44908
rect 129332 44888 129338 44900
rect 131592 44824 131790 44852
rect 128814 44752 128820 44804
rect 128872 44792 128878 44804
rect 131592 44792 131620 44824
rect 128872 44764 131620 44792
rect 128872 44752 128878 44764
rect 131684 44740 131974 44768
rect 131684 44668 131712 44740
rect 131666 44616 131672 44668
rect 131724 44616 131730 44668
rect 128998 44412 129004 44464
rect 129056 44452 129062 44464
rect 132144 44452 132172 44670
rect 132374 44452 132402 44586
rect 129056 44424 132172 44452
rect 132236 44424 132402 44452
rect 132466 44488 132526 44516
rect 129056 44412 129062 44424
rect 43622 44276 43628 44328
rect 43680 44316 43686 44328
rect 132236 44316 132264 44424
rect 43680 44288 132264 44316
rect 132466 44316 132494 44488
rect 132586 44364 132592 44416
rect 132644 44404 132650 44416
rect 132644 44376 132756 44404
rect 132644 44364 132650 44376
rect 132466 44304 132540 44316
rect 132466 44288 132500 44304
rect 43680 44276 43686 44288
rect 132494 44252 132500 44288
rect 132552 44252 132558 44304
rect 132770 44252 132776 44304
rect 132828 44292 132834 44304
rect 132828 44264 132986 44292
rect 132828 44252 132834 44264
rect 43438 44140 43444 44192
rect 43496 44180 43502 44192
rect 131666 44180 131672 44192
rect 43496 44152 131672 44180
rect 43496 44140 43502 44152
rect 131666 44140 131672 44152
rect 131724 44140 131730 44192
rect 132144 44152 133170 44180
rect 131022 44004 131028 44056
rect 131080 44044 131086 44056
rect 132144 44044 132172 44152
rect 131080 44016 132172 44044
rect 131080 44004 131086 44016
rect 440234 43800 440240 43852
rect 440292 43840 440298 43852
rect 441062 43840 441068 43852
rect 440292 43812 441068 43840
rect 440292 43800 440298 43812
rect 441062 43800 441068 43812
rect 441120 43800 441126 43852
rect 187326 42780 187332 42832
rect 187384 42820 187390 42832
rect 255866 42820 255872 42832
rect 187384 42792 255872 42820
rect 187384 42780 187390 42792
rect 255866 42780 255872 42792
rect 255924 42780 255930 42832
rect 307294 42712 307300 42764
rect 307352 42752 307358 42764
rect 431218 42752 431224 42764
rect 307352 42724 431224 42752
rect 307352 42712 307358 42724
rect 431218 42712 431224 42724
rect 431276 42712 431282 42764
rect 441062 42712 441068 42764
rect 441120 42752 441126 42764
rect 449158 42752 449164 42764
rect 441120 42724 449164 42752
rect 441120 42712 441126 42724
rect 449158 42712 449164 42724
rect 449216 42712 449222 42764
rect 453574 42712 453580 42764
rect 453632 42752 453638 42764
rect 464154 42752 464160 42764
rect 453632 42724 464160 42752
rect 453632 42712 453638 42724
rect 464154 42712 464160 42724
rect 464212 42712 464218 42764
rect 310422 42576 310428 42628
rect 310480 42616 310486 42628
rect 427078 42616 427084 42628
rect 310480 42588 427084 42616
rect 310480 42576 310486 42588
rect 427078 42576 427084 42588
rect 427136 42576 427142 42628
rect 441246 42576 441252 42628
rect 441304 42616 441310 42628
rect 446398 42616 446404 42628
rect 441304 42588 446404 42616
rect 441304 42576 441310 42588
rect 446398 42576 446404 42588
rect 446456 42576 446462 42628
rect 454494 42440 454500 42492
rect 454552 42480 454558 42492
rect 463050 42480 463056 42492
rect 454552 42452 463056 42480
rect 454552 42440 454558 42452
rect 463050 42440 463056 42452
rect 463108 42440 463114 42492
rect 404446 42304 404452 42356
rect 404504 42344 404510 42356
rect 405182 42344 405188 42356
rect 404504 42316 405188 42344
rect 404504 42304 404510 42316
rect 405182 42304 405188 42316
rect 405240 42304 405246 42356
rect 420730 42304 420736 42356
rect 420788 42344 420794 42356
rect 426894 42344 426900 42356
rect 420788 42316 426900 42344
rect 420788 42304 420794 42316
rect 426894 42304 426900 42316
rect 426952 42304 426958 42356
rect 661402 42129 661408 42181
rect 661460 42129 661466 42181
rect 427078 41964 427084 42016
rect 427136 42004 427142 42016
rect 427136 41976 427814 42004
rect 427136 41964 427142 41976
rect 427786 41868 427814 41976
rect 431218 41964 431224 42016
rect 431276 42004 431282 42016
rect 441062 42004 441068 42016
rect 431276 41976 441068 42004
rect 431276 41964 431282 41976
rect 441062 41964 441068 41976
rect 441120 41964 441126 42016
rect 446398 41964 446404 42016
rect 446456 42004 446462 42016
rect 454494 42004 454500 42016
rect 446456 41976 454500 42004
rect 446456 41964 446462 41976
rect 454494 41964 454500 41976
rect 454552 41964 454558 42016
rect 441246 41868 441252 41880
rect 427786 41840 441252 41868
rect 441246 41828 441252 41840
rect 441304 41828 441310 41880
rect 449158 41828 449164 41880
rect 449216 41868 449222 41880
rect 453574 41868 453580 41880
rect 449216 41840 453580 41868
rect 449216 41828 449222 41840
rect 453574 41828 453580 41840
rect 453632 41828 453638 41880
rect 404446 41420 404452 41472
rect 404504 41460 404510 41472
rect 420730 41460 420736 41472
rect 404504 41432 420736 41460
rect 404504 41420 404510 41432
rect 420730 41420 420736 41432
rect 420788 41420 420794 41472
rect 426894 41420 426900 41472
rect 426952 41460 426958 41472
rect 459186 41460 459192 41472
rect 426952 41432 459192 41460
rect 426952 41420 426958 41432
rect 459186 41420 459192 41432
rect 459244 41420 459250 41472
<< via1 >>
rect 652024 896996 652076 897048
rect 676036 897064 676088 897116
rect 654784 895772 654836 895824
rect 675852 895772 675904 895824
rect 672724 895636 672776 895688
rect 676036 895636 676088 895688
rect 671068 894412 671120 894464
rect 675852 894412 675904 894464
rect 671896 894276 671948 894328
rect 676036 894276 676088 894328
rect 672908 892984 672960 893036
rect 676036 892984 676088 893036
rect 672540 892848 672592 892900
rect 675852 892848 675904 892900
rect 675024 890332 675076 890384
rect 676036 890332 676088 890384
rect 676220 890128 676272 890180
rect 676864 890128 676916 890180
rect 674656 888904 674708 888956
rect 676036 888904 676088 888956
rect 676220 888700 676272 888752
rect 677048 888700 677100 888752
rect 674380 888496 674432 888548
rect 676036 888496 676088 888548
rect 674196 887272 674248 887324
rect 676036 887272 676088 887324
rect 670884 886864 670936 886916
rect 676036 886864 676088 886916
rect 673092 885640 673144 885692
rect 676036 885640 676088 885692
rect 653404 880472 653456 880524
rect 675392 880336 675444 880388
rect 675024 879588 675076 879640
rect 677048 879452 677100 879504
rect 675944 879316 675996 879368
rect 676864 879316 676916 879368
rect 674748 879180 674800 879232
rect 675760 879044 675812 879096
rect 678244 879044 678296 879096
rect 675208 878772 675260 878824
rect 675392 878772 675444 878824
rect 674932 878160 674984 878212
rect 676404 878568 676456 878620
rect 675944 878432 675996 878484
rect 675208 877752 675260 877804
rect 675484 877208 675536 877260
rect 674840 874148 674892 874200
rect 675300 874148 675352 874200
rect 674380 872108 674432 872160
rect 674840 872108 674892 872160
rect 657544 869388 657596 869440
rect 675024 869388 675076 869440
rect 651472 868844 651524 868896
rect 654784 868844 654836 868896
rect 674196 868708 674248 868760
rect 675300 868708 675352 868760
rect 654140 868028 654192 868080
rect 674840 868028 674892 868080
rect 651472 866600 651524 866652
rect 672724 866600 672776 866652
rect 651380 865172 651432 865224
rect 653404 865172 653456 865224
rect 651472 863812 651524 863864
rect 657544 863812 657596 863864
rect 651472 862452 651524 862504
rect 654140 862452 654192 862504
rect 35808 817096 35860 817148
rect 44824 817096 44876 817148
rect 35624 816960 35676 817012
rect 61384 816960 61436 817012
rect 35808 815736 35860 815788
rect 43076 815736 43128 815788
rect 35440 815600 35492 815652
rect 43444 815600 43496 815652
rect 35624 814376 35676 814428
rect 42892 814376 42944 814428
rect 35808 814240 35860 814292
rect 44180 814240 44232 814292
rect 41328 812812 41380 812864
rect 44456 812812 44508 812864
rect 40960 811384 41012 811436
rect 42616 811384 42668 811436
rect 40684 808596 40736 808648
rect 41788 808596 41840 808648
rect 41144 808052 41196 808104
rect 41604 808052 41656 808104
rect 43444 807916 43496 807968
rect 62948 807916 63000 807968
rect 41144 807304 41196 807356
rect 44640 807304 44692 807356
rect 41328 806080 41380 806132
rect 50344 806080 50396 806132
rect 41144 805944 41196 805996
rect 62672 805944 62724 805996
rect 34520 802544 34572 802596
rect 41788 802544 41840 802596
rect 32404 802408 32456 802460
rect 42708 802408 42760 802460
rect 33784 801184 33836 801236
rect 42616 801184 42668 801236
rect 31024 801048 31076 801100
rect 43444 801048 43496 801100
rect 42432 799076 42484 799128
rect 53104 799008 53156 799060
rect 43628 797648 43680 797700
rect 57244 797648 57296 797700
rect 44640 796288 44692 796340
rect 42432 795608 42484 795660
rect 43628 795608 43680 795660
rect 42248 794996 42300 795048
rect 42248 793772 42300 793824
rect 43168 793772 43220 793824
rect 42616 793500 42668 793552
rect 43444 793500 43496 793552
rect 653404 790780 653456 790832
rect 675392 790780 675444 790832
rect 53104 790712 53156 790764
rect 62212 790712 62264 790764
rect 42432 790576 42484 790628
rect 42156 790372 42208 790424
rect 42248 789760 42300 789812
rect 42248 789488 42300 789540
rect 57244 789148 57296 789200
rect 62120 789148 62172 789200
rect 62120 786632 62172 786684
rect 42524 785612 42576 785664
rect 44824 785136 44876 785188
rect 62120 785136 62172 785188
rect 670608 784252 670660 784304
rect 675116 784252 675168 784304
rect 669228 784116 669280 784168
rect 675392 784116 675444 784168
rect 673736 782620 673788 782672
rect 675116 782620 675168 782672
rect 669044 782484 669096 782536
rect 675300 782484 675352 782536
rect 655520 781056 655572 781108
rect 675024 781056 675076 781108
rect 673920 779968 673972 780020
rect 675116 779968 675168 780020
rect 655060 778336 655112 778388
rect 674932 778336 674984 778388
rect 651472 777588 651524 777640
rect 660304 777588 660356 777640
rect 670424 776976 670476 777028
rect 675300 776976 675352 777028
rect 672724 775616 672776 775668
rect 674932 775616 674984 775668
rect 651472 775548 651524 775600
rect 669964 775548 670016 775600
rect 651380 775276 651432 775328
rect 653404 775276 653456 775328
rect 35808 774188 35860 774240
rect 41696 774188 41748 774240
rect 42064 774188 42116 774240
rect 60004 774188 60056 774240
rect 651472 774120 651524 774172
rect 655520 774120 655572 774172
rect 651472 773780 651524 773832
rect 655060 773780 655112 773832
rect 671436 773372 671488 773424
rect 675300 773372 675352 773424
rect 35808 773304 35860 773356
rect 41696 773304 41748 773356
rect 35808 773100 35860 773152
rect 40776 773100 40828 773152
rect 35532 772964 35584 773016
rect 41696 772964 41748 773016
rect 42064 772964 42116 773016
rect 43168 772964 43220 773016
rect 35348 772828 35400 772880
rect 61384 772828 61436 772880
rect 41696 772692 41748 772744
rect 42064 772692 42116 772744
rect 35808 771808 35860 771860
rect 40224 771808 40276 771860
rect 35624 771536 35676 771588
rect 41052 771604 41104 771656
rect 35808 771400 35860 771452
rect 41696 771400 41748 771452
rect 42064 771400 42116 771452
rect 44180 771400 44232 771452
rect 35808 770448 35860 770500
rect 39856 770448 39908 770500
rect 35624 770176 35676 770228
rect 41512 770176 41564 770228
rect 35808 770040 35860 770092
rect 41696 770040 41748 770092
rect 42064 770040 42116 770092
rect 44548 770040 44600 770092
rect 35808 769156 35860 769208
rect 41696 768952 41748 769004
rect 35532 768816 35584 768868
rect 41236 768816 41288 768868
rect 35808 768680 35860 768732
rect 40040 768680 40092 768732
rect 35808 767320 35860 767372
rect 36544 767320 36596 767372
rect 35808 766028 35860 766080
rect 39764 766028 39816 766080
rect 40040 765280 40092 765332
rect 41696 765280 41748 765332
rect 42064 765144 42116 765196
rect 42524 765144 42576 765196
rect 35808 764804 35860 764856
rect 39396 764804 39448 764856
rect 35808 764532 35860 764584
rect 41696 764600 41748 764652
rect 35624 763444 35676 763496
rect 40960 763444 41012 763496
rect 35808 763172 35860 763224
rect 41696 763104 41748 763156
rect 53104 763172 53156 763224
rect 42432 763036 42484 763088
rect 42064 761880 42116 761932
rect 48964 761880 49016 761932
rect 35808 761812 35860 761864
rect 41696 761812 41748 761864
rect 35164 759772 35216 759824
rect 41696 759772 41748 759824
rect 32404 759636 32456 759688
rect 41604 759636 41656 759688
rect 42064 759500 42116 759552
rect 42432 759500 42484 759552
rect 33784 758276 33836 758328
rect 39212 758276 39264 758328
rect 42248 756032 42300 756084
rect 44732 755488 44784 755540
rect 62948 755488 63000 755540
rect 42248 755420 42300 755472
rect 43628 754876 43680 754928
rect 45008 754876 45060 754928
rect 43996 753516 44048 753568
rect 45376 753516 45428 753568
rect 61384 747260 61436 747312
rect 63040 747260 63092 747312
rect 653404 746580 653456 746632
rect 675392 746580 675444 746632
rect 44824 746512 44876 746564
rect 62120 746512 62172 746564
rect 42800 744064 42852 744116
rect 62120 743860 62172 743912
rect 46204 743724 46256 743776
rect 62120 743724 62172 743776
rect 60004 742364 60056 742416
rect 62120 742364 62172 742416
rect 671804 742160 671856 742212
rect 675392 742160 675444 742212
rect 671620 741140 671672 741192
rect 675116 741140 675168 741192
rect 673552 738624 673604 738676
rect 675392 738624 675444 738676
rect 672264 738420 672316 738472
rect 675116 738420 675168 738472
rect 652024 736856 652076 736908
rect 656164 736856 656216 736908
rect 657544 735564 657596 735616
rect 675300 735700 675352 735752
rect 669596 735564 669648 735616
rect 675116 735564 675168 735616
rect 654784 734136 654836 734188
rect 675116 734204 675168 734256
rect 651472 733388 651524 733440
rect 668584 733388 668636 733440
rect 672080 732708 672132 732760
rect 675300 732708 675352 732760
rect 651472 731416 651524 731468
rect 658924 731416 658976 731468
rect 651380 731076 651432 731128
rect 653404 731076 653456 731128
rect 674932 731076 674984 731128
rect 675116 730872 675168 730924
rect 652668 730668 652720 730720
rect 661684 730668 661736 730720
rect 43628 730260 43680 730312
rect 61384 730260 61436 730312
rect 651472 729988 651524 730040
rect 657544 729988 657596 730040
rect 42248 729308 42300 729360
rect 62948 729308 63000 729360
rect 40960 728764 41012 728816
rect 41696 728832 41748 728884
rect 42064 728832 42116 728884
rect 43076 728832 43128 728884
rect 41144 728628 41196 728680
rect 41696 728628 41748 728680
rect 42064 728628 42116 728680
rect 43444 728628 43496 728680
rect 651472 728492 651524 728544
rect 654784 728492 654836 728544
rect 673092 728288 673144 728340
rect 670884 728084 670936 728136
rect 40868 727404 40920 727456
rect 41696 727404 41748 727456
rect 42064 727404 42116 727456
rect 44364 727404 44416 727456
rect 41328 727268 41380 727320
rect 41696 727268 41748 727320
rect 42064 727268 42116 727320
rect 44640 727268 44692 727320
rect 674564 726724 674616 726776
rect 683396 726724 683448 726776
rect 674748 726520 674800 726572
rect 681004 726520 681056 726572
rect 674380 726384 674432 726436
rect 684040 726384 684092 726436
rect 41328 726180 41380 726232
rect 41696 726180 41748 726232
rect 41144 725908 41196 725960
rect 41604 725908 41656 725960
rect 675300 721692 675352 721744
rect 675300 721216 675352 721268
rect 673920 721012 673972 721064
rect 675300 720808 675352 720860
rect 674472 720468 674524 720520
rect 675300 720468 675352 720520
rect 43628 718972 43680 719024
rect 55864 718972 55916 719024
rect 32404 716796 32456 716848
rect 41696 716796 41748 716848
rect 674288 716456 674340 716508
rect 676036 716456 676088 716508
rect 656164 716252 656216 716304
rect 674012 716252 674064 716304
rect 669964 715708 670016 715760
rect 674012 715708 674064 715760
rect 35164 715640 35216 715692
rect 40408 715640 40460 715692
rect 31668 715436 31720 715488
rect 38016 715436 38068 715488
rect 671068 715300 671120 715352
rect 674012 715300 674064 715352
rect 674288 715028 674340 715080
rect 676036 715028 676088 715080
rect 660304 714960 660356 715012
rect 674012 714960 674064 715012
rect 674288 714892 674340 714944
rect 676036 714892 676088 714944
rect 672448 714824 672500 714876
rect 674012 714824 674064 714876
rect 39304 714756 39356 714808
rect 41604 714756 41656 714808
rect 671896 714484 671948 714536
rect 674012 714484 674064 714536
rect 42064 714008 42116 714060
rect 42616 714008 42668 714060
rect 672632 713668 672684 713720
rect 674012 713668 674064 713720
rect 671068 713192 671120 713244
rect 674012 713192 674064 713244
rect 671896 712376 671948 712428
rect 674012 712376 674064 712428
rect 51724 712104 51776 712156
rect 42248 711084 42300 711136
rect 671436 709996 671488 710048
rect 674012 709996 674064 710048
rect 674288 709724 674340 709776
rect 676036 709724 676088 709776
rect 43628 709316 43680 709368
rect 45284 709316 45336 709368
rect 669044 709316 669096 709368
rect 674012 709316 674064 709368
rect 670608 709180 670660 709232
rect 674012 709180 674064 709232
rect 674288 708704 674340 708756
rect 676036 708704 676088 708756
rect 669228 708228 669280 708280
rect 674012 708228 674064 708280
rect 674472 707140 674524 707192
rect 676036 707140 676088 707192
rect 42432 705508 42484 705560
rect 43444 705508 43496 705560
rect 670424 705304 670476 705356
rect 674012 705304 674064 705356
rect 674288 705304 674340 705356
rect 683120 705304 683172 705356
rect 667848 705168 667900 705220
rect 674012 705168 674064 705220
rect 674288 705168 674340 705220
rect 675852 705168 675904 705220
rect 51724 705100 51776 705152
rect 62120 705100 62172 705152
rect 674288 703876 674340 703928
rect 676036 703876 676088 703928
rect 667020 703808 667072 703860
rect 674012 703808 674064 703860
rect 44180 703740 44232 703792
rect 62120 703740 62172 703792
rect 654784 701156 654836 701208
rect 673736 701156 673788 701208
rect 42708 701020 42760 701072
rect 62948 701020 63000 701072
rect 42064 699184 42116 699236
rect 42524 699184 42576 699236
rect 46204 698232 46256 698284
rect 62212 698232 62264 698284
rect 656532 690208 656584 690260
rect 674012 690208 674064 690260
rect 674472 690004 674524 690056
rect 675116 690004 675168 690056
rect 674932 688984 674984 689036
rect 652760 688780 652812 688832
rect 673000 688780 673052 688832
rect 675116 688780 675168 688832
rect 651472 688644 651524 688696
rect 657544 688644 657596 688696
rect 43444 687488 43496 687540
rect 61384 687488 61436 687540
rect 651472 687216 651524 687268
rect 669964 687216 670016 687268
rect 651472 687012 651524 687064
rect 654784 687012 654836 687064
rect 43444 686468 43496 686520
rect 62948 686468 63000 686520
rect 651656 686468 651708 686520
rect 667204 686468 667256 686520
rect 41328 686264 41380 686316
rect 41696 686264 41748 686316
rect 42064 686264 42116 686316
rect 42800 686264 42852 686316
rect 41144 686060 41196 686112
rect 41696 686060 41748 686112
rect 42064 686060 42116 686112
rect 43076 686060 43128 686112
rect 40960 685856 41012 685908
rect 41696 685856 41748 685908
rect 42064 685856 42116 685908
rect 45100 685856 45152 685908
rect 651472 685516 651524 685568
rect 656532 685516 656584 685568
rect 674288 683952 674340 684004
rect 674656 683952 674708 684004
rect 41328 683408 41380 683460
rect 41696 683408 41748 683460
rect 675484 682524 675536 682576
rect 683212 682524 683264 682576
rect 674748 682388 674800 682440
rect 683488 682388 683540 682440
rect 40776 678580 40828 678632
rect 41696 678580 41748 678632
rect 40776 677696 40828 677748
rect 41604 677696 41656 677748
rect 42432 676200 42484 676252
rect 60004 676200 60056 676252
rect 33048 674092 33100 674144
rect 41420 674092 41472 674144
rect 35164 672732 35216 672784
rect 41604 672732 41656 672784
rect 42616 671304 42668 671356
rect 673552 671304 673604 671356
rect 42616 671168 42668 671220
rect 668584 671100 668636 671152
rect 673552 671100 673604 671152
rect 36544 670964 36596 671016
rect 40500 670964 40552 671016
rect 661684 670692 661736 670744
rect 672448 670556 672500 670608
rect 673368 670556 673420 670608
rect 670240 669604 670292 669656
rect 673368 669604 673420 669656
rect 658924 669468 658976 669520
rect 673552 669468 673604 669520
rect 674840 669468 674892 669520
rect 676496 669468 676548 669520
rect 42432 669332 42484 669384
rect 57244 669332 57296 669384
rect 673552 668652 673604 668704
rect 671068 668516 671120 668568
rect 673552 668516 673604 668568
rect 671068 668108 671120 668160
rect 673552 668108 673604 668160
rect 44548 667904 44600 667956
rect 58624 667904 58676 667956
rect 671436 667904 671488 667956
rect 674840 667020 674892 667072
rect 676496 667020 676548 667072
rect 671896 666884 671948 666936
rect 673552 666884 673604 666936
rect 671896 666544 671948 666596
rect 673552 666544 673604 666596
rect 42248 665796 42300 665848
rect 44548 665796 44600 665848
rect 669596 665252 669648 665304
rect 673552 665252 673604 665304
rect 672264 665116 672316 665168
rect 673368 665116 673420 665168
rect 671712 664368 671764 664420
rect 673552 664368 673604 664420
rect 669412 663892 669464 663944
rect 673552 663892 673604 663944
rect 42616 663756 42668 663808
rect 674840 663756 674892 663808
rect 676036 663756 676088 663808
rect 42616 663552 42668 663604
rect 42248 663416 42300 663468
rect 42800 663416 42852 663468
rect 673552 663348 673604 663400
rect 673920 663348 673972 663400
rect 42248 663008 42300 663060
rect 43996 663008 44048 663060
rect 672080 662396 672132 662448
rect 673920 662396 673972 662448
rect 671252 661580 671304 661632
rect 673920 661580 673972 661632
rect 669228 661104 669280 661156
rect 673920 661104 673972 661156
rect 57244 660900 57296 660952
rect 62120 660900 62172 660952
rect 42156 660492 42208 660544
rect 43628 660492 43680 660544
rect 668860 660084 668912 660136
rect 673920 660084 673972 660136
rect 674840 659812 674892 659864
rect 683120 659812 683172 659864
rect 58624 659540 58676 659592
rect 62120 659540 62172 659592
rect 42156 658996 42208 659048
rect 42616 658996 42668 659048
rect 42524 657500 42576 657552
rect 62120 657500 62172 657552
rect 653404 655528 653456 655580
rect 673920 655528 673972 655580
rect 45468 655460 45520 655512
rect 62120 655460 62172 655512
rect 655520 645872 655572 645924
rect 674012 645872 674064 645924
rect 674564 644580 674616 644632
rect 675300 644580 675352 644632
rect 35808 644444 35860 644496
rect 40132 644444 40184 644496
rect 35808 643492 35860 643544
rect 40592 643492 40644 643544
rect 35532 643220 35584 643272
rect 41696 643288 41748 643340
rect 42064 643288 42116 643340
rect 45100 643288 45152 643340
rect 35348 643084 35400 643136
rect 41696 643084 41748 643136
rect 42064 643084 42116 643136
rect 61384 643084 61436 643136
rect 655336 643084 655388 643136
rect 674012 643084 674064 643136
rect 38568 642472 38620 642524
rect 41696 642472 41748 642524
rect 42064 642336 42116 642388
rect 62948 642336 63000 642388
rect 651472 642336 651524 642388
rect 658924 642336 658976 642388
rect 35808 642132 35860 642184
rect 40316 642132 40368 642184
rect 35440 641860 35492 641912
rect 39948 641860 40000 641912
rect 35624 641724 35676 641776
rect 41696 641724 41748 641776
rect 42064 641724 42116 641776
rect 44364 641724 44416 641776
rect 674748 641044 674800 641096
rect 674748 640840 674800 640892
rect 35808 640704 35860 640756
rect 39948 640704 40000 640756
rect 42064 640500 42116 640552
rect 42984 640500 43036 640552
rect 35532 640432 35584 640484
rect 41696 640432 41748 640484
rect 35348 640296 35400 640348
rect 41696 640296 41748 640348
rect 42064 640296 42116 640348
rect 45468 640296 45520 640348
rect 651472 640296 651524 640348
rect 668584 640296 668636 640348
rect 675208 640228 675260 640280
rect 674840 640160 674892 640212
rect 651380 640092 651432 640144
rect 653404 640092 653456 640144
rect 675024 639888 675076 639940
rect 674840 639752 674892 639804
rect 35808 639140 35860 639192
rect 39304 639072 39356 639124
rect 35808 638936 35860 638988
rect 40040 638936 40092 638988
rect 651656 638868 651708 638920
rect 655336 638868 655388 638920
rect 651472 638732 651524 638784
rect 655520 638732 655572 638784
rect 34428 638188 34480 638240
rect 41696 638188 41748 638240
rect 674748 637712 674800 637764
rect 35808 637576 35860 637628
rect 36544 637576 36596 637628
rect 674748 637576 674800 637628
rect 674288 637440 674340 637492
rect 675484 637440 675536 637492
rect 674748 637032 674800 637084
rect 683212 637032 683264 637084
rect 35624 636828 35676 636880
rect 40316 636828 40368 636880
rect 675484 636828 675536 636880
rect 683396 636828 683448 636880
rect 35808 636692 35860 636744
rect 40868 636624 40920 636676
rect 35808 636352 35860 636404
rect 40500 636352 40552 636404
rect 35532 636216 35584 636268
rect 39120 636148 39172 636200
rect 674932 635468 674984 635520
rect 675668 635468 675720 635520
rect 35808 634788 35860 634840
rect 40500 634788 40552 634840
rect 652024 634040 652076 634092
rect 660304 634040 660356 634092
rect 35808 633836 35860 633888
rect 39764 633700 39816 633752
rect 35808 633428 35860 633480
rect 41512 633428 41564 633480
rect 42064 633428 42116 633480
rect 60188 633428 60240 633480
rect 36544 630572 36596 630624
rect 41604 630504 41656 630556
rect 671528 628736 671580 628788
rect 35164 628532 35216 628584
rect 40500 628532 40552 628584
rect 671344 628396 671396 628448
rect 669964 625948 670016 626000
rect 673552 625948 673604 626000
rect 44180 625812 44232 625864
rect 63132 625812 63184 625864
rect 667204 625676 667256 625728
rect 674012 625676 674064 625728
rect 674748 625676 674800 625728
rect 676496 625676 676548 625728
rect 657544 625132 657596 625184
rect 674012 625132 674064 625184
rect 670240 624996 670292 625048
rect 674012 624996 674064 625048
rect 42248 624656 42300 624708
rect 44180 624656 44232 624708
rect 670240 624656 670292 624708
rect 674012 624656 674064 624708
rect 671436 624316 671488 624368
rect 674012 624316 674064 624368
rect 42248 624044 42300 624096
rect 44364 624044 44416 624096
rect 669412 623840 669464 623892
rect 674012 623840 674064 623892
rect 671068 623500 671120 623552
rect 674012 623500 674064 623552
rect 670424 623024 670476 623076
rect 674012 623024 674064 623076
rect 674380 623024 674432 623076
rect 683396 623024 683448 623076
rect 671896 622684 671948 622736
rect 674012 622684 674064 622736
rect 671436 622208 671488 622260
rect 674012 622208 674064 622260
rect 42248 621664 42300 621716
rect 44180 621664 44232 621716
rect 667664 621596 667716 621648
rect 674012 621596 674064 621648
rect 42248 621528 42300 621580
rect 43996 621528 44048 621580
rect 670884 620644 670936 620696
rect 672540 620644 672592 620696
rect 42248 620372 42300 620424
rect 42708 620372 42760 620424
rect 669044 620372 669096 620424
rect 673644 620372 673696 620424
rect 669780 619828 669832 619880
rect 673644 619828 673696 619880
rect 42248 619624 42300 619676
rect 42892 619624 42944 619676
rect 668216 617924 668268 617976
rect 673644 617924 673696 617976
rect 674288 617516 674340 617568
rect 676220 617516 676272 617568
rect 42248 617312 42300 617364
rect 43076 617312 43128 617364
rect 668400 616836 668452 616888
rect 673644 616836 673696 616888
rect 44180 616768 44232 616820
rect 62120 616768 62172 616820
rect 670608 615476 670660 615528
rect 673644 615476 673696 615528
rect 674288 615476 674340 615528
rect 683120 615476 683172 615528
rect 670608 614864 670660 614916
rect 673644 614864 673696 614916
rect 42708 614116 42760 614168
rect 62120 614116 62172 614168
rect 46204 613368 46256 613420
rect 62120 613368 62172 613420
rect 42248 612348 42300 612400
rect 43812 612620 43864 612672
rect 43996 612212 44048 612264
rect 44732 612212 44784 612264
rect 44088 612076 44140 612128
rect 43875 611940 43927 611992
rect 44272 611668 44324 611720
rect 44916 611532 44968 611584
rect 653404 611328 653456 611380
rect 673644 611328 673696 611380
rect 50160 611260 50212 611312
rect 44318 611124 44370 611176
rect 44732 610716 44784 610768
rect 50160 610104 50212 610156
rect 58624 610104 58676 610156
rect 61384 609968 61436 610020
rect 667664 608608 667716 608660
rect 673184 608608 673236 608660
rect 674288 608336 674340 608388
rect 675484 608336 675536 608388
rect 674288 603236 674340 603288
rect 675116 603236 675168 603288
rect 35808 601672 35860 601724
rect 36544 601672 36596 601724
rect 657544 600448 657596 600500
rect 673828 600380 673880 600432
rect 654784 598952 654836 599004
rect 673184 598952 673236 599004
rect 674472 598952 674524 599004
rect 675300 598952 675352 599004
rect 651472 597524 651524 597576
rect 669964 597524 670016 597576
rect 43076 597388 43128 597440
rect 43076 596980 43128 597032
rect 651472 596164 651524 596216
rect 664444 596164 664496 596216
rect 40132 595756 40184 595808
rect 41696 595756 41748 595808
rect 651656 595484 651708 595536
rect 653404 595484 653456 595536
rect 651472 594804 651524 594856
rect 661684 594804 661736 594856
rect 41328 594736 41380 594788
rect 41696 594736 41748 594788
rect 651472 594668 651524 594720
rect 657544 594668 657596 594720
rect 39948 594260 40000 594312
rect 41604 594260 41656 594312
rect 651472 593240 651524 593292
rect 654784 593240 654836 593292
rect 674288 592628 674340 592680
rect 683396 592628 683448 592680
rect 674840 591472 674892 591524
rect 679624 591472 679676 591524
rect 35624 590792 35676 590844
rect 41696 590724 41748 590776
rect 35808 590656 35860 590708
rect 39672 590656 39724 590708
rect 42064 590656 42116 590708
rect 43260 590656 43312 590708
rect 674656 588548 674708 588600
rect 684040 588548 684092 588600
rect 33048 587120 33100 587172
rect 41512 587120 41564 587172
rect 42248 586236 42300 586288
rect 42616 586236 42668 586288
rect 35164 586100 35216 586152
rect 39396 586032 39448 586084
rect 33784 585896 33836 585948
rect 39764 585896 39816 585948
rect 31024 585760 31076 585812
rect 39212 585760 39264 585812
rect 660304 581000 660356 581052
rect 673184 581000 673236 581052
rect 668584 580252 668636 580304
rect 673184 580252 673236 580304
rect 670240 579980 670292 580032
rect 673184 579980 673236 580032
rect 674380 579708 674432 579760
rect 676220 579708 676272 579760
rect 658924 579640 658976 579692
rect 673184 579640 673236 579692
rect 42248 578960 42300 579012
rect 43260 578960 43312 579012
rect 669412 578892 669464 578944
rect 673184 578892 673236 578944
rect 674472 578416 674524 578468
rect 676220 578416 676272 578468
rect 670792 578212 670844 578264
rect 673184 578212 673236 578264
rect 670240 577600 670292 577652
rect 673184 577600 673236 577652
rect 674380 577532 674432 577584
rect 676220 577532 676272 577584
rect 670424 577396 670476 577448
rect 673184 577396 673236 577448
rect 671436 577124 671488 577176
rect 673184 577124 673236 577176
rect 669412 576852 669464 576904
rect 673184 576852 673236 576904
rect 45100 575424 45152 575476
rect 62120 575424 62172 575476
rect 671620 574540 671672 574592
rect 673920 574540 673972 574592
rect 671988 574268 672040 574320
rect 673920 574268 673972 574320
rect 667480 574064 667532 574116
rect 46940 573996 46992 574048
rect 62120 573996 62172 574048
rect 674380 574064 674432 574116
rect 676220 574064 676272 574116
rect 673920 573860 673972 573912
rect 671804 571548 671856 571600
rect 673920 571548 673972 571600
rect 674564 571548 674616 571600
rect 676036 571548 676088 571600
rect 674380 571412 674432 571464
rect 676220 571412 676272 571464
rect 669596 571344 669648 571396
rect 673920 571344 673972 571396
rect 671344 571072 671396 571124
rect 673920 571072 673972 571124
rect 42064 570936 42116 570988
rect 42616 570936 42668 570988
rect 674840 570460 674892 570512
rect 675484 570460 675536 570512
rect 683120 570460 683172 570512
rect 671988 569916 672040 569968
rect 673920 569916 673972 569968
rect 669780 568556 669832 568608
rect 673920 568556 673972 568608
rect 653404 565836 653456 565888
rect 673920 565836 673972 565888
rect 665088 564408 665140 564460
rect 673920 564408 673972 564460
rect 657820 554752 657872 554804
rect 672724 554752 672776 554804
rect 674656 553460 674708 553512
rect 675300 553460 675352 553512
rect 655152 553392 655204 553444
rect 669596 553392 669648 553444
rect 674472 552916 674524 552968
rect 674932 552984 674984 553036
rect 651472 552644 651524 552696
rect 665824 552644 665876 552696
rect 41328 552032 41380 552084
rect 41696 552032 41748 552084
rect 674472 552032 674524 552084
rect 675116 552032 675168 552084
rect 651472 550604 651524 550656
rect 660304 550604 660356 550656
rect 40960 550400 41012 550452
rect 41696 550400 41748 550452
rect 651380 550332 651432 550384
rect 653404 550332 653456 550384
rect 651656 549856 651708 549908
rect 663064 549856 663116 549908
rect 651472 549176 651524 549228
rect 657820 549176 657872 549228
rect 674932 548836 674984 548888
rect 675300 548836 675352 548888
rect 651472 548768 651524 548820
rect 655152 548768 655204 548820
rect 41328 547884 41380 547936
rect 41696 547884 41748 547936
rect 674288 547340 674340 547392
rect 683212 547340 683264 547392
rect 29644 547136 29696 547188
rect 41696 547136 41748 547188
rect 675576 547136 675628 547188
rect 683396 547136 683448 547188
rect 675208 546592 675260 546644
rect 675576 546592 675628 546644
rect 675392 546456 675444 546508
rect 681004 546456 681056 546508
rect 675116 540948 675168 541000
rect 675576 540948 675628 541000
rect 673552 536120 673604 536172
rect 673920 536120 673972 536172
rect 669964 535916 670016 535968
rect 674012 535916 674064 535968
rect 674288 535848 674340 535900
rect 676036 535848 676088 535900
rect 674288 535644 674340 535696
rect 676220 535644 676272 535696
rect 664444 535440 664496 535492
rect 674012 535440 674064 535492
rect 670976 534964 671028 535016
rect 674012 534964 674064 535016
rect 674288 534896 674340 534948
rect 676036 534896 676088 534948
rect 670792 534692 670844 534744
rect 674012 534692 674064 534744
rect 674288 534624 674340 534676
rect 676496 534624 676548 534676
rect 674288 534488 674340 534540
rect 676220 534488 676272 534540
rect 661684 534080 661736 534132
rect 674012 534080 674064 534132
rect 675484 533332 675536 533384
rect 683580 533332 683632 533384
rect 670240 533264 670292 533316
rect 674012 533264 674064 533316
rect 674288 533196 674340 533248
rect 676036 533196 676088 533248
rect 674288 532788 674340 532840
rect 676036 532788 676088 532840
rect 670792 532720 670844 532772
rect 674012 532720 674064 532772
rect 669412 532516 669464 532568
rect 674012 532516 674064 532568
rect 674288 532448 674340 532500
rect 676036 532448 676088 532500
rect 44824 531972 44876 532024
rect 62120 531972 62172 532024
rect 671620 531972 671672 532024
rect 674012 531972 674064 532024
rect 674288 531972 674340 532024
rect 676036 531972 676088 532024
rect 667664 531836 667716 531888
rect 674012 531836 674064 531888
rect 674288 531768 674340 531820
rect 676220 531768 676272 531820
rect 51724 531224 51776 531276
rect 62304 531224 62356 531276
rect 42708 530884 42760 530936
rect 672172 530884 672224 530936
rect 674012 530884 674064 530936
rect 674288 530816 674340 530868
rect 676036 530816 676088 530868
rect 42156 530680 42208 530732
rect 42248 530272 42300 530324
rect 42892 530272 42944 530324
rect 667296 529932 667348 529984
rect 674012 529932 674064 529984
rect 674288 529932 674340 529984
rect 676036 529932 676088 529984
rect 671160 529388 671212 529440
rect 674012 529388 674064 529440
rect 674288 529320 674340 529372
rect 676036 529320 676088 529372
rect 674288 529184 674340 529236
rect 676220 529184 676272 529236
rect 668400 529116 668452 529168
rect 674012 529116 674064 529168
rect 672356 528844 672408 528896
rect 674012 528844 674064 528896
rect 674288 528776 674340 528828
rect 676036 528776 676088 528828
rect 45192 528572 45244 528624
rect 62120 528572 62172 528624
rect 672540 528028 672592 528080
rect 674012 528028 674064 528080
rect 674288 527960 674340 528012
rect 676036 527960 676088 528012
rect 47584 527076 47636 527128
rect 62120 527076 62172 527128
rect 42064 527008 42116 527060
rect 42708 527008 42760 527060
rect 669044 524560 669096 524612
rect 674012 524560 674064 524612
rect 674288 524560 674340 524612
rect 683120 524560 683172 524612
rect 668584 524424 668636 524476
rect 669044 524424 669096 524476
rect 675484 520208 675536 520260
rect 680360 520208 680412 520260
rect 675668 518780 675720 518832
rect 677876 518780 677928 518832
rect 658464 518168 658516 518220
rect 668584 518168 668636 518220
rect 650644 509872 650696 509924
rect 658464 509872 658516 509924
rect 675116 503616 675168 503668
rect 679624 503616 679676 503668
rect 675300 503480 675352 503532
rect 681004 503480 681056 503532
rect 674840 500896 674892 500948
rect 681188 500896 681240 500948
rect 674288 491648 674340 491700
rect 676036 491648 676088 491700
rect 665824 491580 665876 491632
rect 674012 491580 674064 491632
rect 663064 491444 663116 491496
rect 673828 491444 673880 491496
rect 660304 491308 660356 491360
rect 674012 491308 674064 491360
rect 670976 490900 671028 490952
rect 674012 490900 674064 490952
rect 672540 490696 672592 490748
rect 672908 490696 672960 490748
rect 672448 489608 672500 489660
rect 674012 489608 674064 489660
rect 670792 489268 670844 489320
rect 674012 489268 674064 489320
rect 671620 488452 671672 488504
rect 674012 488452 674064 488504
rect 672632 486004 672684 486056
rect 674012 486004 674064 486056
rect 674288 485868 674340 485920
rect 676036 485868 676088 485920
rect 665088 485800 665140 485852
rect 674012 485800 674064 485852
rect 674288 485120 674340 485172
rect 676036 485120 676088 485172
rect 668768 484372 668820 484424
rect 674012 484372 674064 484424
rect 674472 483964 674524 484016
rect 676036 483964 676088 484016
rect 671804 483148 671856 483200
rect 674012 483148 674064 483200
rect 676220 482944 676272 482996
rect 677416 482944 677468 482996
rect 674656 482332 674708 482384
rect 676036 482332 676088 482384
rect 665180 480360 665232 480412
rect 670424 480360 670476 480412
rect 674012 480360 674064 480412
rect 674288 480360 674340 480412
rect 683120 480360 683172 480412
rect 659660 476144 659712 476196
rect 665180 476144 665232 476196
rect 676036 475124 676088 475176
rect 680360 475124 680412 475176
rect 656164 473424 656216 473476
rect 659660 473424 659712 473476
rect 650828 470568 650880 470620
rect 656164 470568 656216 470620
rect 667020 456560 667072 456612
rect 667848 455948 667900 456000
rect 673368 455812 673420 455864
rect 669228 455608 669280 455660
rect 673276 455336 673328 455388
rect 673388 455200 673440 455252
rect 673506 455200 673558 455252
rect 674288 454860 674340 454912
rect 675852 454860 675904 454912
rect 672080 454792 672132 454844
rect 673046 454588 673098 454640
rect 674288 454588 674340 454640
rect 675484 454588 675536 454640
rect 672816 454452 672868 454504
rect 672954 454316 673006 454368
rect 674288 454316 674340 454368
rect 675668 454316 675720 454368
rect 672264 453908 672316 453960
rect 674288 453908 674340 453960
rect 676036 453908 676088 453960
rect 35808 429156 35860 429208
rect 41696 429156 41748 429208
rect 35808 427932 35860 427984
rect 41696 427932 41748 427984
rect 40960 424328 41012 424380
rect 41696 424328 41748 424380
rect 41144 422356 41196 422408
rect 41604 422356 41656 422408
rect 32036 417392 32088 417444
rect 41696 417392 41748 417444
rect 42064 417256 42116 417308
rect 42616 417256 42668 417308
rect 34520 416032 34572 416084
rect 41696 416032 41748 416084
rect 42248 409776 42300 409828
rect 43168 409776 43220 409828
rect 42248 406988 42300 407040
rect 42616 406988 42668 407040
rect 44732 404268 44784 404320
rect 62120 404268 62172 404320
rect 674564 403248 674616 403300
rect 676220 403248 676272 403300
rect 51448 402908 51500 402960
rect 62120 402908 62172 402960
rect 42432 402228 42484 402280
rect 42984 402228 43036 402280
rect 45192 400256 45244 400308
rect 51080 400188 51132 400240
rect 62120 400188 62172 400240
rect 62120 400052 62172 400104
rect 46388 399440 46440 399492
rect 56048 399440 56100 399492
rect 674932 398828 674984 398880
rect 676036 398828 676088 398880
rect 47768 398760 47820 398812
rect 62120 398760 62172 398812
rect 674564 396040 674616 396092
rect 676036 396040 676088 396092
rect 675208 395700 675260 395752
rect 676220 395700 676272 395752
rect 674380 394272 674432 394324
rect 676220 394272 676272 394324
rect 41328 386384 41380 386436
rect 41696 386384 41748 386436
rect 679624 386724 679676 386776
rect 675484 385976 675536 386028
rect 674840 384752 674892 384804
rect 675392 384752 675444 384804
rect 41328 382236 41380 382288
rect 41696 382236 41748 382288
rect 674380 382168 674432 382220
rect 675116 382168 675168 382220
rect 41328 379720 41380 379772
rect 41512 379720 41564 379772
rect 35808 379516 35860 379568
rect 40408 379584 40460 379636
rect 35808 378156 35860 378208
rect 41696 378156 41748 378208
rect 674380 378088 674432 378140
rect 675116 378088 675168 378140
rect 651472 373940 651524 373992
rect 657544 373940 657596 373992
rect 33968 373260 34020 373312
rect 41696 373260 41748 373312
rect 674656 372512 674708 372564
rect 675300 372512 675352 372564
rect 39304 372036 39356 372088
rect 41696 372036 41748 372088
rect 42064 371900 42116 371952
rect 42708 371900 42760 371952
rect 651472 370948 651524 371000
rect 654784 370948 654836 371000
rect 42432 366800 42484 366852
rect 43076 366800 43128 366852
rect 42248 365848 42300 365900
rect 42708 365848 42760 365900
rect 655520 364964 655572 365016
rect 668584 364964 668636 365016
rect 42340 362856 42392 362908
rect 42708 362856 42760 362908
rect 651012 361564 651064 361616
rect 655520 361564 655572 361616
rect 44640 361496 44692 361548
rect 62120 361496 62172 361548
rect 51080 360136 51132 360188
rect 62120 360136 62172 360188
rect 44640 357416 44692 357468
rect 62120 357416 62172 357468
rect 42248 355988 42300 356040
rect 42892 355988 42944 356040
rect 47768 355988 47820 356040
rect 62120 355988 62172 356040
rect 44640 354492 44692 354544
rect 44732 354288 44784 354340
rect 45468 354560 45520 354612
rect 45468 354084 45520 354136
rect 45468 353812 45520 353864
rect 45303 353676 45355 353728
rect 47952 353404 48004 353456
rect 45422 353132 45474 353184
rect 35808 344564 35860 344616
rect 40040 344564 40092 344616
rect 35532 343748 35584 343800
rect 40040 343748 40092 343800
rect 35808 342252 35860 342304
rect 40224 342252 40276 342304
rect 33048 341368 33100 341420
rect 40224 341368 40276 341420
rect 45468 341368 45520 341420
rect 62212 341368 62264 341420
rect 35808 341164 35860 341216
rect 40224 341164 40276 341216
rect 35624 341028 35676 341080
rect 40040 341028 40092 341080
rect 35532 339600 35584 339652
rect 36544 339600 36596 339652
rect 35808 339464 35860 339516
rect 38844 339464 38896 339516
rect 35808 335316 35860 335368
rect 40224 335316 40276 335368
rect 35624 334228 35676 334280
rect 39396 334228 39448 334280
rect 35808 333956 35860 334008
rect 41696 333956 41748 334008
rect 42064 333956 42116 334008
rect 42984 333956 43036 334008
rect 674472 333888 674524 333940
rect 675116 333888 675168 333940
rect 651380 328244 651432 328296
rect 654784 328244 654836 328296
rect 651380 325592 651432 325644
rect 653404 325592 653456 325644
rect 42248 322872 42300 322924
rect 43168 322872 43220 322924
rect 42248 320220 42300 320272
rect 42616 319948 42668 320000
rect 60372 315936 60424 315988
rect 62120 315936 62172 315988
rect 51080 314712 51132 314764
rect 62120 314712 62172 314764
rect 46388 309068 46440 309120
rect 47768 309068 47820 309120
rect 676220 306348 676272 306400
rect 676864 306348 676916 306400
rect 675852 304920 675904 304972
rect 676404 304920 676456 304972
rect 651380 303492 651432 303544
rect 653404 303492 653456 303544
rect 651472 300772 651524 300824
rect 660304 300772 660356 300824
rect 41144 299616 41196 299668
rect 41604 299616 41656 299668
rect 675852 297032 675904 297084
rect 679624 297032 679676 297084
rect 651932 296760 651984 296812
rect 665824 296692 665876 296744
rect 675484 296352 675536 296404
rect 41328 295604 41380 295656
rect 41696 295604 41748 295656
rect 50528 295332 50580 295384
rect 62120 295332 62172 295384
rect 675484 295196 675536 295248
rect 57244 294040 57296 294092
rect 62120 294040 62172 294092
rect 651472 293972 651524 294024
rect 664444 293972 664496 294024
rect 51908 292544 51960 292596
rect 62120 292544 62172 292596
rect 41144 292204 41196 292256
rect 41604 292204 41656 292256
rect 47584 292136 47636 292188
rect 53472 292136 53524 292188
rect 47768 292000 47820 292052
rect 53656 292000 53708 292052
rect 41236 291252 41288 291304
rect 41696 291252 41748 291304
rect 651472 291184 651524 291236
rect 663064 291184 663116 291236
rect 53288 291116 53340 291168
rect 62120 291116 62172 291168
rect 651380 290368 651432 290420
rect 653404 290368 653456 290420
rect 651472 288396 651524 288448
rect 672172 288396 672224 288448
rect 651472 287036 651524 287088
rect 667572 287036 667624 287088
rect 33784 286288 33836 286340
rect 41696 286288 41748 286340
rect 46388 285676 46440 285728
rect 63040 285676 63092 285728
rect 651472 285676 651524 285728
rect 667388 285676 667440 285728
rect 674472 285608 674524 285660
rect 675116 285608 675168 285660
rect 53656 284928 53708 284980
rect 56324 284928 56376 284980
rect 39304 284724 39356 284776
rect 41696 284724 41748 284776
rect 42064 284656 42116 284708
rect 42616 284656 42668 284708
rect 60372 284384 60424 284436
rect 62120 284384 62172 284436
rect 651472 284316 651524 284368
rect 672356 284316 672408 284368
rect 47768 282888 47820 282940
rect 62120 282888 62172 282940
rect 651472 282140 651524 282192
rect 666560 282140 666612 282192
rect 53288 281528 53340 281580
rect 62120 281528 62172 281580
rect 58808 280168 58860 280220
rect 62120 280168 62172 280220
rect 651472 280168 651524 280220
rect 667204 280168 667256 280220
rect 62580 278672 62632 278724
rect 671344 278672 671396 278724
rect 63408 278536 63460 278588
rect 671712 278536 671764 278588
rect 56048 278400 56100 278452
rect 651012 278400 651064 278452
rect 51724 278264 51776 278316
rect 635004 278264 635056 278316
rect 47952 278128 48004 278180
rect 637764 278128 637816 278180
rect 64144 277992 64196 278044
rect 667940 277992 667992 278044
rect 53472 277856 53524 277908
rect 56324 277720 56376 277772
rect 69664 277856 69716 277908
rect 629484 277856 629536 277908
rect 650828 277856 650880 277908
rect 64328 277584 64380 277636
rect 650644 277720 650696 277772
rect 69664 277448 69716 277500
rect 629484 277448 629536 277500
rect 636200 277584 636252 277636
rect 42248 277312 42300 277364
rect 42800 277312 42852 277364
rect 482836 277312 482888 277364
rect 557540 277312 557592 277364
rect 487988 277176 488040 277228
rect 565820 277176 565872 277228
rect 497924 277040 497976 277092
rect 579988 277040 580040 277092
rect 511632 276904 511684 276956
rect 600136 276904 600188 276956
rect 514484 276768 514536 276820
rect 603632 276768 603684 276820
rect 518716 276632 518768 276684
rect 609612 276632 609664 276684
rect 479984 276496 480036 276548
rect 555240 276496 555292 276548
rect 477040 276360 477092 276412
rect 550456 276360 550508 276412
rect 471612 276224 471664 276276
rect 543372 276224 543424 276276
rect 107200 275952 107252 276004
rect 163504 275952 163556 276004
rect 167552 275952 167604 276004
rect 178868 275952 178920 276004
rect 185216 275952 185268 276004
rect 221280 275952 221332 276004
rect 232504 275952 232556 276004
rect 239220 275952 239272 276004
rect 410800 275952 410852 276004
rect 455880 275952 455932 276004
rect 456064 275952 456116 276004
rect 509056 275952 509108 276004
rect 513196 275952 513248 276004
rect 601332 275952 601384 276004
rect 139124 275816 139176 275868
rect 174268 275816 174320 275868
rect 178132 275816 178184 275868
rect 216680 275816 216732 275868
rect 224224 275816 224276 275868
rect 232688 275816 232740 275868
rect 236092 275816 236144 275868
rect 250444 275816 250496 275868
rect 286876 275816 286928 275868
rect 291844 275816 291896 275868
rect 430212 275816 430264 275868
rect 484308 275816 484360 275868
rect 490564 275816 490616 275868
rect 505560 275816 505612 275868
rect 522764 275816 522816 275868
rect 615500 275816 615552 275868
rect 260932 275748 260984 275800
rect 266360 275748 266412 275800
rect 93032 275680 93084 275732
rect 152832 275680 152884 275732
rect 160468 275680 160520 275732
rect 199568 275680 199620 275732
rect 217140 275680 217192 275732
rect 224224 275680 224276 275732
rect 229008 275680 229060 275732
rect 243544 275680 243596 275732
rect 250260 275680 250312 275732
rect 259368 275680 259420 275732
rect 284576 275680 284628 275732
rect 290096 275680 290148 275732
rect 416412 275680 416464 275732
rect 462964 275680 463016 275732
rect 463148 275680 463200 275732
rect 516232 275680 516284 275732
rect 528192 275680 528244 275732
rect 622584 275680 622636 275732
rect 76472 275544 76524 275596
rect 86224 275544 86276 275596
rect 90732 275544 90784 275596
rect 154764 275544 154816 275596
rect 171048 275544 171100 275596
rect 211620 275544 211672 275596
rect 218336 275544 218388 275596
rect 233884 275544 233936 275596
rect 239588 275544 239640 275596
rect 255964 275544 256016 275596
rect 257344 275544 257396 275596
rect 262312 275544 262364 275596
rect 266820 275544 266872 275596
rect 276480 275544 276532 275596
rect 363880 275544 363932 275596
rect 388536 275544 388588 275596
rect 445024 275544 445076 275596
rect 498476 275544 498528 275596
rect 498844 275544 498896 275596
rect 512644 275544 512696 275596
rect 516784 275544 516836 275596
rect 526812 275544 526864 275596
rect 532332 275544 532384 275596
rect 629668 275544 629720 275596
rect 277492 275476 277544 275528
rect 285128 275476 285180 275528
rect 100116 275408 100168 275460
rect 71780 275272 71832 275324
rect 141056 275272 141108 275324
rect 156880 275408 156932 275460
rect 159456 275272 159508 275324
rect 163964 275408 164016 275460
rect 206376 275408 206428 275460
rect 221924 275408 221976 275460
rect 243728 275408 243780 275460
rect 256148 275408 256200 275460
rect 200764 275272 200816 275324
rect 214840 275272 214892 275324
rect 239404 275272 239456 275324
rect 243176 275272 243228 275324
rect 256700 275272 256752 275324
rect 358636 275408 358688 275460
rect 381452 275408 381504 275460
rect 386052 275408 386104 275460
rect 420460 275408 420512 275460
rect 435640 275408 435692 275460
rect 485044 275408 485096 275460
rect 485228 275408 485280 275460
rect 530400 275408 530452 275460
rect 537668 275408 537720 275460
rect 636752 275408 636804 275460
rect 269212 275340 269264 275392
rect 274640 275340 274692 275392
rect 276296 275272 276348 275324
rect 283104 275272 283156 275324
rect 285680 275272 285732 275324
rect 291292 275272 291344 275324
rect 291660 275272 291712 275324
rect 295340 275272 295392 275324
rect 299940 275272 299992 275324
rect 301136 275272 301188 275324
rect 326436 275272 326488 275324
rect 335360 275272 335412 275324
rect 371056 275272 371108 275324
rect 399208 275272 399260 275324
rect 418804 275272 418856 275324
rect 466552 275272 466604 275324
rect 467564 275272 467616 275324
rect 537484 275272 537536 275324
rect 542268 275272 542320 275324
rect 643836 275272 643888 275324
rect 270132 275204 270184 275256
rect 96620 275136 96672 275188
rect 149612 275136 149664 275188
rect 153384 275136 153436 275188
rect 169024 275136 169076 275188
rect 190000 275136 190052 275188
rect 222936 275136 222988 275188
rect 292856 275136 292908 275188
rect 295800 275136 295852 275188
rect 298744 275136 298796 275188
rect 300032 275136 300084 275188
rect 427084 275136 427136 275188
rect 477224 275136 477276 275188
rect 485044 275136 485096 275188
rect 491392 275136 491444 275188
rect 507492 275136 507544 275188
rect 594248 275136 594300 275188
rect 263232 275068 263284 275120
rect 273260 275068 273312 275120
rect 136824 275000 136876 275052
rect 137652 275000 137704 275052
rect 146208 275000 146260 275052
rect 185308 275000 185360 275052
rect 288072 275000 288124 275052
rect 292856 275000 292908 275052
rect 420552 275000 420604 275052
rect 470140 275000 470192 275052
rect 484308 275000 484360 275052
rect 485228 275000 485280 275052
rect 503444 275000 503496 275052
rect 587072 275000 587124 275052
rect 81256 274932 81308 274984
rect 293960 274932 294012 274984
rect 297180 274932 297232 274984
rect 145288 274864 145340 274916
rect 149796 274864 149848 274916
rect 189080 274864 189132 274916
rect 289268 274864 289320 274916
rect 292672 274864 292724 274916
rect 473084 274864 473136 274916
rect 544568 274864 544620 274916
rect 296352 274796 296404 274848
rect 298376 274796 298428 274848
rect 128544 274728 128596 274780
rect 168288 274728 168340 274780
rect 207756 274728 207808 274780
rect 210700 274728 210752 274780
rect 476764 274728 476816 274780
rect 523316 274728 523368 274780
rect 523684 274728 523736 274780
rect 533896 274728 533948 274780
rect 534724 274728 534776 274780
rect 540980 274728 541032 274780
rect 74172 274660 74224 274712
rect 76840 274660 76892 274712
rect 85948 274660 86000 274712
rect 90364 274660 90416 274712
rect 103704 274660 103756 274712
rect 104808 274660 104860 274712
rect 110788 274660 110840 274712
rect 111708 274660 111760 274712
rect 253848 274660 253900 274712
rect 256884 274660 256936 274712
rect 275100 274660 275152 274712
rect 278320 274660 278372 274712
rect 283380 274660 283432 274712
rect 289176 274660 289228 274712
rect 290464 274660 290516 274712
rect 294144 274660 294196 274712
rect 295156 274660 295208 274712
rect 296812 274660 296864 274712
rect 297548 274660 297600 274712
rect 299480 274660 299532 274712
rect 303436 274660 303488 274712
rect 303988 274660 304040 274712
rect 321192 274660 321244 274712
rect 328276 274660 328328 274712
rect 114376 274592 114428 274644
rect 171600 274592 171652 274644
rect 179328 274592 179380 274644
rect 214564 274592 214616 274644
rect 409788 274592 409840 274644
rect 453580 274592 453632 274644
rect 457444 274592 457496 274644
rect 480720 274592 480772 274644
rect 486792 274592 486844 274644
rect 563428 274592 563480 274644
rect 101312 274456 101364 274508
rect 160928 274456 160980 274508
rect 168748 274456 168800 274508
rect 208400 274456 208452 274508
rect 381544 274456 381596 274508
rect 392124 274456 392176 274508
rect 413836 274456 413888 274508
rect 460664 274456 460716 274508
rect 463240 274456 463292 274508
rect 484308 274456 484360 274508
rect 488356 274456 488408 274508
rect 567016 274456 567068 274508
rect 95424 274320 95476 274372
rect 157616 274320 157668 274372
rect 159272 274320 159324 274372
rect 202328 274320 202380 274372
rect 223120 274320 223172 274372
rect 247224 274320 247276 274372
rect 369124 274320 369176 274372
rect 387340 274320 387392 274372
rect 419080 274320 419132 274372
rect 467748 274320 467800 274372
rect 506204 274320 506256 274372
rect 591856 274320 591908 274372
rect 331864 274252 331916 274304
rect 337752 274252 337804 274304
rect 67088 274184 67140 274236
rect 130384 274184 130436 274236
rect 130844 274184 130896 274236
rect 182456 274184 182508 274236
rect 193496 274184 193548 274236
rect 226432 274184 226484 274236
rect 239220 274184 239272 274236
rect 253940 274184 253992 274236
rect 359464 274184 359516 274236
rect 380256 274184 380308 274236
rect 388996 274184 389048 274236
rect 425152 274184 425204 274236
rect 425704 274184 425756 274236
rect 474832 274184 474884 274236
rect 511816 274184 511868 274236
rect 598940 274184 598992 274236
rect 77668 274048 77720 274100
rect 144920 274048 144972 274100
rect 154488 274048 154540 274100
rect 198096 274048 198148 274100
rect 210056 274048 210108 274100
rect 237840 274048 237892 274100
rect 249064 274048 249116 274100
rect 265256 274048 265308 274100
rect 266360 274048 266412 274100
rect 273536 274048 273588 274100
rect 278596 274048 278648 274100
rect 285864 274048 285916 274100
rect 337752 274048 337804 274100
rect 351920 274048 351972 274100
rect 353944 274048 353996 274100
rect 369584 274048 369636 274100
rect 373264 274048 373316 274100
rect 400312 274048 400364 274100
rect 401508 274048 401560 274100
rect 442908 274048 442960 274100
rect 451188 274048 451240 274100
rect 513840 274048 513892 274100
rect 536748 274048 536800 274100
rect 634360 274048 634412 274100
rect 69388 273912 69440 273964
rect 139400 273912 139452 273964
rect 148600 273912 148652 273964
rect 194784 273912 194836 273964
rect 208860 273912 208912 273964
rect 237472 273912 237524 273964
rect 238484 273912 238536 273964
rect 88340 273776 88392 273828
rect 119344 273776 119396 273828
rect 120264 273776 120316 273828
rect 175280 273776 175332 273828
rect 192392 273776 192444 273828
rect 224960 273776 225012 273828
rect 271512 273912 271564 273964
rect 280344 273912 280396 273964
rect 322756 273912 322808 273964
rect 330576 273912 330628 273964
rect 335268 273912 335320 273964
rect 348332 273912 348384 273964
rect 350356 273912 350408 273964
rect 368480 273912 368532 273964
rect 377772 273912 377824 273964
rect 408592 273912 408644 273964
rect 422116 273912 422168 273964
rect 472440 273912 472492 273964
rect 474648 273912 474700 273964
rect 545764 273912 545816 273964
rect 545948 273912 546000 273964
rect 639144 273912 639196 273964
rect 258080 273776 258132 273828
rect 259368 273776 259420 273828
rect 266360 273776 266412 273828
rect 397000 273776 397052 273828
rect 435824 273776 435876 273828
rect 438124 273776 438176 273828
rect 473636 273776 473688 273828
rect 481364 273776 481416 273828
rect 556344 273776 556396 273828
rect 556804 273776 556856 273828
rect 590660 273776 590712 273828
rect 119068 273640 119120 273692
rect 173256 273640 173308 273692
rect 447600 273640 447652 273692
rect 481916 273640 481968 273692
rect 484216 273640 484268 273692
rect 559932 273640 559984 273692
rect 132040 273504 132092 273556
rect 153844 273504 153896 273556
rect 440884 273504 440936 273556
rect 471244 273504 471296 273556
rect 476028 273504 476080 273556
rect 549260 273504 549312 273556
rect 549904 273504 549956 273556
rect 583576 273504 583628 273556
rect 145288 273368 145340 273420
rect 147864 273368 147916 273420
rect 478696 273368 478748 273420
rect 552848 273368 552900 273420
rect 327724 273232 327776 273284
rect 329472 273232 329524 273284
rect 42432 273164 42484 273216
rect 43260 273164 43312 273216
rect 108396 273164 108448 273216
rect 165896 273164 165948 273216
rect 186412 273164 186464 273216
rect 218704 273164 218756 273216
rect 362776 273164 362828 273216
rect 385868 273164 385920 273216
rect 400036 273164 400088 273216
rect 439320 273164 439372 273216
rect 444012 273164 444064 273216
rect 503168 273164 503220 273216
rect 504180 273164 504232 273216
rect 511448 273164 511500 273216
rect 102508 273028 102560 273080
rect 162860 273028 162912 273080
rect 172244 273028 172296 273080
rect 209780 273028 209832 273080
rect 219532 273028 219584 273080
rect 244556 273028 244608 273080
rect 280988 273028 281040 273080
rect 286324 273028 286376 273080
rect 361212 273028 361264 273080
rect 384948 273028 385000 273080
rect 385684 273028 385736 273080
rect 395620 273028 395672 273080
rect 404176 273028 404228 273080
rect 446496 273028 446548 273080
rect 446864 273028 446916 273080
rect 507952 273028 508004 273080
rect 509700 273028 509752 273080
rect 515220 273164 515272 273216
rect 515404 273164 515456 273216
rect 519728 273164 519780 273216
rect 521476 273164 521528 273216
rect 614304 273164 614356 273216
rect 513840 273028 513892 273080
rect 518532 273028 518584 273080
rect 94228 272892 94280 272944
rect 155960 272892 156012 272944
rect 166356 272892 166408 272944
rect 207296 272892 207348 272944
rect 211252 272892 211304 272944
rect 220084 272892 220136 272944
rect 220728 272892 220780 272944
rect 245752 272892 245804 272944
rect 247868 272892 247920 272944
rect 264244 272892 264296 272944
rect 333796 272892 333848 272944
rect 345940 272892 345992 272944
rect 348424 272892 348476 272944
rect 362500 272892 362552 272944
rect 365444 272892 365496 272944
rect 390928 272892 390980 272944
rect 405556 272892 405608 272944
rect 448796 272892 448848 272944
rect 455328 272892 455380 272944
rect 461400 272892 461452 272944
rect 82452 272756 82504 272808
rect 148416 272756 148468 272808
rect 155684 272756 155736 272808
rect 200120 272756 200172 272808
rect 205364 272756 205416 272808
rect 234804 272756 234856 272808
rect 245384 272756 245436 272808
rect 72976 272620 73028 272672
rect 142160 272620 142212 272672
rect 142712 272620 142764 272672
rect 145564 272620 145616 272672
rect 147404 272620 147456 272672
rect 193220 272620 193272 272672
rect 197084 272620 197136 272672
rect 229100 272620 229152 272672
rect 233700 272620 233752 272672
rect 254400 272620 254452 272672
rect 262312 272756 262364 272808
rect 270960 272756 271012 272808
rect 274272 272756 274324 272808
rect 282920 272756 282972 272808
rect 325332 272756 325384 272808
rect 332968 272756 333020 272808
rect 344652 272756 344704 272808
rect 361396 272756 361448 272808
rect 362224 272756 362276 272808
rect 370320 272756 370372 272808
rect 370504 272756 370556 272808
rect 396816 272756 396868 272808
rect 406844 272756 406896 272808
rect 449992 272756 450044 272808
rect 452292 272756 452344 272808
rect 515036 272892 515088 272944
rect 515220 272892 515272 272944
rect 569408 273028 569460 273080
rect 532516 272892 532568 272944
rect 262680 272620 262732 272672
rect 264428 272620 264480 272672
rect 276020 272620 276072 272672
rect 324044 272620 324096 272672
rect 331404 272620 331456 272672
rect 332324 272620 332376 272672
rect 343640 272620 343692 272672
rect 346216 272620 346268 272672
rect 363696 272620 363748 272672
rect 376116 272620 376168 272672
rect 406292 272620 406344 272672
rect 412272 272620 412324 272672
rect 456800 272620 456852 272672
rect 457168 272620 457220 272672
rect 461032 272620 461084 272672
rect 461400 272620 461452 272672
rect 513840 272756 513892 272808
rect 514024 272756 514076 272808
rect 525616 272756 525668 272808
rect 529848 272756 529900 272808
rect 532884 272756 532936 272808
rect 533712 272756 533764 272808
rect 538680 272756 538732 272808
rect 539048 272892 539100 272944
rect 624976 272892 625028 272944
rect 628472 272756 628524 272808
rect 461860 272620 461912 272672
rect 466414 272620 466466 272672
rect 522120 272620 522172 272672
rect 526812 272620 526864 272672
rect 621388 272620 621440 272672
rect 65892 272484 65944 272536
rect 136824 272484 136876 272536
rect 137928 272484 137980 272536
rect 116676 272348 116728 272400
rect 172520 272348 172572 272400
rect 181720 272484 181772 272536
rect 186964 272484 187016 272536
rect 195888 272484 195940 272536
rect 227904 272484 227956 272536
rect 228088 272484 228140 272536
rect 249064 272484 249116 272536
rect 254952 272484 255004 272536
rect 269304 272484 269356 272536
rect 270316 272484 270368 272536
rect 280528 272484 280580 272536
rect 329748 272484 329800 272536
rect 338856 272484 338908 272536
rect 339224 272484 339276 272536
rect 354220 272484 354272 272536
rect 354496 272484 354548 272536
rect 375564 272484 375616 272536
rect 379428 272484 379480 272536
rect 410984 272484 411036 272536
rect 416596 272484 416648 272536
rect 463700 272484 463752 272536
rect 470554 272484 470606 272536
rect 470692 272484 470744 272536
rect 532700 272484 532752 272536
rect 532884 272484 532936 272536
rect 538496 272484 538548 272536
rect 538680 272484 538732 272536
rect 632060 272892 632112 272944
rect 187700 272348 187752 272400
rect 194968 272348 195020 272400
rect 227168 272348 227220 272400
rect 318708 272348 318760 272400
rect 324688 272348 324740 272400
rect 395988 272348 396040 272400
rect 434628 272348 434680 272400
rect 449716 272348 449768 272400
rect 504180 272348 504232 272400
rect 504364 272348 504416 272400
rect 514024 272348 514076 272400
rect 517428 272348 517480 272400
rect 600964 272348 601016 272400
rect 601148 272348 601200 272400
rect 635556 272756 635608 272808
rect 634084 272620 634136 272672
rect 640340 272620 640392 272672
rect 127348 272212 127400 272264
rect 179880 272212 179932 272264
rect 189080 272212 189132 272264
rect 196440 272212 196492 272264
rect 391848 272212 391900 272264
rect 428740 272212 428792 272264
rect 450544 272212 450596 272264
rect 510252 272212 510304 272264
rect 520096 272212 520148 272264
rect 610716 272212 610768 272264
rect 145104 272076 145156 272128
rect 192392 272076 192444 272128
rect 384948 272076 385000 272128
rect 418068 272076 418120 272128
rect 428464 272076 428516 272128
rect 470554 272076 470606 272128
rect 470784 272076 470836 272128
rect 124956 271940 125008 271992
rect 151084 271940 151136 271992
rect 431684 271940 431736 271992
rect 480168 271940 480220 271992
rect 480536 272076 480588 272128
rect 547512 272076 547564 272128
rect 547696 272076 547748 272128
rect 504364 271940 504416 271992
rect 504548 271940 504600 271992
rect 562324 271940 562376 271992
rect 600964 272076 601016 272128
rect 607220 272076 607272 272128
rect 601148 271940 601200 271992
rect 106004 271804 106056 271856
rect 164976 271804 165028 271856
rect 174268 271804 174320 271856
rect 189264 271804 189316 271856
rect 202972 271804 203024 271856
rect 233240 271804 233292 271856
rect 274640 271804 274692 271856
rect 279240 271804 279292 271856
rect 355324 271804 355376 271856
rect 356612 271804 356664 271856
rect 375288 271804 375340 271856
rect 403900 271804 403952 271856
rect 433156 271804 433208 271856
rect 480168 271804 480220 271856
rect 480444 271804 480496 271856
rect 484860 271804 484912 271856
rect 97816 271668 97868 271720
rect 158812 271668 158864 271720
rect 169852 271668 169904 271720
rect 209964 271668 210016 271720
rect 225420 271668 225472 271720
rect 228364 271668 228416 271720
rect 351184 271668 351236 271720
rect 366088 271668 366140 271720
rect 382004 271668 382056 271720
rect 414572 271668 414624 271720
rect 430396 271668 430448 271720
rect 483572 271668 483624 271720
rect 485044 271668 485096 271720
rect 501420 271804 501472 271856
rect 496544 271668 496596 271720
rect 578516 271804 578568 271856
rect 578884 271804 578936 271856
rect 604828 271804 604880 271856
rect 504548 271668 504600 271720
rect 585968 271668 586020 271720
rect 87144 271532 87196 271584
rect 152004 271532 152056 271584
rect 165160 271532 165212 271584
rect 205640 271532 205692 271584
rect 215944 271532 215996 271584
rect 242072 271532 242124 271584
rect 337936 271532 337988 271584
rect 350724 271532 350776 271584
rect 360844 271532 360896 271584
rect 377588 271532 377640 271584
rect 387708 271532 387760 271584
rect 421656 271532 421708 271584
rect 437204 271532 437256 271584
rect 493692 271532 493744 271584
rect 499304 271532 499356 271584
rect 582380 271532 582432 271584
rect 583024 271532 583076 271584
rect 611636 271532 611688 271584
rect 612004 271532 612056 271584
rect 618996 271532 619048 271584
rect 75368 271396 75420 271448
rect 142712 271396 142764 271448
rect 162676 271396 162728 271448
rect 204720 271396 204772 271448
rect 213644 271396 213696 271448
rect 240416 271396 240468 271448
rect 240784 271396 240836 271448
rect 259644 271396 259696 271448
rect 260104 271396 260156 271448
rect 272616 271396 272668 271448
rect 325516 271396 325568 271448
rect 334164 271396 334216 271448
rect 347688 271396 347740 271448
rect 364892 271396 364944 271448
rect 366364 271396 366416 271448
rect 383844 271396 383896 271448
rect 384764 271396 384816 271448
rect 419264 271396 419316 271448
rect 420184 271396 420236 271448
rect 431132 271396 431184 271448
rect 439964 271396 440016 271448
rect 497280 271396 497332 271448
rect 501972 271396 502024 271448
rect 504548 271396 504600 271448
rect 505008 271396 505060 271448
rect 589464 271396 589516 271448
rect 589924 271396 589976 271448
rect 633256 271396 633308 271448
rect 76840 271260 76892 271312
rect 143540 271260 143592 271312
rect 152188 271260 152240 271312
rect 197360 271260 197412 271312
rect 198280 271260 198332 271312
rect 229560 271260 229612 271312
rect 235264 271260 235316 271312
rect 255320 271260 255372 271312
rect 256700 271260 256752 271312
rect 261024 271260 261076 271312
rect 262036 271260 262088 271312
rect 274640 271260 274692 271312
rect 329564 271260 329616 271312
rect 340052 271260 340104 271312
rect 340604 271260 340656 271312
rect 355140 271260 355192 271312
rect 357164 271260 357216 271312
rect 379060 271260 379112 271312
rect 390284 271260 390336 271312
rect 426348 271260 426400 271312
rect 68192 271124 68244 271176
rect 138480 271124 138532 271176
rect 141516 271124 141568 271176
rect 189080 271124 189132 271176
rect 191196 271124 191248 271176
rect 225144 271124 225196 271176
rect 230204 271124 230256 271176
rect 252008 271124 252060 271176
rect 268016 271124 268068 271176
rect 278780 271124 278832 271176
rect 279792 271124 279844 271176
rect 287060 271124 287112 271176
rect 331128 271124 331180 271176
rect 342444 271124 342496 271176
rect 343548 271124 343600 271176
rect 360200 271124 360252 271176
rect 364156 271124 364208 271176
rect 389732 271124 389784 271176
rect 394332 271124 394384 271176
rect 432236 271260 432288 271312
rect 442908 271260 442960 271312
rect 500868 271260 500920 271312
rect 507676 271260 507728 271312
rect 593052 271260 593104 271312
rect 598204 271260 598256 271312
rect 645032 271260 645084 271312
rect 113456 270988 113508 271040
rect 169944 270988 169996 271040
rect 187424 270988 187476 271040
rect 215944 270988 215996 271040
rect 251456 270988 251508 271040
rect 266912 270988 266964 271040
rect 417424 270988 417476 271040
rect 437940 271124 437992 271176
rect 441344 271124 441396 271176
rect 445024 271124 445076 271176
rect 445668 271124 445720 271176
rect 503996 271124 504048 271176
rect 524052 271124 524104 271176
rect 617340 271124 617392 271176
rect 617524 271124 617576 271176
rect 626080 271124 626132 271176
rect 427452 270988 427504 271040
rect 479156 270988 479208 271040
rect 480260 270988 480312 271040
rect 486608 270988 486660 271040
rect 495072 270988 495124 271040
rect 575296 270988 575348 271040
rect 123760 270852 123812 270904
rect 177488 270852 177540 270904
rect 407764 270852 407816 270904
rect 440516 270852 440568 270904
rect 449164 270852 449216 270904
rect 490196 270852 490248 270904
rect 492588 270852 492640 270904
rect 571708 270852 571760 270904
rect 134432 270716 134484 270768
rect 185124 270716 185176 270768
rect 321376 270716 321428 270768
rect 327080 270716 327132 270768
rect 414664 270716 414716 270768
rect 450820 270716 450872 270768
rect 486976 270716 487028 270768
rect 564624 270716 564676 270768
rect 567844 270716 567896 270768
rect 597744 270716 597796 270768
rect 121460 270580 121512 270632
rect 168104 270580 168156 270632
rect 403624 270580 403676 270632
rect 433432 270580 433484 270632
rect 453304 270580 453356 270632
rect 487804 270580 487856 270632
rect 489644 270580 489696 270632
rect 568212 270580 568264 270632
rect 84108 270444 84160 270496
rect 137468 270444 137520 270496
rect 137652 270444 137704 270496
rect 186136 270444 186188 270496
rect 200764 270444 200816 270496
rect 201868 270444 201920 270496
rect 206836 270444 206888 270496
rect 235816 270444 235868 270496
rect 278320 270444 278372 270496
rect 283840 270444 283892 270496
rect 400864 270444 400916 270496
rect 441620 270444 441672 270496
rect 456432 270444 456484 270496
rect 520280 270444 520332 270496
rect 523132 270444 523184 270496
rect 532884 270444 532936 270496
rect 78864 270308 78916 270360
rect 132500 270308 132552 270360
rect 133788 270308 133840 270360
rect 183652 270308 183704 270360
rect 185308 270308 185360 270360
rect 194416 270308 194468 270360
rect 199936 270308 199988 270360
rect 230848 270308 230900 270360
rect 232688 270308 232740 270360
rect 248236 270308 248288 270360
rect 283104 270308 283156 270360
rect 284668 270308 284720 270360
rect 355048 270308 355100 270360
rect 376944 270308 376996 270360
rect 379704 270308 379756 270360
rect 404360 270308 404412 270360
rect 415032 270308 415084 270360
rect 461216 270308 461268 270360
rect 461400 270308 461452 270360
rect 111984 270172 112036 270224
rect 168748 270172 168800 270224
rect 184848 270172 184900 270224
rect 219348 270172 219400 270224
rect 244372 270172 244424 270224
rect 262312 270172 262364 270224
rect 334348 270172 334400 270224
rect 346400 270172 346452 270224
rect 372252 270172 372304 270224
rect 397460 270172 397512 270224
rect 409604 270172 409656 270224
rect 454040 270172 454092 270224
rect 458824 270172 458876 270224
rect 524420 270172 524472 270224
rect 525616 270308 525668 270360
rect 619640 270444 619692 270496
rect 533528 270308 533580 270360
rect 626540 270308 626592 270360
rect 527180 270172 527232 270224
rect 528376 270172 528428 270224
rect 623964 270172 624016 270224
rect 89628 270036 89680 270088
rect 153016 270036 153068 270088
rect 176568 270036 176620 270088
rect 211160 270036 211212 270088
rect 212448 270036 212500 270088
rect 239956 270036 240008 270088
rect 241888 270036 241940 270088
rect 260656 270036 260708 270088
rect 266176 270036 266228 270088
rect 277216 270036 277268 270088
rect 345296 270036 345348 270088
rect 358820 270036 358872 270088
rect 366640 270036 366692 270088
rect 393320 270036 393372 270088
rect 394700 270036 394752 270088
rect 408776 270036 408828 270088
rect 412456 270036 412508 270088
rect 458180 270036 458232 270088
rect 463516 270036 463568 270088
rect 530768 270036 530820 270088
rect 530952 270036 531004 270088
rect 533160 270036 533212 270088
rect 85488 269900 85540 269952
rect 149428 269900 149480 269952
rect 152832 269900 152884 269952
rect 157156 269900 157208 269952
rect 173808 269900 173860 269952
rect 212632 269900 212684 269952
rect 226616 269900 226668 269952
rect 249892 269900 249944 269952
rect 256884 269900 256936 269952
rect 268936 269900 268988 269952
rect 330208 269900 330260 269952
rect 340880 269900 340932 269952
rect 341800 269900 341852 269952
rect 357440 269900 357492 269952
rect 359188 269900 359240 269952
rect 382280 269900 382332 269952
rect 383016 269900 383068 269952
rect 411260 269900 411312 269952
rect 419632 269900 419684 269952
rect 467932 269900 467984 269952
rect 468484 269900 468536 269952
rect 538312 270036 538364 270088
rect 533988 269900 534040 269952
rect 630680 270036 630732 270088
rect 540520 269900 540572 269952
rect 640524 269900 640576 269952
rect 70584 269764 70636 269816
rect 79324 269764 79376 269816
rect 80060 269764 80112 269816
rect 146392 269764 146444 269816
rect 158628 269764 158680 269816
rect 201040 269764 201092 269816
rect 201684 269764 201736 269816
rect 232504 269764 232556 269816
rect 237288 269764 237340 269816
rect 257344 269764 257396 269816
rect 258540 269764 258592 269816
rect 272248 269764 272300 269816
rect 273076 269764 273128 269816
rect 282184 269764 282236 269816
rect 326896 269764 326948 269816
rect 335544 269764 335596 269816
rect 336004 269764 336056 269816
rect 349160 269764 349212 269816
rect 351736 269764 351788 269816
rect 371240 269764 371292 269816
rect 376576 269764 376628 269816
rect 407120 269764 407172 269816
rect 417148 269764 417200 269816
rect 465080 269764 465132 269816
rect 466000 269764 466052 269816
rect 530400 269764 530452 269816
rect 122748 269628 122800 269680
rect 176200 269628 176252 269680
rect 183468 269628 183520 269680
rect 205456 269628 205508 269680
rect 392032 269628 392084 269680
rect 401692 269628 401744 269680
rect 404360 269628 404412 269680
rect 423680 269628 423732 269680
rect 423864 269628 423916 269680
rect 451372 269628 451424 269680
rect 453580 269628 453632 269680
rect 509240 269628 509292 269680
rect 538496 269764 538548 269816
rect 538680 269764 538732 269816
rect 541164 269764 541216 269816
rect 541348 269764 541400 269816
rect 637580 269764 637632 269816
rect 129648 269492 129700 269544
rect 181168 269492 181220 269544
rect 204168 269492 204220 269544
rect 223488 269492 223540 269544
rect 398748 269492 398800 269544
rect 412640 269492 412692 269544
rect 424600 269492 424652 269544
rect 475016 269492 475068 269544
rect 495256 269492 495308 269544
rect 532884 269628 532936 269680
rect 616420 269628 616472 269680
rect 509884 269492 509936 269544
rect 596180 269492 596232 269544
rect 126888 269356 126940 269408
rect 178684 269356 178736 269408
rect 408408 269356 408460 269408
rect 426532 269356 426584 269408
rect 441620 269356 441672 269408
rect 458456 269356 458508 269408
rect 470968 269356 471020 269408
rect 538312 269356 538364 269408
rect 538496 269356 538548 269408
rect 575480 269356 575532 269408
rect 143908 269220 143960 269272
rect 191104 269220 191156 269272
rect 282736 269220 282788 269272
rect 288808 269220 288860 269272
rect 401692 269220 401744 269272
rect 416780 269220 416832 269272
rect 474280 269220 474332 269272
rect 546500 269152 546552 269204
rect 319444 269084 319496 269136
rect 325700 269084 325752 269136
rect 118608 269016 118660 269068
rect 174544 269016 174596 269068
rect 175096 269016 175148 269068
rect 177672 269016 177724 269068
rect 273260 269016 273312 269068
rect 275560 269016 275612 269068
rect 433708 269016 433760 269068
rect 488540 269016 488592 269068
rect 493324 269016 493376 269068
rect 574100 269016 574152 269068
rect 115848 268880 115900 268932
rect 171232 268880 171284 268932
rect 382372 268880 382424 268932
rect 415400 268880 415452 268932
rect 436560 268880 436612 268932
rect 491668 268880 491720 268932
rect 498292 268880 498344 268932
rect 581000 268880 581052 268932
rect 110328 268744 110380 268796
rect 167920 268744 167972 268796
rect 168288 268744 168340 268796
rect 181996 268744 182048 268796
rect 188896 268744 188948 268796
rect 190460 268744 190512 268796
rect 200580 268744 200632 268796
rect 231308 268744 231360 268796
rect 387340 268744 387392 268796
rect 422300 268744 422352 268796
rect 438676 268744 438728 268796
rect 495440 268744 495492 268796
rect 500776 268744 500828 268796
rect 583760 268744 583812 268796
rect 104992 268608 105044 268660
rect 163780 268608 163832 268660
rect 176936 268608 176988 268660
rect 215116 268608 215168 268660
rect 224224 268608 224276 268660
rect 243268 268608 243320 268660
rect 352564 268608 352616 268660
rect 372620 268608 372672 268660
rect 393688 268608 393740 268660
rect 429200 268608 429252 268660
rect 441160 268608 441212 268660
rect 499580 268608 499632 268660
rect 503260 268608 503312 268660
rect 587900 268608 587952 268660
rect 99288 268472 99340 268524
rect 160468 268472 160520 268524
rect 180616 268472 180668 268524
rect 217600 268472 217652 268524
rect 231676 268472 231728 268524
rect 253204 268472 253256 268524
rect 338488 268472 338540 268524
rect 352104 268472 352156 268524
rect 367468 268472 367520 268524
rect 393504 268472 393556 268524
rect 397276 268472 397328 268524
rect 436100 268472 436152 268524
rect 446128 268472 446180 268524
rect 506480 268472 506532 268524
rect 508228 268472 508280 268524
rect 594800 268472 594852 268524
rect 92388 268336 92440 268388
rect 155500 268336 155552 268388
rect 161572 268336 161624 268388
rect 203524 268336 203576 268388
rect 210700 268336 210752 268388
rect 236644 268336 236696 268388
rect 252652 268336 252704 268388
rect 268108 268336 268160 268388
rect 348792 268336 348844 268388
rect 367100 268336 367152 268388
rect 372436 268336 372488 268388
rect 400496 268336 400548 268388
rect 402244 268336 402296 268388
rect 443092 268336 443144 268388
rect 461860 268336 461912 268388
rect 528560 268336 528612 268388
rect 541348 268336 541400 268388
rect 641720 268336 641772 268388
rect 135628 268200 135680 268252
rect 140136 268200 140188 268252
rect 140688 268200 140740 268252
rect 188620 268200 188672 268252
rect 416228 268200 416280 268252
rect 447140 268200 447192 268252
rect 448428 268200 448480 268252
rect 494060 268200 494112 268252
rect 495808 268200 495860 268252
rect 576860 268200 576912 268252
rect 151728 268064 151780 268116
rect 196072 268064 196124 268116
rect 422300 268064 422352 268116
rect 444380 268064 444432 268116
rect 527180 268064 527232 268116
rect 607404 268064 607456 268116
rect 490840 267928 490892 267980
rect 569960 267928 570012 267980
rect 276480 267724 276532 267776
rect 278044 267724 278096 267776
rect 119344 267656 119396 267708
rect 153476 267656 153528 267708
rect 153844 267656 153896 267708
rect 184480 267656 184532 267708
rect 365812 267656 365864 267708
rect 381544 267656 381596 267708
rect 388168 267656 388220 267708
rect 404360 267656 404412 267708
rect 408040 267656 408092 267708
rect 423864 267656 423916 267708
rect 445300 267656 445352 267708
rect 490564 267656 490616 267708
rect 509884 267656 509936 267708
rect 567844 267656 567896 267708
rect 111708 267520 111760 267572
rect 168564 267520 168616 267572
rect 169024 267520 169076 267572
rect 199384 267520 199436 267572
rect 215944 267520 215996 267572
rect 222568 267520 222620 267572
rect 371608 267520 371660 267572
rect 373264 267520 373316 267572
rect 390652 267520 390704 267572
rect 408408 267520 408460 267572
rect 421288 267520 421340 267572
rect 440884 267520 440936 267572
rect 447784 267520 447836 267572
rect 456064 267520 456116 267572
rect 460204 267520 460256 267572
rect 516784 267520 516836 267572
rect 519820 267520 519872 267572
rect 583024 267520 583076 267572
rect 86224 267384 86276 267436
rect 144736 267384 144788 267436
rect 145564 267384 145616 267436
rect 191932 267384 191984 267436
rect 199568 267384 199620 267436
rect 204352 267384 204404 267436
rect 205456 267384 205508 267436
rect 218428 267384 218480 267436
rect 233884 267384 233936 267436
rect 104808 267248 104860 267300
rect 164608 267248 164660 267300
rect 186964 267248 187016 267300
rect 219256 267248 219308 267300
rect 223488 267248 223540 267300
rect 234160 267248 234212 267300
rect 243544 267384 243596 267436
rect 251548 267384 251600 267436
rect 315304 267384 315356 267436
rect 319168 267384 319220 267436
rect 340972 267384 341024 267436
rect 355324 267384 355376 267436
rect 362500 267384 362552 267436
rect 369124 267384 369176 267436
rect 244096 267248 244148 267300
rect 321928 267248 321980 267300
rect 327724 267248 327776 267300
rect 350908 267248 350960 267300
rect 362224 267248 362276 267300
rect 90364 267112 90416 267164
rect 151360 267112 151412 267164
rect 168104 267112 168156 267164
rect 177028 267112 177080 267164
rect 177672 267112 177724 267164
rect 214288 267112 214340 267164
rect 220084 267112 220136 267164
rect 239128 267112 239180 267164
rect 246948 267112 247000 267164
rect 263968 267112 264020 267164
rect 312820 267112 312872 267164
rect 316040 267112 316092 267164
rect 360016 267112 360068 267164
rect 366364 267112 366416 267164
rect 79324 266976 79376 267028
rect 140136 266976 140188 267028
rect 186964 266976 187016 267028
rect 190460 266976 190512 267028
rect 224224 266976 224276 267028
rect 228364 266976 228416 267028
rect 140596 266840 140648 266892
rect 137468 266704 137520 266756
rect 150532 266840 150584 266892
rect 159456 266840 159508 266892
rect 162124 266840 162176 266892
rect 178868 266840 178920 266892
rect 209320 266840 209372 266892
rect 218704 266840 218756 266892
rect 220912 266840 220964 266892
rect 249064 266976 249116 267028
rect 250720 266976 250772 267028
rect 255964 266976 256016 267028
rect 259000 266976 259052 267028
rect 286324 266976 286376 267028
rect 287980 266976 288032 267028
rect 314476 266976 314528 267028
rect 318984 266976 319036 267028
rect 353392 266976 353444 267028
rect 374460 267384 374512 267436
rect 380716 267384 380768 267436
rect 398748 267384 398800 267436
rect 403072 267384 403124 267436
rect 422300 267384 422352 267436
rect 428740 267384 428792 267436
rect 447600 267384 447652 267436
rect 450268 267384 450320 267436
rect 498844 267384 498896 267436
rect 514852 267384 514904 267436
rect 578884 267384 578936 267436
rect 373264 267248 373316 267300
rect 392032 267248 392084 267300
rect 398104 267248 398156 267300
rect 417424 267248 417476 267300
rect 436744 267248 436796 267300
rect 457444 267248 457496 267300
rect 459376 267248 459428 267300
rect 460848 267248 460900 267300
rect 465172 267248 465224 267300
rect 523684 267248 523736 267300
rect 524788 267248 524840 267300
rect 612004 267248 612056 267300
rect 249064 266840 249116 266892
rect 332692 266840 332744 266892
rect 343824 266840 343876 266892
rect 368296 266840 368348 266892
rect 385684 267112 385736 267164
rect 393136 267112 393188 267164
rect 420184 267112 420236 267164
rect 432880 267112 432932 267164
rect 453304 267112 453356 267164
rect 455144 267112 455196 267164
rect 515404 267112 515456 267164
rect 517244 267112 517296 267164
rect 527180 267112 527232 267164
rect 529664 267112 529716 267164
rect 617524 267112 617576 267164
rect 383200 266976 383252 267028
rect 401692 266976 401744 267028
rect 413008 266976 413060 267028
rect 470140 266976 470192 267028
rect 534724 266976 534776 267028
rect 535552 266976 535604 267028
rect 536748 266976 536800 267028
rect 539692 266976 539744 267028
rect 634084 266976 634136 267028
rect 378232 266840 378284 266892
rect 394700 266840 394752 266892
rect 404728 266840 404780 266892
rect 416228 266840 416280 266892
rect 422944 266840 422996 266892
rect 438124 266840 438176 266892
rect 441620 266840 441672 266892
rect 442724 266840 442776 266892
rect 485044 266840 485096 266892
rect 499948 266840 500000 266892
rect 507860 266840 507912 266892
rect 534724 266840 534776 266892
rect 589924 266840 589976 266892
rect 316960 266772 317012 266824
rect 321560 266772 321612 266824
rect 151084 266704 151136 266756
rect 179512 266704 179564 266756
rect 394792 266704 394844 266756
rect 403624 266704 403676 266756
rect 407212 266704 407264 266756
rect 414664 266704 414716 266756
rect 308680 266636 308732 266688
rect 310520 266636 310572 266688
rect 313648 266636 313700 266688
rect 317420 266636 317472 266688
rect 317788 266636 317840 266688
rect 322940 266636 322992 266688
rect 347504 266636 347556 266688
rect 351184 266636 351236 266688
rect 427912 266636 427964 266688
rect 436744 266636 436796 266688
rect 449164 266704 449216 266756
rect 457720 266704 457772 266756
rect 476764 266704 476816 266756
rect 485044 266704 485096 266756
rect 130384 266568 130436 266620
rect 138112 266568 138164 266620
rect 149612 266568 149664 266620
rect 159640 266568 159692 266620
rect 399760 266568 399812 266620
rect 407764 266568 407816 266620
rect 310336 266500 310388 266552
rect 311900 266500 311952 266552
rect 312268 266500 312320 266552
rect 314660 266500 314712 266552
rect 316132 266500 316184 266552
rect 320180 266500 320232 266552
rect 327724 266500 327776 266552
rect 331864 266500 331916 266552
rect 345112 266500 345164 266552
rect 348424 266500 348476 266552
rect 350080 266500 350132 266552
rect 353944 266500 353996 266552
rect 355876 266500 355928 266552
rect 360844 266500 360896 266552
rect 369952 266500 370004 266552
rect 372252 266500 372304 266552
rect 374920 266500 374972 266552
rect 379704 266500 379756 266552
rect 423772 266500 423824 266552
rect 425704 266500 425756 266552
rect 426256 266500 426308 266552
rect 428464 266500 428516 266552
rect 434536 266500 434588 266552
rect 452752 266568 452804 266620
rect 462964 266568 463016 266620
rect 490012 266704 490064 266756
rect 509700 266704 509752 266756
rect 510712 266704 510764 266756
rect 511816 266704 511868 266756
rect 512368 266704 512420 266756
rect 513196 266704 513248 266756
rect 516508 266704 516560 266756
rect 517428 266704 517480 266756
rect 518992 266704 519044 266756
rect 520096 266704 520148 266756
rect 527272 266704 527324 266756
rect 528192 266704 528244 266756
rect 528928 266704 528980 266756
rect 529848 266704 529900 266756
rect 531412 266704 531464 266756
rect 532516 266704 532568 266756
rect 533068 266704 533120 266756
rect 533988 266704 534040 266756
rect 543004 266704 543056 266756
rect 598204 266704 598256 266756
rect 501604 266568 501656 266620
rect 504824 266568 504876 266620
rect 556804 266568 556856 266620
rect 437848 266500 437900 266552
rect 448428 266500 448480 266552
rect 132500 266432 132552 266484
rect 147220 266432 147272 266484
rect 491668 266432 491720 266484
rect 492588 266432 492640 266484
rect 494152 266432 494204 266484
rect 495072 266432 495124 266484
rect 502432 266432 502484 266484
rect 503444 266432 503496 266484
rect 504088 266432 504140 266484
rect 505008 266432 505060 266484
rect 506572 266432 506624 266484
rect 507676 266432 507728 266484
rect 507860 266432 507912 266484
rect 549904 266432 549956 266484
rect 163504 266364 163556 266416
rect 167092 266364 167144 266416
rect 168564 266364 168616 266416
rect 169576 266364 169628 266416
rect 211160 266364 211212 266416
rect 213460 266364 213512 266416
rect 214564 266364 214616 266416
rect 215944 266364 215996 266416
rect 239404 266364 239456 266416
rect 241612 266364 241664 266416
rect 243728 266364 243780 266416
rect 246580 266364 246632 266416
rect 250444 266364 250496 266416
rect 256516 266364 256568 266416
rect 300952 266364 301004 266416
rect 302056 266364 302108 266416
rect 303712 266364 303764 266416
rect 304540 266364 304592 266416
rect 307852 266364 307904 266416
rect 309140 266364 309192 266416
rect 309508 266364 309560 266416
rect 310704 266364 310756 266416
rect 311164 266364 311216 266416
rect 313280 266364 313332 266416
rect 320272 266364 320324 266416
rect 321376 266364 321428 266416
rect 324412 266364 324464 266416
rect 325332 266364 325384 266416
rect 328552 266364 328604 266416
rect 329748 266364 329800 266416
rect 336832 266364 336884 266416
rect 337936 266364 337988 266416
rect 342628 266364 342680 266416
rect 345296 266364 345348 266416
rect 346768 266364 346820 266416
rect 347688 266364 347740 266416
rect 349252 266364 349304 266416
rect 350356 266364 350408 266416
rect 357532 266364 357584 266416
rect 359464 266364 359516 266416
rect 361672 266364 361724 266416
rect 362776 266364 362828 266416
rect 369124 266364 369176 266416
rect 370504 266364 370556 266416
rect 374092 266364 374144 266416
rect 375288 266364 375340 266416
rect 379888 266364 379940 266416
rect 383016 266364 383068 266416
rect 384028 266364 384080 266416
rect 384948 266364 385000 266416
rect 386512 266364 386564 266416
rect 387708 266364 387760 266416
rect 392308 266364 392360 266416
rect 393688 266364 393740 266416
rect 398932 266364 398984 266416
rect 400036 266364 400088 266416
rect 408868 266364 408920 266416
rect 409788 266364 409840 266416
rect 411352 266364 411404 266416
rect 412272 266364 412324 266416
rect 415492 266364 415544 266416
rect 416412 266364 416464 266416
rect 417976 266364 418028 266416
rect 418804 266364 418856 266416
rect 425428 266364 425480 266416
rect 427084 266364 427136 266416
rect 429568 266364 429620 266416
rect 430396 266364 430448 266416
rect 432052 266364 432104 266416
rect 433156 266364 433208 266416
rect 440332 266364 440384 266416
rect 441344 266364 441396 266416
rect 441988 266364 442040 266416
rect 442908 266364 442960 266416
rect 444472 266364 444524 266416
rect 445668 266364 445720 266416
rect 448612 266364 448664 266416
rect 450544 266364 450596 266416
rect 454408 266364 454460 266416
rect 455328 266364 455380 266416
rect 473452 266364 473504 266416
rect 474648 266364 474700 266416
rect 475108 266364 475160 266416
rect 479524 266364 479576 266416
rect 481732 266364 481784 266416
rect 482836 266364 482888 266416
rect 483388 266364 483440 266416
rect 484216 266364 484268 266416
rect 485872 266364 485924 266416
rect 486792 266364 486844 266416
rect 487160 266296 487212 266348
rect 557724 266296 557776 266348
rect 484216 266160 484268 266212
rect 560300 266160 560352 266212
rect 482560 266024 482612 266076
rect 487160 266024 487212 266076
rect 492496 266024 492548 266076
rect 572720 266024 572772 266076
rect 513196 265888 513248 265940
rect 601700 265888 601752 265940
rect 515680 265752 515732 265804
rect 605840 265752 605892 265804
rect 189080 265616 189132 265668
rect 189908 265616 189960 265668
rect 209780 265616 209832 265668
rect 210700 265616 210752 265668
rect 224960 265616 225012 265668
rect 225604 265616 225656 265668
rect 280344 265616 280396 265668
rect 280988 265616 281040 265668
rect 292672 265616 292724 265668
rect 293500 265616 293552 265668
rect 296812 265616 296864 265668
rect 297548 265616 297600 265668
rect 520648 265616 520700 265668
rect 612740 265616 612792 265668
rect 479248 265480 479300 265532
rect 553400 265480 553452 265532
rect 477592 265344 477644 265396
rect 550640 265344 550692 265396
rect 469312 265208 469364 265260
rect 539968 265208 540020 265260
rect 466828 265072 466880 265124
rect 535736 265072 535788 265124
rect 58624 264324 58676 264376
rect 668124 264324 668176 264376
rect 46204 264188 46256 264240
rect 669228 264188 669280 264240
rect 570604 261468 570656 261520
rect 645860 261468 645912 261520
rect 554412 260856 554464 260908
rect 568580 260856 568632 260908
rect 554320 259428 554372 259480
rect 563704 259428 563756 259480
rect 675852 258748 675904 258800
rect 676404 258748 676456 258800
rect 35808 256912 35860 256964
rect 39488 256912 39540 256964
rect 35624 256708 35676 256760
rect 41696 256708 41748 256760
rect 42064 256708 42116 256760
rect 43352 256708 43404 256760
rect 553952 256708 554004 256760
rect 560944 256708 560996 256760
rect 554504 255552 554556 255604
rect 558184 255552 558236 255604
rect 35808 255416 35860 255468
rect 40224 255416 40276 255468
rect 51724 254532 51776 254584
rect 62396 254532 62448 254584
rect 35624 252696 35676 252748
rect 40684 252696 40736 252748
rect 35808 252560 35860 252612
rect 41328 252560 41380 252612
rect 554412 252560 554464 252612
rect 562324 252560 562376 252612
rect 35808 251200 35860 251252
rect 39304 251200 39356 251252
rect 554136 251200 554188 251252
rect 556804 251200 556856 251252
rect 35624 250044 35676 250096
rect 40132 250044 40184 250096
rect 35808 249772 35860 249824
rect 41696 249772 41748 249824
rect 42064 249772 42116 249824
rect 42984 249772 43036 249824
rect 674932 249704 674984 249756
rect 675484 249704 675536 249756
rect 674932 249160 674984 249212
rect 674932 249024 674984 249076
rect 35808 247256 35860 247308
rect 39856 247256 39908 247308
rect 559564 246304 559616 246356
rect 647240 246304 647292 246356
rect 553860 245624 553912 245676
rect 596824 245624 596876 245676
rect 674840 245420 674892 245472
rect 675208 245420 675260 245472
rect 553492 244264 553544 244316
rect 555424 244264 555476 244316
rect 39304 242700 39356 242752
rect 41696 242700 41748 242752
rect 42064 242632 42116 242684
rect 42524 242632 42576 242684
rect 34428 242156 34480 242208
rect 41696 242156 41748 242208
rect 576124 242156 576176 242208
rect 648620 242156 648672 242208
rect 553676 241476 553728 241528
rect 629944 241476 629996 241528
rect 554504 240116 554556 240168
rect 577504 240116 577556 240168
rect 554320 238688 554372 238740
rect 576124 238688 576176 238740
rect 672264 236988 672316 237040
rect 671252 236852 671304 236904
rect 553768 236784 553820 236836
rect 559564 236784 559616 236836
rect 672954 236648 673006 236700
rect 671712 236444 671764 236496
rect 673184 236444 673236 236496
rect 671068 235900 671120 235952
rect 673414 235832 673466 235884
rect 672080 235696 672132 235748
rect 673184 235492 673236 235544
rect 673000 235016 673052 235068
rect 673460 234812 673512 234864
rect 674088 234676 674140 234728
rect 554412 234540 554464 234592
rect 570604 234540 570656 234592
rect 669780 234540 669832 234592
rect 669596 234132 669648 234184
rect 675852 233996 675904 234048
rect 678244 233996 678296 234048
rect 652392 233860 652444 233912
rect 670884 233928 670936 233980
rect 671372 233724 671424 233776
rect 674104 233724 674156 233776
rect 672264 233248 672316 233300
rect 673184 233248 673236 233300
rect 670884 233180 670936 233232
rect 672080 233180 672132 233232
rect 673460 233180 673512 233232
rect 674288 233180 674340 233232
rect 670332 233044 670384 233096
rect 673000 233044 673052 233096
rect 663064 232636 663116 232688
rect 674104 232636 674156 232688
rect 675852 232636 675904 232688
rect 683212 232636 683264 232688
rect 653404 232500 653456 232552
rect 676036 232500 676088 232552
rect 683396 232500 683448 232552
rect 674104 232364 674156 232416
rect 666284 231548 666336 231600
rect 674840 231548 674892 231600
rect 134984 231412 135036 231464
rect 137652 231412 137704 231464
rect 61384 231276 61436 231328
rect 668860 231276 668912 231328
rect 92388 231140 92440 231192
rect 170772 231140 170824 231192
rect 665088 231140 665140 231192
rect 128268 231004 128320 231056
rect 195888 231004 195940 231056
rect 666468 230936 666520 230988
rect 104808 230868 104860 230920
rect 179144 230868 179196 230920
rect 674840 230800 674892 230852
rect 118608 230732 118660 230784
rect 188160 230732 188212 230784
rect 94504 230596 94556 230648
rect 171416 230596 171468 230648
rect 194416 230596 194468 230648
rect 196900 230596 196952 230648
rect 672080 230596 672132 230648
rect 439320 230528 439372 230580
rect 137652 230460 137704 230512
rect 201040 230460 201092 230512
rect 42156 230392 42208 230444
rect 43260 230392 43312 230444
rect 133788 230392 133840 230444
rect 137468 230392 137520 230444
rect 213092 230392 213144 230444
rect 261576 230392 261628 230444
rect 311992 230392 312044 230444
rect 313096 230392 313148 230444
rect 374644 230392 374696 230444
rect 376208 230392 376260 230444
rect 433432 230392 433484 230444
rect 434168 230392 434220 230444
rect 440700 230392 440752 230444
rect 441896 230392 441948 230444
rect 443460 230392 443512 230444
rect 451556 230392 451608 230444
rect 453304 230392 453356 230444
rect 532516 230392 532568 230444
rect 538312 230392 538364 230444
rect 673276 230392 673328 230444
rect 387432 230324 387484 230376
rect 388444 230324 388496 230376
rect 398104 230324 398156 230376
rect 399392 230324 399444 230376
rect 436100 230324 436152 230376
rect 436744 230324 436796 230376
rect 438676 230324 438728 230376
rect 439320 230324 439372 230376
rect 443828 230324 443880 230376
rect 444932 230324 444984 230376
rect 455420 230324 455472 230376
rect 457168 230324 457220 230376
rect 463792 230324 463844 230376
rect 465724 230324 465776 230376
rect 470876 230324 470928 230376
rect 471888 230324 471940 230376
rect 476028 230324 476080 230376
rect 478604 230324 478656 230376
rect 493416 230324 493468 230376
rect 496360 230324 496412 230376
rect 497280 230324 497332 230376
rect 498108 230324 498160 230376
rect 510804 230324 510856 230376
rect 511908 230324 511960 230376
rect 521108 230324 521160 230376
rect 526444 230324 526496 230376
rect 530124 230324 530176 230376
rect 531136 230324 531188 230376
rect 126888 230256 126940 230308
rect 194416 230256 194468 230308
rect 194876 230256 194928 230308
rect 195428 230256 195480 230308
rect 195612 230256 195664 230308
rect 204904 230256 204956 230308
rect 206284 230256 206336 230308
rect 256424 230256 256476 230308
rect 256608 230256 256660 230308
rect 297640 230256 297692 230308
rect 297824 230256 297876 230308
rect 323400 230256 323452 230308
rect 444472 230188 444524 230240
rect 447600 230188 447652 230240
rect 452844 230188 452896 230240
rect 454316 230188 454368 230240
rect 468300 230188 468352 230240
rect 469128 230188 469180 230240
rect 487620 230188 487672 230240
rect 488448 230188 488500 230240
rect 95240 230120 95292 230172
rect 165988 230120 166040 230172
rect 166264 230120 166316 230172
rect 185584 230120 185636 230172
rect 186044 230120 186096 230172
rect 235816 230120 235868 230172
rect 240324 230120 240376 230172
rect 282184 230120 282236 230172
rect 282644 230120 282696 230172
rect 307944 230120 307996 230172
rect 308128 230120 308180 230172
rect 334992 230120 335044 230172
rect 335176 230120 335228 230172
rect 350448 230120 350500 230172
rect 454132 230052 454184 230104
rect 455328 230052 455380 230104
rect 82084 229984 82136 230036
rect 86224 229984 86276 230036
rect 137284 229984 137336 230036
rect 137468 229984 137520 230036
rect 195060 229984 195112 230036
rect 195428 229984 195480 230036
rect 215208 229984 215260 230036
rect 230480 229984 230532 230036
rect 277032 229984 277084 230036
rect 277216 229984 277268 230036
rect 302792 229984 302844 230036
rect 303252 229984 303304 230036
rect 329840 229984 329892 230036
rect 330944 229984 330996 230036
rect 355600 229984 355652 230036
rect 448336 229984 448388 230036
rect 448980 229984 449032 230036
rect 484400 229984 484452 230036
rect 495164 230188 495216 230240
rect 511448 230188 511500 230240
rect 517520 230188 517572 230240
rect 530768 230188 530820 230240
rect 539600 230256 539652 230308
rect 673460 230188 673512 230240
rect 532700 230120 532752 230172
rect 547144 230120 547196 230172
rect 491484 230052 491536 230104
rect 492496 230052 492548 230104
rect 528836 230052 528888 230104
rect 532516 230052 532568 230104
rect 560944 230052 560996 230104
rect 568120 230052 568172 230104
rect 517244 229984 517296 230036
rect 524604 229984 524656 230036
rect 534632 229984 534684 230036
rect 550548 229984 550600 230036
rect 674104 229984 674156 230036
rect 453488 229916 453540 229968
rect 455788 229916 455840 229968
rect 151728 229848 151780 229900
rect 151912 229848 151964 229900
rect 166264 229848 166316 229900
rect 68284 229712 68336 229764
rect 144460 229712 144512 229764
rect 144828 229712 144880 229764
rect 146300 229712 146352 229764
rect 137284 229576 137336 229628
rect 154028 229712 154080 229764
rect 154212 229712 154264 229764
rect 161388 229712 161440 229764
rect 151176 229576 151228 229628
rect 161756 229712 161808 229764
rect 163964 229712 164016 229764
rect 225512 229848 225564 229900
rect 225696 229848 225748 229900
rect 271880 229848 271932 229900
rect 275652 229848 275704 229900
rect 311992 229848 312044 229900
rect 312636 229848 312688 229900
rect 340144 229848 340196 229900
rect 345664 229848 345716 229900
rect 360752 229848 360804 229900
rect 361212 229848 361264 229900
rect 378784 229848 378836 229900
rect 449624 229848 449676 229900
rect 450544 229848 450596 229900
rect 467012 229848 467064 229900
rect 474004 229848 474056 229900
rect 476672 229848 476724 229900
rect 481640 229848 481692 229900
rect 481824 229848 481876 229900
rect 493600 229848 493652 229900
rect 495992 229848 496044 229900
rect 506388 229848 506440 229900
rect 507584 229848 507636 229900
rect 516784 229848 516836 229900
rect 519176 229848 519228 229900
rect 528560 229848 528612 229900
rect 536564 229848 536616 229900
rect 559564 229848 559616 229900
rect 674104 229780 674156 229832
rect 173716 229712 173768 229764
rect 175924 229712 175976 229764
rect 176384 229712 176436 229764
rect 185400 229712 185452 229764
rect 185584 229712 185636 229764
rect 194876 229712 194928 229764
rect 195060 229712 195112 229764
rect 202328 229712 202380 229764
rect 204904 229712 204956 229764
rect 246120 229712 246172 229764
rect 246488 229712 246540 229764
rect 287336 229712 287388 229764
rect 287704 229712 287756 229764
rect 318248 229712 318300 229764
rect 161756 229576 161808 229628
rect 220360 229576 220412 229628
rect 102140 229440 102192 229492
rect 145656 229440 145708 229492
rect 146024 229372 146076 229424
rect 150992 229508 151044 229560
rect 151774 229440 151826 229492
rect 210056 229440 210108 229492
rect 220452 229440 220504 229492
rect 251272 229576 251324 229628
rect 251732 229576 251784 229628
rect 292488 229576 292540 229628
rect 318064 229576 318116 229628
rect 345296 229712 345348 229764
rect 351736 229712 351788 229764
rect 371056 229712 371108 229764
rect 377680 229712 377732 229764
rect 389088 229712 389140 229764
rect 399852 229712 399904 229764
rect 409696 229712 409748 229764
rect 410892 229712 410944 229764
rect 417424 229712 417476 229764
rect 457352 229712 457404 229764
rect 463884 229712 463936 229764
rect 465448 229712 465500 229764
rect 467472 229712 467524 229764
rect 469588 229712 469640 229764
rect 476764 229712 476816 229764
rect 479248 229712 479300 229764
rect 489920 229712 489972 229764
rect 492128 229712 492180 229764
rect 507124 229712 507176 229764
rect 523040 229712 523092 229764
rect 534724 229712 534776 229764
rect 538496 229712 538548 229764
rect 566832 229712 566884 229764
rect 663708 229712 663760 229764
rect 672080 229712 672132 229764
rect 509516 229644 509568 229696
rect 515496 229644 515548 229696
rect 388628 229576 388680 229628
rect 398748 229576 398800 229628
rect 526904 229576 526956 229628
rect 536104 229576 536156 229628
rect 673368 229576 673420 229628
rect 449256 229508 449308 229560
rect 451924 229508 451976 229560
rect 148324 229372 148376 229424
rect 151636 229372 151688 229424
rect 110328 229304 110380 229356
rect 145840 229304 145892 229356
rect 123484 229168 123536 229220
rect 153384 229304 153436 229356
rect 153844 229304 153896 229356
rect 157800 229304 157852 229356
rect 157984 229304 158036 229356
rect 163688 229304 163740 229356
rect 164240 229304 164292 229356
rect 169116 229304 169168 229356
rect 170956 229304 171008 229356
rect 230664 229304 230716 229356
rect 413836 229304 413888 229356
rect 420000 229304 420052 229356
rect 472164 229304 472216 229356
rect 472992 229304 473044 229356
rect 674104 229304 674156 229356
rect 446404 229236 446456 229288
rect 448612 229236 448664 229288
rect 450268 229236 450320 229288
rect 451740 229236 451792 229288
rect 495348 229236 495400 229288
rect 500224 229236 500276 229288
rect 505652 229236 505704 229288
rect 510620 229236 510672 229288
rect 513380 229236 513432 229288
rect 519176 229236 519228 229288
rect 660948 229236 661000 229288
rect 666284 229236 666336 229288
rect 151912 229168 151964 229220
rect 155960 229168 156012 229220
rect 157248 229168 157300 229220
rect 161296 229168 161348 229220
rect 161480 229168 161532 229220
rect 173716 229168 173768 229220
rect 173900 229168 173952 229220
rect 174820 229168 174872 229220
rect 175924 229168 175976 229220
rect 180432 229168 180484 229220
rect 183376 229168 183428 229220
rect 240968 229168 241020 229220
rect 423496 229100 423548 229152
rect 427728 229100 427780 229152
rect 441252 229100 441304 229152
rect 442080 229100 442132 229152
rect 450912 229100 450964 229152
rect 452752 229100 452804 229152
rect 503720 229100 503772 229152
rect 509884 229100 509936 229152
rect 515312 229100 515364 229152
rect 520924 229100 520976 229152
rect 524972 229100 525024 229152
rect 529940 229100 529992 229152
rect 662328 229100 662380 229152
rect 666468 229100 666520 229152
rect 673552 229100 673604 229152
rect 100668 229032 100720 229084
rect 174636 229032 174688 229084
rect 174820 229032 174872 229084
rect 179788 229032 179840 229084
rect 180064 229032 180116 229084
rect 185584 229032 185636 229084
rect 189724 229032 189776 229084
rect 106188 228896 106240 228948
rect 173900 228896 173952 228948
rect 93584 228760 93636 228812
rect 161434 228760 161486 228812
rect 161572 228760 161624 228812
rect 166540 228760 166592 228812
rect 184940 228896 184992 228948
rect 185400 228896 185452 228948
rect 190092 228896 190144 228948
rect 192852 229032 192904 229084
rect 195244 229032 195296 229084
rect 201408 229032 201460 229084
rect 252560 229032 252612 229084
rect 255228 229032 255280 229084
rect 295708 229032 295760 229084
rect 305552 229032 305604 229084
rect 315672 229032 315724 229084
rect 326896 229032 326948 229084
rect 351092 229032 351144 229084
rect 195244 228896 195296 228948
rect 195428 228896 195480 228948
rect 246764 228896 246816 228948
rect 248236 228896 248288 228948
rect 291844 228896 291896 228948
rect 302148 228896 302200 228948
rect 331220 228896 331272 228948
rect 506388 228896 506440 228948
rect 512736 228896 512788 228948
rect 526444 228896 526496 228948
rect 544016 228896 544068 228948
rect 176108 228760 176160 228812
rect 231308 228760 231360 228812
rect 238576 228760 238628 228812
rect 282828 228760 282880 228812
rect 291844 228760 291896 228812
rect 300216 228760 300268 228812
rect 300676 228760 300728 228812
rect 330484 228760 330536 228812
rect 376024 228760 376076 228812
rect 387800 228760 387852 228812
rect 478880 228760 478932 228812
rect 490380 228760 490432 228812
rect 499856 228760 499908 228812
rect 518164 228760 518216 228812
rect 518532 228760 518584 228812
rect 541532 228760 541584 228812
rect 67548 228624 67600 228676
rect 146208 228624 146260 228676
rect 61384 228488 61436 228540
rect 57244 228352 57296 228404
rect 136824 228352 136876 228404
rect 137376 228488 137428 228540
rect 165988 228624 166040 228676
rect 181444 228624 181496 228676
rect 181628 228624 181680 228676
rect 185400 228624 185452 228676
rect 185584 228624 185636 228676
rect 226156 228624 226208 228676
rect 226340 228624 226392 228676
rect 272524 228624 272576 228676
rect 296628 228624 296680 228676
rect 329196 228624 329248 228676
rect 336464 228624 336516 228676
rect 358820 228624 358872 228676
rect 359924 228624 359976 228676
rect 376852 228624 376904 228676
rect 485688 228624 485740 228676
rect 498292 228624 498344 228676
rect 498568 228624 498620 228676
rect 515772 228624 515824 228676
rect 517888 228624 517940 228676
rect 539416 228624 539468 228676
rect 539600 228624 539652 228676
rect 556988 228624 557040 228676
rect 147128 228488 147180 228540
rect 200120 228488 200172 228540
rect 200304 228488 200356 228540
rect 221004 228488 221056 228540
rect 112996 228216 113048 228268
rect 137192 228216 137244 228268
rect 139308 228352 139360 228404
rect 143080 228216 143132 228268
rect 143448 228216 143500 228268
rect 146024 228216 146076 228268
rect 146208 228216 146260 228268
rect 148876 228216 148928 228268
rect 153476 228352 153528 228404
rect 154212 228352 154264 228404
rect 154396 228352 154448 228404
rect 215852 228352 215904 228404
rect 216404 228352 216456 228404
rect 264796 228488 264848 228540
rect 272524 228488 272576 228540
rect 309876 228488 309928 228540
rect 313832 228488 313884 228540
rect 320824 228488 320876 228540
rect 325424 228488 325476 228540
rect 349160 228488 349212 228540
rect 350448 228488 350500 228540
rect 369124 228488 369176 228540
rect 371056 228488 371108 228540
rect 385224 228488 385276 228540
rect 386052 228488 386104 228540
rect 397460 228488 397512 228540
rect 224776 228352 224828 228404
rect 273812 228352 273864 228404
rect 285588 228352 285640 228404
rect 318892 228352 318944 228404
rect 330484 228352 330536 228404
rect 354956 228352 355008 228404
rect 355324 228352 355376 228404
rect 372988 228352 373040 228404
rect 373448 228352 373500 228404
rect 387156 228352 387208 228404
rect 390008 228352 390060 228404
rect 400036 228352 400088 228404
rect 205548 228216 205600 228268
rect 205732 228216 205784 228268
rect 257068 228216 257120 228268
rect 257620 228216 257672 228268
rect 296352 228216 296404 228268
rect 407764 228488 407816 228540
rect 409788 228488 409840 228540
rect 415492 228488 415544 228540
rect 485044 228488 485096 228540
rect 498660 228488 498712 228540
rect 502432 228488 502484 228540
rect 521108 228488 521160 228540
rect 527548 228488 527600 228540
rect 553308 228488 553360 228540
rect 556804 228488 556856 228540
rect 570604 228488 570656 228540
rect 402796 228352 402848 228404
rect 411628 228352 411680 228404
rect 474464 228352 474516 228404
rect 484492 228352 484544 228404
rect 490196 228352 490248 228404
rect 505192 228352 505244 228404
rect 512092 228352 512144 228404
rect 532976 228352 533028 228404
rect 537208 228352 537260 228404
rect 565636 228352 565688 228404
rect 539416 228216 539468 228268
rect 540796 228216 540848 228268
rect 119988 228080 120040 228132
rect 181260 228080 181312 228132
rect 181444 228080 181496 228132
rect 126704 227944 126756 227996
rect 192852 227944 192904 227996
rect 195244 228080 195296 228132
rect 239036 228080 239088 228132
rect 246304 228080 246356 228132
rect 253848 228080 253900 228132
rect 268936 228080 268988 228132
rect 306012 228080 306064 228132
rect 400128 228080 400180 228132
rect 415032 228012 415084 228064
rect 421932 228012 421984 228064
rect 200304 227944 200356 227996
rect 210424 227944 210476 227996
rect 238392 227944 238444 227996
rect 416688 227876 416740 227928
rect 420644 227876 420696 227928
rect 447048 227876 447100 227928
rect 450544 227876 450596 227928
rect 88248 227808 88300 227860
rect 95240 227808 95292 227860
rect 133512 227808 133564 227860
rect 136640 227808 136692 227860
rect 136824 227808 136876 227860
rect 141148 227808 141200 227860
rect 141516 227808 141568 227860
rect 200488 227808 200540 227860
rect 200672 227808 200724 227860
rect 210240 227808 210292 227860
rect 409052 227740 409104 227792
rect 410340 227740 410392 227792
rect 411904 227740 411956 227792
rect 413560 227740 413612 227792
rect 420644 227740 420696 227792
rect 423864 227740 423916 227792
rect 471520 227740 471572 227792
rect 479524 227740 479576 227792
rect 662052 227740 662104 227792
rect 663892 227740 663944 227792
rect 42432 227672 42484 227724
rect 43076 227672 43128 227724
rect 64788 227672 64840 227724
rect 110328 227672 110380 227724
rect 110512 227672 110564 227724
rect 182364 227672 182416 227724
rect 185400 227672 185452 227724
rect 192668 227672 192720 227724
rect 60648 227536 60700 227588
rect 102140 227536 102192 227588
rect 103428 227536 103480 227588
rect 175372 227536 175424 227588
rect 181536 227536 181588 227588
rect 96436 227400 96488 227452
rect 170772 227400 170824 227452
rect 171094 227400 171146 227452
rect 175924 227468 175976 227520
rect 185584 227400 185636 227452
rect 186136 227536 186188 227588
rect 214380 227672 214432 227724
rect 214748 227672 214800 227724
rect 262220 227672 262272 227724
rect 277032 227672 277084 227724
rect 311808 227672 311860 227724
rect 465908 227604 465960 227656
rect 469864 227604 469916 227656
rect 200212 227536 200264 227588
rect 251916 227536 251968 227588
rect 259276 227536 259328 227588
rect 298284 227536 298336 227588
rect 301504 227536 301556 227588
rect 308588 227536 308640 227588
rect 524604 227536 524656 227588
rect 539968 227536 540020 227588
rect 219900 227400 219952 227452
rect 220084 227400 220136 227452
rect 241612 227400 241664 227452
rect 257804 227400 257856 227452
rect 299572 227400 299624 227452
rect 304908 227400 304960 227452
rect 333704 227400 333756 227452
rect 333888 227400 333940 227452
rect 356244 227400 356296 227452
rect 357072 227400 357124 227452
rect 374276 227400 374328 227452
rect 514024 227400 514076 227452
rect 535736 227400 535788 227452
rect 538312 227400 538364 227452
rect 556068 227400 556120 227452
rect 89628 227264 89680 227316
rect 161434 227264 161486 227316
rect 161572 227264 161624 227316
rect 176752 227264 176804 227316
rect 228732 227264 228784 227316
rect 235816 227264 235868 227316
rect 280252 227264 280304 227316
rect 306196 227264 306248 227316
rect 336924 227264 336976 227316
rect 340696 227264 340748 227316
rect 361396 227264 361448 227316
rect 382096 227264 382148 227316
rect 392952 227264 393004 227316
rect 63040 227128 63092 227180
rect 144828 227128 144880 227180
rect 150072 227128 150124 227180
rect 213368 227128 213420 227180
rect 214380 227128 214432 227180
rect 220084 227128 220136 227180
rect 220268 227128 220320 227180
rect 223580 227128 223632 227180
rect 56508 226992 56560 227044
rect 142436 226992 142488 227044
rect 143264 226992 143316 227044
rect 208124 226992 208176 227044
rect 122748 226856 122800 226908
rect 185400 226856 185452 226908
rect 185584 226856 185636 226908
rect 218428 226992 218480 227044
rect 262864 227128 262916 227180
rect 263508 227128 263560 227180
rect 277216 227128 277268 227180
rect 281356 227128 281408 227180
rect 317604 227128 317656 227180
rect 322848 227128 322900 227180
rect 349804 227128 349856 227180
rect 355876 227128 355928 227180
rect 375564 227128 375616 227180
rect 376668 227128 376720 227180
rect 389732 227128 389784 227180
rect 393136 227128 393188 227180
rect 402612 227264 402664 227316
rect 494704 227264 494756 227316
rect 402244 227128 402296 227180
rect 408408 227128 408460 227180
rect 478604 227128 478656 227180
rect 486792 227128 486844 227180
rect 489552 227128 489604 227180
rect 504180 227128 504232 227180
rect 213828 226856 213880 226908
rect 228916 226992 228968 227044
rect 271236 226992 271288 227044
rect 271788 226992 271840 227044
rect 301504 226992 301556 227044
rect 310428 226992 310480 227044
rect 338212 226992 338264 227044
rect 338672 226992 338724 227044
rect 360108 226992 360160 227044
rect 362776 226992 362828 227044
rect 379428 226992 379480 227044
rect 391848 226992 391900 227044
rect 403532 226992 403584 227044
rect 412548 226992 412600 227044
rect 419356 226992 419408 227044
rect 486976 226992 487028 227044
rect 500960 226992 501012 227044
rect 220268 226856 220320 226908
rect 267372 226856 267424 226908
rect 293776 226856 293828 226908
rect 324964 226856 325016 226908
rect 510620 227264 510672 227316
rect 524420 227264 524472 227316
rect 526260 227264 526312 227316
rect 550916 227264 550968 227316
rect 506204 227128 506256 227180
rect 525984 227128 526036 227180
rect 533344 227128 533396 227180
rect 560944 227128 560996 227180
rect 505008 226992 505060 227044
rect 523040 226992 523092 227044
rect 523684 226992 523736 227044
rect 548340 226992 548392 227044
rect 555424 226992 555476 227044
rect 633716 226992 633768 227044
rect 668584 226924 668636 226976
rect 672816 226992 672868 227044
rect 510988 226856 511040 226908
rect 676036 226788 676088 226840
rect 678244 226788 678296 226840
rect 117228 226720 117280 226772
rect 187516 226720 187568 226772
rect 190000 226720 190052 226772
rect 233884 226720 233936 226772
rect 249616 226720 249668 226772
rect 290556 226720 290608 226772
rect 243452 226652 243504 226704
rect 248696 226652 248748 226704
rect 129556 226584 129608 226636
rect 197360 226584 197412 226636
rect 203524 226584 203576 226636
rect 136548 226448 136600 226500
rect 141608 226448 141660 226500
rect 142252 226448 142304 226500
rect 202972 226448 203024 226500
rect 212172 226448 212224 226500
rect 214748 226448 214800 226500
rect 219348 226584 219400 226636
rect 220268 226584 220320 226636
rect 222936 226584 222988 226636
rect 231032 226584 231084 226636
rect 243268 226584 243320 226636
rect 264244 226516 264296 226568
rect 269304 226516 269356 226568
rect 673092 226516 673144 226568
rect 221832 226448 221884 226500
rect 228916 226448 228968 226500
rect 351092 226448 351144 226500
rect 353024 226448 353076 226500
rect 403992 226448 404044 226500
rect 412272 226448 412324 226500
rect 474740 226448 474792 226500
rect 482744 226448 482796 226500
rect 141792 226380 141844 226432
rect 142114 226380 142166 226432
rect 271144 226380 271196 226432
rect 279608 226380 279660 226432
rect 672724 226380 672776 226432
rect 350264 226312 350316 226364
rect 351736 226312 351788 226364
rect 388536 226312 388588 226364
rect 391664 226312 391716 226364
rect 407764 226312 407816 226364
rect 408684 226312 408736 226364
rect 481640 226312 481692 226364
rect 487804 226312 487856 226364
rect 122564 226244 122616 226296
rect 193956 226244 194008 226296
rect 194140 226244 194192 226296
rect 244188 226244 244240 226296
rect 286324 226244 286376 226296
rect 289912 226244 289964 226296
rect 291016 226244 291068 226296
rect 322112 226244 322164 226296
rect 458640 226244 458692 226296
rect 462964 226244 463016 226296
rect 127624 226108 127676 226160
rect 142114 226108 142166 226160
rect 142252 226108 142304 226160
rect 203708 226108 203760 226160
rect 203892 226108 203944 226160
rect 72424 225972 72476 226024
rect 147588 225972 147640 226024
rect 147772 225972 147824 226024
rect 149796 225972 149848 226024
rect 151912 225972 151964 226024
rect 214380 225972 214432 226024
rect 214748 226108 214800 226160
rect 259644 226108 259696 226160
rect 261852 226108 261904 226160
rect 300860 226108 300912 226160
rect 309048 226108 309100 226160
rect 336280 226108 336332 226160
rect 528560 226108 528612 226160
rect 543004 226108 543056 226160
rect 672604 226108 672656 226160
rect 220084 225972 220136 226024
rect 220268 225972 220320 226024
rect 266084 225972 266136 226024
rect 267004 225972 267056 226024
rect 274456 225972 274508 226024
rect 278412 225972 278464 226024
rect 313280 225972 313332 226024
rect 321376 225972 321428 226024
rect 346584 225972 346636 226024
rect 352932 225972 352984 226024
rect 371700 225972 371752 226024
rect 498108 225972 498160 226024
rect 514300 225972 514352 226024
rect 516600 225972 516652 226024
rect 538680 225972 538732 226024
rect 672494 225904 672546 225956
rect 83464 225836 83516 225888
rect 163044 225836 163096 225888
rect 193588 225836 193640 225888
rect 194140 225836 194192 225888
rect 198004 225836 198056 225888
rect 203892 225836 203944 225888
rect 204904 225836 204956 225888
rect 231492 225836 231544 225888
rect 249340 225836 249392 225888
rect 252468 225836 252520 225888
rect 293132 225836 293184 225888
rect 296444 225836 296496 225888
rect 327908 225836 327960 225888
rect 329748 225836 329800 225888
rect 353668 225836 353720 225888
rect 354588 225836 354640 225888
rect 372344 225836 372396 225888
rect 373816 225836 373868 225888
rect 377680 225836 377732 225888
rect 377864 225836 377916 225888
rect 390376 225836 390428 225888
rect 394332 225836 394384 225888
rect 403256 225836 403308 225888
rect 483756 225836 483808 225888
rect 497280 225836 497332 225888
rect 501144 225836 501196 225888
rect 519268 225836 519320 225888
rect 521752 225836 521804 225888
rect 545764 225836 545816 225888
rect 558184 225836 558236 225888
rect 571984 225836 572036 225888
rect 76564 225700 76616 225752
rect 151728 225700 151780 225752
rect 151912 225700 151964 225752
rect 154304 225700 154356 225752
rect 66168 225564 66220 225616
rect 142114 225564 142166 225616
rect 142252 225564 142304 225616
rect 184296 225700 184348 225752
rect 184480 225700 184532 225752
rect 212540 225700 212592 225752
rect 215208 225700 215260 225752
rect 154672 225564 154724 225616
rect 217140 225564 217192 225616
rect 220084 225700 220136 225752
rect 237288 225700 237340 225752
rect 240324 225700 240376 225752
rect 255044 225700 255096 225752
rect 296996 225700 297048 225752
rect 315672 225700 315724 225752
rect 344652 225700 344704 225752
rect 347044 225700 347096 225752
rect 367836 225700 367888 225752
rect 371792 225700 371844 225752
rect 382740 225700 382792 225752
rect 382924 225700 382976 225752
rect 396172 225700 396224 225752
rect 488908 225700 488960 225752
rect 503628 225700 503680 225752
rect 508872 225700 508924 225752
rect 529204 225700 529256 225752
rect 535920 225700 535972 225752
rect 563980 225700 564032 225752
rect 672380 225700 672432 225752
rect 672264 225632 672316 225684
rect 220268 225564 220320 225616
rect 222016 225564 222068 225616
rect 269948 225564 270000 225616
rect 270224 225564 270276 225616
rect 282644 225564 282696 225616
rect 284116 225564 284168 225616
rect 320180 225564 320232 225616
rect 332232 225564 332284 225616
rect 357532 225564 357584 225616
rect 372528 225564 372580 225616
rect 387432 225564 387484 225616
rect 390192 225564 390244 225616
rect 401968 225564 402020 225616
rect 410984 225564 411036 225616
rect 416136 225564 416188 225616
rect 467656 225564 467708 225616
rect 476580 225564 476632 225616
rect 477316 225564 477368 225616
rect 488816 225564 488868 225616
rect 494060 225564 494112 225616
rect 509700 225564 509752 225616
rect 510160 225564 510212 225616
rect 531044 225564 531096 225616
rect 531412 225564 531464 225616
rect 558276 225564 558328 225616
rect 110144 225428 110196 225480
rect 127624 225428 127676 225480
rect 125232 225292 125284 225344
rect 196164 225428 196216 225480
rect 196348 225428 196400 225480
rect 204904 225428 204956 225480
rect 208124 225428 208176 225480
rect 257436 225428 257488 225480
rect 463148 225360 463200 225412
rect 467288 225360 467340 225412
rect 672156 225360 672208 225412
rect 129372 225292 129424 225344
rect 199108 225292 199160 225344
rect 203708 225292 203760 225344
rect 209412 225292 209464 225344
rect 209688 225292 209740 225344
rect 214748 225292 214800 225344
rect 231492 225292 231544 225344
rect 236460 225292 236512 225344
rect 241152 225292 241204 225344
rect 286692 225292 286744 225344
rect 135168 225156 135220 225208
rect 204260 225156 204312 225208
rect 242716 225156 242768 225208
rect 285404 225156 285456 225208
rect 132408 225020 132460 225072
rect 201684 225020 201736 225072
rect 202236 225020 202288 225072
rect 254492 225020 254544 225072
rect 297272 224952 297324 225004
rect 305368 224952 305420 225004
rect 327724 224952 327776 225004
rect 332048 224952 332100 225004
rect 369124 224952 369176 225004
rect 373632 224952 373684 225004
rect 404176 224952 404228 225004
rect 410616 224952 410668 225004
rect 416504 224952 416556 225004
rect 422208 224952 422260 225004
rect 493600 224952 493652 225004
rect 494704 224952 494756 225004
rect 495164 224952 495216 225004
rect 567016 225088 567068 225140
rect 571432 225088 571484 225140
rect 563704 224952 563756 225004
rect 672034 225224 672086 225276
rect 96252 224884 96304 224936
rect 173348 224884 173400 224936
rect 174912 224884 174964 224936
rect 181352 224884 181404 224936
rect 181996 224884 182048 224936
rect 102048 224748 102100 224800
rect 178500 224748 178552 224800
rect 178776 224748 178828 224800
rect 185400 224748 185452 224800
rect 185768 224884 185820 224936
rect 195244 224884 195296 224936
rect 195428 224884 195480 224936
rect 242900 224884 242952 224936
rect 266176 224884 266228 224936
rect 460572 224884 460624 224936
rect 463148 224884 463200 224936
rect 630864 224952 630916 225004
rect 658188 224952 658240 225004
rect 568948 224884 569000 224936
rect 303436 224816 303488 224868
rect 610992 224816 611044 224868
rect 614948 224816 615000 224868
rect 204536 224748 204588 224800
rect 204720 224748 204772 224800
rect 79968 224612 80020 224664
rect 160468 224612 160520 224664
rect 162768 224612 162820 224664
rect 223856 224612 223908 224664
rect 224224 224748 224276 224800
rect 230020 224748 230072 224800
rect 232964 224748 233016 224800
rect 237748 224748 237800 224800
rect 245292 224748 245344 224800
rect 287980 224748 288032 224800
rect 311532 224748 311584 224800
rect 338856 224748 338908 224800
rect 462504 224748 462556 224800
rect 469312 224748 469364 224800
rect 506940 224748 506992 224800
rect 526720 224748 526772 224800
rect 529940 224748 529992 224800
rect 534540 224748 534592 224800
rect 224408 224612 224460 224664
rect 224592 224612 224644 224664
rect 270592 224612 270644 224664
rect 274272 224612 274324 224664
rect 312452 224612 312504 224664
rect 319812 224612 319864 224664
rect 345940 224612 345992 224664
rect 346216 224612 346268 224664
rect 366548 224680 366600 224732
rect 505192 224612 505244 224664
rect 557356 224748 557408 224800
rect 535276 224612 535328 224664
rect 562140 224748 562192 224800
rect 562324 224748 562376 224800
rect 567016 224748 567068 224800
rect 567844 224748 567896 224800
rect 610808 224748 610860 224800
rect 668492 224680 668544 224732
rect 557816 224612 557868 224664
rect 610440 224612 610492 224664
rect 610624 224612 610676 224664
rect 616052 224612 616104 224664
rect 671820 224680 671872 224732
rect 85488 224476 85540 224528
rect 165620 224476 165672 224528
rect 181352 224476 181404 224528
rect 235172 224476 235224 224528
rect 251088 224476 251140 224528
rect 294420 224476 294472 224528
rect 319996 224476 320048 224528
rect 347228 224476 347280 224528
rect 363512 224476 363564 224528
rect 368480 224476 368532 224528
rect 387708 224476 387760 224528
rect 397828 224476 397880 224528
rect 456064 224476 456116 224528
rect 459744 224476 459796 224528
rect 491300 224476 491352 224528
rect 506112 224476 506164 224528
rect 515956 224476 516008 224528
rect 530860 224476 530912 224528
rect 73712 224340 73764 224392
rect 88984 224340 89036 224392
rect 89444 224340 89496 224392
rect 167828 224340 167880 224392
rect 168288 224340 168340 224392
rect 224224 224340 224276 224392
rect 224408 224340 224460 224392
rect 232964 224340 233016 224392
rect 233148 224340 233200 224392
rect 277676 224340 277728 224392
rect 299296 224340 299348 224392
rect 331772 224340 331824 224392
rect 335176 224340 335228 224392
rect 356888 224340 356940 224392
rect 361212 224340 361264 224392
rect 377496 224340 377548 224392
rect 379244 224340 379296 224392
rect 393596 224340 393648 224392
rect 480536 224340 480588 224392
rect 492772 224340 492824 224392
rect 499212 224340 499264 224392
rect 516784 224340 516836 224392
rect 520464 224340 520516 224392
rect 544108 224476 544160 224528
rect 544292 224476 544344 224528
rect 549996 224476 550048 224528
rect 550364 224476 550416 224528
rect 551192 224476 551244 224528
rect 557172 224476 557224 224528
rect 426440 224272 426492 224324
rect 426992 224272 427044 224324
rect 68928 224068 68980 224120
rect 151636 224204 151688 224256
rect 151774 224204 151826 224256
rect 155316 224204 155368 224256
rect 165528 224204 165580 224256
rect 227444 224204 227496 224256
rect 231676 224204 231728 224256
rect 278964 224204 279016 224256
rect 290832 224204 290884 224256
rect 323676 224204 323728 224256
rect 323952 224204 324004 224256
rect 334992 224204 335044 224256
rect 339408 224204 339460 224256
rect 88984 224068 89036 224120
rect 142114 224068 142166 224120
rect 142252 224068 142304 224120
rect 194600 224068 194652 224120
rect 195244 224068 195296 224120
rect 204720 224068 204772 224120
rect 204904 224068 204956 224120
rect 250628 224068 250680 224120
rect 275100 224068 275152 224120
rect 311164 224068 311216 224120
rect 358084 224204 358136 224256
rect 362960 224204 363012 224256
rect 366732 224204 366784 224256
rect 381636 224204 381688 224256
rect 394516 224204 394568 224256
rect 404544 224204 404596 224256
rect 405556 224204 405608 224256
rect 414204 224204 414256 224256
rect 427912 224204 427964 224256
rect 428740 224204 428792 224256
rect 470232 224204 470284 224256
rect 480444 224204 480496 224256
rect 486608 224204 486660 224256
rect 500408 224204 500460 224256
rect 504364 224204 504416 224256
rect 523500 224204 523552 224256
rect 525616 224204 525668 224256
rect 550640 224340 550692 224392
rect 550824 224340 550876 224392
rect 625252 224476 625304 224528
rect 667756 224408 667808 224460
rect 557816 224340 557868 224392
rect 625436 224340 625488 224392
rect 532700 224204 532752 224256
rect 619640 224204 619692 224256
rect 651288 224204 651340 224256
rect 658188 224204 658240 224256
rect 362316 224068 362368 224120
rect 377404 224068 377456 224120
rect 385868 224068 385920 224120
rect 519084 224068 519136 224120
rect 530676 224068 530728 224120
rect 530860 224068 530912 224120
rect 534356 224068 534408 224120
rect 534540 224068 534592 224120
rect 543740 224068 543792 224120
rect 667020 224068 667072 224120
rect 543924 224000 543976 224052
rect 545028 224000 545080 224052
rect 623780 224000 623832 224052
rect 671482 224068 671534 224120
rect 106004 223932 106056 223984
rect 181076 223932 181128 223984
rect 201224 223932 201276 223984
rect 255780 223932 255832 223984
rect 286692 223932 286744 223984
rect 319536 223932 319588 223984
rect 667756 223932 667808 223984
rect 279424 223864 279476 223916
rect 284760 223864 284812 223916
rect 509700 223864 509752 223916
rect 510160 223864 510212 223916
rect 610624 223864 610676 223916
rect 610808 223864 610860 223916
rect 622676 223864 622728 223916
rect 108672 223796 108724 223848
rect 183836 223796 183888 223848
rect 184848 223796 184900 223848
rect 112812 223660 112864 223712
rect 185952 223660 186004 223712
rect 186964 223796 187016 223848
rect 217784 223796 217836 223848
rect 228732 223796 228784 223848
rect 274916 223796 274968 223848
rect 524420 223728 524472 223780
rect 525064 223728 525116 223780
rect 532700 223728 532752 223780
rect 195428 223660 195480 223712
rect 195888 223660 195940 223712
rect 204904 223660 204956 223712
rect 238024 223660 238076 223712
rect 266728 223660 266780 223712
rect 319628 223660 319680 223712
rect 319996 223660 320048 223712
rect 530676 223592 530728 223644
rect 535000 223728 535052 223780
rect 621572 223728 621624 223780
rect 534356 223592 534408 223644
rect 538312 223592 538364 223644
rect 539968 223592 540020 223644
rect 567844 223592 567896 223644
rect 568304 223592 568356 223644
rect 628748 223592 628800 223644
rect 670424 223592 670476 223644
rect 78588 223524 78640 223576
rect 154028 223524 154080 223576
rect 154212 223524 154264 223576
rect 161940 223524 161992 223576
rect 162124 223524 162176 223576
rect 186596 223524 186648 223576
rect 187332 223524 187384 223576
rect 242256 223524 242308 223576
rect 250904 223524 250956 223576
rect 291200 223524 291252 223576
rect 297916 223524 297968 223576
rect 303252 223524 303304 223576
rect 307668 223524 307720 223576
rect 335636 223524 335688 223576
rect 406752 223524 406804 223576
rect 414848 223524 414900 223576
rect 454868 223524 454920 223576
rect 460480 223524 460532 223576
rect 473452 223524 473504 223576
rect 475568 223524 475620 223576
rect 75828 223388 75880 223440
rect 154948 223388 155000 223440
rect 155500 223388 155552 223440
rect 159180 223388 159232 223440
rect 159364 223388 159416 223440
rect 181812 223388 181864 223440
rect 184020 223388 184072 223440
rect 239680 223388 239732 223440
rect 244096 223388 244148 223440
rect 286048 223388 286100 223440
rect 304724 223388 304776 223440
rect 308128 223388 308180 223440
rect 312912 223388 312964 223440
rect 342076 223456 342128 223508
rect 666652 223456 666704 223508
rect 342812 223388 342864 223440
rect 347872 223388 347924 223440
rect 517520 223388 517572 223440
rect 531504 223388 531556 223440
rect 534724 223388 534776 223440
rect 547420 223388 547472 223440
rect 561956 223388 562008 223440
rect 568764 223388 568816 223440
rect 336004 223320 336056 223372
rect 342260 223320 342312 223372
rect 66904 223252 66956 223304
rect 146668 223252 146720 223304
rect 147312 223252 147364 223304
rect 176660 223252 176712 223304
rect 188896 223252 188948 223304
rect 245108 223252 245160 223304
rect 246856 223252 246908 223304
rect 288624 223252 288676 223304
rect 289728 223252 289780 223304
rect 297732 223252 297784 223304
rect 299112 223252 299164 223304
rect 328552 223252 328604 223304
rect 347228 223252 347280 223304
rect 357900 223252 357952 223304
rect 483112 223252 483164 223304
rect 496084 223252 496136 223304
rect 503352 223252 503404 223304
rect 69572 223116 69624 223168
rect 149520 223116 149572 223168
rect 71412 222980 71464 223032
rect 152096 223116 152148 223168
rect 154396 223116 154448 223168
rect 216220 223116 216272 223168
rect 241336 223116 241388 223168
rect 283472 223116 283524 223168
rect 288256 223116 288308 223168
rect 321100 223116 321152 223168
rect 344652 223116 344704 223168
rect 364616 223116 364668 223168
rect 365536 223116 365588 223168
rect 379612 223116 379664 223168
rect 380072 223116 380124 223168
rect 386512 223116 386564 223168
rect 488632 223116 488684 223168
rect 503168 223116 503220 223168
rect 508228 223116 508280 223168
rect 514668 223252 514720 223304
rect 536288 223252 536340 223304
rect 554044 223252 554096 223304
rect 562508 223252 562560 223304
rect 566832 223252 566884 223304
rect 568304 223252 568356 223304
rect 586980 223252 587032 223304
rect 593972 223252 594024 223304
rect 153660 222980 153712 223032
rect 155500 222980 155552 223032
rect 155684 222980 155736 223032
rect 219532 222980 219584 223032
rect 230204 222980 230256 223032
rect 275468 222980 275520 223032
rect 278596 222980 278648 223032
rect 315028 222980 315080 223032
rect 316684 222980 316736 223032
rect 327264 222980 327316 223032
rect 328092 222980 328144 223032
rect 351460 222980 351512 223032
rect 353944 222980 353996 223032
rect 365904 222980 365956 223032
rect 366916 222980 366968 223032
rect 383844 222980 383896 223032
rect 384212 222980 384264 223032
rect 393964 222980 394016 223032
rect 493048 222980 493100 223032
rect 508504 222980 508556 223032
rect 521752 223116 521804 223168
rect 532056 223116 532108 223168
rect 559012 223116 559064 223168
rect 559840 223116 559892 223168
rect 567660 223116 567712 223168
rect 527824 222980 527876 223032
rect 529480 222980 529532 223032
rect 555700 222980 555752 223032
rect 559380 222980 559432 223032
rect 568304 222980 568356 223032
rect 587164 222980 587216 223032
rect 620652 223116 620704 223168
rect 667020 223116 667072 223168
rect 617340 222980 617392 223032
rect 625620 222980 625672 223032
rect 62764 222844 62816 222896
rect 141976 222844 142028 222896
rect 142160 222844 142212 222896
rect 144000 222844 144052 222896
rect 146024 222844 146076 222896
rect 211988 222844 212040 222896
rect 215944 222844 215996 222896
rect 233332 222844 233384 222896
rect 234528 222844 234580 222896
rect 281540 222844 281592 222896
rect 282460 222844 282512 222896
rect 316316 222844 316368 222896
rect 324136 222844 324188 222896
rect 348516 222844 348568 222896
rect 349068 222844 349120 222896
rect 367192 222844 367244 222896
rect 368388 222844 368440 222896
rect 382372 222844 382424 222896
rect 383476 222844 383528 222896
rect 394884 222844 394936 222896
rect 395804 222844 395856 222896
rect 406476 222844 406528 222896
rect 420828 222844 420880 222896
rect 425152 222844 425204 222896
rect 459928 222844 459980 222896
rect 467104 222844 467156 222896
rect 467472 222844 467524 222896
rect 473728 222844 473780 222896
rect 479892 222844 479944 222896
rect 491944 222844 491996 222896
rect 500776 222844 500828 222896
rect 517520 222844 517572 222896
rect 519820 222844 519872 222896
rect 542360 222844 542412 222896
rect 543832 222844 543884 222896
rect 552480 222844 552532 222896
rect 562324 222844 562376 222896
rect 562508 222844 562560 222896
rect 632704 222844 632756 222896
rect 81348 222708 81400 222760
rect 153660 222708 153712 222760
rect 154028 222708 154080 222760
rect 156972 222708 157024 222760
rect 166264 222708 166316 222760
rect 192024 222708 192076 222760
rect 194508 222708 194560 222760
rect 247408 222708 247460 222760
rect 264796 222708 264848 222760
rect 304356 222708 304408 222760
rect 482744 222708 482796 222760
rect 586980 222708 587032 222760
rect 587164 222708 587216 222760
rect 99288 222572 99340 222624
rect 175740 222572 175792 222624
rect 197176 222572 197228 222624
rect 249984 222572 250036 222624
rect 557540 222572 557592 222624
rect 559840 222572 559892 222624
rect 562324 222572 562376 222624
rect 617340 222572 617392 222624
rect 620468 222708 620520 222760
rect 627092 222708 627144 222760
rect 629852 222572 629904 222624
rect 175924 222504 175976 222556
rect 87972 222436 88024 222488
rect 164976 222436 165028 222488
rect 207480 222436 207532 222488
rect 207664 222436 207716 222488
rect 258356 222436 258408 222488
rect 489920 222436 489972 222488
rect 491116 222436 491168 222488
rect 172152 222368 172204 222420
rect 85304 222300 85356 222352
rect 154212 222300 154264 222352
rect 199752 222300 199804 222352
rect 211804 222300 211856 222352
rect 228088 222300 228140 222352
rect 287888 222300 287940 222352
rect 295064 222300 295116 222352
rect 484492 222300 484544 222352
rect 504364 222436 504416 222488
rect 523684 222436 523736 222488
rect 529848 222436 529900 222488
rect 619916 222436 619968 222488
rect 118424 222164 118476 222216
rect 141976 222164 142028 222216
rect 142160 222164 142212 222216
rect 191012 222164 191064 222216
rect 568304 222300 568356 222352
rect 568764 222300 568816 222352
rect 627920 222300 627972 222352
rect 504364 222164 504416 222216
rect 523684 222164 523736 222216
rect 559380 222164 559432 222216
rect 567660 222164 567712 222216
rect 620468 222164 620520 222216
rect 620652 222164 620704 222216
rect 631508 222164 631560 222216
rect 160836 222096 160888 222148
rect 166080 222096 166132 222148
rect 97908 221960 97960 222012
rect 172704 222096 172756 222148
rect 174084 222096 174136 222148
rect 191472 222096 191524 222148
rect 247592 222096 247644 222148
rect 258080 222096 258132 222148
rect 263692 222096 263744 222148
rect 270040 222096 270092 222148
rect 306380 222096 306432 222148
rect 310704 222096 310756 222148
rect 312636 222096 312688 222148
rect 331404 222096 331456 222148
rect 353760 222096 353812 222148
rect 424968 222096 425020 222148
rect 429292 222096 429344 222148
rect 452568 222096 452620 222148
rect 455604 222096 455656 222148
rect 462136 222096 462188 222148
rect 468760 222096 468812 222148
rect 471888 222096 471940 222148
rect 477868 222096 477920 222148
rect 559564 222096 559616 222148
rect 564808 222096 564860 222148
rect 167000 221960 167052 222012
rect 169760 221960 169812 222012
rect 171784 221960 171836 222012
rect 178960 221960 179012 222012
rect 495164 222028 495216 222080
rect 497740 222028 497792 222080
rect 515496 222028 515548 222080
rect 529848 222028 529900 222080
rect 533988 222028 534040 222080
rect 559380 222028 559432 222080
rect 592040 222028 592092 222080
rect 596640 222028 596692 222080
rect 596824 222028 596876 222080
rect 605012 222028 605064 222080
rect 231860 221960 231912 222012
rect 233700 221960 233752 222012
rect 277952 221960 278004 222012
rect 280068 221960 280120 222012
rect 314016 221960 314068 222012
rect 318248 221960 318300 222012
rect 343824 221960 343876 222012
rect 367652 221960 367704 222012
rect 380256 221960 380308 222012
rect 536104 221892 536156 221944
rect 543694 221892 543746 221944
rect 557172 221892 557224 221944
rect 608600 221892 608652 221944
rect 104532 221824 104584 221876
rect 176292 221824 176344 221876
rect 80520 221688 80572 221740
rect 86224 221688 86276 221740
rect 94688 221688 94740 221740
rect 161434 221688 161486 221740
rect 161572 221688 161624 221740
rect 167184 221688 167236 221740
rect 167460 221688 167512 221740
rect 171416 221688 171468 221740
rect 171600 221688 171652 221740
rect 182640 221824 182692 221876
rect 182824 221824 182876 221876
rect 240140 221824 240192 221876
rect 263324 221824 263376 221876
rect 301228 221824 301280 221876
rect 301412 221824 301464 221876
rect 310888 221824 310940 221876
rect 313188 221824 313240 221876
rect 340420 221824 340472 221876
rect 351276 221824 351328 221876
rect 369308 221824 369360 221876
rect 509884 221824 509936 221876
rect 522672 221824 522724 221876
rect 546592 221824 546644 221876
rect 547144 221824 547196 221876
rect 556804 221824 556856 221876
rect 178960 221688 179012 221740
rect 232228 221688 232280 221740
rect 239220 221688 239272 221740
rect 283656 221688 283708 221740
rect 303252 221688 303304 221740
rect 332784 221688 332836 221740
rect 357164 221688 357216 221740
rect 374644 221688 374696 221740
rect 391020 221688 391072 221740
rect 400312 221688 400364 221740
rect 475844 221688 475896 221740
rect 486148 221688 486200 221740
rect 496268 221688 496320 221740
rect 513564 221688 513616 221740
rect 522856 221688 522908 221740
rect 549260 221688 549312 221740
rect 606668 221688 606720 221740
rect 59360 221552 59412 221604
rect 138296 221552 138348 221604
rect 138480 221552 138532 221604
rect 140780 221552 140832 221604
rect 140964 221552 141016 221604
rect 205916 221552 205968 221604
rect 208400 221552 208452 221604
rect 260840 221552 260892 221604
rect 261024 221552 261076 221604
rect 301780 221552 301832 221604
rect 308864 221552 308916 221604
rect 339684 221552 339736 221604
rect 341340 221552 341392 221604
rect 361764 221552 361816 221604
rect 369492 221552 369544 221604
rect 384028 221552 384080 221604
rect 384396 221552 384448 221604
rect 395160 221552 395212 221604
rect 400772 221552 400824 221604
rect 405740 221552 405792 221604
rect 480812 221552 480864 221604
rect 492956 221552 493008 221604
rect 497464 221552 497516 221604
rect 515128 221552 515180 221604
rect 524236 221552 524288 221604
rect 73896 221416 73948 221468
rect 82084 221416 82136 221468
rect 86316 221416 86368 221468
rect 91284 221280 91336 221332
rect 118148 221280 118200 221332
rect 127440 221280 127492 221332
rect 161434 221280 161486 221332
rect 161756 221416 161808 221468
rect 164424 221280 164476 221332
rect 171600 221280 171652 221332
rect 171968 221416 172020 221468
rect 226524 221416 226576 221468
rect 227904 221416 227956 221468
rect 276112 221416 276164 221468
rect 292488 221416 292540 221468
rect 326252 221416 326304 221468
rect 342168 221416 342220 221468
rect 364800 221416 364852 221468
rect 375288 221416 375340 221468
rect 390744 221416 390796 221468
rect 396816 221416 396868 221468
rect 407304 221416 407356 221468
rect 408408 221416 408460 221468
rect 416872 221416 416924 221468
rect 468944 221416 468996 221468
rect 476212 221416 476264 221468
rect 483756 221416 483808 221468
rect 533252 221416 533304 221468
rect 533620 221552 533672 221604
rect 601976 221552 602028 221604
rect 193312 221280 193364 221332
rect 204168 221280 204220 221332
rect 252744 221280 252796 221332
rect 266820 221280 266872 221332
rect 303804 221280 303856 221332
rect 523500 221280 523552 221332
rect 533160 221280 533212 221332
rect 538680 221348 538732 221400
rect 543648 221212 543700 221264
rect 543832 221212 543884 221264
rect 548524 221212 548576 221264
rect 597008 221416 597060 221468
rect 633440 221416 633492 221468
rect 548892 221348 548944 221400
rect 596824 221348 596876 221400
rect 669780 221348 669832 221400
rect 604644 221212 604696 221264
rect 111156 221008 111208 221060
rect 118148 221008 118200 221060
rect 124404 221008 124456 221060
rect 127256 221008 127308 221060
rect 127440 221008 127492 221060
rect 166080 221144 166132 221196
rect 221280 221144 221332 221196
rect 222752 221144 222804 221196
rect 268292 221144 268344 221196
rect 521108 221076 521160 221128
rect 591948 221076 592000 221128
rect 592132 221076 592184 221128
rect 600412 221076 600464 221128
rect 669780 221076 669832 221128
rect 127900 221008 127952 221060
rect 146392 221008 146444 221060
rect 206468 221008 206520 221060
rect 219808 221008 219860 221060
rect 263048 221008 263100 221060
rect 83004 220872 83056 220924
rect 142114 220872 142166 220924
rect 142252 220872 142304 220924
rect 145564 220872 145616 220924
rect 525984 220940 526036 220992
rect 601792 220940 601844 220992
rect 161434 220872 161486 220924
rect 161572 220872 161624 220924
rect 222292 220872 222344 220924
rect 282644 220872 282696 220924
rect 287704 220872 287756 220924
rect 456708 220872 456760 220924
rect 253848 220804 253900 220856
rect 258632 220804 258684 220856
rect 418344 220804 418396 220856
rect 424048 220804 424100 220856
rect 466092 220872 466144 220924
rect 471428 220872 471480 220924
rect 669412 220872 669464 220924
rect 462136 220804 462188 220856
rect 517520 220804 517572 220856
rect 518532 220804 518584 220856
rect 592040 220804 592092 220856
rect 596916 220804 596968 220856
rect 600688 220804 600740 220856
rect 114284 220736 114336 220788
rect 145840 220736 145892 220788
rect 146944 220736 146996 220788
rect 177212 220736 177264 220788
rect 177396 220736 177448 220788
rect 181260 220736 181312 220788
rect 181444 220736 181496 220788
rect 190368 220736 190420 220788
rect 190552 220736 190604 220788
rect 236644 220736 236696 220788
rect 242624 220736 242676 220788
rect 246488 220736 246540 220788
rect 260196 220736 260248 220788
rect 298560 220736 298612 220788
rect 302424 220736 302476 220788
rect 334072 220736 334124 220788
rect 385224 220736 385276 220788
rect 388720 220736 388772 220788
rect 414204 220736 414256 220788
rect 418160 220736 418212 220788
rect 455328 220736 455380 220788
rect 458824 220736 458876 220788
rect 465724 220736 465776 220788
rect 469588 220736 469640 220788
rect 474004 220736 474056 220788
rect 475384 220736 475436 220788
rect 476764 220736 476816 220788
rect 478696 220736 478748 220788
rect 511816 220736 511868 220788
rect 101220 220600 101272 220652
rect 175096 220600 175148 220652
rect 175280 220600 175332 220652
rect 224224 220600 224276 220652
rect 253572 220600 253624 220652
rect 293316 220600 293368 220652
rect 294972 220600 295024 220652
rect 325884 220600 325936 220652
rect 357900 220600 357952 220652
rect 374460 220600 374512 220652
rect 500224 220600 500276 220652
rect 511816 220600 511868 220652
rect 332692 220532 332744 220584
rect 337200 220532 337252 220584
rect 69756 220464 69808 220516
rect 136916 220464 136968 220516
rect 137100 220464 137152 220516
rect 146944 220464 146996 220516
rect 147128 220464 147180 220516
rect 208584 220464 208636 220516
rect 210516 220464 210568 220516
rect 259920 220464 259972 220516
rect 267648 220464 267700 220516
rect 306840 220464 306892 220516
rect 338028 220464 338080 220516
rect 359004 220464 359056 220516
rect 469128 220464 469180 220516
rect 474556 220464 474608 220516
rect 488448 220464 488500 220516
rect 501880 220464 501932 220516
rect 543648 220668 543700 220720
rect 549076 220668 549128 220720
rect 520924 220600 520976 220652
rect 537484 220600 537536 220652
rect 551008 220600 551060 220652
rect 554228 220600 554280 220652
rect 555700 220600 555752 220652
rect 562876 220600 562928 220652
rect 563060 220600 563112 220652
rect 587348 220600 587400 220652
rect 587532 220600 587584 220652
rect 596732 220736 596784 220788
rect 669412 220736 669464 220788
rect 669872 220736 669924 220788
rect 670240 220736 670292 220788
rect 538312 220532 538364 220584
rect 543832 220532 543884 220584
rect 531688 220464 531740 220516
rect 73068 220328 73120 220380
rect 145656 220328 145708 220380
rect 145840 220328 145892 220380
rect 153476 220328 153528 220380
rect 154396 220328 154448 220380
rect 214104 220328 214156 220380
rect 214288 220328 214340 220380
rect 79692 220192 79744 220244
rect 158904 220192 158956 220244
rect 164148 220192 164200 220244
rect 223672 220192 223724 220244
rect 224408 220328 224460 220380
rect 267924 220328 267976 220380
rect 273444 220328 273496 220380
rect 309232 220328 309284 220380
rect 314844 220328 314896 220380
rect 341064 220328 341116 220380
rect 342996 220328 343048 220380
rect 363328 220328 363380 220380
rect 472992 220328 473044 220380
rect 481180 220328 481232 220380
rect 496452 220328 496504 220380
rect 509332 220328 509384 220380
rect 516968 220328 517020 220380
rect 527548 220328 527600 220380
rect 531228 220328 531280 220380
rect 556528 220464 556580 220516
rect 234160 220192 234212 220244
rect 237012 220192 237064 220244
rect 280436 220192 280488 220244
rect 283380 220192 283432 220244
rect 316500 220192 316552 220244
rect 321652 220192 321704 220244
rect 324504 220192 324556 220244
rect 76380 220056 76432 220108
rect 156144 220056 156196 220108
rect 157524 220056 157576 220108
rect 214104 220056 214156 220108
rect 107844 219920 107896 219972
rect 114284 219920 114336 219972
rect 114468 219920 114520 219972
rect 121092 219784 121144 219836
rect 127624 219920 127676 219972
rect 181444 219920 181496 219972
rect 181628 219920 181680 219972
rect 214288 219920 214340 219972
rect 137100 219784 137152 219836
rect 127624 219648 127676 219700
rect 131028 219648 131080 219700
rect 197636 219784 197688 219836
rect 197820 219784 197872 219836
rect 244280 220056 244332 220108
rect 244464 220056 244516 220108
rect 288532 220056 288584 220108
rect 288716 220056 288768 220108
rect 136916 219512 136968 219564
rect 144644 219648 144696 219700
rect 144828 219648 144880 219700
rect 146760 219648 146812 219700
rect 137652 219512 137704 219564
rect 203156 219648 203208 219700
rect 203892 219648 203944 219700
rect 254768 219920 254820 219972
rect 316500 220056 316552 220108
rect 342628 220192 342680 220244
rect 348792 220192 348844 220244
rect 369952 220192 370004 220244
rect 370504 220192 370556 220244
rect 381084 220192 381136 220244
rect 388720 220192 388772 220244
rect 400956 220192 401008 220244
rect 432236 220192 432288 220244
rect 434812 220192 434864 220244
rect 459468 220192 459520 220244
rect 465448 220192 465500 220244
rect 473176 220192 473228 220244
rect 482008 220192 482060 220244
rect 482928 220192 482980 220244
rect 495256 220192 495308 220244
rect 501328 220192 501380 220244
rect 520188 220192 520240 220244
rect 528376 220192 528428 220244
rect 554044 220328 554096 220380
rect 554228 220328 554280 220380
rect 562140 220464 562192 220516
rect 558276 220328 558328 220380
rect 561772 220328 561824 220380
rect 566832 220328 566884 220380
rect 567292 220328 567344 220380
rect 568580 220464 568632 220516
rect 569776 220464 569828 220516
rect 572674 220464 572726 220516
rect 610532 220464 610584 220516
rect 572352 220328 572404 220380
rect 574744 220328 574796 220380
rect 611452 220328 611504 220380
rect 548708 220192 548760 220244
rect 562876 220192 562928 220244
rect 608968 220192 609020 220244
rect 325608 220056 325660 220108
rect 352104 220056 352156 220108
rect 358820 220056 358872 220108
rect 378324 220056 378376 220108
rect 379428 220056 379480 220108
rect 392124 220056 392176 220108
rect 395988 220056 396040 220108
rect 404728 220056 404780 220108
rect 421656 220056 421708 220108
rect 426808 220056 426860 220108
rect 478328 220056 478380 220108
rect 489460 220056 489512 220108
rect 492496 220056 492548 220108
rect 506848 220056 506900 220108
rect 513104 220056 513156 220108
rect 534172 220056 534224 220108
rect 538128 220056 538180 220108
rect 561772 220056 561824 220108
rect 587348 220056 587400 220108
rect 608784 220056 608836 220108
rect 562140 219988 562192 220040
rect 322388 219920 322440 219972
rect 503628 219852 503680 219904
rect 586980 219852 587032 219904
rect 607312 219852 607364 219904
rect 217140 219784 217192 219836
rect 265164 219784 265216 219836
rect 220452 219648 220504 219700
rect 224408 219648 224460 219700
rect 227076 219648 227128 219700
rect 272708 219648 272760 219700
rect 464988 219580 465040 219632
rect 472072 219580 472124 219632
rect 527548 219580 527600 219632
rect 548708 219716 548760 219768
rect 548892 219716 548944 219768
rect 595628 219716 595680 219768
rect 540796 219580 540848 219632
rect 606024 219716 606076 219768
rect 147588 219512 147640 219564
rect 211344 219512 211396 219564
rect 214104 219512 214156 219564
rect 218704 219512 218756 219564
rect 224224 219512 224276 219564
rect 229284 219512 229336 219564
rect 405924 219444 405976 219496
rect 412732 219444 412784 219496
rect 70584 219376 70636 219428
rect 117596 219376 117648 219428
rect 117780 219376 117832 219428
rect 118700 219376 118752 219428
rect 131856 219376 131908 219428
rect 132408 219376 132460 219428
rect 132592 219376 132644 219428
rect 168932 219376 168984 219428
rect 169116 219376 169168 219428
rect 169576 219376 169628 219428
rect 169760 219376 169812 219428
rect 172152 219376 172204 219428
rect 172428 219376 172480 219428
rect 173164 219376 173216 219428
rect 178224 219376 178276 219428
rect 178776 219376 178828 219428
rect 181628 219376 181680 219428
rect 182088 219376 182140 219428
rect 182272 219376 182324 219428
rect 184480 219376 184532 219428
rect 185676 219376 185728 219428
rect 186136 219376 186188 219428
rect 186274 219376 186326 219428
rect 215944 219376 215996 219428
rect 219624 219376 219676 219428
rect 261208 219376 261260 219428
rect 262680 219376 262732 219428
rect 263600 219376 263652 219428
rect 272340 219376 272392 219428
rect 301412 219376 301464 219428
rect 308220 219376 308272 219428
rect 309140 219376 309192 219428
rect 314016 219376 314068 219428
rect 330300 219376 330352 219428
rect 333704 219376 333756 219428
rect 347228 219376 347280 219428
rect 349620 219376 349672 219428
rect 350540 219376 350592 219428
rect 352104 219376 352156 219428
rect 355324 219376 355376 219428
rect 362040 219376 362092 219428
rect 367652 219376 367704 219428
rect 380256 219376 380308 219428
rect 384212 219376 384264 219428
rect 399300 219376 399352 219428
rect 400220 219376 400272 219428
rect 415860 219376 415912 219428
rect 416780 219376 416832 219428
rect 417516 219376 417568 219428
rect 421012 219444 421064 219496
rect 432052 219512 432104 219564
rect 501144 219512 501196 219564
rect 428280 219376 428332 219428
rect 582380 219444 582432 219496
rect 620100 219580 620152 219632
rect 93768 219240 93820 219292
rect 94412 219240 94464 219292
rect 117964 219240 118016 219292
rect 159364 219240 159416 219292
rect 162492 219240 162544 219292
rect 171600 219240 171652 219292
rect 64604 219104 64656 219156
rect 66904 219104 66956 219156
rect 83832 219104 83884 219156
rect 157984 219104 158036 219156
rect 165804 219104 165856 219156
rect 180064 219240 180116 219292
rect 181444 219240 181496 219292
rect 190000 219240 190052 219292
rect 190644 219240 190696 219292
rect 194876 219240 194928 219292
rect 195060 219240 195112 219292
rect 224040 219240 224092 219292
rect 237840 219240 237892 219292
rect 239220 219240 239272 219292
rect 239496 219240 239548 219292
rect 272892 219240 272944 219292
rect 285864 219240 285916 219292
rect 313832 219240 313884 219292
rect 419172 219240 419224 219292
rect 422668 219240 422720 219292
rect 536196 219240 536248 219292
rect 536656 219240 536708 219292
rect 171968 219104 172020 219156
rect 175924 219104 175976 219156
rect 62304 218968 62356 219020
rect 72424 218968 72476 219020
rect 77208 218968 77260 219020
rect 150624 218968 150676 219020
rect 152372 218968 152424 219020
rect 153844 218968 153896 219020
rect 154028 218968 154080 219020
rect 160192 218968 160244 219020
rect 161480 218968 161532 219020
rect 166264 218968 166316 219020
rect 169760 218968 169812 219020
rect 207848 219104 207900 219156
rect 208860 219104 208912 219156
rect 209688 219104 209740 219156
rect 211344 219104 211396 219156
rect 217324 219104 217376 219156
rect 218796 219104 218848 219156
rect 219348 219104 219400 219156
rect 224224 219104 224276 219156
rect 253388 219104 253440 219156
rect 261208 219104 261260 219156
rect 264244 219104 264296 219156
rect 264428 219104 264480 219156
rect 267004 219104 267056 219156
rect 272708 219104 272760 219156
rect 179052 218968 179104 219020
rect 196256 218968 196308 219020
rect 200212 218968 200264 219020
rect 204168 218968 204220 219020
rect 204720 218968 204772 219020
rect 246304 218968 246356 219020
rect 252744 218968 252796 219020
rect 282184 218968 282236 219020
rect 295800 219104 295852 219156
rect 296720 219104 296772 219156
rect 320640 219104 320692 219156
rect 342812 219104 342864 219156
rect 343824 219104 343876 219156
rect 353944 219104 353996 219156
rect 363696 219104 363748 219156
rect 370504 219104 370556 219156
rect 542544 219104 542596 219156
rect 543004 219104 543056 219156
rect 548892 219240 548944 219292
rect 557356 219240 557408 219292
rect 562048 219308 562100 219360
rect 297272 218968 297324 219020
rect 307392 218968 307444 219020
rect 59820 218832 59872 218884
rect 139952 218832 140004 218884
rect 142252 218832 142304 218884
rect 146944 218832 146996 218884
rect 150900 218832 150952 218884
rect 154396 218832 154448 218884
rect 159824 218832 159876 218884
rect 203524 218832 203576 218884
rect 206468 218832 206520 218884
rect 253848 218832 253900 218884
rect 259092 218832 259144 218884
rect 58992 218696 59044 218748
rect 145104 218696 145156 218748
rect 146760 218696 146812 218748
rect 180524 218696 180576 218748
rect 180708 218696 180760 218748
rect 185952 218696 186004 218748
rect 186504 218696 186556 218748
rect 195060 218696 195112 218748
rect 195612 218696 195664 218748
rect 198004 218696 198056 218748
rect 198280 218696 198332 218748
rect 243452 218696 243504 218748
rect 253204 218696 253256 218748
rect 286324 218696 286376 218748
rect 291660 218832 291712 218884
rect 291844 218696 291896 218748
rect 300492 218832 300544 218884
rect 327724 218832 327776 218884
rect 330300 218968 330352 219020
rect 336004 218968 336056 219020
rect 337200 218968 337252 219020
rect 345664 218968 345716 219020
rect 347228 218968 347280 219020
rect 363512 218968 363564 219020
rect 368664 218968 368716 219020
rect 377404 218968 377456 219020
rect 332692 218832 332744 218884
rect 340512 218832 340564 218884
rect 358084 218832 358136 218884
rect 376944 218832 376996 218884
rect 382740 218832 382792 218884
rect 383476 218832 383528 218884
rect 386880 218968 386932 219020
rect 398104 218968 398156 219020
rect 388536 218832 388588 218884
rect 402612 218832 402664 218884
rect 409052 218832 409104 218884
rect 411720 218832 411772 218884
rect 412548 218832 412600 218884
rect 512736 218832 512788 218884
rect 561312 219104 561364 219156
rect 572536 219308 572588 219360
rect 572674 219240 572726 219292
rect 595628 219308 595680 219360
rect 607496 219444 607548 219496
rect 586980 219172 587032 219224
rect 597560 219172 597612 219224
rect 548708 218968 548760 219020
rect 574560 219104 574612 219156
rect 321652 218696 321704 218748
rect 327264 218696 327316 218748
rect 351092 218696 351144 218748
rect 353760 218696 353812 218748
rect 369124 218696 369176 218748
rect 370320 218696 370372 218748
rect 380072 218696 380124 218748
rect 383568 218696 383620 218748
rect 396264 218696 396316 218748
rect 412548 218696 412600 218748
rect 417148 218696 417200 218748
rect 482744 218696 482796 218748
rect 485320 218696 485372 218748
rect 500408 218696 500460 218748
rect 508044 218696 508096 218748
rect 517704 218696 517756 218748
rect 518164 218696 518216 218748
rect 520004 218696 520056 218748
rect 547420 218832 547472 218884
rect 563152 218968 563204 219020
rect 563336 218968 563388 219020
rect 563520 218968 563572 219020
rect 572352 218968 572404 219020
rect 572674 218968 572726 219020
rect 603080 218968 603132 219020
rect 562600 218832 562652 218884
rect 562968 218832 563020 218884
rect 563336 218832 563388 218884
rect 614120 218832 614172 218884
rect 537484 218696 537536 218748
rect 107016 218560 107068 218612
rect 117964 218560 118016 218612
rect 118148 218560 118200 218612
rect 162124 218560 162176 218612
rect 166632 218560 166684 218612
rect 169760 218560 169812 218612
rect 169944 218560 169996 218612
rect 170956 218560 171008 218612
rect 171600 218560 171652 218612
rect 181076 218560 181128 218612
rect 182364 218560 182416 218612
rect 189724 218560 189776 218612
rect 192852 218560 192904 218612
rect 100392 218288 100444 218340
rect 142252 218424 142304 218476
rect 142436 218424 142488 218476
rect 150440 218424 150492 218476
rect 150624 218424 150676 218476
rect 152372 218424 152424 218476
rect 152556 218424 152608 218476
rect 153108 218424 153160 218476
rect 153384 218424 153436 218476
rect 154028 218424 154080 218476
rect 155040 218424 155092 218476
rect 155684 218424 155736 218476
rect 156696 218424 156748 218476
rect 157248 218424 157300 218476
rect 159180 218424 159232 218476
rect 160008 218424 160060 218476
rect 160192 218424 160244 218476
rect 186964 218424 187016 218476
rect 189816 218424 189868 218476
rect 195244 218424 195296 218476
rect 198096 218560 198148 218612
rect 200212 218560 200264 218612
rect 200396 218560 200448 218612
rect 210332 218560 210384 218612
rect 213000 218560 213052 218612
rect 224224 218560 224276 218612
rect 225972 218560 226024 218612
rect 264428 218560 264480 218612
rect 265992 218560 266044 218612
rect 272708 218560 272760 218612
rect 272892 218560 272944 218612
rect 279424 218560 279476 218612
rect 198280 218424 198332 218476
rect 199752 218424 199804 218476
rect 204720 218424 204772 218476
rect 113640 218288 113692 218340
rect 118148 218288 118200 218340
rect 120264 218288 120316 218340
rect 161480 218288 161532 218340
rect 161664 218288 161716 218340
rect 162768 218288 162820 218340
rect 163320 218288 163372 218340
rect 163964 218288 164016 218340
rect 164976 218288 165028 218340
rect 165528 218288 165580 218340
rect 170772 218288 170824 218340
rect 175280 218288 175332 218340
rect 175740 218288 175792 218340
rect 181444 218288 181496 218340
rect 192024 218288 192076 218340
rect 193588 218288 193640 218340
rect 196440 218288 196492 218340
rect 209688 218288 209740 218340
rect 213184 218288 213236 218340
rect 216312 218424 216364 218476
rect 217324 218424 217376 218476
rect 219808 218424 219860 218476
rect 224040 218424 224092 218476
rect 231032 218424 231084 218476
rect 238024 218424 238076 218476
rect 55680 218152 55732 218204
rect 56508 218152 56560 218204
rect 57428 218152 57480 218204
rect 61384 218152 61436 218204
rect 66444 218152 66496 218204
rect 67548 218152 67600 218204
rect 68100 218152 68152 218204
rect 69572 218152 69624 218204
rect 75552 218152 75604 218204
rect 76564 218152 76616 218204
rect 97080 218152 97132 218204
rect 56508 218016 56560 218068
rect 57244 218016 57296 218068
rect 58164 218016 58216 218068
rect 59360 218016 59412 218068
rect 61476 218016 61528 218068
rect 62764 218016 62816 218068
rect 63960 218016 64012 218068
rect 64788 218016 64840 218068
rect 65616 218016 65668 218068
rect 66168 218016 66220 218068
rect 67272 218016 67324 218068
rect 68284 218016 68336 218068
rect 72240 218016 72292 218068
rect 73712 218016 73764 218068
rect 74724 218016 74776 218068
rect 75828 218016 75880 218068
rect 78036 218016 78088 218068
rect 78588 218016 78640 218068
rect 78864 218016 78916 218068
rect 79968 218016 80020 218068
rect 82176 218016 82228 218068
rect 83464 218016 83516 218068
rect 84660 218016 84712 218068
rect 85304 218016 85356 218068
rect 87144 218016 87196 218068
rect 88248 218016 88300 218068
rect 88800 218016 88852 218068
rect 89444 218016 89496 218068
rect 92940 218016 92992 218068
rect 93584 218016 93636 218068
rect 95424 218016 95476 218068
rect 96252 218016 96304 218068
rect 98736 218016 98788 218068
rect 99288 218016 99340 218068
rect 99564 218016 99616 218068
rect 100668 218016 100720 218068
rect 117596 218152 117648 218204
rect 123392 218152 123444 218204
rect 123576 218152 123628 218204
rect 102876 218084 102928 218136
rect 103428 218084 103480 218136
rect 103704 218016 103756 218068
rect 104808 218016 104860 218068
rect 105360 218016 105412 218068
rect 106004 218016 106056 218068
rect 109500 218016 109552 218068
rect 110420 218016 110472 218068
rect 111984 218016 112036 218068
rect 112812 218016 112864 218068
rect 116124 218016 116176 218068
rect 117228 218016 117280 218068
rect 119436 218016 119488 218068
rect 119988 218016 120040 218068
rect 121920 218016 121972 218068
rect 122564 218016 122616 218068
rect 126060 218016 126112 218068
rect 126704 218016 126756 218068
rect 127716 218016 127768 218068
rect 128268 218016 128320 218068
rect 128544 218016 128596 218068
rect 129372 218016 129424 218068
rect 130200 218016 130252 218068
rect 132500 218016 132552 218068
rect 132684 218016 132736 218068
rect 133512 218016 133564 218068
rect 135996 218016 136048 218068
rect 136548 218016 136600 218068
rect 136916 218152 136968 218204
rect 137284 218016 137336 218068
rect 140136 218016 140188 218068
rect 142436 218016 142488 218068
rect 142620 218016 142672 218068
rect 143264 218016 143316 218068
rect 144276 218016 144328 218068
rect 144828 218016 144880 218068
rect 145104 218016 145156 218068
rect 145932 218016 145984 218068
rect 148416 218016 148468 218068
rect 148876 218016 148928 218068
rect 149244 218016 149296 218068
rect 150072 218016 150124 218068
rect 150440 218152 150492 218204
rect 171416 218152 171468 218204
rect 179328 218152 179380 218204
rect 179880 218152 179932 218204
rect 200396 218152 200448 218204
rect 200580 218152 200632 218204
rect 201500 218152 201552 218204
rect 204720 218152 204772 218204
rect 207664 218152 207716 218204
rect 207848 218152 207900 218204
rect 211804 218152 211856 218204
rect 232872 218288 232924 218340
rect 271144 218424 271196 218476
rect 279240 218424 279292 218476
rect 305552 218560 305604 218612
rect 398472 218560 398524 218612
rect 407764 218560 407816 218612
rect 429936 218560 429988 218612
rect 432696 218560 432748 218612
rect 469864 218560 469916 218612
rect 471244 218560 471296 218612
rect 475568 218560 475620 218612
rect 482836 218560 482888 218612
rect 507676 218560 507728 218612
rect 548708 218560 548760 218612
rect 548892 218560 548944 218612
rect 562600 218560 562652 218612
rect 598112 218696 598164 218748
rect 564164 218560 564216 218612
rect 572536 218560 572588 218612
rect 572674 218560 572726 218612
rect 610716 218560 610768 218612
rect 282184 218424 282236 218476
rect 287888 218424 287940 218476
rect 294144 218424 294196 218476
rect 316684 218424 316736 218476
rect 502800 218424 502852 218476
rect 503168 218424 503220 218476
rect 507860 218424 507912 218476
rect 508044 218424 508096 218476
rect 604460 218424 604512 218476
rect 458180 218356 458232 218408
rect 246120 218288 246172 218340
rect 253204 218288 253256 218340
rect 253388 218288 253440 218340
rect 258080 218288 258132 218340
rect 426624 218288 426676 218340
rect 429568 218288 429620 218340
rect 434904 218288 434956 218340
rect 436652 218288 436704 218340
rect 450728 218288 450780 218340
rect 453856 218288 453908 218340
rect 461308 218288 461360 218340
rect 497464 218288 497516 218340
rect 595996 218288 596048 218340
rect 217968 218152 218020 218204
rect 222752 218152 222804 218204
rect 222936 218152 222988 218204
rect 225604 218152 225656 218204
rect 241980 218152 242032 218204
rect 242900 218152 242952 218204
rect 249432 218152 249484 218204
rect 251732 218152 251784 218204
rect 328920 218152 328972 218204
rect 330484 218152 330536 218204
rect 365352 218152 365404 218204
rect 371792 218152 371844 218204
rect 374460 218152 374512 218204
rect 376024 218152 376076 218204
rect 381912 218152 381964 218204
rect 382924 218152 382976 218204
rect 401784 218152 401836 218204
rect 402796 218152 402848 218204
rect 407580 218152 407632 218204
rect 411904 218152 411956 218204
rect 422484 218152 422536 218204
rect 425428 218152 425480 218204
rect 425796 218152 425848 218204
rect 428464 218152 428516 218204
rect 433248 218152 433300 218204
rect 435272 218152 435324 218204
rect 461952 218152 462004 218204
rect 466276 218152 466328 218204
rect 491944 218152 491996 218204
rect 502248 218152 502300 218204
rect 507124 218152 507176 218204
rect 507676 218152 507728 218204
rect 507860 218152 507912 218204
rect 563060 218152 563112 218204
rect 572674 218152 572726 218204
rect 173256 218016 173308 218068
rect 186228 218016 186280 218068
rect 188160 218016 188212 218068
rect 188896 218016 188948 218068
rect 174268 217880 174320 217932
rect 188896 217880 188948 217932
rect 192024 218016 192076 218068
rect 192300 218016 192352 218068
rect 193036 218016 193088 218068
rect 193956 218016 194008 218068
rect 194508 218016 194560 218068
rect 194784 218016 194836 218068
rect 195888 218016 195940 218068
rect 198924 218016 198976 218068
rect 200028 218016 200080 218068
rect 203064 218016 203116 218068
rect 206284 218016 206336 218068
rect 207204 218016 207256 218068
rect 208124 218016 208176 218068
rect 214656 218016 214708 218068
rect 215208 218016 215260 218068
rect 215484 218016 215536 218068
rect 216128 218016 216180 218068
rect 220084 218016 220136 218068
rect 221280 218016 221332 218068
rect 221832 218016 221884 218068
rect 223764 218016 223816 218068
rect 224592 218016 224644 218068
rect 225420 218016 225472 218068
rect 226156 218016 226208 218068
rect 229560 218016 229612 218068
rect 230480 218016 230532 218068
rect 231216 218016 231268 218068
rect 231676 218016 231728 218068
rect 232044 218016 232096 218068
rect 233148 218016 233200 218068
rect 235356 218016 235408 218068
rect 235816 218016 235868 218068
rect 236184 218016 236236 218068
rect 237288 218016 237340 218068
rect 240324 218016 240376 218068
rect 241336 218016 241388 218068
rect 243636 218016 243688 218068
rect 244096 218016 244148 218068
rect 247776 218016 247828 218068
rect 248236 218016 248288 218068
rect 248604 218016 248656 218068
rect 249616 218016 249668 218068
rect 250260 218016 250312 218068
rect 250904 218016 250956 218068
rect 251916 218016 251968 218068
rect 252468 218016 252520 218068
rect 254400 218016 254452 218068
rect 255044 218016 255096 218068
rect 256056 218016 256108 218068
rect 256516 218016 256568 218068
rect 256884 218016 256936 218068
rect 257528 218016 257580 218068
rect 258540 218016 258592 218068
rect 259276 218016 259328 218068
rect 264336 218016 264388 218068
rect 264796 218016 264848 218068
rect 265164 218016 265216 218068
rect 266176 218016 266228 218068
rect 268476 218016 268528 218068
rect 268936 218016 268988 218068
rect 269304 218016 269356 218068
rect 270224 218016 270276 218068
rect 270960 218016 271012 218068
rect 272524 218016 272576 218068
rect 276756 218016 276808 218068
rect 277216 218016 277268 218068
rect 277584 218016 277636 218068
rect 278596 218016 278648 218068
rect 280896 218016 280948 218068
rect 281448 218016 281500 218068
rect 281724 218016 281776 218068
rect 282460 218016 282512 218068
rect 285036 218016 285088 218068
rect 285496 218016 285548 218068
rect 287520 218016 287572 218068
rect 288716 218016 288768 218068
rect 289176 218016 289228 218068
rect 289728 218016 289780 218068
rect 290004 218016 290056 218068
rect 291108 218016 291160 218068
rect 293316 218016 293368 218068
rect 293776 218016 293828 218068
rect 297456 218016 297508 218068
rect 297916 218016 297968 218068
rect 298284 218016 298336 218068
rect 299112 218016 299164 218068
rect 299940 218016 299992 218068
rect 300676 218016 300728 218068
rect 301596 218016 301648 218068
rect 302148 218016 302200 218068
rect 304080 218016 304132 218068
rect 304724 218016 304776 218068
rect 305736 218016 305788 218068
rect 306196 218016 306248 218068
rect 306564 218016 306616 218068
rect 307668 218016 307720 218068
rect 309876 218016 309928 218068
rect 310428 218016 310480 218068
rect 312360 218016 312412 218068
rect 312912 218016 312964 218068
rect 317328 218016 317380 218068
rect 317972 218016 318024 218068
rect 318984 218016 319036 218068
rect 319628 218016 319680 218068
rect 322296 218016 322348 218068
rect 322848 218016 322900 218068
rect 323124 218016 323176 218068
rect 324136 218016 324188 218068
rect 324780 218016 324832 218068
rect 325424 218016 325476 218068
rect 326436 218016 326488 218068
rect 326896 218016 326948 218068
rect 330576 218016 330628 218068
rect 331036 218016 331088 218068
rect 333060 218016 333112 218068
rect 333888 218016 333940 218068
rect 334716 218016 334768 218068
rect 335176 218016 335228 218068
rect 335544 218016 335596 218068
rect 338672 218016 338724 218068
rect 338856 218016 338908 218068
rect 339408 218016 339460 218068
rect 339684 218016 339736 218068
rect 340696 218016 340748 218068
rect 345480 218016 345532 218068
rect 347044 218016 347096 218068
rect 347964 218016 348016 218068
rect 349068 218016 349120 218068
rect 355416 218016 355468 218068
rect 355876 218016 355928 218068
rect 356244 218016 356296 218068
rect 356980 218016 357032 218068
rect 359556 218016 359608 218068
rect 360108 218016 360160 218068
rect 360384 218016 360436 218068
rect 361028 218016 361080 218068
rect 364524 218016 364576 218068
rect 365536 218016 365588 218068
rect 366180 218016 366232 218068
rect 366732 218016 366784 218068
rect 367836 218016 367888 218068
rect 368388 218016 368440 218068
rect 371976 218016 372028 218068
rect 372528 218016 372580 218068
rect 372804 218016 372856 218068
rect 373448 218016 373500 218068
rect 376116 218016 376168 218068
rect 376668 218016 376720 218068
rect 378600 218016 378652 218068
rect 379244 218016 379296 218068
rect 381084 218016 381136 218068
rect 382096 218016 382148 218068
rect 389364 218016 389416 218068
rect 390008 218016 390060 218068
rect 392676 218016 392728 218068
rect 393136 218016 393188 218068
rect 393504 218016 393556 218068
rect 394516 218016 394568 218068
rect 395160 218016 395212 218068
rect 395804 218016 395856 218068
rect 397644 218016 397696 218068
rect 400772 218016 400824 218068
rect 400956 218016 401008 218068
rect 402244 218016 402296 218068
rect 403440 218016 403492 218068
rect 403992 218016 404044 218068
rect 405096 218016 405148 218068
rect 405556 218016 405608 218068
rect 409236 218016 409288 218068
rect 409788 218016 409840 218068
rect 410064 218016 410116 218068
rect 410708 218016 410760 218068
rect 413376 218016 413428 218068
rect 413836 218016 413888 218068
rect 420000 218016 420052 218068
rect 420920 218016 420972 218068
rect 424140 218016 424192 218068
rect 426992 218016 427044 218068
rect 427452 218016 427504 218068
rect 427912 218016 427964 218068
rect 429108 218016 429160 218068
rect 430580 218016 430632 218068
rect 432420 218016 432472 218068
rect 433708 218016 433760 218068
rect 435732 218016 435784 218068
rect 436284 218016 436336 218068
rect 436560 218016 436612 218068
rect 437480 218016 437532 218068
rect 438216 218016 438268 218068
rect 438860 218016 438912 218068
rect 439872 218016 439924 218068
rect 440332 218016 440384 218068
rect 453304 218016 453356 218068
rect 455420 218016 455472 218068
rect 455604 218016 455656 218068
rect 457168 218016 457220 218068
rect 463148 218016 463200 218068
rect 464620 218016 464672 218068
rect 467288 218016 467340 218068
rect 467932 218016 467984 218068
rect 471428 218016 471480 218068
rect 472900 218016 472952 218068
rect 490380 218016 490432 218068
rect 497004 218016 497056 218068
rect 497464 218016 497516 218068
rect 563336 217948 563388 218000
rect 572352 217948 572404 218000
rect 612280 217948 612332 218000
rect 644940 218016 644992 218068
rect 653588 218016 653640 218068
rect 614488 217948 614540 218000
rect 523040 217812 523092 217864
rect 524236 217812 524288 217864
rect 533436 217676 533488 217728
rect 604000 217812 604052 217864
rect 116952 217540 117004 217592
rect 189172 217540 189224 217592
rect 530952 217540 531004 217592
rect 603448 217676 603500 217728
rect 604460 217676 604512 217728
rect 614304 217676 614356 217728
rect 542360 217540 542412 217592
rect 543280 217540 543332 217592
rect 606208 217540 606260 217592
rect 614120 217540 614172 217592
rect 626632 217540 626684 217592
rect 115296 217404 115348 217456
rect 187976 217404 188028 217456
rect 527824 217404 527876 217456
rect 528468 217404 528520 217456
rect 596916 217404 596968 217456
rect 603080 217404 603132 217456
rect 628288 217404 628340 217456
rect 90410 217200 90462 217252
rect 168564 217268 168616 217320
rect 506112 217268 506164 217320
rect 436100 217200 436152 217252
rect 437342 217200 437394 217252
rect 447140 217200 447192 217252
rect 448106 217200 448158 217252
rect 469312 217200 469364 217252
rect 470462 217200 470514 217252
rect 498200 217200 498252 217252
rect 499442 217200 499494 217252
rect 508550 217132 508602 217184
rect 563060 217132 563112 217184
rect 563336 217268 563388 217320
rect 571984 217268 572036 217320
rect 597928 217268 597980 217320
rect 598112 217268 598164 217320
rect 622400 217268 622452 217320
rect 572674 217132 572726 217184
rect 596548 217132 596600 217184
rect 596916 217132 596968 217184
rect 603080 217132 603132 217184
rect 498614 217064 498666 217116
rect 574192 216996 574244 217048
rect 610072 216996 610124 217048
rect 596364 216860 596416 216912
rect 596548 216860 596600 216912
rect 598480 216860 598532 216912
rect 595996 216724 596048 216776
rect 613384 216860 613436 216912
rect 610716 216724 610768 216776
rect 615684 216724 615736 216776
rect 646320 216044 646372 216096
rect 654784 216044 654836 216096
rect 649632 215908 649684 215960
rect 659108 215908 659160 215960
rect 675852 215364 675904 215416
rect 676956 215364 677008 215416
rect 574744 214820 574796 214872
rect 616880 214820 616932 214872
rect 574376 214684 574428 214736
rect 623320 214684 623372 214736
rect 574560 214548 574612 214600
rect 601792 214412 601844 214464
rect 602344 214412 602396 214464
rect 607312 214548 607364 214600
rect 607864 214548 607916 214600
rect 608784 214548 608836 214600
rect 609520 214548 609572 214600
rect 618260 214548 618312 214600
rect 618904 214548 618956 214600
rect 619916 214548 619968 214600
rect 620560 214548 620612 214600
rect 623964 214548 624016 214600
rect 624424 214412 624476 214464
rect 625436 214548 625488 214600
rect 626080 214548 626132 214600
rect 630036 214548 630088 214600
rect 632888 214548 632940 214600
rect 648252 214548 648304 214600
rect 664444 214548 664496 214600
rect 664812 214548 664864 214600
rect 666008 214548 666060 214600
rect 629392 214412 629444 214464
rect 35808 213936 35860 213988
rect 41696 213936 41748 213988
rect 646044 213868 646096 213920
rect 646504 213868 646556 213920
rect 653220 213868 653272 213920
rect 656164 213868 656216 213920
rect 645492 213732 645544 213784
rect 649816 213732 649868 213784
rect 654140 213732 654192 213784
rect 654784 213732 654836 213784
rect 663156 213732 663208 213784
rect 665824 213732 665876 213784
rect 654600 213256 654652 213308
rect 657544 213256 657596 213308
rect 673736 213256 673788 213308
rect 575480 213188 575532 213240
rect 594800 213188 594852 213240
rect 643836 213188 643888 213240
rect 653404 213188 653456 213240
rect 600688 213120 600740 213172
rect 601240 213120 601292 213172
rect 632704 212984 632756 213036
rect 634360 212984 634412 213036
rect 664260 212984 664312 213036
rect 665088 212984 665140 213036
rect 673552 213188 673604 213240
rect 673552 213052 673604 213104
rect 673736 212916 673788 212968
rect 658188 212848 658240 212900
rect 658924 212848 658976 212900
rect 650460 212712 650512 212764
rect 651288 212712 651340 212764
rect 35808 212644 35860 212696
rect 39580 212644 39632 212696
rect 591304 212644 591356 212696
rect 639880 212644 639932 212696
rect 659568 212644 659620 212696
rect 662420 212644 662472 212696
rect 592684 212508 592736 212560
rect 641720 212508 641772 212560
rect 656532 212508 656584 212560
rect 657912 212508 657964 212560
rect 578516 211148 578568 211200
rect 580908 211148 580960 211200
rect 600412 210400 600464 210452
rect 601010 210400 601062 210452
rect 35808 209924 35860 209976
rect 40132 209924 40184 209976
rect 579528 209788 579580 209840
rect 582288 209788 582340 209840
rect 35624 208632 35676 208684
rect 39764 208632 39816 208684
rect 581644 208564 581696 208616
rect 632152 209516 632204 209568
rect 652024 209516 652076 209568
rect 667020 209040 667072 209092
rect 35808 208360 35860 208412
rect 40040 208360 40092 208412
rect 578884 208292 578936 208344
rect 589464 208292 589516 208344
rect 35808 207136 35860 207188
rect 40132 207136 40184 207188
rect 580908 206864 580960 206916
rect 589464 206864 589516 206916
rect 35808 205776 35860 205828
rect 40224 205776 40276 205828
rect 579528 205776 579580 205828
rect 581000 205776 581052 205828
rect 582288 205504 582340 205556
rect 589464 205504 589516 205556
rect 35808 204416 35860 204468
rect 41512 204416 41564 204468
rect 35624 204280 35676 204332
rect 41696 204280 41748 204332
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 35808 202852 35860 202904
rect 37924 202852 37976 202904
rect 578332 202852 578384 202904
rect 580264 202852 580316 202904
rect 581000 202784 581052 202836
rect 589464 202784 589516 202836
rect 578792 200132 578844 200184
rect 590384 200132 590436 200184
rect 580264 199996 580316 200048
rect 589464 199996 589516 200048
rect 579528 198704 579580 198756
rect 589464 198704 589516 198756
rect 578516 195984 578568 196036
rect 589280 195984 589332 196036
rect 579528 194556 579580 194608
rect 589464 194556 589516 194608
rect 579528 191836 579580 191888
rect 589464 191836 589516 191888
rect 579528 190476 579580 190528
rect 590568 190476 590620 190528
rect 579528 187688 579580 187740
rect 589464 187688 589516 187740
rect 42432 187416 42484 187468
rect 43260 187416 43312 187468
rect 579528 186260 579580 186312
rect 589648 186260 589700 186312
rect 579528 184832 579580 184884
rect 589464 184832 589516 184884
rect 669228 184832 669280 184884
rect 670700 184832 670752 184884
rect 42156 183472 42208 183524
rect 42984 183472 43036 183524
rect 579528 182112 579580 182164
rect 589464 182112 589516 182164
rect 578792 180752 578844 180804
rect 590568 180752 590620 180804
rect 578792 178032 578844 178084
rect 589464 178032 589516 178084
rect 668216 177964 668268 178016
rect 670792 177964 670844 178016
rect 579528 177896 579580 177948
rect 589648 177896 589700 177948
rect 579988 175244 580040 175296
rect 589464 175312 589516 175364
rect 667940 174700 667992 174752
rect 669596 174700 669648 174752
rect 578424 174496 578476 174548
rect 589648 174496 589700 174548
rect 578240 172864 578292 172916
rect 579988 172864 580040 172916
rect 580908 172524 580960 172576
rect 589464 172524 589516 172576
rect 580264 171096 580316 171148
rect 589464 171096 589516 171148
rect 578700 169736 578752 169788
rect 580908 169736 580960 169788
rect 667940 169668 667992 169720
rect 669780 169668 669832 169720
rect 582380 168376 582432 168428
rect 589464 168376 589516 168428
rect 578240 167288 578292 167340
rect 580264 167288 580316 167340
rect 579988 167016 580040 167068
rect 589464 167016 589516 167068
rect 579528 166268 579580 166320
rect 589648 166268 589700 166320
rect 579344 165180 579396 165232
rect 582380 165180 582432 165232
rect 668032 164908 668084 164960
rect 670332 164908 670384 164960
rect 582472 164228 582524 164280
rect 589464 164228 589516 164280
rect 578240 163616 578292 163668
rect 579988 163616 580040 163668
rect 675852 163208 675904 163260
rect 679624 163208 679676 163260
rect 580908 162868 580960 162920
rect 589464 162868 589516 162920
rect 676036 162732 676088 162784
rect 681004 162732 681056 162784
rect 578424 162664 578476 162716
rect 582472 162664 582524 162716
rect 580540 161440 580592 161492
rect 589464 161440 589516 161492
rect 580724 160080 580776 160132
rect 589464 160080 589516 160132
rect 668216 160012 668268 160064
rect 670792 160012 670844 160064
rect 578884 158720 578936 158772
rect 580908 158720 580960 158772
rect 585784 158720 585836 158772
rect 589464 158720 589516 158772
rect 587164 157360 587216 157412
rect 589280 157360 589332 157412
rect 668216 155116 668268 155168
rect 670792 155116 670844 155168
rect 578332 154776 578384 154828
rect 580540 154776 580592 154828
rect 584404 154572 584456 154624
rect 589464 154572 589516 154624
rect 583024 153212 583076 153264
rect 589464 153212 589516 153264
rect 578240 152736 578292 152788
rect 580724 152736 580776 152788
rect 580264 151784 580316 151836
rect 589464 151784 589516 151836
rect 578884 150560 578936 150612
rect 585784 150560 585836 150612
rect 585140 149064 585192 149116
rect 589464 149064 589516 149116
rect 579528 148316 579580 148368
rect 587164 148316 587216 148368
rect 578884 146276 578936 146328
rect 585140 146276 585192 146328
rect 668768 146004 668820 146056
rect 670792 146004 670844 146056
rect 584772 144916 584824 144968
rect 589464 144916 589516 144968
rect 579252 144644 579304 144696
rect 584404 144644 584456 144696
rect 585968 143556 586020 143608
rect 589464 143556 589516 143608
rect 579528 143420 579580 143472
rect 583024 143420 583076 143472
rect 587164 142400 587216 142452
rect 589832 142400 589884 142452
rect 580448 140768 580500 140820
rect 589464 140768 589516 140820
rect 578608 140700 578660 140752
rect 580264 140700 580316 140752
rect 583024 139408 583076 139460
rect 589464 139408 589516 139460
rect 578608 139272 578660 139324
rect 589924 139272 589976 139324
rect 579528 138660 579580 138712
rect 588544 138660 588596 138712
rect 579068 137300 579120 137352
rect 584772 137300 584824 137352
rect 584588 136620 584640 136672
rect 589464 136620 589516 136672
rect 580264 134512 580316 134564
rect 589464 134512 589516 134564
rect 667940 133764 667992 133816
rect 669964 133764 670016 133816
rect 585784 132472 585836 132524
rect 589464 132472 589516 132524
rect 581828 131248 581880 131300
rect 589464 131248 589516 131300
rect 578884 131112 578936 131164
rect 585968 131112 586020 131164
rect 668676 130636 668728 130688
rect 670792 130636 670844 130688
rect 667940 129548 667992 129600
rect 670148 129548 670200 129600
rect 583208 129140 583260 129192
rect 590384 129140 590436 129192
rect 579528 129004 579580 129056
rect 587164 129004 587216 129056
rect 579068 126964 579120 127016
rect 589464 126964 589516 127016
rect 578332 125604 578384 125656
rect 580448 125604 580500 125656
rect 580448 124176 580500 124228
rect 589464 124176 589516 124228
rect 578424 123564 578476 123616
rect 583024 123564 583076 123616
rect 584404 122816 584456 122868
rect 589464 122816 589516 122868
rect 578884 122136 578936 122188
rect 584588 122136 584640 122188
rect 580632 122000 580684 122052
rect 589924 122000 589976 122052
rect 675852 120028 675904 120080
rect 676404 120028 676456 120080
rect 587348 118668 587400 118720
rect 590016 118668 590068 118720
rect 578516 118396 578568 118448
rect 580264 118396 580316 118448
rect 579528 116900 579580 116952
rect 583208 116900 583260 116952
rect 586152 115948 586204 116000
rect 589464 115948 589516 116000
rect 583208 115200 583260 115252
rect 589648 115200 589700 115252
rect 579252 114452 579304 114504
rect 581644 114452 581696 114504
rect 583024 113160 583076 113212
rect 589464 113160 589516 113212
rect 668124 112888 668176 112940
rect 670148 112888 670200 112940
rect 579528 112820 579580 112872
rect 585784 112820 585836 112872
rect 585968 112412 586020 112464
rect 590108 112412 590160 112464
rect 581644 110440 581696 110492
rect 589464 110440 589516 110492
rect 579344 110100 579396 110152
rect 581828 110100 581880 110152
rect 584588 109012 584640 109064
rect 589280 109012 589332 109064
rect 578332 108672 578384 108724
rect 580632 108672 580684 108724
rect 668400 107992 668452 108044
rect 670792 107992 670844 108044
rect 578884 107584 578936 107636
rect 589464 107652 589516 107704
rect 587164 106292 587216 106344
rect 589832 106292 589884 106344
rect 580264 104864 580316 104916
rect 589464 104864 589516 104916
rect 667940 104524 667992 104576
rect 669964 104524 670016 104576
rect 579528 103436 579580 103488
rect 588544 103436 588596 103488
rect 579528 101804 579580 101856
rect 584404 101804 584456 101856
rect 584404 100104 584456 100156
rect 589464 100104 589516 100156
rect 579068 99356 579120 99408
rect 586152 99356 586204 99408
rect 622308 99288 622360 99340
rect 630772 99288 630824 99340
rect 578608 99220 578660 99272
rect 580448 99220 580500 99272
rect 623688 99152 623740 99204
rect 633440 99152 633492 99204
rect 577504 99084 577556 99136
rect 595260 99084 595312 99136
rect 625068 99016 625120 99068
rect 636292 99016 636344 99068
rect 628288 98880 628340 98932
rect 642180 98880 642232 98932
rect 629024 98744 629076 98796
rect 643652 98744 643704 98796
rect 647148 98608 647200 98660
rect 661960 98608 662012 98660
rect 630496 98472 630548 98524
rect 646596 98472 646648 98524
rect 631048 98200 631100 98252
rect 640708 98132 640760 98184
rect 578332 97928 578384 97980
rect 587348 97928 587400 97980
rect 620192 97928 620244 97980
rect 626264 97928 626316 97980
rect 629760 97928 629812 97980
rect 645308 97996 645360 98048
rect 659200 97928 659252 97980
rect 663892 97928 663944 97980
rect 618720 97792 618772 97844
rect 625804 97792 625856 97844
rect 627552 97792 627604 97844
rect 631048 97792 631100 97844
rect 634176 97792 634228 97844
rect 650552 97792 650604 97844
rect 655428 97792 655480 97844
rect 634728 97656 634780 97708
rect 650184 97656 650236 97708
rect 651840 97656 651892 97708
rect 659568 97656 659620 97708
rect 659936 97792 659988 97844
rect 665180 97792 665232 97844
rect 662512 97656 662564 97708
rect 621664 97520 621716 97572
rect 629300 97520 629352 97572
rect 631968 97520 632020 97572
rect 647516 97520 647568 97572
rect 650368 97452 650420 97504
rect 658280 97452 658332 97504
rect 612648 97384 612700 97436
rect 618904 97384 618956 97436
rect 623136 97384 623188 97436
rect 632060 97384 632112 97436
rect 633256 97384 633308 97436
rect 648620 97384 648672 97436
rect 658096 97316 658148 97368
rect 663064 97316 663116 97368
rect 605472 97248 605524 97300
rect 611912 97248 611964 97300
rect 626080 97248 626132 97300
rect 637764 97248 637816 97300
rect 644296 97248 644348 97300
rect 626816 97112 626868 97164
rect 639236 97112 639288 97164
rect 643008 97112 643060 97164
rect 624608 96976 624660 97028
rect 635004 96976 635056 97028
rect 635556 96976 635608 97028
rect 647700 96976 647752 97028
rect 598940 96908 598992 96960
rect 599676 96908 599728 96960
rect 606208 96908 606260 96960
rect 607128 96908 607180 96960
rect 615776 96908 615828 96960
rect 616788 96908 616840 96960
rect 612096 96840 612148 96892
rect 612648 96840 612700 96892
rect 617248 96840 617300 96892
rect 618168 96840 618220 96892
rect 632704 96840 632756 96892
rect 648252 96840 648304 96892
rect 653956 96840 654008 96892
rect 654600 96840 654652 96892
rect 654784 96840 654836 96892
rect 655428 96840 655480 96892
rect 656808 97180 656860 97232
rect 661408 97180 661460 97232
rect 658832 97044 658884 97096
rect 656716 96908 656768 96960
rect 660120 96908 660172 96960
rect 660120 96772 660172 96824
rect 610624 96704 610676 96756
rect 611268 96704 611320 96756
rect 640524 96568 640576 96620
rect 647884 96704 647936 96756
rect 645768 96568 645820 96620
rect 656348 96568 656400 96620
rect 639052 96432 639104 96484
rect 645124 96432 645176 96484
rect 646412 96432 646464 96484
rect 652024 96432 652076 96484
rect 652576 96432 652628 96484
rect 665548 96432 665600 96484
rect 631232 96296 631284 96348
rect 647148 96296 647200 96348
rect 648896 96296 648948 96348
rect 664168 96296 664220 96348
rect 637580 96160 637632 96212
rect 660672 96160 660724 96212
rect 611084 96024 611136 96076
rect 622124 96024 622176 96076
rect 649908 96024 649960 96076
rect 663708 96024 663760 96076
rect 644940 95956 644992 96008
rect 649080 95956 649132 96008
rect 607680 95888 607732 95940
rect 624976 95888 625028 95940
rect 643468 95820 643520 95872
rect 649264 95820 649316 95872
rect 665364 95888 665416 95940
rect 638592 95684 638644 95736
rect 647332 95684 647384 95736
rect 647884 95684 647936 95736
rect 653312 95616 653364 95668
rect 664352 95616 664404 95668
rect 640064 95548 640116 95600
rect 647884 95548 647936 95600
rect 641536 95412 641588 95464
rect 645124 95412 645176 95464
rect 651840 95412 651892 95464
rect 649908 95276 649960 95328
rect 620928 95140 620980 95192
rect 626448 95140 626500 95192
rect 647700 95140 647752 95192
rect 648804 95140 648856 95192
rect 579528 95004 579580 95056
rect 583208 95004 583260 95056
rect 616512 95004 616564 95056
rect 623044 95004 623096 95056
rect 609152 94460 609204 94512
rect 620284 94460 620336 94512
rect 619548 93780 619600 93832
rect 626448 93780 626500 93832
rect 651288 93508 651340 93560
rect 655428 93508 655480 93560
rect 578516 93440 578568 93492
rect 585968 93440 586020 93492
rect 649080 93236 649132 93288
rect 656164 93236 656216 93288
rect 611268 93100 611320 93152
rect 619272 93100 619324 93152
rect 606944 92828 606996 92880
rect 610072 92828 610124 92880
rect 648620 92488 648672 92540
rect 650000 92488 650052 92540
rect 617984 92420 618036 92472
rect 626448 92420 626500 92472
rect 647332 92352 647384 92404
rect 654324 92352 654376 92404
rect 579344 91060 579396 91112
rect 584588 91060 584640 91112
rect 618168 90992 618220 91044
rect 626448 90992 626500 91044
rect 651840 90652 651892 90704
rect 655428 90652 655480 90704
rect 623044 89632 623096 89684
rect 626448 89564 626500 89616
rect 585140 88952 585192 89004
rect 589924 88952 589976 89004
rect 649724 88748 649776 88800
rect 658556 88748 658608 88800
rect 662328 88748 662380 88800
rect 663892 88748 663944 88800
rect 656348 88612 656400 88664
rect 657452 88612 657504 88664
rect 610072 88272 610124 88324
rect 626448 88272 626500 88324
rect 655244 88272 655296 88324
rect 658464 88272 658516 88324
rect 622124 88136 622176 88188
rect 626264 88136 626316 88188
rect 579528 88068 579580 88120
rect 585140 88068 585192 88120
rect 648436 86980 648488 87032
rect 662512 86980 662564 87032
rect 656716 86844 656768 86896
rect 659568 86844 659620 86896
rect 649264 86708 649316 86760
rect 661408 86708 661460 86760
rect 647884 86572 647936 86624
rect 660120 86572 660172 86624
rect 656164 86436 656216 86488
rect 660672 86436 660724 86488
rect 619272 86300 619324 86352
rect 626448 86300 626500 86352
rect 652024 86300 652076 86352
rect 657176 86300 657228 86352
rect 620284 85484 620336 85536
rect 626448 85484 626500 85536
rect 609888 85348 609940 85400
rect 625344 85280 625396 85332
rect 579160 84124 579212 84176
rect 581644 84124 581696 84176
rect 608508 84124 608560 84176
rect 625804 84124 625856 84176
rect 579068 82356 579120 82408
rect 583024 82356 583076 82408
rect 579528 82084 579580 82136
rect 587164 82084 587216 82136
rect 628748 80928 628800 80980
rect 642456 80928 642508 80980
rect 612648 80792 612700 80844
rect 647424 80792 647476 80844
rect 595444 80656 595496 80708
rect 636752 80656 636804 80708
rect 629208 79976 629260 80028
rect 633440 79976 633492 80028
rect 613752 79432 613804 79484
rect 645952 79432 646004 79484
rect 579068 79296 579120 79348
rect 588728 79296 588780 79348
rect 613936 79296 613988 79348
rect 646504 79296 646556 79348
rect 633440 78072 633492 78124
rect 645308 78072 645360 78124
rect 631048 77936 631100 77988
rect 643100 77936 643152 77988
rect 628472 77732 628524 77784
rect 632796 77732 632848 77784
rect 625804 77256 625856 77308
rect 631048 77256 631100 77308
rect 616788 76644 616840 76696
rect 646320 76644 646372 76696
rect 612004 76508 612056 76560
rect 662420 76508 662472 76560
rect 578240 75828 578292 75880
rect 580264 75828 580316 75880
rect 618904 75420 618956 75472
rect 648620 75420 648672 75472
rect 615408 75284 615460 75336
rect 646872 75284 646924 75336
rect 607128 75148 607180 75200
rect 646136 75148 646188 75200
rect 578884 72428 578936 72480
rect 601700 72428 601752 72480
rect 579068 71340 579120 71392
rect 584404 71340 584456 71392
rect 580264 68280 580316 68332
rect 604460 68280 604512 68332
rect 577504 59984 577556 60036
rect 603080 59984 603132 60036
rect 576124 58624 576176 58676
rect 601884 58624 601936 58676
rect 574928 57196 574980 57248
rect 600504 57196 600556 57248
rect 574560 55972 574612 56024
rect 598940 55972 598992 56024
rect 574744 55836 574796 55888
rect 600320 55836 600372 55888
rect 596456 55156 596508 55208
rect 597652 55020 597704 55072
rect 597928 54884 597980 54936
rect 463240 53592 463292 53644
rect 464068 53592 464120 53644
rect 464252 53592 464304 53644
rect 459468 53456 459520 53508
rect 599124 54748 599176 54800
rect 624424 54612 624476 54664
rect 625804 54476 625856 54528
rect 596180 54340 596232 54392
rect 465264 53592 465316 53644
rect 465448 53592 465500 53644
rect 464988 53456 465040 53508
rect 581644 54204 581696 54256
rect 574744 54068 574796 54120
rect 466368 53592 466420 53644
rect 467104 53592 467156 53644
rect 471060 53592 471112 53644
rect 574560 53932 574612 53984
rect 463056 53320 463108 53372
rect 574928 53796 574980 53848
rect 50528 53184 50580 53236
rect 130384 53184 130436 53236
rect 463240 53184 463292 53236
rect 463792 53184 463844 53236
rect 312360 53116 312412 53168
rect 313740 53116 313792 53168
rect 316316 53116 316368 53168
rect 317696 53116 317748 53168
rect 48964 53048 49016 53100
rect 130568 53048 130620 53100
rect 463608 53048 463660 53100
rect 464252 53048 464304 53100
rect 465448 53048 465500 53100
rect 466368 53048 466420 53100
rect 461308 52912 461360 52964
rect 471060 52912 471112 52964
rect 461906 52776 461958 52828
rect 467104 52776 467156 52828
rect 47584 51960 47636 52012
rect 130752 51960 130804 52012
rect 50344 51824 50396 51876
rect 129004 51824 129056 51876
rect 129648 51824 129700 51876
rect 591304 51824 591356 51876
rect 128820 51688 128872 51740
rect 592684 51688 592736 51740
rect 318340 50464 318392 50516
rect 458180 50464 458232 50516
rect 46204 50328 46256 50380
rect 131028 50328 131080 50380
rect 314016 50328 314068 50380
rect 458364 50328 458416 50380
rect 522948 50328 523000 50380
rect 544016 50328 544068 50380
rect 49148 49104 49200 49156
rect 129280 49104 129332 49156
rect 45468 48968 45520 49020
rect 129464 48968 129516 49020
rect 130568 46044 130620 46096
rect 132316 46044 132368 46096
rect 130752 45500 130804 45552
rect 132592 45500 132644 45552
rect 129464 45364 129516 45416
rect 129648 45024 129700 45076
rect 129280 44888 129332 44940
rect 128820 44752 128872 44804
rect 131672 44616 131724 44668
rect 129004 44412 129056 44464
rect 43628 44276 43680 44328
rect 132592 44364 132644 44416
rect 132500 44252 132552 44304
rect 132776 44252 132828 44304
rect 43444 44140 43496 44192
rect 131672 44140 131724 44192
rect 131028 44004 131080 44056
rect 440240 43800 440292 43852
rect 441068 43800 441120 43852
rect 187332 42780 187384 42832
rect 255872 42780 255924 42832
rect 307300 42712 307352 42764
rect 431224 42712 431276 42764
rect 441068 42712 441120 42764
rect 449164 42712 449216 42764
rect 453580 42712 453632 42764
rect 464160 42712 464212 42764
rect 310428 42576 310480 42628
rect 427084 42576 427136 42628
rect 441252 42576 441304 42628
rect 446404 42576 446456 42628
rect 454500 42440 454552 42492
rect 463056 42440 463108 42492
rect 404452 42304 404504 42356
rect 405188 42304 405240 42356
rect 420736 42304 420788 42356
rect 426900 42304 426952 42356
rect 661408 42129 661460 42181
rect 427084 41964 427136 42016
rect 431224 41964 431276 42016
rect 441068 41964 441120 42016
rect 446404 41964 446456 42016
rect 454500 41964 454552 42016
rect 441252 41828 441304 41880
rect 449164 41828 449216 41880
rect 453580 41828 453632 41880
rect 404452 41420 404504 41472
rect 420736 41420 420788 41472
rect 426900 41420 426952 41472
rect 459192 41420 459244 41472
<< metal2 >>
rect 703694 897668 703722 897804
rect 704154 897668 704182 897804
rect 704614 897668 704642 897804
rect 705074 897668 705102 897804
rect 705534 897668 705562 897804
rect 705994 897668 706022 897804
rect 706454 897668 706482 897804
rect 706914 897668 706942 897804
rect 707374 897668 707402 897804
rect 707834 897668 707862 897804
rect 708294 897668 708322 897804
rect 708754 897668 708782 897804
rect 709214 897668 709242 897804
rect 676034 897152 676090 897161
rect 676034 897087 676036 897096
rect 676088 897087 676090 897096
rect 676036 897058 676088 897064
rect 652024 897048 652076 897054
rect 652024 896990 652076 896996
rect 651472 868896 651524 868902
rect 651472 868838 651524 868844
rect 651484 868601 651512 868838
rect 651470 868592 651526 868601
rect 651470 868527 651526 868536
rect 652036 867649 652064 896990
rect 675850 896744 675906 896753
rect 675850 896679 675906 896688
rect 675864 895830 675892 896679
rect 676034 896336 676090 896345
rect 676034 896271 676090 896280
rect 654784 895824 654836 895830
rect 654784 895766 654836 895772
rect 675852 895824 675904 895830
rect 675852 895766 675904 895772
rect 653404 880524 653456 880530
rect 653404 880466 653456 880472
rect 652022 867640 652078 867649
rect 652022 867575 652078 867584
rect 651472 866652 651524 866658
rect 651472 866594 651524 866600
rect 651484 866289 651512 866594
rect 651470 866280 651526 866289
rect 651470 866215 651526 866224
rect 653416 865230 653444 880466
rect 654796 868902 654824 895766
rect 676048 895694 676076 896271
rect 672724 895688 672776 895694
rect 672724 895630 672776 895636
rect 676036 895688 676088 895694
rect 676036 895630 676088 895636
rect 671068 894464 671120 894470
rect 671068 894406 671120 894412
rect 670884 886916 670936 886922
rect 670884 886858 670936 886864
rect 657544 869440 657596 869446
rect 657544 869382 657596 869388
rect 654784 868896 654836 868902
rect 654784 868838 654836 868844
rect 654140 868080 654192 868086
rect 654140 868022 654192 868028
rect 651380 865224 651432 865230
rect 651378 865192 651380 865201
rect 653404 865224 653456 865230
rect 651432 865192 651434 865201
rect 653404 865166 653456 865172
rect 651378 865127 651434 865136
rect 651472 863864 651524 863870
rect 651470 863832 651472 863841
rect 651524 863832 651526 863841
rect 651470 863767 651526 863776
rect 654152 862510 654180 868022
rect 657556 863870 657584 869382
rect 657544 863864 657596 863870
rect 657544 863806 657596 863812
rect 651472 862504 651524 862510
rect 651472 862446 651524 862452
rect 654140 862504 654192 862510
rect 654140 862446 654192 862452
rect 651484 862345 651512 862446
rect 651470 862336 651526 862345
rect 651470 862271 651526 862280
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35622 818000 35678 818009
rect 35622 817935 35678 817944
rect 35636 817018 35664 817935
rect 35806 817320 35862 817329
rect 35806 817255 35862 817264
rect 35820 817154 35848 817255
rect 35808 817148 35860 817154
rect 35808 817090 35860 817096
rect 44824 817148 44876 817154
rect 44824 817090 44876 817096
rect 35624 817012 35676 817018
rect 35624 816954 35676 816960
rect 35438 816912 35494 816921
rect 35438 816847 35494 816856
rect 35452 815658 35480 816847
rect 35806 816096 35862 816105
rect 35806 816031 35862 816040
rect 35820 815794 35848 816031
rect 35808 815788 35860 815794
rect 35808 815730 35860 815736
rect 43076 815788 43128 815794
rect 43076 815730 43128 815736
rect 35440 815652 35492 815658
rect 35440 815594 35492 815600
rect 35622 815280 35678 815289
rect 35622 815215 35678 815224
rect 35636 814434 35664 815215
rect 35806 814464 35862 814473
rect 35624 814428 35676 814434
rect 35806 814399 35862 814408
rect 42892 814428 42944 814434
rect 35624 814370 35676 814376
rect 35820 814298 35848 814399
rect 42892 814370 42944 814376
rect 35808 814292 35860 814298
rect 35808 814234 35860 814240
rect 42904 814214 42932 814370
rect 42904 814186 43024 814214
rect 41326 813648 41382 813657
rect 41326 813583 41382 813592
rect 41340 812870 41368 813583
rect 41328 812864 41380 812870
rect 40958 812832 41014 812841
rect 41328 812806 41380 812812
rect 40958 812767 41014 812776
rect 32402 811608 32458 811617
rect 32402 811543 32458 811552
rect 31022 809976 31078 809985
rect 31022 809911 31078 809920
rect 31036 801106 31064 809911
rect 32416 802466 32444 811543
rect 40972 811442 41000 812767
rect 41142 812424 41198 812433
rect 41142 812359 41198 812368
rect 40960 811436 41012 811442
rect 40960 811378 41012 811384
rect 34518 811200 34574 811209
rect 34518 811135 34574 811144
rect 33782 809568 33838 809577
rect 33782 809503 33838 809512
rect 32404 802460 32456 802466
rect 32404 802402 32456 802408
rect 33796 801242 33824 809503
rect 34532 802602 34560 811135
rect 40958 808752 41014 808761
rect 40958 808687 41014 808696
rect 40684 808648 40736 808654
rect 40684 808590 40736 808596
rect 34520 802596 34572 802602
rect 34520 802538 34572 802544
rect 33784 801236 33836 801242
rect 33784 801178 33836 801184
rect 31024 801100 31076 801106
rect 31024 801042 31076 801048
rect 40696 800601 40724 808590
rect 40972 805225 41000 808687
rect 41156 808110 41184 812359
rect 42616 811436 42668 811442
rect 42616 811378 42668 811384
rect 41970 810792 42026 810801
rect 41970 810727 42026 810736
rect 41786 809160 41842 809169
rect 41786 809095 41842 809104
rect 41800 808654 41828 809095
rect 41788 808648 41840 808654
rect 41788 808590 41840 808596
rect 41144 808104 41196 808110
rect 41144 808046 41196 808052
rect 41604 808104 41656 808110
rect 41604 808046 41656 808052
rect 41142 807936 41198 807945
rect 41142 807871 41198 807880
rect 41156 807362 41184 807871
rect 41144 807356 41196 807362
rect 41144 807298 41196 807304
rect 41142 806712 41198 806721
rect 41142 806647 41198 806656
rect 41156 806002 41184 806647
rect 41326 806304 41382 806313
rect 41326 806239 41382 806248
rect 41340 806138 41368 806239
rect 41328 806132 41380 806138
rect 41328 806074 41380 806080
rect 41144 805996 41196 806002
rect 41144 805938 41196 805944
rect 40958 805216 41014 805225
rect 40958 805151 41014 805160
rect 41616 804681 41644 808046
rect 41984 805633 42012 810727
rect 42154 810384 42210 810393
rect 42154 810319 42210 810328
rect 41970 805624 42026 805633
rect 41970 805559 42026 805568
rect 42168 804953 42196 810319
rect 42154 804944 42210 804953
rect 42154 804879 42210 804888
rect 41602 804672 41658 804681
rect 41602 804607 41658 804616
rect 42628 804554 42656 811378
rect 42996 804554 43024 814186
rect 42260 804526 42656 804554
rect 42904 804526 43024 804554
rect 41788 802596 41840 802602
rect 41788 802538 41840 802544
rect 40682 800592 40738 800601
rect 40682 800527 40738 800536
rect 41800 800329 41828 802538
rect 41786 800320 41842 800329
rect 41786 800255 41842 800264
rect 41786 799912 41842 799921
rect 41786 799847 41842 799856
rect 41800 799445 41828 799847
rect 42260 797619 42288 804526
rect 42708 802460 42760 802466
rect 42708 802402 42760 802408
rect 42720 801794 42748 802402
rect 42720 801766 42840 801794
rect 42616 801236 42668 801242
rect 42616 801178 42668 801184
rect 42432 799128 42484 799134
rect 42432 799070 42484 799076
rect 42182 797591 42288 797619
rect 42444 796974 42472 799070
rect 42628 798946 42656 801178
rect 42182 796946 42472 796974
rect 42536 798918 42656 798946
rect 42536 795779 42564 798918
rect 42182 795751 42564 795779
rect 42432 795660 42484 795666
rect 42432 795602 42484 795608
rect 42444 795138 42472 795602
rect 42182 795110 42472 795138
rect 42248 795048 42300 795054
rect 42248 794990 42300 794996
rect 42260 794894 42288 794990
rect 42260 794866 42380 794894
rect 42352 794594 42380 794866
rect 42182 794566 42380 794594
rect 41786 794472 41842 794481
rect 41786 794407 41842 794416
rect 41800 793900 41828 794407
rect 42248 793824 42300 793830
rect 42168 793772 42248 793778
rect 42168 793766 42300 793772
rect 42168 793750 42288 793766
rect 42168 793288 42196 793750
rect 42812 793642 42840 801766
rect 42260 793614 42840 793642
rect 42260 792758 42288 793614
rect 42616 793552 42668 793558
rect 42430 793520 42486 793529
rect 42616 793494 42668 793500
rect 42430 793455 42486 793464
rect 42182 792730 42288 792758
rect 42246 792024 42302 792033
rect 42246 791959 42302 791968
rect 42260 790514 42288 791959
rect 42444 790634 42472 793455
rect 42432 790628 42484 790634
rect 42432 790570 42484 790576
rect 42260 790486 42380 790514
rect 42156 790424 42208 790430
rect 42156 790366 42208 790372
rect 42168 790228 42196 790366
rect 42352 790242 42380 790486
rect 42260 790214 42380 790242
rect 42260 789818 42288 790214
rect 42248 789812 42300 789818
rect 42248 789754 42300 789760
rect 42628 789698 42656 793494
rect 42168 789670 42656 789698
rect 42168 789616 42196 789670
rect 42522 789576 42578 789585
rect 42248 789540 42300 789546
rect 42522 789511 42578 789520
rect 42248 789482 42300 789488
rect 42260 789290 42288 789482
rect 42536 789426 42564 789511
rect 42168 789262 42288 789290
rect 42444 789398 42564 789426
rect 42168 788936 42196 789262
rect 42246 788896 42302 788905
rect 42246 788831 42302 788840
rect 41878 788624 41934 788633
rect 41878 788559 41934 788568
rect 41892 788392 41920 788559
rect 42260 786570 42288 788831
rect 42182 786542 42288 786570
rect 42444 785958 42472 789398
rect 42614 789304 42670 789313
rect 42614 789239 42670 789248
rect 42168 785890 42196 785944
rect 42260 785930 42472 785958
rect 42260 785890 42288 785930
rect 42168 785862 42288 785890
rect 42628 785754 42656 789239
rect 42352 785726 42656 785754
rect 42352 785278 42380 785726
rect 42524 785664 42576 785670
rect 42524 785606 42576 785612
rect 42182 785250 42380 785278
rect 42536 785234 42564 785606
rect 42444 785206 42564 785234
rect 42444 784734 42472 785206
rect 42182 784706 42472 784734
rect 42904 779714 42932 804526
rect 43088 794894 43116 815730
rect 43444 815652 43496 815658
rect 43444 815594 43496 815600
rect 43258 808344 43314 808353
rect 43258 808279 43314 808288
rect 43272 794894 43300 808279
rect 43456 807974 43484 815594
rect 44180 814292 44232 814298
rect 44180 814234 44232 814240
rect 43444 807968 43496 807974
rect 43444 807910 43496 807916
rect 43810 807528 43866 807537
rect 43810 807463 43866 807472
rect 43444 801100 43496 801106
rect 43444 801042 43496 801048
rect 42996 794866 43116 794894
rect 43180 794866 43300 794894
rect 42996 785234 43024 794866
rect 43180 793830 43208 794866
rect 43168 793824 43220 793830
rect 43168 793766 43220 793772
rect 43456 793558 43484 801042
rect 43628 797700 43680 797706
rect 43628 797642 43680 797648
rect 43640 795666 43668 797642
rect 43628 795660 43680 795666
rect 43628 795602 43680 795608
rect 43444 793552 43496 793558
rect 43444 793494 43496 793500
rect 42996 785206 43208 785234
rect 42812 779686 42932 779714
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 774752 35862 774761
rect 35806 774687 35862 774696
rect 35820 774246 35848 774687
rect 35808 774240 35860 774246
rect 35808 774182 35860 774188
rect 41696 774240 41748 774246
rect 42064 774240 42116 774246
rect 41748 774188 42064 774194
rect 41696 774182 42116 774188
rect 41708 774166 42104 774182
rect 35346 773936 35402 773945
rect 35346 773871 35402 773880
rect 35360 772886 35388 773871
rect 35530 773528 35586 773537
rect 35530 773463 35586 773472
rect 35806 773528 35862 773537
rect 35806 773463 35862 773472
rect 41694 773528 41750 773537
rect 41694 773463 41750 773472
rect 35544 773022 35572 773463
rect 35820 773362 35848 773463
rect 41708 773362 41736 773463
rect 35808 773356 35860 773362
rect 35808 773298 35860 773304
rect 41696 773356 41748 773362
rect 41696 773298 41748 773304
rect 35808 773152 35860 773158
rect 35806 773120 35808 773129
rect 40776 773152 40828 773158
rect 35860 773120 35862 773129
rect 35806 773055 35862 773064
rect 40774 773120 40776 773129
rect 40828 773120 40830 773129
rect 40774 773055 40830 773064
rect 35532 773016 35584 773022
rect 35532 772958 35584 772964
rect 41696 773016 41748 773022
rect 42064 773016 42116 773022
rect 41748 772964 42064 772970
rect 41696 772958 42116 772964
rect 41708 772942 42104 772958
rect 35348 772880 35400 772886
rect 35348 772822 35400 772828
rect 41696 772744 41748 772750
rect 42064 772744 42116 772750
rect 41748 772692 42064 772698
rect 41696 772686 42116 772692
rect 41708 772670 42104 772686
rect 35806 772304 35862 772313
rect 35806 772239 35862 772248
rect 35622 771896 35678 771905
rect 35820 771866 35848 772239
rect 42812 771905 42840 779686
rect 42982 773120 43038 773129
rect 42982 773055 43038 773064
rect 40222 771896 40278 771905
rect 35622 771831 35678 771840
rect 35808 771860 35860 771866
rect 35636 771594 35664 771831
rect 40222 771831 40224 771840
rect 35808 771802 35860 771808
rect 40276 771831 40278 771840
rect 42798 771896 42854 771905
rect 42798 771831 42854 771840
rect 40224 771802 40276 771808
rect 41052 771656 41104 771662
rect 41052 771598 41104 771604
rect 35624 771588 35676 771594
rect 35624 771530 35676 771536
rect 41064 771497 41092 771598
rect 35806 771488 35862 771497
rect 35806 771423 35808 771432
rect 35860 771423 35862 771432
rect 41050 771488 41106 771497
rect 41708 771458 42104 771474
rect 41050 771423 41106 771432
rect 41696 771452 42116 771458
rect 35808 771394 35860 771400
rect 41748 771446 42064 771452
rect 41696 771394 41748 771400
rect 42064 771394 42116 771400
rect 35806 771080 35862 771089
rect 35806 771015 35862 771024
rect 41510 771080 41566 771089
rect 41510 771015 41566 771024
rect 35622 770672 35678 770681
rect 35622 770607 35678 770616
rect 35636 770234 35664 770607
rect 35820 770506 35848 771015
rect 35808 770500 35860 770506
rect 35808 770442 35860 770448
rect 39856 770500 39908 770506
rect 39856 770442 39908 770448
rect 39868 770273 39896 770442
rect 35806 770264 35862 770273
rect 35624 770228 35676 770234
rect 35806 770199 35862 770208
rect 39854 770264 39910 770273
rect 41524 770234 41552 771015
rect 39854 770199 39910 770208
rect 41512 770228 41564 770234
rect 35624 770170 35676 770176
rect 35820 770098 35848 770199
rect 41512 770170 41564 770176
rect 41708 770098 42104 770114
rect 35808 770092 35860 770098
rect 35808 770034 35860 770040
rect 41696 770092 42116 770098
rect 41748 770086 42064 770092
rect 41696 770034 41748 770040
rect 42064 770034 42116 770040
rect 35806 769448 35862 769457
rect 35806 769383 35862 769392
rect 35820 769214 35848 769383
rect 35808 769208 35860 769214
rect 35808 769150 35860 769156
rect 35530 769040 35586 769049
rect 35530 768975 35586 768984
rect 35806 769040 35862 769049
rect 35806 768975 35862 768984
rect 41696 769004 41748 769010
rect 35544 768874 35572 768975
rect 35532 768868 35584 768874
rect 35532 768810 35584 768816
rect 35820 768738 35848 768975
rect 41696 768946 41748 768952
rect 41236 768868 41288 768874
rect 41236 768810 41288 768816
rect 35808 768732 35860 768738
rect 35808 768674 35860 768680
rect 40040 768732 40092 768738
rect 40040 768674 40092 768680
rect 35162 768224 35218 768233
rect 35162 768159 35218 768168
rect 32402 767816 32458 767825
rect 32402 767751 32458 767760
rect 32416 759694 32444 767751
rect 33782 767000 33838 767009
rect 33782 766935 33838 766944
rect 32404 759688 32456 759694
rect 32404 759630 32456 759636
rect 33796 758334 33824 766935
rect 35176 759830 35204 768159
rect 35806 767408 35862 767417
rect 35806 767343 35808 767352
rect 35860 767343 35862 767352
rect 36544 767372 36596 767378
rect 35808 767314 35860 767320
rect 36544 767314 36596 767320
rect 35806 766592 35862 766601
rect 35806 766527 35862 766536
rect 35820 766086 35848 766527
rect 35808 766080 35860 766086
rect 35808 766022 35860 766028
rect 35806 765776 35862 765785
rect 35806 765711 35862 765720
rect 35820 764862 35848 765711
rect 35808 764856 35860 764862
rect 35808 764798 35860 764804
rect 35808 764584 35860 764590
rect 35806 764552 35808 764561
rect 35860 764552 35862 764561
rect 35806 764487 35862 764496
rect 35622 764144 35678 764153
rect 35622 764079 35678 764088
rect 35636 763502 35664 764079
rect 35806 763736 35862 763745
rect 35806 763671 35862 763680
rect 35624 763496 35676 763502
rect 35624 763438 35676 763444
rect 35820 763230 35848 763671
rect 35808 763224 35860 763230
rect 35808 763166 35860 763172
rect 35806 762920 35862 762929
rect 35806 762855 35862 762864
rect 35820 761870 35848 762855
rect 35808 761864 35860 761870
rect 35808 761806 35860 761812
rect 35164 759824 35216 759830
rect 35164 759766 35216 759772
rect 33784 758328 33836 758334
rect 33784 758270 33836 758276
rect 36556 757761 36584 767314
rect 39764 766080 39816 766086
rect 39764 766022 39816 766028
rect 39776 765785 39804 766022
rect 39762 765776 39818 765785
rect 39762 765711 39818 765720
rect 40052 765338 40080 768674
rect 41248 767417 41276 768810
rect 41234 767408 41290 767417
rect 41234 767343 41290 767352
rect 41708 765914 41736 768946
rect 41708 765886 42288 765914
rect 40040 765332 40092 765338
rect 40040 765274 40092 765280
rect 41696 765332 41748 765338
rect 41696 765274 41748 765280
rect 41708 765218 41736 765274
rect 41708 765202 42104 765218
rect 41708 765196 42116 765202
rect 41708 765190 42064 765196
rect 42064 765138 42116 765144
rect 39396 764856 39448 764862
rect 39396 764798 39448 764804
rect 39408 764561 39436 764798
rect 41696 764652 41748 764658
rect 41696 764594 41748 764600
rect 39394 764552 39450 764561
rect 39394 764487 39450 764496
rect 41708 763745 41736 764594
rect 41694 763736 41750 763745
rect 41694 763671 41750 763680
rect 40960 763496 41012 763502
rect 40960 763438 41012 763444
rect 40972 763337 41000 763438
rect 40958 763328 41014 763337
rect 40958 763263 41014 763272
rect 41696 763156 41748 763162
rect 41696 763098 41748 763104
rect 41708 762929 41736 763098
rect 41694 762920 41750 762929
rect 41694 762855 41750 762864
rect 42064 761932 42116 761938
rect 42064 761874 42116 761880
rect 41696 761864 41748 761870
rect 42076 761818 42104 761874
rect 41748 761812 42104 761818
rect 41696 761806 42104 761812
rect 41708 761790 42104 761806
rect 41696 759824 41748 759830
rect 41748 759784 42104 759812
rect 41696 759766 41748 759772
rect 41604 759688 41656 759694
rect 41656 759636 41828 759642
rect 41604 759630 41828 759636
rect 41616 759614 41828 759630
rect 39212 758328 39264 758334
rect 39212 758270 39264 758276
rect 36542 757752 36598 757761
rect 36542 757687 36598 757696
rect 39224 757353 39252 758270
rect 39210 757344 39266 757353
rect 39210 757279 39266 757288
rect 41800 757081 41828 759614
rect 42076 759558 42104 759784
rect 42064 759552 42116 759558
rect 42064 759494 42116 759500
rect 41786 757072 41842 757081
rect 41786 757007 41842 757016
rect 41878 756664 41934 756673
rect 41878 756599 41934 756608
rect 41892 756226 41920 756599
rect 42260 756090 42288 765886
rect 42524 765196 42576 765202
rect 42524 765138 42576 765144
rect 42536 763154 42564 765138
rect 42536 763126 42840 763154
rect 42432 763088 42484 763094
rect 42432 763030 42484 763036
rect 42444 762929 42472 763030
rect 42430 762920 42486 762929
rect 42430 762855 42486 762864
rect 42432 759552 42484 759558
rect 42484 759500 42564 759506
rect 42432 759494 42564 759500
rect 42444 759478 42564 759494
rect 42248 756084 42300 756090
rect 42248 756026 42300 756032
rect 42338 755848 42394 755857
rect 42338 755783 42394 755792
rect 42352 755562 42380 755783
rect 42352 755534 42472 755562
rect 42248 755472 42300 755478
rect 42248 755414 42300 755420
rect 42260 754406 42288 755414
rect 42182 754378 42288 754406
rect 42062 754080 42118 754089
rect 42062 754015 42118 754024
rect 42076 753780 42104 754015
rect 42154 752992 42210 753001
rect 42154 752927 42210 752936
rect 42168 752556 42196 752927
rect 42076 751777 42104 751944
rect 42062 751768 42118 751777
rect 42062 751703 42118 751712
rect 42168 751233 42196 751369
rect 42154 751224 42210 751233
rect 42154 751159 42210 751168
rect 42154 750952 42210 750961
rect 42154 750887 42210 750896
rect 42168 750720 42196 750887
rect 42444 750122 42472 755534
rect 42168 749986 42196 750108
rect 42260 750094 42472 750122
rect 42260 749986 42288 750094
rect 42168 749958 42288 749986
rect 42536 749578 42564 759478
rect 42812 755154 42840 763126
rect 42444 749550 42564 749578
rect 42628 755126 42840 755154
rect 42444 749543 42472 749550
rect 42182 749515 42472 749543
rect 42062 749184 42118 749193
rect 42118 749142 42288 749170
rect 42062 749119 42118 749128
rect 42260 747062 42288 749142
rect 42182 747034 42288 747062
rect 41786 746872 41842 746881
rect 41786 746807 41842 746816
rect 41800 746401 41828 746807
rect 42628 746415 42656 755126
rect 42798 755032 42854 755041
rect 42798 754967 42854 754976
rect 42812 753494 42840 754967
rect 42260 746387 42656 746415
rect 42720 753466 42840 753494
rect 42062 746056 42118 746065
rect 42062 745991 42118 746000
rect 42076 745756 42104 745991
rect 42260 745634 42288 746387
rect 42720 746065 42748 753466
rect 42706 746056 42762 746065
rect 42706 745991 42762 746000
rect 42168 745606 42288 745634
rect 42168 745212 42196 745606
rect 42430 745376 42486 745385
rect 42430 745311 42486 745320
rect 42246 744832 42302 744841
rect 42246 744767 42302 744776
rect 42260 743730 42288 744767
rect 42168 743702 42288 743730
rect 42168 743376 42196 743702
rect 42168 742750 42288 742778
rect 42168 742696 42196 742750
rect 42260 742710 42288 742750
rect 42444 742710 42472 745311
rect 42614 745104 42670 745113
rect 42614 745039 42670 745048
rect 42260 742682 42472 742710
rect 42628 742098 42656 745039
rect 42800 744116 42852 744122
rect 42800 744058 42852 744064
rect 42812 744002 42840 744058
rect 42182 742070 42656 742098
rect 42720 743974 42840 744002
rect 42720 741690 42748 743974
rect 42536 741662 42748 741690
rect 42536 741554 42564 741662
rect 42182 741526 42564 741554
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 42246 730552 42302 730561
rect 42246 730487 42302 730496
rect 40958 729736 41014 729745
rect 40958 729671 41014 729680
rect 40972 728822 41000 729671
rect 42260 729366 42288 730487
rect 42996 730153 43024 773055
rect 43180 773022 43208 785206
rect 43168 773016 43220 773022
rect 43168 772958 43220 772964
rect 43442 771488 43498 771497
rect 43442 771423 43498 771432
rect 43258 763328 43314 763337
rect 43258 763263 43314 763272
rect 42982 730144 43038 730153
rect 42982 730079 43038 730088
rect 42248 729360 42300 729366
rect 41142 729328 41198 729337
rect 42248 729302 42300 729308
rect 41142 729263 41198 729272
rect 40960 728816 41012 728822
rect 40960 728758 41012 728764
rect 40866 728682 40922 728691
rect 41156 728686 41184 729263
rect 42890 728920 42946 728929
rect 41708 728890 42104 728906
rect 41696 728884 42116 728890
rect 41748 728878 42064 728884
rect 41696 728826 41748 728832
rect 42890 728855 42946 728864
rect 43076 728884 43128 728890
rect 42064 728826 42116 728832
rect 40866 728617 40922 728626
rect 41144 728680 41196 728686
rect 41144 728622 41196 728628
rect 41696 728680 41748 728686
rect 42064 728680 42116 728686
rect 41748 728640 42064 728668
rect 41696 728622 41748 728628
rect 42064 728622 42116 728628
rect 40880 727462 40908 728617
rect 40868 727456 40920 727462
rect 40868 727398 40920 727404
rect 41326 727458 41382 727467
rect 41326 727393 41382 727402
rect 41696 727456 41748 727462
rect 42064 727456 42116 727462
rect 41748 727416 42064 727444
rect 41696 727398 41748 727404
rect 42064 727398 42116 727404
rect 41340 727326 41368 727393
rect 41328 727320 41380 727326
rect 41328 727262 41380 727268
rect 41696 727320 41748 727326
rect 42064 727320 42116 727326
rect 41748 727280 42064 727308
rect 41696 727262 41748 727268
rect 42064 727262 42116 727268
rect 41142 726880 41198 726889
rect 41142 726815 41198 726824
rect 40958 726234 41014 726243
rect 40958 726169 41014 726178
rect 40774 725656 40830 725665
rect 40774 725591 40830 725600
rect 32402 725248 32458 725257
rect 32402 725183 32458 725192
rect 31666 724024 31722 724033
rect 31666 723959 31722 723968
rect 31680 715494 31708 723959
rect 32416 716854 32444 725183
rect 35162 724840 35218 724849
rect 35162 724775 35218 724784
rect 32404 716848 32456 716854
rect 32404 716790 32456 716796
rect 35176 715698 35204 724775
rect 37278 724432 37334 724441
rect 37278 724367 37334 724376
rect 37292 716961 37320 724367
rect 39302 723208 39358 723217
rect 39302 723143 39358 723152
rect 37278 716952 37334 716961
rect 37278 716887 37334 716896
rect 35164 715692 35216 715698
rect 35164 715634 35216 715640
rect 31668 715488 31720 715494
rect 31668 715430 31720 715436
rect 38016 715488 38068 715494
rect 38016 715430 38068 715436
rect 38028 714513 38056 715430
rect 39316 714814 39344 723143
rect 40788 719273 40816 725591
rect 40972 723058 41000 726169
rect 41156 725966 41184 726815
rect 41326 726234 41382 726243
rect 41326 726169 41382 726178
rect 41696 726232 41748 726238
rect 41748 726180 42196 726186
rect 41696 726174 42196 726180
rect 41708 726158 42196 726174
rect 41144 725960 41196 725966
rect 41144 725902 41196 725908
rect 41604 725960 41656 725966
rect 41604 725902 41656 725908
rect 41616 725778 41644 725902
rect 41786 725792 41842 725801
rect 41616 725750 41786 725778
rect 41786 725727 41842 725736
rect 41786 723072 41842 723081
rect 40972 723030 41786 723058
rect 41786 723007 41842 723016
rect 41786 722392 41842 722401
rect 41786 722327 41842 722336
rect 40774 719264 40830 719273
rect 40774 719199 40830 719208
rect 41800 718593 41828 722327
rect 41970 721984 42026 721993
rect 41970 721919 42026 721928
rect 41786 718584 41842 718593
rect 41786 718519 41842 718528
rect 41984 718321 42012 721919
rect 41970 718312 42026 718321
rect 41970 718247 42026 718256
rect 41696 716848 41748 716854
rect 41748 716796 41920 716802
rect 41696 716790 41920 716796
rect 41708 716774 41920 716790
rect 40408 715692 40460 715698
rect 40408 715634 40460 715640
rect 40420 714921 40448 715634
rect 40406 714912 40462 714921
rect 40406 714847 40462 714856
rect 39304 714808 39356 714814
rect 39304 714750 39356 714756
rect 41604 714808 41656 714814
rect 41656 714756 41828 714762
rect 41604 714750 41828 714756
rect 41616 714734 41828 714750
rect 38014 714504 38070 714513
rect 38014 714439 38070 714448
rect 41800 713969 41828 714734
rect 41892 714082 41920 716774
rect 42168 716530 42196 726158
rect 42706 719264 42762 719273
rect 42706 719199 42762 719208
rect 42168 716502 42472 716530
rect 42154 714912 42210 714921
rect 42154 714847 42210 714856
rect 42168 714241 42196 714847
rect 42154 714232 42210 714241
rect 42154 714167 42210 714176
rect 41892 714066 42104 714082
rect 41892 714060 42116 714066
rect 41892 714054 42064 714060
rect 42064 714002 42116 714008
rect 41786 713960 41842 713969
rect 41786 713895 41842 713904
rect 42154 713552 42210 713561
rect 42154 713487 42210 713496
rect 42168 713048 42196 713487
rect 42444 713474 42472 716502
rect 42720 714877 42748 719199
rect 42706 714868 42762 714877
rect 42706 714803 42762 714812
rect 42616 714060 42668 714066
rect 42616 714002 42668 714008
rect 42628 713474 42656 714002
rect 42352 713446 42472 713474
rect 42536 713446 42656 713474
rect 42352 712314 42380 713446
rect 42260 712286 42380 712314
rect 42260 711226 42288 712286
rect 42536 712042 42564 713446
rect 42536 712014 42656 712042
rect 42182 711198 42288 711226
rect 42248 711136 42300 711142
rect 42248 711078 42300 711084
rect 42260 710575 42288 711078
rect 42628 710575 42656 712014
rect 42182 710547 42288 710575
rect 42536 710547 42656 710575
rect 42246 710424 42302 710433
rect 42246 710359 42302 710368
rect 42260 709390 42288 710359
rect 42182 709362 42288 709390
rect 42246 709200 42302 709209
rect 42246 709135 42302 709144
rect 42062 708928 42118 708937
rect 42062 708863 42118 708872
rect 42076 708696 42104 708863
rect 42062 708384 42118 708393
rect 42062 708319 42118 708328
rect 42076 708152 42104 708319
rect 41984 707441 42012 707540
rect 41970 707432 42026 707441
rect 42260 707418 42288 709135
rect 41970 707367 42026 707376
rect 42168 707390 42288 707418
rect 42168 706860 42196 707390
rect 42536 706330 42564 710547
rect 42706 710016 42762 710025
rect 42706 709951 42762 709960
rect 42182 706302 42564 706330
rect 42430 706208 42486 706217
rect 42486 706166 42656 706194
rect 42430 706143 42486 706152
rect 42432 705560 42484 705566
rect 42432 705502 42484 705508
rect 41970 704304 42026 704313
rect 41970 704239 42026 704248
rect 41984 703868 42012 704239
rect 42444 703202 42472 705502
rect 42182 703174 42472 703202
rect 42628 702658 42656 706166
rect 42352 702630 42656 702658
rect 42352 702590 42380 702630
rect 42168 702522 42196 702576
rect 42260 702562 42380 702590
rect 42260 702522 42288 702562
rect 42168 702494 42288 702522
rect 42720 702250 42748 709951
rect 42904 706194 42932 728855
rect 43076 728826 43128 728832
rect 43088 714854 43116 728826
rect 43088 714826 43208 714854
rect 42812 706166 42932 706194
rect 42812 705922 42840 706166
rect 42812 705894 42932 705922
rect 41984 702222 42748 702250
rect 41984 702032 42012 702222
rect 42246 701856 42302 701865
rect 42246 701791 42302 701800
rect 41786 700496 41842 700505
rect 41786 700431 41842 700440
rect 41800 700165 41828 700431
rect 42260 699938 42288 701791
rect 42522 701584 42578 701593
rect 42522 701519 42578 701528
rect 42168 699910 42288 699938
rect 42168 699516 42196 699910
rect 42536 699242 42564 701519
rect 42708 701072 42760 701078
rect 42708 701014 42760 701020
rect 42064 699236 42116 699242
rect 42064 699178 42116 699184
rect 42524 699236 42576 699242
rect 42524 699178 42576 699184
rect 42076 698904 42104 699178
rect 42720 698339 42748 701014
rect 42182 698311 42748 698339
rect 42904 698294 42932 705894
rect 43180 705194 43208 714826
rect 42812 698266 42932 698294
rect 43088 705166 43208 705194
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 41142 686896 41198 686905
rect 41142 686831 41198 686840
rect 40958 686488 41014 686497
rect 40958 686423 41014 686432
rect 40774 685910 40830 685919
rect 40972 685914 41000 686423
rect 41156 686118 41184 686831
rect 42812 686322 42840 698266
rect 41328 686316 41380 686322
rect 41328 686258 41380 686264
rect 41696 686316 41748 686322
rect 42064 686316 42116 686322
rect 41748 686276 42064 686304
rect 41696 686258 41748 686264
rect 42064 686258 42116 686264
rect 42800 686316 42852 686322
rect 42800 686258 42852 686264
rect 41144 686112 41196 686118
rect 41144 686054 41196 686060
rect 41340 685919 41368 686258
rect 43088 686118 43116 705166
rect 41696 686112 41748 686118
rect 42064 686112 42116 686118
rect 41748 686072 42064 686100
rect 41696 686054 41748 686060
rect 42064 686054 42116 686060
rect 43076 686112 43128 686118
rect 43076 686054 43128 686060
rect 40774 685845 40830 685854
rect 40960 685908 41012 685914
rect 40960 685850 41012 685856
rect 41326 685910 41382 685919
rect 41326 685845 41382 685854
rect 41696 685908 41748 685914
rect 42064 685908 42116 685914
rect 41748 685868 42064 685896
rect 41696 685850 41748 685856
rect 42064 685850 42116 685856
rect 35162 682000 35218 682009
rect 35162 681935 35218 681944
rect 33046 681592 33102 681601
rect 33046 681527 33102 681536
rect 33060 674150 33088 681527
rect 33782 681184 33838 681193
rect 33782 681119 33838 681128
rect 33048 674144 33100 674150
rect 33048 674086 33100 674092
rect 33796 672761 33824 681119
rect 35176 672790 35204 681935
rect 36542 680776 36598 680785
rect 36542 680711 36598 680720
rect 35164 672784 35216 672790
rect 33782 672752 33838 672761
rect 35164 672726 35216 672732
rect 33782 672687 33838 672696
rect 36556 671022 36584 680711
rect 40788 678638 40816 685845
rect 42982 684176 43038 684185
rect 42982 684111 43038 684120
rect 41326 683462 41382 683471
rect 41326 683397 41382 683406
rect 41696 683460 41748 683466
rect 41696 683402 41748 683408
rect 40958 682816 41014 682825
rect 40958 682751 41014 682760
rect 40972 678974 41000 682751
rect 41708 678974 41736 683402
rect 42614 682408 42670 682417
rect 42614 682343 42670 682352
rect 40972 678946 41368 678974
rect 41708 678946 42288 678974
rect 41340 678858 41368 678946
rect 41786 678872 41842 678881
rect 41340 678830 41786 678858
rect 41786 678807 41842 678816
rect 40776 678632 40828 678638
rect 41696 678632 41748 678638
rect 40776 678574 40828 678580
rect 41694 678600 41696 678609
rect 41748 678600 41750 678609
rect 41694 678535 41750 678544
rect 41786 678328 41842 678337
rect 41616 678286 41786 678314
rect 40774 677750 40830 677759
rect 41616 677754 41644 678286
rect 41786 678263 41842 678272
rect 40774 677685 40830 677694
rect 41604 677748 41656 677754
rect 41604 677690 41656 677696
rect 41420 674144 41472 674150
rect 41420 674086 41472 674092
rect 36544 671016 36596 671022
rect 40500 671016 40552 671022
rect 36544 670958 36596 670964
rect 40498 670984 40500 670993
rect 41432 670993 41460 674086
rect 41604 672784 41656 672790
rect 41604 672726 41656 672732
rect 41616 671129 41644 672726
rect 41602 671120 41658 671129
rect 41602 671055 41658 671064
rect 40552 670984 40554 670993
rect 40498 670919 40554 670928
rect 41418 670984 41474 670993
rect 41418 670919 41474 670928
rect 41786 670304 41842 670313
rect 41786 670239 41842 670248
rect 41800 669868 41828 670239
rect 42168 667978 42196 668032
rect 42260 667978 42288 678946
rect 42430 677104 42486 677113
rect 42430 677039 42486 677048
rect 42444 676258 42472 677039
rect 42432 676252 42484 676258
rect 42432 676194 42484 676200
rect 42628 671362 42656 682343
rect 42798 679960 42854 679969
rect 42798 679895 42854 679904
rect 42812 671537 42840 679895
rect 42798 671528 42854 671537
rect 42798 671463 42854 671472
rect 42616 671356 42668 671362
rect 42616 671298 42668 671304
rect 42616 671220 42668 671226
rect 42616 671162 42668 671168
rect 42432 669384 42484 669390
rect 42432 669326 42484 669332
rect 42168 667950 42288 667978
rect 42444 667706 42472 669326
rect 42628 669314 42656 671162
rect 42798 671120 42854 671129
rect 42798 671055 42854 671064
rect 42812 670834 42840 671055
rect 42812 670806 42932 670834
rect 42628 669286 42748 669314
rect 42168 667678 42472 667706
rect 42168 667352 42196 667678
rect 42338 667448 42394 667457
rect 42338 667383 42394 667392
rect 42154 666632 42210 666641
rect 42154 666567 42210 666576
rect 42168 666165 42196 666567
rect 42352 666554 42380 667383
rect 42720 666554 42748 669286
rect 42352 666526 42472 666554
rect 42248 665848 42300 665854
rect 42248 665790 42300 665796
rect 42260 665530 42288 665790
rect 42182 665502 42288 665530
rect 42062 665408 42118 665417
rect 42118 665366 42288 665394
rect 42062 665343 42118 665352
rect 41786 665136 41842 665145
rect 41786 665071 41842 665080
rect 41800 664972 41828 665071
rect 42062 664592 42118 664601
rect 42062 664527 42118 664536
rect 42076 664325 42104 664527
rect 42260 663694 42288 665366
rect 42444 663762 42472 666526
rect 42536 666526 42748 666554
rect 42536 663898 42564 666526
rect 42536 663870 42656 663898
rect 42628 663814 42656 663870
rect 42182 663666 42288 663694
rect 42352 663734 42472 663762
rect 42616 663808 42668 663814
rect 42616 663750 42668 663756
rect 42352 663626 42380 663734
rect 42352 663598 42472 663626
rect 42248 663468 42300 663474
rect 42248 663410 42300 663416
rect 42260 663150 42288 663410
rect 42182 663122 42288 663150
rect 42248 663060 42300 663066
rect 42248 663002 42300 663008
rect 42260 660770 42288 663002
rect 42168 660742 42288 660770
rect 42168 660620 42196 660742
rect 42156 660544 42208 660550
rect 42156 660486 42208 660492
rect 42168 660008 42196 660486
rect 42444 659371 42472 663598
rect 42616 663604 42668 663610
rect 42616 663546 42668 663552
rect 42182 659343 42472 659371
rect 42628 659054 42656 663546
rect 42904 663490 42932 670806
rect 42812 663474 42932 663490
rect 42800 663468 42932 663474
rect 42852 663462 42932 663468
rect 42800 663410 42852 663416
rect 42156 659048 42208 659054
rect 42156 658990 42208 658996
rect 42616 659048 42668 659054
rect 42616 658990 42668 658996
rect 42168 658784 42196 658990
rect 42522 658608 42578 658617
rect 42352 658566 42522 658594
rect 41800 658430 42288 658458
rect 41800 658345 41828 658430
rect 41786 658336 41842 658345
rect 41786 658271 41842 658280
rect 41786 657248 41842 657257
rect 41786 657183 41842 657192
rect 41800 656948 41828 657183
rect 42260 656350 42288 658430
rect 42182 656322 42288 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42352 655670 42380 658566
rect 42522 658543 42578 658552
rect 42524 657552 42576 657558
rect 42524 657494 42576 657500
rect 42260 655642 42380 655670
rect 42536 655126 42564 657494
rect 42182 655098 42564 655126
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 35820 644502 35848 644671
rect 35808 644496 35860 644502
rect 35808 644438 35860 644444
rect 40132 644496 40184 644502
rect 40132 644438 40184 644444
rect 38566 644328 38622 644337
rect 38566 644263 38622 644272
rect 35346 643920 35402 643929
rect 35346 643855 35402 643864
rect 35360 643142 35388 643855
rect 35808 643544 35860 643550
rect 35530 643512 35586 643521
rect 35530 643447 35586 643456
rect 35806 643512 35808 643521
rect 35860 643512 35862 643521
rect 35806 643447 35862 643456
rect 35544 643278 35572 643447
rect 35532 643272 35584 643278
rect 35532 643214 35584 643220
rect 35348 643136 35400 643142
rect 35348 643078 35400 643084
rect 35438 642696 35494 642705
rect 35438 642631 35494 642640
rect 35806 642696 35862 642705
rect 35806 642631 35862 642640
rect 35452 641918 35480 642631
rect 35622 642288 35678 642297
rect 35622 642223 35678 642232
rect 35440 641912 35492 641918
rect 35440 641854 35492 641860
rect 35636 641782 35664 642223
rect 35820 642190 35848 642631
rect 38580 642530 38608 644263
rect 38568 642524 38620 642530
rect 38568 642466 38620 642472
rect 39946 642288 40002 642297
rect 39946 642223 40002 642232
rect 35808 642184 35860 642190
rect 35808 642126 35860 642132
rect 39960 641918 39988 642223
rect 39948 641912 40000 641918
rect 39948 641854 40000 641860
rect 35624 641776 35676 641782
rect 35624 641718 35676 641724
rect 40144 641481 40172 644438
rect 40592 643544 40644 643550
rect 40592 643486 40644 643492
rect 40316 642184 40368 642190
rect 40316 642126 40368 642132
rect 35346 641472 35402 641481
rect 35346 641407 35402 641416
rect 40130 641472 40186 641481
rect 40130 641407 40186 641416
rect 35360 640354 35388 641407
rect 35530 641064 35586 641073
rect 35530 640999 35586 641008
rect 35806 641064 35862 641073
rect 35806 640999 35862 641008
rect 35544 640490 35572 640999
rect 35820 640762 35848 640999
rect 35808 640756 35860 640762
rect 35808 640698 35860 640704
rect 39948 640756 40000 640762
rect 39948 640698 40000 640704
rect 35532 640484 35584 640490
rect 35532 640426 35584 640432
rect 35348 640348 35400 640354
rect 35348 640290 35400 640296
rect 39960 640257 39988 640698
rect 39946 640248 40002 640257
rect 39946 640183 40002 640192
rect 40328 639849 40356 642126
rect 40604 641073 40632 643486
rect 41708 643346 42104 643362
rect 41696 643340 42116 643346
rect 41748 643334 42064 643340
rect 41696 643282 41748 643288
rect 42064 643282 42116 643288
rect 41696 643136 41748 643142
rect 42064 643136 42116 643142
rect 41748 643084 42064 643090
rect 41696 643078 42116 643084
rect 41708 643062 42104 643078
rect 41696 642524 41748 642530
rect 41748 642484 42104 642512
rect 41696 642466 41748 642472
rect 42076 642394 42104 642484
rect 42064 642388 42116 642394
rect 42064 642330 42116 642336
rect 41696 641776 41748 641782
rect 42064 641776 42116 641782
rect 41748 641724 42064 641730
rect 41696 641718 42116 641724
rect 41708 641702 42104 641718
rect 40590 641064 40646 641073
rect 40590 640999 40646 641008
rect 42996 640558 43024 684111
rect 42064 640552 42116 640558
rect 41708 640500 42064 640506
rect 41708 640494 42116 640500
rect 42984 640552 43036 640558
rect 42984 640494 43036 640500
rect 41708 640490 42104 640494
rect 41696 640484 42104 640490
rect 41748 640478 42104 640484
rect 41696 640426 41748 640432
rect 41696 640348 41748 640354
rect 42064 640348 42116 640354
rect 41748 640306 42064 640334
rect 41696 640290 41748 640296
rect 42064 640290 42116 640296
rect 34426 639840 34482 639849
rect 34426 639775 34482 639784
rect 40314 639840 40370 639849
rect 40314 639775 40370 639784
rect 34440 638246 34468 639775
rect 35806 639432 35862 639441
rect 35806 639367 35862 639376
rect 35820 639198 35848 639367
rect 35808 639192 35860 639198
rect 35808 639134 35860 639140
rect 39304 639124 39356 639130
rect 39304 639066 39356 639072
rect 35806 639024 35862 639033
rect 35806 638959 35808 638968
rect 35860 638959 35862 638968
rect 35808 638930 35860 638936
rect 35622 638616 35678 638625
rect 35622 638551 35678 638560
rect 34428 638240 34480 638246
rect 34428 638182 34480 638188
rect 32402 637800 32458 637809
rect 32402 637735 32458 637744
rect 32416 629921 32444 637735
rect 35162 637392 35218 637401
rect 35162 637327 35218 637336
rect 32402 629912 32458 629921
rect 32402 629847 32458 629856
rect 35176 628590 35204 637327
rect 35636 636886 35664 638551
rect 35806 638208 35862 638217
rect 35806 638143 35862 638152
rect 35820 637634 35848 638143
rect 35808 637628 35860 637634
rect 35808 637570 35860 637576
rect 36544 637628 36596 637634
rect 36544 637570 36596 637576
rect 35806 636984 35862 636993
rect 35806 636919 35862 636928
rect 35624 636880 35676 636886
rect 35624 636822 35676 636828
rect 35820 636750 35848 636919
rect 35808 636744 35860 636750
rect 35808 636686 35860 636692
rect 35530 636576 35586 636585
rect 35530 636511 35586 636520
rect 35806 636576 35862 636585
rect 35806 636511 35862 636520
rect 35544 636274 35572 636511
rect 35820 636410 35848 636511
rect 35808 636404 35860 636410
rect 35808 636346 35860 636352
rect 35532 636268 35584 636274
rect 35532 636210 35584 636216
rect 35806 635760 35862 635769
rect 35806 635695 35862 635704
rect 35820 634846 35848 635695
rect 35808 634840 35860 634846
rect 35808 634782 35860 634788
rect 35806 634536 35862 634545
rect 35806 634471 35862 634480
rect 35820 633894 35848 634471
rect 35808 633888 35860 633894
rect 35808 633830 35860 633836
rect 35806 633720 35862 633729
rect 35806 633655 35862 633664
rect 35820 633486 35848 633655
rect 35808 633480 35860 633486
rect 35808 633422 35860 633428
rect 36556 630630 36584 637570
rect 39120 636200 39172 636206
rect 39118 636168 39120 636177
rect 39172 636168 39174 636177
rect 39118 636103 39174 636112
rect 36544 630624 36596 630630
rect 36544 630566 36596 630572
rect 39316 629241 39344 639066
rect 40040 638988 40092 638994
rect 40040 638930 40092 638936
rect 39764 633752 39816 633758
rect 39762 633720 39764 633729
rect 39816 633720 39818 633729
rect 39762 633655 39818 633664
rect 40052 630329 40080 638930
rect 41696 638240 41748 638246
rect 41696 638182 41748 638188
rect 40316 636880 40368 636886
rect 40316 636822 40368 636828
rect 40328 634545 40356 636822
rect 40868 636676 40920 636682
rect 40868 636618 40920 636624
rect 40500 636404 40552 636410
rect 40500 636346 40552 636352
rect 40512 635769 40540 636346
rect 40498 635760 40554 635769
rect 40498 635695 40554 635704
rect 40500 634840 40552 634846
rect 40500 634782 40552 634788
rect 40314 634536 40370 634545
rect 40314 634471 40370 634480
rect 40512 630601 40540 634782
rect 40880 632369 40908 636618
rect 41512 633480 41564 633486
rect 41512 633422 41564 633428
rect 41524 633321 41552 633422
rect 41510 633312 41566 633321
rect 41510 633247 41566 633256
rect 40866 632360 40922 632369
rect 40866 632295 40922 632304
rect 41708 630674 41736 638182
rect 42706 634536 42762 634545
rect 42706 634471 42762 634480
rect 42064 633480 42116 633486
rect 42064 633422 42116 633428
rect 42076 633321 42104 633422
rect 42062 633312 42118 633321
rect 42062 633247 42118 633256
rect 41708 630646 41920 630674
rect 40498 630592 40554 630601
rect 40498 630527 40554 630536
rect 41604 630556 41656 630562
rect 41604 630498 41656 630504
rect 41616 630442 41644 630498
rect 41616 630414 41828 630442
rect 40038 630320 40094 630329
rect 40038 630255 40094 630264
rect 39302 629232 39358 629241
rect 39302 629167 39358 629176
rect 35164 628584 35216 628590
rect 35164 628526 35216 628532
rect 40500 628584 40552 628590
rect 40500 628526 40552 628532
rect 40512 628425 40540 628526
rect 40498 628416 40554 628425
rect 40498 628351 40554 628360
rect 41800 627473 41828 630414
rect 41892 628266 41920 630646
rect 42522 630320 42578 630329
rect 42522 630255 42578 630264
rect 42338 628416 42394 628425
rect 42338 628351 42394 628360
rect 41892 628238 42288 628266
rect 41786 627464 41842 627473
rect 41786 627399 41842 627408
rect 41786 627192 41842 627201
rect 41786 627127 41842 627136
rect 41800 626620 41828 627127
rect 42260 625274 42288 628238
rect 42168 625246 42288 625274
rect 42168 624784 42196 625246
rect 42352 625002 42380 628351
rect 42352 624974 42472 625002
rect 42248 624708 42300 624714
rect 42248 624650 42300 624656
rect 42260 624186 42288 624650
rect 42182 624158 42288 624186
rect 42248 624096 42300 624102
rect 42248 624038 42300 624044
rect 42260 623098 42288 624038
rect 42168 623070 42288 623098
rect 42168 622948 42196 623070
rect 42182 622322 42288 622350
rect 41786 622024 41842 622033
rect 41786 621959 41842 621968
rect 41800 621792 41828 621959
rect 42260 621722 42288 622322
rect 42248 621716 42300 621722
rect 42248 621658 42300 621664
rect 42248 621580 42300 621586
rect 42248 621522 42300 621528
rect 42260 621126 42288 621522
rect 42182 621098 42288 621126
rect 41786 620800 41842 620809
rect 41786 620735 41842 620744
rect 41800 620500 41828 620735
rect 42248 620424 42300 620430
rect 42248 620366 42300 620372
rect 42260 620242 42288 620366
rect 42076 620214 42288 620242
rect 42076 619956 42104 620214
rect 42248 619676 42300 619682
rect 42248 619618 42300 619624
rect 42260 617454 42288 619618
rect 42182 617426 42288 617454
rect 42248 617364 42300 617370
rect 42248 617306 42300 617312
rect 42260 617250 42288 617306
rect 42076 617222 42288 617250
rect 42076 616828 42104 617222
rect 42444 616298 42472 624974
rect 42536 620242 42564 630255
rect 42720 620430 42748 634471
rect 43074 632360 43130 632369
rect 43074 632295 43130 632304
rect 42890 630592 42946 630601
rect 42890 630527 42946 630536
rect 42708 620424 42760 620430
rect 42708 620366 42760 620372
rect 42536 620214 42748 620242
rect 42168 616270 42472 616298
rect 42168 616148 42196 616270
rect 41878 616040 41934 616049
rect 41934 615998 42288 616026
rect 41878 615975 41934 615984
rect 42062 615904 42118 615913
rect 42062 615839 42118 615848
rect 42076 615604 42104 615839
rect 42260 614122 42288 615998
rect 42720 615913 42748 620214
rect 42904 619682 42932 630527
rect 42892 619676 42944 619682
rect 42892 619618 42944 619624
rect 43088 617370 43116 632295
rect 43076 617364 43128 617370
rect 43076 617306 43128 617312
rect 42706 615904 42762 615913
rect 42706 615839 42762 615848
rect 42614 615496 42670 615505
rect 42614 615431 42670 615440
rect 42628 615346 42656 615431
rect 42168 614094 42288 614122
rect 42536 615318 42656 615346
rect 42168 613768 42196 614094
rect 41878 613456 41934 613465
rect 41878 613391 41934 613400
rect 41892 613121 41920 613391
rect 42536 612490 42564 615318
rect 42708 614168 42760 614174
rect 42708 614110 42760 614116
rect 42182 612462 42564 612490
rect 42248 612400 42300 612406
rect 42246 612368 42248 612377
rect 42300 612368 42302 612377
rect 42246 612303 42302 612312
rect 42720 612082 42748 614110
rect 43272 612241 43300 763263
rect 43456 728686 43484 771423
rect 43628 754928 43680 754934
rect 43628 754870 43680 754876
rect 43640 753001 43668 754870
rect 43626 752992 43682 753001
rect 43626 752927 43682 752936
rect 43626 731368 43682 731377
rect 43626 731303 43682 731312
rect 43640 730318 43668 731303
rect 43628 730312 43680 730318
rect 43628 730254 43680 730260
rect 43444 728680 43496 728686
rect 43444 728622 43496 728628
rect 43442 723616 43498 723625
rect 43442 723551 43498 723560
rect 43456 705566 43484 723551
rect 43626 720352 43682 720361
rect 43626 720287 43682 720296
rect 43640 719030 43668 720287
rect 43628 719024 43680 719030
rect 43628 718966 43680 718972
rect 43628 709368 43680 709374
rect 43628 709310 43680 709316
rect 43640 707441 43668 709310
rect 43626 707432 43682 707441
rect 43626 707367 43682 707376
rect 43444 705560 43496 705566
rect 43444 705502 43496 705508
rect 43442 688120 43498 688129
rect 43442 688055 43498 688064
rect 43456 687546 43484 688055
rect 43444 687540 43496 687546
rect 43444 687482 43496 687488
rect 43442 687304 43498 687313
rect 43442 687239 43498 687248
rect 43456 686526 43484 687239
rect 43444 686520 43496 686526
rect 43444 686462 43496 686468
rect 43626 680368 43682 680377
rect 43626 680303 43682 680312
rect 43442 677920 43498 677929
rect 43442 677855 43498 677864
rect 43456 630674 43484 677855
rect 43640 660550 43668 680303
rect 43628 660544 43680 660550
rect 43628 660486 43680 660492
rect 43626 633720 43682 633729
rect 43626 633655 43682 633664
rect 43456 630646 43576 630674
rect 43258 612232 43314 612241
rect 43258 612167 43314 612176
rect 42536 612054 42748 612082
rect 42536 611946 42564 612054
rect 42182 611918 42564 611946
rect 43548 611266 43576 630646
rect 43640 612354 43668 633655
rect 43824 612678 43852 807463
rect 44192 771458 44220 814234
rect 44456 812864 44508 812870
rect 44456 812806 44508 812812
rect 44180 771452 44232 771458
rect 44180 771394 44232 771400
rect 44468 771089 44496 812806
rect 44640 807356 44692 807362
rect 44640 807298 44692 807304
rect 44652 796346 44680 807298
rect 44640 796340 44692 796346
rect 44640 796282 44692 796288
rect 44836 785194 44864 817090
rect 61384 817012 61436 817018
rect 61384 816954 61436 816960
rect 50344 806132 50396 806138
rect 50344 806074 50396 806080
rect 44824 785188 44876 785194
rect 44824 785130 44876 785136
rect 46202 773528 46258 773537
rect 46202 773463 46258 773472
rect 44454 771080 44510 771089
rect 44454 771015 44510 771024
rect 44270 770264 44326 770273
rect 44270 770199 44326 770208
rect 43996 753568 44048 753574
rect 43996 753510 44048 753516
rect 44008 751233 44036 753510
rect 43994 751224 44050 751233
rect 43994 751159 44050 751168
rect 44284 736934 44312 770199
rect 44548 770092 44600 770098
rect 44548 770034 44600 770040
rect 44284 736906 44404 736934
rect 44178 728104 44234 728113
rect 44178 728039 44234 728048
rect 44192 724514 44220 728039
rect 44376 727462 44404 736906
rect 44560 727705 44588 770034
rect 45006 765776 45062 765785
rect 45006 765711 45062 765720
rect 44732 755540 44784 755546
rect 44732 755482 44784 755488
rect 44744 754089 44772 755482
rect 45020 754934 45048 765711
rect 45190 764552 45246 764561
rect 45190 764487 45246 764496
rect 45008 754928 45060 754934
rect 45008 754870 45060 754876
rect 44730 754080 44786 754089
rect 44730 754015 44786 754024
rect 44822 751768 44878 751777
rect 44822 751703 44878 751712
rect 44836 746570 44864 751703
rect 45204 750961 45232 764487
rect 45374 763736 45430 763745
rect 45374 763671 45430 763680
rect 45388 753574 45416 763671
rect 45376 753568 45428 753574
rect 45376 753510 45428 753516
rect 45190 750952 45246 750961
rect 45190 750887 45246 750896
rect 44824 746564 44876 746570
rect 44824 746506 44876 746512
rect 46216 743782 46244 773463
rect 48964 761932 49016 761938
rect 48964 761874 49016 761880
rect 46204 743776 46256 743782
rect 46204 743718 46256 743724
rect 46202 730960 46258 730969
rect 46202 730895 46258 730904
rect 44546 727696 44602 727705
rect 44546 727631 44602 727640
rect 44364 727456 44416 727462
rect 44364 727398 44416 727404
rect 44640 727320 44692 727326
rect 44640 727262 44692 727268
rect 44192 724486 44404 724514
rect 44178 721576 44234 721585
rect 44178 721511 44234 721520
rect 44192 709050 44220 721511
rect 44008 709022 44220 709050
rect 44008 708393 44036 709022
rect 44178 708928 44234 708937
rect 44178 708863 44234 708872
rect 43994 708384 44050 708393
rect 43994 708319 44050 708328
rect 44192 703798 44220 708863
rect 44180 703792 44232 703798
rect 44180 703734 44232 703740
rect 44376 685273 44404 724486
rect 44362 685264 44418 685273
rect 44362 685199 44418 685208
rect 44362 684856 44418 684865
rect 44362 684791 44418 684800
rect 44178 679552 44234 679561
rect 44178 679487 44234 679496
rect 43994 679144 44050 679153
rect 43994 679079 44050 679088
rect 44008 663066 44036 679079
rect 44192 664601 44220 679487
rect 44178 664592 44234 664601
rect 44178 664527 44234 664536
rect 43996 663060 44048 663066
rect 43996 663002 44048 663008
rect 44376 641782 44404 684791
rect 44652 684457 44680 727262
rect 45282 722800 45338 722809
rect 45282 722735 45338 722744
rect 44914 721168 44970 721177
rect 44914 721103 44970 721112
rect 44638 684448 44694 684457
rect 44638 684383 44694 684392
rect 44548 667956 44600 667962
rect 44548 667898 44600 667904
rect 44560 665854 44588 667898
rect 44548 665848 44600 665854
rect 44548 665790 44600 665796
rect 44364 641776 44416 641782
rect 44364 641718 44416 641724
rect 44546 641064 44602 641073
rect 44546 640999 44602 641008
rect 44362 636168 44418 636177
rect 44362 636103 44418 636112
rect 43994 635760 44050 635769
rect 43994 635695 44050 635704
rect 44008 621586 44036 635695
rect 44180 625864 44232 625870
rect 44180 625806 44232 625812
rect 44192 624714 44220 625806
rect 44180 624708 44232 624714
rect 44180 624650 44232 624656
rect 44376 624102 44404 636103
rect 44364 624096 44416 624102
rect 44364 624038 44416 624044
rect 44180 621716 44232 621722
rect 44180 621658 44232 621664
rect 43996 621580 44048 621586
rect 43996 621522 44048 621528
rect 44192 616826 44220 621658
rect 44180 616820 44232 616826
rect 44180 616762 44232 616768
rect 43812 612672 43864 612678
rect 43812 612614 43864 612620
rect 43640 612326 44036 612354
rect 44008 612270 44036 612326
rect 43996 612264 44048 612270
rect 43873 612232 43929 612241
rect 43996 612206 44048 612212
rect 43873 612167 43929 612176
rect 43887 611998 43915 612167
rect 44088 612128 44140 612134
rect 44088 612070 44140 612076
rect 43875 611992 43927 611998
rect 43875 611934 43927 611940
rect 44100 611425 44128 612070
rect 44272 611720 44324 611726
rect 44270 611688 44272 611697
rect 44324 611688 44326 611697
rect 44270 611623 44326 611632
rect 44086 611416 44142 611425
rect 44086 611351 44142 611360
rect 43548 611238 44358 611266
rect 44330 611182 44358 611238
rect 44318 611176 44370 611182
rect 44318 611118 44370 611124
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 40314 602032 40370 602041
rect 40314 601967 40370 601976
rect 35806 601760 35862 601769
rect 35806 601695 35808 601704
rect 35860 601695 35862 601704
rect 36544 601724 36596 601730
rect 35808 601666 35860 601672
rect 36544 601666 36596 601672
rect 35162 595810 35218 595819
rect 35162 595745 35218 595754
rect 33046 595232 33102 595241
rect 33046 595167 33102 595176
rect 31022 594416 31078 594425
rect 31022 594351 31078 594360
rect 31036 585818 31064 594351
rect 33060 587178 33088 595167
rect 33782 593600 33838 593609
rect 33782 593535 33838 593544
rect 33048 587172 33100 587178
rect 33048 587114 33100 587120
rect 33796 585954 33824 593535
rect 35176 586158 35204 595745
rect 35622 591968 35678 591977
rect 35622 591903 35678 591912
rect 35636 590850 35664 591903
rect 35806 591560 35862 591569
rect 35806 591495 35862 591504
rect 35624 590844 35676 590850
rect 35624 590786 35676 590792
rect 35820 590714 35848 591495
rect 35808 590708 35860 590714
rect 35808 590650 35860 590656
rect 36556 589665 36584 601666
rect 39946 601352 40002 601361
rect 39946 601287 40002 601296
rect 37922 594824 37978 594833
rect 37922 594759 37978 594768
rect 36542 589656 36598 589665
rect 36542 589591 36598 589600
rect 35164 586152 35216 586158
rect 35164 586094 35216 586100
rect 33784 585948 33836 585954
rect 33784 585890 33836 585896
rect 31024 585812 31076 585818
rect 31024 585754 31076 585760
rect 37936 585177 37964 594759
rect 39960 594318 39988 601287
rect 40130 600944 40186 600953
rect 40130 600879 40186 600888
rect 40144 595814 40172 600879
rect 40132 595808 40184 595814
rect 40132 595750 40184 595756
rect 39948 594312 40000 594318
rect 39948 594254 40000 594260
rect 40328 592034 40356 601967
rect 44560 600545 44588 640999
rect 44732 612264 44784 612270
rect 44732 612206 44784 612212
rect 44744 610774 44772 612206
rect 44928 611590 44956 721103
rect 45296 709374 45324 722735
rect 45284 709368 45336 709374
rect 45284 709310 45336 709316
rect 46216 698290 46244 730895
rect 46204 698284 46256 698290
rect 46204 698226 46256 698232
rect 45466 687712 45522 687721
rect 45466 687647 45522 687656
rect 45100 685908 45152 685914
rect 45100 685850 45152 685856
rect 45112 643346 45140 685850
rect 45282 678600 45338 678609
rect 45282 678535 45338 678544
rect 45100 643340 45152 643346
rect 45100 643282 45152 643288
rect 45296 642297 45324 678535
rect 45480 655518 45508 687647
rect 45468 655512 45520 655518
rect 45468 655454 45520 655460
rect 45282 642288 45338 642297
rect 45282 642223 45338 642232
rect 46202 641472 46258 641481
rect 46202 641407 46258 641416
rect 45468 640348 45520 640354
rect 45468 640290 45520 640296
rect 45282 640248 45338 640257
rect 45282 640183 45338 640192
rect 45098 639840 45154 639849
rect 45098 639775 45154 639784
rect 44916 611584 44968 611590
rect 44916 611526 44968 611532
rect 44732 610768 44784 610774
rect 44732 610710 44784 610716
rect 44546 600536 44602 600545
rect 44546 600471 44602 600480
rect 44638 600128 44694 600137
rect 44638 600063 44694 600072
rect 43074 597680 43130 597689
rect 43074 597615 43130 597624
rect 43088 597446 43116 597615
rect 43076 597440 43128 597446
rect 43076 597382 43128 597388
rect 43076 597032 43128 597038
rect 42798 597000 42854 597009
rect 43076 596974 43128 596980
rect 42798 596935 42854 596944
rect 42430 596864 42486 596873
rect 42430 596799 42486 596808
rect 40958 596218 41014 596227
rect 40958 596153 41014 596162
rect 40972 592090 41000 596153
rect 41326 595810 41382 595819
rect 41696 595808 41748 595814
rect 41326 595745 41382 595754
rect 41694 595776 41696 595785
rect 41748 595776 41750 595785
rect 41340 594794 41368 595745
rect 41694 595711 41750 595720
rect 41328 594788 41380 594794
rect 41328 594730 41380 594736
rect 41696 594788 41748 594794
rect 41696 594730 41748 594736
rect 41708 594402 41736 594730
rect 41708 594374 42012 594402
rect 41604 594312 41656 594318
rect 41786 594280 41842 594289
rect 41656 594260 41786 594266
rect 41604 594254 41786 594260
rect 41616 594238 41786 594254
rect 41786 594215 41842 594224
rect 41694 592104 41750 592113
rect 40972 592062 41694 592090
rect 41694 592039 41750 592048
rect 41984 592034 42012 594374
rect 40328 592006 40448 592034
rect 41984 592006 42288 592034
rect 39672 590708 39724 590714
rect 39672 590650 39724 590656
rect 39684 589393 39712 590650
rect 39670 589384 39726 589393
rect 39670 589319 39726 589328
rect 39394 586120 39450 586129
rect 39394 586055 39396 586064
rect 39448 586055 39450 586064
rect 39396 586026 39448 586032
rect 39764 585948 39816 585954
rect 39764 585890 39816 585896
rect 39212 585812 39264 585818
rect 39212 585754 39264 585760
rect 37922 585168 37978 585177
rect 37922 585103 37978 585112
rect 39224 584905 39252 585754
rect 39210 584896 39266 584905
rect 39210 584831 39266 584840
rect 39776 584633 39804 585890
rect 40420 585721 40448 592006
rect 41696 590776 41748 590782
rect 41748 590724 42104 590730
rect 41696 590718 42104 590724
rect 41708 590714 42104 590718
rect 41708 590708 42116 590714
rect 41708 590702 42064 590708
rect 42064 590650 42116 590656
rect 41512 587172 41564 587178
rect 41512 587114 41564 587120
rect 40406 585712 40462 585721
rect 40406 585647 40462 585656
rect 41524 585290 41552 587114
rect 42260 586294 42288 592006
rect 42248 586288 42300 586294
rect 42248 586230 42300 586236
rect 41524 585262 42288 585290
rect 39762 584624 39818 584633
rect 39762 584559 39818 584568
rect 42260 583930 42288 585262
rect 42168 583902 42288 583930
rect 42168 583440 42196 583902
rect 42444 581618 42472 596799
rect 42812 592034 42840 596935
rect 42812 592006 42932 592034
rect 42616 586288 42668 586294
rect 42536 586236 42616 586242
rect 42536 586230 42668 586236
rect 42536 586214 42656 586230
rect 42536 585970 42564 586214
rect 42706 586120 42762 586129
rect 42706 586055 42762 586064
rect 42536 585942 42656 585970
rect 42182 581590 42472 581618
rect 42182 580947 42288 580975
rect 42260 580281 42288 580947
rect 41786 580272 41842 580281
rect 41786 580207 41842 580216
rect 42246 580272 42302 580281
rect 42246 580207 42302 580216
rect 41800 579768 41828 580207
rect 42430 580000 42486 580009
rect 42430 579935 42486 579944
rect 42444 579465 42472 579935
rect 42430 579456 42486 579465
rect 42430 579391 42486 579400
rect 42338 579184 42394 579193
rect 42182 579128 42338 579135
rect 42182 579119 42394 579128
rect 42182 579107 42380 579119
rect 42248 579012 42300 579018
rect 42248 578954 42300 578960
rect 42260 578626 42288 578954
rect 42168 578598 42288 578626
rect 42168 578544 42196 578598
rect 42338 578368 42394 578377
rect 42628 578354 42656 585942
rect 42394 578326 42656 578354
rect 42338 578303 42394 578312
rect 42062 578096 42118 578105
rect 42720 578082 42748 586055
rect 42904 582374 42932 592006
rect 42062 578031 42118 578040
rect 42352 578054 42748 578082
rect 42812 582346 42932 582374
rect 42076 577932 42104 578031
rect 41786 577824 41842 577833
rect 41786 577759 41842 577768
rect 41800 577281 41828 577759
rect 42352 576858 42380 578054
rect 42168 576830 42380 576858
rect 42168 576708 42196 576830
rect 41786 574696 41842 574705
rect 41786 574631 41842 574640
rect 41800 574260 41828 574631
rect 42614 574016 42670 574025
rect 42614 573951 42670 573960
rect 41800 573481 41828 573580
rect 41786 573472 41842 573481
rect 41786 573407 41842 573416
rect 42154 573472 42210 573481
rect 42154 573407 42210 573416
rect 42168 572968 42196 573407
rect 42062 572656 42118 572665
rect 42062 572591 42118 572600
rect 42076 572424 42104 572591
rect 42062 571568 42118 571577
rect 42062 571503 42118 571512
rect 42076 571282 42104 571503
rect 42430 571432 42486 571441
rect 42430 571367 42486 571376
rect 42076 571254 42380 571282
rect 42064 570988 42116 570994
rect 42064 570930 42116 570936
rect 42076 570588 42104 570930
rect 41786 570208 41842 570217
rect 41786 570143 41842 570152
rect 41800 569908 41828 570143
rect 42352 569310 42380 571254
rect 42168 569242 42196 569296
rect 42260 569282 42380 569310
rect 42260 569242 42288 569282
rect 42168 569214 42288 569242
rect 42444 568766 42472 571367
rect 42628 570994 42656 573951
rect 42616 570988 42668 570994
rect 42616 570930 42668 570936
rect 42168 568698 42196 568752
rect 42260 568738 42472 568766
rect 42260 568698 42288 568738
rect 42168 568670 42288 568698
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 40958 558104 41014 558113
rect 40958 558039 41014 558048
rect 37922 553408 37978 553417
rect 37922 553343 37978 553352
rect 29642 551984 29698 551993
rect 29642 551919 29698 551928
rect 29656 547194 29684 551919
rect 29644 547188 29696 547194
rect 29644 547130 29696 547136
rect 37936 542337 37964 553343
rect 40972 550458 41000 558039
rect 42812 555665 42840 582346
rect 42798 555656 42854 555665
rect 42798 555591 42854 555600
rect 43088 554849 43116 596974
rect 44362 593192 44418 593201
rect 44362 593127 44418 593136
rect 43260 590708 43312 590714
rect 43260 590650 43312 590656
rect 43272 579018 43300 590650
rect 43442 589384 43498 589393
rect 43442 589319 43498 589328
rect 43260 579012 43312 579018
rect 43260 578954 43312 578960
rect 43074 554840 43130 554849
rect 43074 554775 43130 554784
rect 43166 554432 43222 554441
rect 43166 554367 43222 554376
rect 41326 553408 41382 553417
rect 41156 553366 41326 553394
rect 40960 550452 41012 550458
rect 40960 550394 41012 550400
rect 40774 549944 40830 549953
rect 40774 549879 40830 549888
rect 40788 545601 40816 549879
rect 41156 545873 41184 553366
rect 41326 553343 41382 553352
rect 41326 552392 41382 552401
rect 41326 552327 41382 552336
rect 41340 552090 41368 552327
rect 41328 552084 41380 552090
rect 41328 552026 41380 552032
rect 41696 552084 41748 552090
rect 41696 552026 41748 552032
rect 41708 551857 41736 552026
rect 41694 551848 41750 551857
rect 41694 551783 41750 551792
rect 42982 551168 43038 551177
rect 42982 551103 43038 551112
rect 41708 550458 42012 550474
rect 41696 550452 42012 550458
rect 41748 550446 42012 550452
rect 41696 550394 41748 550400
rect 41984 550202 42012 550446
rect 42154 550216 42210 550225
rect 41984 550174 42154 550202
rect 42154 550151 42210 550160
rect 42798 549128 42854 549137
rect 42798 549063 42854 549072
rect 41326 548312 41382 548321
rect 41326 548247 41382 548256
rect 41340 547942 41368 548247
rect 41328 547936 41380 547942
rect 41328 547878 41380 547884
rect 41696 547936 41748 547942
rect 41696 547878 41748 547884
rect 41708 547777 41736 547878
rect 41694 547768 41750 547777
rect 41694 547703 41750 547712
rect 41696 547188 41748 547194
rect 41696 547130 41748 547136
rect 41142 545864 41198 545873
rect 41142 545799 41198 545808
rect 40774 545592 40830 545601
rect 40774 545527 40830 545536
rect 41708 543734 41736 547130
rect 42338 545864 42394 545873
rect 42338 545799 42394 545808
rect 41708 543706 42288 543734
rect 37922 542328 37978 542337
rect 37922 542263 37978 542272
rect 42260 540274 42288 543706
rect 42182 540246 42288 540274
rect 42352 538438 42380 545799
rect 42614 539608 42670 539617
rect 42614 539543 42670 539552
rect 42168 538370 42196 538424
rect 42260 538410 42380 538438
rect 42260 538370 42288 538410
rect 42168 538342 42288 538370
rect 42430 538248 42486 538257
rect 42430 538183 42486 538192
rect 42076 537441 42104 537744
rect 42062 537432 42118 537441
rect 42062 537367 42118 537376
rect 42062 537024 42118 537033
rect 42062 536959 42118 536968
rect 42076 536588 42104 536959
rect 42444 535922 42472 538183
rect 42628 537033 42656 539543
rect 42614 537024 42670 537033
rect 42614 536959 42670 536968
rect 42812 536874 42840 549063
rect 42996 540974 43024 551103
rect 42182 535894 42472 535922
rect 42536 536846 42840 536874
rect 42904 540946 43024 540974
rect 42062 535664 42118 535673
rect 42062 535599 42118 535608
rect 42076 535364 42104 535599
rect 41786 535256 41842 535265
rect 41786 535191 41842 535200
rect 41800 534752 41828 535191
rect 42536 534086 42564 536846
rect 42706 536752 42762 536761
rect 42706 536687 42762 536696
rect 42720 535673 42748 536687
rect 42706 535664 42762 535673
rect 42706 535599 42762 535608
rect 42182 534058 42564 534086
rect 42430 533896 42486 533905
rect 42430 533831 42486 533840
rect 42444 533542 42472 533831
rect 42182 533514 42472 533542
rect 42246 533352 42302 533361
rect 42246 533287 42302 533296
rect 42260 531059 42288 533287
rect 42706 532808 42762 532817
rect 42706 532743 42762 532752
rect 42430 531720 42486 531729
rect 42430 531655 42486 531664
rect 42182 531031 42288 531059
rect 42156 530732 42208 530738
rect 42156 530674 42208 530680
rect 42168 530400 42196 530674
rect 42248 530324 42300 530330
rect 42248 530266 42300 530272
rect 42260 529771 42288 530266
rect 42182 529743 42288 529771
rect 42444 529219 42472 531655
rect 42720 530942 42748 532743
rect 42708 530936 42760 530942
rect 42708 530878 42760 530884
rect 42614 530768 42670 530777
rect 42614 530703 42670 530712
rect 42182 529191 42472 529219
rect 42628 529122 42656 530703
rect 42904 530330 42932 540946
rect 42892 530324 42944 530330
rect 42892 530266 42944 530272
rect 42798 529816 42854 529825
rect 42260 529094 42656 529122
rect 42720 529760 42798 529771
rect 42720 529751 42854 529760
rect 42720 529743 42840 529751
rect 42260 527762 42288 529094
rect 42430 529000 42486 529009
rect 42430 528935 42486 528944
rect 42168 527734 42288 527762
rect 42168 527340 42196 527734
rect 42064 527060 42116 527066
rect 42064 527002 42116 527008
rect 42076 526728 42104 527002
rect 42444 526091 42472 528935
rect 42720 527066 42748 529743
rect 42708 527060 42760 527066
rect 42708 527002 42760 527008
rect 42614 526824 42670 526833
rect 42614 526759 42670 526768
rect 42182 526063 42472 526091
rect 42168 525558 42288 525586
rect 42168 525504 42196 525558
rect 42260 525518 42288 525558
rect 42628 525518 42656 526759
rect 42260 525490 42656 525518
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 35806 430128 35862 430137
rect 35806 430063 35862 430072
rect 35820 429214 35848 430063
rect 35808 429208 35860 429214
rect 35808 429150 35860 429156
rect 41696 429208 41748 429214
rect 41748 429156 42196 429162
rect 41696 429150 42196 429156
rect 41708 429134 42196 429150
rect 35806 428496 35862 428505
rect 35806 428431 35862 428440
rect 35820 427990 35848 428431
rect 35808 427984 35860 427990
rect 35808 427926 35860 427932
rect 41696 427984 41748 427990
rect 41696 427926 41748 427932
rect 41708 427666 41736 427926
rect 41708 427638 42012 427666
rect 41984 426465 42012 427638
rect 42168 427145 42196 429134
rect 43180 427417 43208 554367
rect 43166 427408 43222 427417
rect 43166 427343 43222 427352
rect 42154 427136 42210 427145
rect 42154 427071 42210 427080
rect 41142 426456 41198 426465
rect 41142 426391 41198 426400
rect 41970 426456 42026 426465
rect 41970 426391 42026 426400
rect 42798 426456 42854 426465
rect 42798 426391 42854 426400
rect 40958 426048 41014 426057
rect 40958 425983 41014 425992
rect 39302 425640 39358 425649
rect 39302 425575 39358 425584
rect 32034 424824 32090 424833
rect 32034 424759 32090 424768
rect 32048 417450 32076 424759
rect 34518 424416 34574 424425
rect 34518 424351 34574 424360
rect 33782 424008 33838 424017
rect 33782 423943 33838 423952
rect 32036 417444 32088 417450
rect 32036 417386 32088 417392
rect 33796 414633 33824 423943
rect 34532 416090 34560 424351
rect 34520 416084 34572 416090
rect 34520 416026 34572 416032
rect 39316 415313 39344 425575
rect 40972 424386 41000 425983
rect 41156 424538 41184 426391
rect 41156 424510 41460 424538
rect 40960 424380 41012 424386
rect 40960 424322 41012 424328
rect 41142 423600 41198 423609
rect 41432 423586 41460 424510
rect 41696 424380 41748 424386
rect 41748 424340 42012 424368
rect 41696 424322 41748 424328
rect 41786 423600 41842 423609
rect 41432 423558 41786 423586
rect 41142 423535 41198 423544
rect 41786 423535 41842 423544
rect 41156 422414 41184 423535
rect 41144 422408 41196 422414
rect 41144 422350 41196 422356
rect 41604 422408 41656 422414
rect 41656 422385 41828 422396
rect 41656 422376 41842 422385
rect 41656 422368 41786 422376
rect 41604 422350 41656 422356
rect 41786 422311 41842 422320
rect 41786 421968 41842 421977
rect 41616 421926 41786 421954
rect 41616 418713 41644 421926
rect 41786 421903 41842 421912
rect 41786 421560 41842 421569
rect 41786 421495 41842 421504
rect 41602 418704 41658 418713
rect 41602 418639 41658 418648
rect 41800 418441 41828 421495
rect 41786 418432 41842 418441
rect 41786 418367 41842 418376
rect 41984 418154 42012 424340
rect 41984 418126 42380 418154
rect 41696 417444 41748 417450
rect 41696 417386 41748 417392
rect 41708 417330 41736 417386
rect 41708 417314 42104 417330
rect 41708 417308 42116 417314
rect 41708 417302 42064 417308
rect 42064 417250 42116 417256
rect 41696 416084 41748 416090
rect 41696 416026 41748 416032
rect 41708 415970 41736 416026
rect 41708 415942 42288 415970
rect 39302 415304 39358 415313
rect 39302 415239 39358 415248
rect 33782 414624 33838 414633
rect 33782 414559 33838 414568
rect 42260 413114 42288 415942
rect 42168 413086 42288 413114
rect 42168 412624 42196 413086
rect 42352 412634 42380 418126
rect 42616 417308 42668 417314
rect 42616 417250 42668 417256
rect 42260 412606 42380 412634
rect 42260 411346 42288 412606
rect 42168 411318 42288 411346
rect 42168 410788 42196 411318
rect 42182 410162 42472 410190
rect 42248 409828 42300 409834
rect 42248 409770 42300 409776
rect 42260 408966 42288 409770
rect 42182 408938 42288 408966
rect 42168 408218 42196 408340
rect 42168 408190 42288 408218
rect 42062 408096 42118 408105
rect 42062 408031 42118 408040
rect 42076 407796 42104 408031
rect 42260 407130 42288 408190
rect 42444 407289 42472 410162
rect 42430 407280 42486 407289
rect 42430 407215 42486 407224
rect 41800 407017 41828 407116
rect 42260 407102 42472 407130
rect 42248 407040 42300 407046
rect 41786 407008 41842 407017
rect 42248 406982 42300 406988
rect 41786 406943 41842 406952
rect 41786 406736 41842 406745
rect 41786 406671 41842 406680
rect 41800 406504 41828 406671
rect 42260 406042 42288 406982
rect 42168 406014 42288 406042
rect 42168 405929 42196 406014
rect 42444 404977 42472 407102
rect 42628 407046 42656 417250
rect 42616 407040 42668 407046
rect 42616 406982 42668 406988
rect 42430 404968 42486 404977
rect 42430 404903 42486 404912
rect 42246 404560 42302 404569
rect 42246 404495 42302 404504
rect 42260 403458 42288 404495
rect 42182 403430 42288 403458
rect 42338 402928 42394 402937
rect 42168 402886 42338 402914
rect 42168 402801 42196 402886
rect 42338 402863 42394 402872
rect 42246 402520 42302 402529
rect 42246 402455 42302 402464
rect 42260 402166 42288 402455
rect 42432 402280 42484 402286
rect 42432 402222 42484 402228
rect 42182 402138 42288 402166
rect 42444 401622 42472 402222
rect 42182 401594 42472 401622
rect 41786 400072 41842 400081
rect 41786 400007 41842 400016
rect 41800 399772 41828 400007
rect 41786 399392 41842 399401
rect 41786 399327 41842 399336
rect 41800 399121 41828 399327
rect 41970 398848 42026 398857
rect 41970 398783 42026 398792
rect 41984 398480 42012 398783
rect 42168 395729 42196 397936
rect 42154 395720 42210 395729
rect 42154 395655 42210 395664
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41326 387152 41382 387161
rect 41326 387087 41382 387096
rect 41142 386744 41198 386753
rect 41142 386679 41198 386688
rect 41156 385937 41184 386679
rect 41340 386442 41368 387087
rect 41328 386436 41380 386442
rect 41328 386378 41380 386384
rect 41696 386436 41748 386442
rect 41748 386396 41920 386424
rect 41696 386378 41748 386384
rect 40958 385928 41014 385937
rect 40958 385863 41014 385872
rect 41142 385928 41198 385937
rect 41142 385863 41198 385872
rect 40972 382265 41000 385863
rect 41142 383072 41198 383081
rect 41142 383007 41198 383016
rect 40038 382256 40094 382265
rect 40038 382191 40094 382200
rect 40958 382256 41014 382265
rect 40958 382191 41014 382200
rect 35438 381848 35494 381857
rect 35438 381783 35494 381792
rect 33966 381032 34022 381041
rect 33966 380967 34022 380976
rect 33980 373318 34008 380967
rect 35452 374649 35480 381783
rect 39302 381440 39358 381449
rect 39302 381375 39358 381384
rect 35808 379568 35860 379574
rect 35808 379510 35860 379516
rect 35820 379409 35848 379510
rect 35806 379400 35862 379409
rect 35806 379335 35862 379344
rect 35808 378208 35860 378214
rect 35806 378176 35808 378185
rect 35860 378176 35862 378185
rect 35806 378111 35862 378120
rect 35806 376544 35862 376553
rect 35806 376479 35862 376488
rect 35820 376145 35848 376479
rect 35806 376136 35862 376145
rect 35806 376071 35862 376080
rect 35438 374640 35494 374649
rect 35438 374575 35494 374584
rect 33968 373312 34020 373318
rect 33968 373254 34020 373260
rect 39316 372094 39344 381375
rect 40052 379409 40080 382191
rect 41156 381857 41184 383007
rect 41326 382664 41382 382673
rect 41326 382599 41382 382608
rect 41340 382294 41368 382599
rect 41328 382288 41380 382294
rect 41328 382230 41380 382236
rect 41696 382288 41748 382294
rect 41696 382230 41748 382236
rect 41142 381848 41198 381857
rect 41142 381783 41198 381792
rect 41326 379808 41382 379817
rect 41326 379743 41328 379752
rect 41380 379743 41382 379752
rect 41510 379808 41566 379817
rect 41510 379743 41512 379752
rect 41328 379714 41380 379720
rect 41564 379743 41566 379752
rect 41512 379714 41564 379720
rect 40408 379636 40460 379642
rect 40408 379578 40460 379584
rect 40038 379400 40094 379409
rect 40038 379335 40094 379344
rect 40420 376961 40448 379578
rect 41708 379514 41736 382230
rect 41892 381585 41920 386396
rect 42812 385665 42840 426391
rect 42982 425232 43038 425241
rect 42982 425167 43038 425176
rect 42996 402286 43024 425167
rect 43166 422784 43222 422793
rect 43166 422719 43222 422728
rect 43180 409834 43208 422719
rect 43168 409828 43220 409834
rect 43168 409770 43220 409776
rect 42984 402280 43036 402286
rect 42984 402222 43036 402228
rect 42798 385656 42854 385665
rect 42798 385591 42854 385600
rect 43258 385248 43314 385257
rect 43258 385183 43314 385192
rect 41878 381576 41934 381585
rect 41878 381511 41934 381520
rect 42890 380760 42946 380769
rect 42890 380695 42946 380704
rect 41708 379486 42380 379514
rect 41696 378208 41748 378214
rect 41694 378176 41696 378185
rect 41748 378176 41750 378185
rect 41694 378111 41750 378120
rect 40406 376952 40462 376961
rect 40406 376887 40462 376896
rect 41696 373312 41748 373318
rect 41748 373260 42288 373266
rect 41696 373254 42288 373260
rect 41708 373238 42288 373254
rect 39304 372088 39356 372094
rect 39304 372030 39356 372036
rect 41696 372088 41748 372094
rect 41748 372036 42104 372042
rect 41696 372030 42104 372036
rect 41708 372014 42104 372030
rect 42076 371958 42104 372014
rect 42064 371952 42116 371958
rect 42064 371894 42116 371900
rect 42260 369458 42288 373238
rect 42182 369430 42288 369458
rect 42352 367622 42380 379486
rect 42708 371952 42760 371958
rect 42708 371894 42760 371900
rect 42182 367594 42380 367622
rect 42182 366947 42288 366975
rect 42260 365906 42288 366947
rect 42432 366852 42484 366858
rect 42432 366794 42484 366800
rect 42248 365900 42300 365906
rect 42248 365842 42300 365848
rect 42444 365786 42472 366794
rect 42720 366602 42748 371894
rect 42182 365758 42472 365786
rect 42536 366574 42748 366602
rect 42182 365107 42288 365135
rect 41786 364848 41842 364857
rect 41786 364783 41842 364792
rect 41800 364548 41828 364783
rect 42260 364334 42288 365107
rect 42260 364306 42380 364334
rect 41786 364168 41842 364177
rect 41786 364103 41842 364112
rect 41800 363936 41828 364103
rect 42154 363624 42210 363633
rect 42154 363559 42210 363568
rect 42168 363256 42196 363559
rect 42352 362914 42380 364306
rect 42340 362908 42392 362914
rect 42340 362850 42392 362856
rect 42168 362766 42288 362794
rect 42168 362712 42196 362766
rect 42260 362726 42288 362766
rect 42536 362726 42564 366574
rect 42708 365900 42760 365906
rect 42708 365842 42760 365848
rect 42720 363089 42748 365842
rect 42706 363080 42762 363089
rect 42706 363015 42762 363024
rect 42708 362908 42760 362914
rect 42708 362850 42760 362856
rect 42260 362698 42564 362726
rect 42720 362273 42748 362850
rect 42706 362264 42762 362273
rect 42706 362199 42762 362208
rect 41800 360097 41828 360264
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 42154 359952 42210 359961
rect 42154 359887 42210 359896
rect 42168 359584 42196 359887
rect 42430 359000 42486 359009
rect 42182 358958 42430 358986
rect 42430 358935 42486 358944
rect 41878 358728 41934 358737
rect 41878 358663 41934 358672
rect 41892 358428 41920 358663
rect 41786 356960 41842 356969
rect 41786 356895 41842 356904
rect 41800 356592 41828 356895
rect 42904 356046 42932 380695
rect 43074 376952 43130 376961
rect 43074 376887 43130 376896
rect 43088 366858 43116 376887
rect 43076 366852 43128 366858
rect 43076 366794 43128 366800
rect 42248 356040 42300 356046
rect 42892 356040 42944 356046
rect 42248 355982 42300 355988
rect 42430 356008 42486 356017
rect 42260 355926 42288 355982
rect 42892 355982 42944 355988
rect 42430 355943 42486 355952
rect 42182 355898 42288 355926
rect 41878 355736 41934 355745
rect 41878 355671 41934 355680
rect 41892 355300 41920 355671
rect 42444 354739 42472 355943
rect 42182 354711 42472 354739
rect 43272 345545 43300 385183
rect 43456 354793 43484 589319
rect 44376 578105 44404 593127
rect 44362 578096 44418 578105
rect 44362 578031 44418 578040
rect 44652 558793 44680 600063
rect 45112 599729 45140 639775
rect 45098 599720 45154 599729
rect 45098 599655 45154 599664
rect 44914 599312 44970 599321
rect 44914 599247 44970 599256
rect 44638 558784 44694 558793
rect 44638 558719 44694 558728
rect 44928 556481 44956 599247
rect 45296 598097 45324 640183
rect 45480 598913 45508 640290
rect 46216 613426 46244 641407
rect 46204 613420 46256 613426
rect 46204 613362 46256 613368
rect 46202 611688 46258 611697
rect 46202 611623 46258 611632
rect 45466 598904 45522 598913
rect 45466 598839 45522 598848
rect 45282 598088 45338 598097
rect 45282 598023 45338 598032
rect 45098 580272 45154 580281
rect 45098 580207 45154 580216
rect 45112 575482 45140 580207
rect 45100 575476 45152 575482
rect 45100 575418 45152 575424
rect 45098 556880 45154 556889
rect 45098 556815 45154 556824
rect 44914 556472 44970 556481
rect 44914 556407 44970 556416
rect 44638 556064 44694 556073
rect 44638 555999 44694 556008
rect 44362 555248 44418 555257
rect 44362 555183 44418 555192
rect 43994 551848 44050 551857
rect 43994 551783 44050 551792
rect 43810 550760 43866 550769
rect 43810 550695 43866 550704
rect 43626 547768 43682 547777
rect 43626 547703 43682 547712
rect 43442 354784 43498 354793
rect 43442 354719 43498 354728
rect 43640 354113 43668 547703
rect 43824 532817 43852 550695
rect 44008 533905 44036 551783
rect 44178 548720 44234 548729
rect 44178 548655 44234 548664
rect 44192 536897 44220 548655
rect 44178 536888 44234 536897
rect 44178 536823 44234 536832
rect 43994 533896 44050 533905
rect 43994 533831 44050 533840
rect 43810 532808 43866 532817
rect 43810 532743 43866 532752
rect 44376 428097 44404 555183
rect 44652 428913 44680 555999
rect 44822 550488 44878 550497
rect 44822 550423 44878 550432
rect 44836 539617 44864 550423
rect 45112 543734 45140 556815
rect 45282 551576 45338 551585
rect 45282 551511 45338 551520
rect 45020 543706 45140 543734
rect 44822 539608 44878 539617
rect 44822 539543 44878 539552
rect 44822 537432 44878 537441
rect 44822 537367 44878 537376
rect 44836 532030 44864 537367
rect 44824 532024 44876 532030
rect 44824 531966 44876 531972
rect 45020 429729 45048 543706
rect 45296 529825 45324 551511
rect 45282 529816 45338 529825
rect 45282 529751 45338 529760
rect 45192 528624 45244 528630
rect 45192 528566 45244 528572
rect 45204 527241 45232 528566
rect 45190 527232 45246 527241
rect 45190 527167 45246 527176
rect 45282 430944 45338 430953
rect 45282 430879 45338 430888
rect 45006 429720 45062 429729
rect 45006 429655 45062 429664
rect 45098 429312 45154 429321
rect 45098 429247 45154 429256
rect 44638 428904 44694 428913
rect 44638 428839 44694 428848
rect 44362 428088 44418 428097
rect 44362 428023 44418 428032
rect 44362 427680 44418 427689
rect 44362 427615 44418 427624
rect 44178 426864 44234 426873
rect 44178 426799 44234 426808
rect 43810 422376 43866 422385
rect 43810 422311 43866 422320
rect 43824 402529 43852 422311
rect 43994 421152 44050 421161
rect 43994 421087 44050 421096
rect 44008 408105 44036 421087
rect 43994 408096 44050 408105
rect 43994 408031 44050 408040
rect 43810 402520 43866 402529
rect 43810 402455 43866 402464
rect 44192 384033 44220 426799
rect 44376 384849 44404 427615
rect 44546 423192 44602 423201
rect 44546 423127 44602 423136
rect 44560 402937 44588 423127
rect 44730 407280 44786 407289
rect 44730 407215 44786 407224
rect 44744 404326 44772 407215
rect 44732 404320 44784 404326
rect 44732 404262 44784 404268
rect 45112 402974 45140 429247
rect 45296 412634 45324 430879
rect 45466 420744 45522 420753
rect 45466 420679 45522 420688
rect 45480 412634 45508 420679
rect 45020 402946 45140 402974
rect 45204 412606 45324 412634
rect 45388 412606 45508 412634
rect 44546 402928 44602 402937
rect 44546 402863 44602 402872
rect 45020 400194 45048 402946
rect 45204 400314 45232 412606
rect 45192 400308 45244 400314
rect 45192 400250 45244 400256
rect 45020 400166 45140 400194
rect 45112 386481 45140 400166
rect 45098 386472 45154 386481
rect 45098 386407 45154 386416
rect 44362 384840 44418 384849
rect 44362 384775 44418 384784
rect 45190 384432 45246 384441
rect 45190 384367 45246 384376
rect 45204 384282 45232 384367
rect 45204 384254 45324 384282
rect 44178 384024 44234 384033
rect 44178 383959 44234 383968
rect 45098 383616 45154 383625
rect 45098 383551 45154 383560
rect 44914 382256 44970 382265
rect 44914 382191 44970 382200
rect 44638 380352 44694 380361
rect 44638 380287 44694 380296
rect 43810 379808 43866 379817
rect 43810 379743 43866 379752
rect 43824 359961 43852 379743
rect 43994 378176 44050 378185
rect 43994 378111 44050 378120
rect 44008 363633 44036 378111
rect 44270 377496 44326 377505
rect 44270 377431 44326 377440
rect 43994 363624 44050 363633
rect 43994 363559 44050 363568
rect 44284 360194 44312 377431
rect 44652 364334 44680 380287
rect 44192 360166 44312 360194
rect 44468 364306 44680 364334
rect 43810 359952 43866 359961
rect 43810 359887 43866 359896
rect 43626 354104 43682 354113
rect 43626 354039 43682 354048
rect 44192 353161 44220 360166
rect 44468 359009 44496 364306
rect 44638 363080 44694 363089
rect 44638 363015 44694 363024
rect 44652 361554 44680 363015
rect 44640 361548 44692 361554
rect 44640 361490 44692 361496
rect 44454 359000 44510 359009
rect 44454 358935 44510 358944
rect 44640 357468 44692 357474
rect 44640 357410 44692 357416
rect 44652 356017 44680 357410
rect 44638 356008 44694 356017
rect 44638 355943 44694 355952
rect 44454 354784 44510 354793
rect 44454 354719 44510 354728
rect 44468 354362 44496 354719
rect 44640 354544 44692 354550
rect 44638 354512 44640 354521
rect 44692 354512 44694 354521
rect 44638 354447 44694 354456
rect 44468 354346 44772 354362
rect 44468 354340 44784 354346
rect 44468 354334 44732 354340
rect 44732 354282 44784 354288
rect 44178 353152 44234 353161
rect 44178 353087 44234 353096
rect 40222 345536 40278 345545
rect 40222 345471 40278 345480
rect 43258 345536 43314 345545
rect 43258 345471 43314 345480
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 35808 344616 35860 344622
rect 35808 344558 35860 344564
rect 40040 344616 40092 344622
rect 40040 344558 40092 344564
rect 35820 344321 35848 344558
rect 40052 344321 40080 344558
rect 35530 344312 35586 344321
rect 35530 344247 35586 344256
rect 35806 344312 35862 344321
rect 35806 344247 35862 344256
rect 40038 344312 40094 344321
rect 40038 344247 40094 344256
rect 35544 343806 35572 344247
rect 35532 343800 35584 343806
rect 35532 343742 35584 343748
rect 40040 343800 40092 343806
rect 40040 343742 40092 343748
rect 33046 343496 33102 343505
rect 33046 343431 33102 343440
rect 33060 341426 33088 343431
rect 35808 342304 35860 342310
rect 35806 342272 35808 342281
rect 35860 342272 35862 342281
rect 35806 342207 35862 342216
rect 40052 341873 40080 343742
rect 40236 342310 40264 345471
rect 44928 343369 44956 382191
rect 44914 343360 44970 343369
rect 44914 343295 44970 343304
rect 40224 342304 40276 342310
rect 40224 342246 40276 342252
rect 40038 341864 40094 341873
rect 40038 341799 40094 341808
rect 35622 341456 35678 341465
rect 33048 341420 33100 341426
rect 35622 341391 35678 341400
rect 40222 341456 40278 341465
rect 40222 341391 40224 341400
rect 33048 341362 33100 341368
rect 35636 341086 35664 341391
rect 40276 341391 40278 341400
rect 40224 341362 40276 341368
rect 35808 341216 35860 341222
rect 35808 341158 35860 341164
rect 40224 341216 40276 341222
rect 40224 341158 40276 341164
rect 35624 341080 35676 341086
rect 35820 341057 35848 341158
rect 40040 341080 40092 341086
rect 35624 341022 35676 341028
rect 35806 341048 35862 341057
rect 35806 340983 35862 340992
rect 39854 341048 39910 341057
rect 40236 341057 40264 341158
rect 45112 341057 45140 383551
rect 45296 369854 45324 384254
rect 45204 369826 45324 369854
rect 45204 345014 45232 369826
rect 45388 360194 45416 412606
rect 45296 360166 45416 360194
rect 45296 353734 45324 360166
rect 45468 354612 45520 354618
rect 45468 354554 45520 354560
rect 45480 354385 45508 354554
rect 45466 354376 45522 354385
rect 45466 354311 45522 354320
rect 45468 354136 45520 354142
rect 45466 354104 45468 354113
rect 45520 354104 45522 354113
rect 45466 354039 45522 354048
rect 45468 353864 45520 353870
rect 45468 353806 45520 353812
rect 45296 353728 45355 353734
rect 45296 353676 45303 353728
rect 45296 353670 45355 353676
rect 45296 353654 45343 353670
rect 45480 353433 45508 353806
rect 45466 353424 45522 353433
rect 45466 353359 45522 353368
rect 45422 353184 45474 353190
rect 45420 353152 45422 353161
rect 45474 353152 45476 353161
rect 45420 353087 45476 353096
rect 45204 344986 45324 345014
rect 40040 341022 40092 341028
rect 40222 341048 40278 341057
rect 39854 340983 39910 340992
rect 39868 339833 39896 340983
rect 40052 340649 40080 341022
rect 40222 340983 40278 340992
rect 45098 341048 45154 341057
rect 45098 340983 45154 340992
rect 45296 340649 45324 344986
rect 45466 341456 45522 341465
rect 45466 341391 45468 341400
rect 45520 341391 45522 341400
rect 45468 341362 45520 341368
rect 40038 340640 40094 340649
rect 40038 340575 40094 340584
rect 45282 340640 45338 340649
rect 45282 340575 45338 340584
rect 35530 339824 35586 339833
rect 35530 339759 35586 339768
rect 35806 339824 35862 339833
rect 35806 339759 35862 339768
rect 39854 339824 39910 339833
rect 39854 339759 39910 339768
rect 35544 339658 35572 339759
rect 35532 339652 35584 339658
rect 35532 339594 35584 339600
rect 35820 339522 35848 339759
rect 36544 339652 36596 339658
rect 36544 339594 36596 339600
rect 35808 339516 35860 339522
rect 35808 339458 35860 339464
rect 35162 338600 35218 338609
rect 35162 338535 35218 338544
rect 35176 331809 35204 338535
rect 35806 336152 35862 336161
rect 35806 336087 35862 336096
rect 35820 335374 35848 336087
rect 35808 335368 35860 335374
rect 35808 335310 35860 335316
rect 35622 334928 35678 334937
rect 35622 334863 35678 334872
rect 35636 334286 35664 334863
rect 35806 334520 35862 334529
rect 35806 334455 35862 334464
rect 35624 334280 35676 334286
rect 35624 334222 35676 334228
rect 35820 334014 35848 334455
rect 35808 334008 35860 334014
rect 35808 333950 35860 333956
rect 36556 332897 36584 339594
rect 38844 339516 38896 339522
rect 38844 339458 38896 339464
rect 38856 336569 38884 339458
rect 45650 338464 45706 338473
rect 45650 338399 45706 338408
rect 45466 336832 45522 336841
rect 45466 336767 45522 336776
rect 38842 336560 38898 336569
rect 38842 336495 38898 336504
rect 40224 335368 40276 335374
rect 40224 335310 40276 335316
rect 40236 334529 40264 335310
rect 43994 334656 44050 334665
rect 43994 334591 44050 334600
rect 40222 334520 40278 334529
rect 40222 334455 40278 334464
rect 43166 334520 43222 334529
rect 43166 334455 43222 334464
rect 39396 334280 39448 334286
rect 39396 334222 39448 334228
rect 36542 332888 36598 332897
rect 36542 332823 36598 332832
rect 39408 332489 39436 334222
rect 41696 334008 41748 334014
rect 42064 334008 42116 334014
rect 41748 333956 42064 333962
rect 41696 333950 42116 333956
rect 42984 334008 43036 334014
rect 42984 333950 43036 333956
rect 41708 333934 42104 333950
rect 39394 332480 39450 332489
rect 39394 332415 39450 332424
rect 42798 332480 42854 332489
rect 42798 332415 42854 332424
rect 35162 331800 35218 331809
rect 35162 331735 35218 331744
rect 42168 325938 42196 326264
rect 42168 325910 42288 325938
rect 41786 324864 41842 324873
rect 41786 324799 41842 324808
rect 41800 324428 41828 324799
rect 42260 324329 42288 325910
rect 42246 324320 42302 324329
rect 42246 324255 42302 324264
rect 42182 323734 42472 323762
rect 42248 322924 42300 322930
rect 42248 322866 42300 322872
rect 42260 322810 42288 322866
rect 42076 322782 42288 322810
rect 42076 322592 42104 322782
rect 42182 321898 42288 321926
rect 42076 321201 42104 321368
rect 41786 321192 41842 321201
rect 41786 321127 41842 321136
rect 42062 321192 42118 321201
rect 42062 321127 42118 321136
rect 41800 320725 41828 321127
rect 42260 320278 42288 321898
rect 42444 320793 42472 323734
rect 42430 320784 42486 320793
rect 42430 320719 42486 320728
rect 42248 320272 42300 320278
rect 42248 320214 42300 320220
rect 42812 320090 42840 332415
rect 42996 321201 43024 333950
rect 43180 322930 43208 334455
rect 43168 322924 43220 322930
rect 43168 322866 43220 322872
rect 42982 321192 43038 321201
rect 42982 321127 43038 321136
rect 42182 320062 42840 320090
rect 42616 320000 42668 320006
rect 42616 319942 42668 319948
rect 42182 319518 42472 319546
rect 42444 319161 42472 319518
rect 42628 319433 42656 319942
rect 42614 319424 42670 319433
rect 42614 319359 42670 319368
rect 42430 319152 42486 319161
rect 42430 319087 42486 319096
rect 41786 317384 41842 317393
rect 41786 317319 41842 317328
rect 41800 317045 41828 317319
rect 42182 316390 42472 316418
rect 41786 316024 41842 316033
rect 41786 315959 41842 315968
rect 41800 315757 41828 315959
rect 41786 315616 41842 315625
rect 41786 315551 41842 315560
rect 41800 315180 41828 315551
rect 42444 314673 42472 316390
rect 42430 314664 42486 314673
rect 42430 314599 42486 314608
rect 41786 313712 41842 313721
rect 41786 313647 41842 313656
rect 41800 313344 41828 313647
rect 42430 312760 42486 312769
rect 42182 312718 42430 312746
rect 42430 312695 42486 312704
rect 42168 312174 42288 312202
rect 42168 312052 42196 312174
rect 42260 312066 42288 312174
rect 42260 312038 42472 312066
rect 42076 310457 42104 311508
rect 42062 310448 42118 310457
rect 42062 310383 42118 310392
rect 42444 310185 42472 312038
rect 42430 310176 42486 310185
rect 42430 310111 42486 310120
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41142 300520 41198 300529
rect 41142 300455 41198 300464
rect 41156 299674 41184 300455
rect 42890 299704 42946 299713
rect 41144 299668 41196 299674
rect 41144 299610 41196 299616
rect 41604 299668 41656 299674
rect 41656 299628 41828 299656
rect 42890 299639 42946 299648
rect 41604 299610 41656 299616
rect 41800 299474 41828 299628
rect 41800 299446 42012 299474
rect 41984 297401 42012 299446
rect 41970 297392 42026 297401
rect 41970 297327 42026 297336
rect 41326 296440 41382 296449
rect 41326 296375 41382 296384
rect 40958 296032 41014 296041
rect 40958 295967 41014 295976
rect 39302 295624 39358 295633
rect 39302 295559 39358 295568
rect 33782 294808 33838 294817
rect 33782 294743 33838 294752
rect 33796 286346 33824 294743
rect 37922 294400 37978 294409
rect 37922 294335 37978 294344
rect 33784 286340 33836 286346
rect 33784 286282 33836 286288
rect 37936 284345 37964 294335
rect 39316 284782 39344 295559
rect 40972 293026 41000 295967
rect 41340 295662 41368 296375
rect 41328 295656 41380 295662
rect 41328 295598 41380 295604
rect 41696 295656 41748 295662
rect 41696 295598 41748 295604
rect 41142 295216 41198 295225
rect 41142 295151 41198 295160
rect 41156 293026 41184 295151
rect 40972 292998 41092 293026
rect 41156 292998 41276 293026
rect 41064 292890 41092 292998
rect 41064 292862 41184 292890
rect 41156 292262 41184 292862
rect 41248 292574 41276 292998
rect 41708 292574 41736 295598
rect 42706 292768 42762 292777
rect 42706 292703 42762 292712
rect 41248 292546 41368 292574
rect 41708 292546 42472 292574
rect 41340 292482 41368 292546
rect 41340 292454 41552 292482
rect 41524 292346 41552 292454
rect 41524 292318 42380 292346
rect 41144 292256 41196 292262
rect 41144 292198 41196 292204
rect 41604 292256 41656 292262
rect 41786 292224 41842 292233
rect 41656 292204 41786 292210
rect 41604 292198 41786 292204
rect 41616 292182 41786 292198
rect 41786 292159 41842 292168
rect 41234 291544 41290 291553
rect 41234 291479 41290 291488
rect 41248 291310 41276 291479
rect 41236 291304 41288 291310
rect 41236 291246 41288 291252
rect 41696 291304 41748 291310
rect 41748 291281 42012 291292
rect 41748 291272 42026 291281
rect 41748 291264 41970 291272
rect 41696 291246 41748 291252
rect 41970 291207 42026 291216
rect 41786 290320 41842 290329
rect 41786 290255 41842 290264
rect 41800 289241 41828 290255
rect 41786 289232 41842 289241
rect 41786 289167 41842 289176
rect 41696 286340 41748 286346
rect 41696 286282 41748 286288
rect 41708 286226 41736 286282
rect 41708 286198 42288 286226
rect 39304 284776 39356 284782
rect 39304 284718 39356 284724
rect 41696 284776 41748 284782
rect 41748 284724 42104 284730
rect 41696 284718 42104 284724
rect 41708 284714 42104 284718
rect 41708 284708 42116 284714
rect 41708 284702 42064 284708
rect 42064 284650 42116 284656
rect 37922 284336 37978 284345
rect 37922 284271 37978 284280
rect 42260 283059 42288 286198
rect 42352 284458 42380 292318
rect 42444 289814 42472 292546
rect 42720 289814 42748 292703
rect 42444 289786 42564 289814
rect 42720 289786 42840 289814
rect 42536 284889 42564 289786
rect 42522 284880 42578 284889
rect 42522 284815 42578 284824
rect 42616 284708 42668 284714
rect 42616 284650 42668 284656
rect 42352 284430 42564 284458
rect 42182 283031 42288 283059
rect 41786 282296 41842 282305
rect 41786 282231 41842 282240
rect 41800 281860 41828 282231
rect 42154 281752 42210 281761
rect 42154 281687 42210 281696
rect 42168 281180 42196 281687
rect 42168 280265 42196 280568
rect 42154 280256 42210 280265
rect 42154 280191 42210 280200
rect 42536 280154 42564 284430
rect 42444 280126 42564 280154
rect 42154 279712 42210 279721
rect 42154 279647 42210 279656
rect 42168 279344 42196 279647
rect 42182 278718 42380 278746
rect 42062 278488 42118 278497
rect 42062 278423 42118 278432
rect 42076 278188 42104 278423
rect 42154 277944 42210 277953
rect 42154 277879 42210 277888
rect 42168 277508 42196 277879
rect 42352 277794 42380 278718
rect 42260 277766 42380 277794
rect 42260 277370 42288 277766
rect 42248 277364 42300 277370
rect 42248 277306 42300 277312
rect 41786 277128 41842 277137
rect 41786 277063 41842 277072
rect 41800 276896 41828 277063
rect 42444 276366 42472 280126
rect 42168 276298 42196 276352
rect 42260 276338 42472 276366
rect 42260 276298 42288 276338
rect 42168 276270 42288 276298
rect 41786 274272 41842 274281
rect 41786 274207 41842 274216
rect 41800 273836 41828 274207
rect 42168 273057 42196 273224
rect 42432 273216 42484 273222
rect 42432 273158 42484 273164
rect 42154 273048 42210 273057
rect 42154 272983 42210 272992
rect 42444 272558 42472 273158
rect 42182 272530 42472 272558
rect 42628 272014 42656 284650
rect 42812 277953 42840 289786
rect 42904 287722 42932 299639
rect 43166 293992 43222 294001
rect 43166 293927 43222 293936
rect 42904 287694 43024 287722
rect 42798 277944 42854 277953
rect 42798 277879 42854 277888
rect 42800 277364 42852 277370
rect 42800 277306 42852 277312
rect 42812 275913 42840 277306
rect 42798 275904 42854 275913
rect 42798 275839 42854 275848
rect 42996 273254 43024 287694
rect 43180 282914 43208 293927
rect 43442 293176 43498 293185
rect 43442 293111 43498 293120
rect 43180 282886 43300 282914
rect 42182 271986 42656 272014
rect 42812 273226 43024 273254
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 41800 270164 41828 270399
rect 41786 269784 41842 269793
rect 41786 269719 41842 269728
rect 41800 269521 41828 269719
rect 41970 269104 42026 269113
rect 41970 269039 42026 269048
rect 41984 268872 42012 269039
rect 42168 266257 42196 268328
rect 42154 266248 42210 266257
rect 42154 266183 42210 266192
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 42812 257145 42840 273226
rect 43272 273222 43300 282886
rect 43456 279721 43484 293111
rect 43626 291272 43682 291281
rect 43626 291207 43682 291216
rect 43442 279712 43498 279721
rect 43442 279647 43498 279656
rect 43640 278497 43668 291207
rect 43626 278488 43682 278497
rect 43626 278423 43682 278432
rect 43442 273864 43498 273873
rect 43442 273799 43498 273808
rect 43260 273216 43312 273222
rect 43260 273158 43312 273164
rect 43456 263594 43484 273799
rect 43364 263566 43484 263594
rect 35622 257136 35678 257145
rect 35622 257071 35678 257080
rect 39486 257136 39542 257145
rect 39486 257071 39542 257080
rect 42798 257136 42854 257145
rect 42798 257071 42854 257080
rect 35636 256766 35664 257071
rect 39500 256970 39528 257071
rect 35808 256964 35860 256970
rect 35808 256906 35860 256912
rect 39488 256964 39540 256970
rect 39488 256906 39540 256912
rect 35624 256760 35676 256766
rect 35820 256737 35848 256906
rect 43364 256766 43392 263566
rect 41696 256760 41748 256766
rect 35624 256702 35676 256708
rect 35806 256728 35862 256737
rect 42064 256760 42116 256766
rect 41748 256708 42064 256714
rect 41696 256702 42116 256708
rect 43352 256760 43404 256766
rect 43352 256702 43404 256708
rect 41708 256686 42104 256702
rect 35806 256663 35862 256672
rect 35806 256320 35862 256329
rect 35806 256255 35862 256264
rect 35820 255474 35848 256255
rect 35808 255468 35860 255474
rect 35808 255410 35860 255416
rect 40224 255468 40276 255474
rect 40224 255410 40276 255416
rect 40236 253473 40264 255410
rect 35622 253464 35678 253473
rect 35622 253399 35678 253408
rect 40222 253464 40278 253473
rect 40222 253399 40278 253408
rect 42798 253464 42854 253473
rect 42798 253399 42854 253408
rect 35636 252754 35664 253399
rect 35806 253056 35862 253065
rect 35806 252991 35862 253000
rect 35624 252748 35676 252754
rect 35624 252690 35676 252696
rect 35820 252618 35848 252991
rect 40684 252748 40736 252754
rect 40684 252690 40736 252696
rect 35808 252612 35860 252618
rect 35808 252554 35860 252560
rect 35806 252240 35862 252249
rect 35806 252175 35862 252184
rect 35820 251258 35848 252175
rect 35808 251252 35860 251258
rect 35808 251194 35860 251200
rect 39304 251252 39356 251258
rect 39304 251194 39356 251200
rect 35622 250608 35678 250617
rect 35622 250543 35678 250552
rect 35636 250102 35664 250543
rect 35806 250200 35862 250209
rect 35806 250135 35862 250144
rect 35624 250096 35676 250102
rect 35624 250038 35676 250044
rect 35820 249830 35848 250135
rect 35808 249824 35860 249830
rect 35808 249766 35860 249772
rect 35806 247752 35862 247761
rect 35806 247687 35862 247696
rect 35820 247314 35848 247687
rect 35808 247308 35860 247314
rect 35808 247250 35860 247256
rect 34426 246936 34482 246945
rect 34426 246871 34482 246880
rect 34440 242214 34468 246871
rect 39316 242758 39344 251194
rect 40132 250096 40184 250102
rect 40132 250038 40184 250044
rect 39856 247308 39908 247314
rect 39856 247250 39908 247256
rect 39868 244089 39896 247250
rect 40144 245721 40172 250038
rect 40130 245712 40186 245721
rect 40130 245647 40186 245656
rect 39854 244080 39910 244089
rect 39854 244015 39910 244024
rect 39304 242752 39356 242758
rect 39304 242694 39356 242700
rect 34428 242208 34480 242214
rect 34428 242150 34480 242156
rect 40696 240961 40724 252690
rect 41328 252612 41380 252618
rect 41328 252554 41380 252560
rect 41340 248414 41368 252554
rect 41696 249824 41748 249830
rect 42064 249824 42116 249830
rect 41748 249772 42064 249778
rect 41696 249766 42116 249772
rect 41708 249750 42104 249766
rect 41340 248386 41460 248414
rect 41432 244274 41460 248386
rect 41432 244246 42380 244274
rect 41696 242752 41748 242758
rect 41748 242700 42104 242706
rect 41696 242694 42104 242700
rect 41708 242690 42104 242694
rect 41708 242684 42116 242690
rect 41708 242678 42064 242684
rect 42064 242626 42116 242632
rect 41696 242208 41748 242214
rect 41748 242156 42288 242162
rect 41696 242150 42288 242156
rect 41708 242134 42288 242150
rect 40682 240952 40738 240961
rect 40682 240887 40738 240896
rect 42062 240136 42118 240145
rect 42062 240071 42118 240080
rect 42076 239836 42104 240071
rect 42260 238663 42288 242134
rect 42182 238635 42288 238663
rect 42352 238014 42380 244246
rect 42524 242684 42576 242690
rect 42524 242626 42576 242632
rect 42536 238105 42564 242626
rect 42522 238096 42578 238105
rect 42522 238031 42578 238040
rect 42182 237986 42380 238014
rect 41786 236600 41842 236609
rect 41786 236535 41842 236544
rect 41800 236164 41828 236535
rect 42430 235920 42486 235929
rect 42430 235855 42486 235864
rect 42444 234983 42472 235855
rect 42182 234955 42472 234983
rect 41786 234696 41842 234705
rect 41786 234631 41842 234640
rect 41800 234328 41828 234631
rect 42430 234560 42486 234569
rect 42430 234495 42486 234504
rect 42444 233695 42472 234495
rect 42182 233667 42472 233695
rect 42168 233158 42288 233186
rect 42168 233104 42196 233158
rect 42260 233118 42288 233158
rect 42260 233090 42472 233118
rect 42444 232257 42472 233090
rect 42430 232248 42486 232257
rect 42430 232183 42486 232192
rect 42430 231840 42486 231849
rect 42430 231775 42486 231784
rect 42444 230670 42472 231775
rect 42182 230642 42472 230670
rect 42156 230444 42208 230450
rect 42156 230386 42208 230392
rect 42168 229976 42196 230386
rect 42430 229392 42486 229401
rect 42182 229350 42430 229378
rect 42430 229327 42486 229336
rect 41970 228984 42026 228993
rect 41970 228919 42026 228928
rect 41984 228820 42012 228919
rect 42432 227724 42484 227730
rect 42432 227666 42484 227672
rect 42444 226998 42472 227666
rect 42168 226930 42196 226984
rect 42260 226970 42472 226998
rect 42260 226930 42288 226970
rect 42168 226902 42288 226930
rect 42154 226672 42210 226681
rect 42154 226607 42210 226616
rect 42168 226304 42196 226607
rect 42430 225720 42486 225729
rect 42182 225678 42430 225706
rect 42430 225655 42486 225664
rect 41694 224496 41750 224505
rect 41694 224431 41750 224440
rect 35530 217968 35586 217977
rect 35530 217903 35586 217912
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 35544 214713 35572 217903
rect 35530 214704 35586 214713
rect 35530 214639 35586 214648
rect 35806 214704 35862 214713
rect 35806 214639 35862 214648
rect 35820 213994 35848 214639
rect 41708 213994 41736 224431
rect 42168 223553 42196 225148
rect 42154 223544 42210 223553
rect 42154 223479 42210 223488
rect 35808 213988 35860 213994
rect 35808 213930 35860 213936
rect 41696 213988 41748 213994
rect 41696 213930 41748 213936
rect 42812 213489 42840 253399
rect 42984 249824 43036 249830
rect 42984 249766 43036 249772
rect 42996 244274 43024 249766
rect 43626 245712 43682 245721
rect 43626 245647 43682 245656
rect 42996 244246 43300 244274
rect 43074 240952 43130 240961
rect 43074 240887 43130 240896
rect 43088 227730 43116 240887
rect 43272 230450 43300 244246
rect 43442 244080 43498 244089
rect 43442 244015 43498 244024
rect 43260 230444 43312 230450
rect 43260 230386 43312 230392
rect 43076 227724 43128 227730
rect 43076 227666 43128 227672
rect 43456 215294 43484 244015
rect 43640 229401 43668 245647
rect 44008 231033 44036 334591
rect 44822 334112 44878 334121
rect 44822 334047 44878 334056
rect 44270 298072 44326 298081
rect 44270 298007 44326 298016
rect 44284 255241 44312 298007
rect 44546 297120 44602 297129
rect 44546 297055 44602 297064
rect 44270 255232 44326 255241
rect 44270 255167 44326 255176
rect 44178 254824 44234 254833
rect 44178 254759 44234 254768
rect 43994 231024 44050 231033
rect 43994 230959 44050 230968
rect 43626 229392 43682 229401
rect 43626 229327 43682 229336
rect 43456 215266 43576 215294
rect 35806 213480 35862 213489
rect 35806 213415 35862 213424
rect 39578 213480 39634 213489
rect 39578 213415 39634 213424
rect 42798 213480 42854 213489
rect 42798 213415 42854 213424
rect 35820 212702 35848 213415
rect 39592 212702 39620 213415
rect 35808 212696 35860 212702
rect 35808 212638 35860 212644
rect 39580 212696 39632 212702
rect 39580 212638 39632 212644
rect 43548 212534 43576 215266
rect 43456 212506 43576 212534
rect 35806 210216 35862 210225
rect 35806 210151 35862 210160
rect 35820 209982 35848 210151
rect 35808 209976 35860 209982
rect 35808 209918 35860 209924
rect 40132 209976 40184 209982
rect 40132 209918 40184 209924
rect 40144 209409 40172 209918
rect 35622 209400 35678 209409
rect 35622 209335 35678 209344
rect 40130 209400 40186 209409
rect 40130 209335 40186 209344
rect 42982 209400 43038 209409
rect 42982 209335 43038 209344
rect 35636 208690 35664 209335
rect 35806 208992 35862 209001
rect 35806 208927 35862 208936
rect 35624 208684 35676 208690
rect 35624 208626 35676 208632
rect 35820 208418 35848 208927
rect 39764 208684 39816 208690
rect 39764 208626 39816 208632
rect 35808 208412 35860 208418
rect 35808 208354 35860 208360
rect 39776 207777 39804 208626
rect 40040 208412 40092 208418
rect 40040 208354 40092 208360
rect 40052 208185 40080 208354
rect 40038 208176 40094 208185
rect 40038 208111 40094 208120
rect 35806 207768 35862 207777
rect 35806 207703 35862 207712
rect 39762 207768 39818 207777
rect 39762 207703 39818 207712
rect 35820 207194 35848 207703
rect 35808 207188 35860 207194
rect 35808 207130 35860 207136
rect 40132 207188 40184 207194
rect 40132 207130 40184 207136
rect 40144 206961 40172 207130
rect 40130 206952 40186 206961
rect 40130 206887 40186 206896
rect 42798 206952 42854 206961
rect 42798 206887 42854 206896
rect 35806 206136 35862 206145
rect 35806 206071 35862 206080
rect 35820 205834 35848 206071
rect 35808 205828 35860 205834
rect 35808 205770 35860 205776
rect 40224 205828 40276 205834
rect 40224 205770 40276 205776
rect 40236 204921 40264 205770
rect 35622 204912 35678 204921
rect 35622 204847 35678 204856
rect 40222 204912 40278 204921
rect 40222 204847 40278 204856
rect 35636 204338 35664 204847
rect 35806 204504 35862 204513
rect 35806 204439 35808 204448
rect 35860 204439 35862 204448
rect 41512 204468 41564 204474
rect 35808 204410 35860 204416
rect 41512 204410 41564 204416
rect 35624 204332 35676 204338
rect 35624 204274 35676 204280
rect 41524 203697 41552 204410
rect 41696 204332 41748 204338
rect 41696 204274 41748 204280
rect 41708 204105 41736 204274
rect 41694 204096 41750 204105
rect 41694 204031 41750 204040
rect 35806 203688 35862 203697
rect 35806 203623 35862 203632
rect 41510 203688 41566 203697
rect 41510 203623 41566 203632
rect 35820 202910 35848 203623
rect 35808 202904 35860 202910
rect 35808 202846 35860 202852
rect 37924 202904 37976 202910
rect 37924 202846 37976 202852
rect 37936 198801 37964 202846
rect 37922 198792 37978 198801
rect 37922 198727 37978 198736
rect 42430 197296 42486 197305
rect 42430 197231 42486 197240
rect 42444 196670 42472 197231
rect 42182 196642 42472 196670
rect 41970 195800 42026 195809
rect 41970 195735 42026 195744
rect 41984 195432 42012 195735
rect 41786 195256 41842 195265
rect 41786 195191 41842 195200
rect 41800 194820 41828 195191
rect 42246 194984 42302 194993
rect 42246 194919 42302 194928
rect 41786 193488 41842 193497
rect 41786 193423 41842 193432
rect 41800 192984 41828 193423
rect 42076 191593 42104 191760
rect 42062 191584 42118 191593
rect 42062 191519 42118 191528
rect 42168 191026 42196 191148
rect 42260 191026 42288 194919
rect 42168 190998 42288 191026
rect 42430 190496 42486 190505
rect 42182 190454 42430 190482
rect 42430 190431 42486 190440
rect 42182 189910 42472 189938
rect 42444 187649 42472 189910
rect 42430 187640 42486 187649
rect 42430 187575 42486 187584
rect 42432 187468 42484 187474
rect 42182 187431 42432 187459
rect 42432 187410 42484 187416
rect 42430 186824 42486 186833
rect 42182 186782 42430 186810
rect 42430 186759 42486 186768
rect 41786 186416 41842 186425
rect 41786 186351 41842 186360
rect 41800 186184 41828 186351
rect 41786 186008 41842 186017
rect 41786 185943 41842 185952
rect 41800 185605 41828 185943
rect 42168 183530 42196 183765
rect 42156 183524 42208 183530
rect 42156 183466 42208 183472
rect 42812 183274 42840 206887
rect 42996 183530 43024 209335
rect 43258 204912 43314 204921
rect 43258 204847 43314 204856
rect 43272 187474 43300 204847
rect 43260 187468 43312 187474
rect 43260 187410 43312 187416
rect 42984 183524 43036 183530
rect 42984 183466 43036 183472
rect 42536 183246 42840 183274
rect 42536 183138 42564 183246
rect 42182 183110 42564 183138
rect 42430 183016 42486 183025
rect 42430 182951 42486 182960
rect 42444 182491 42472 182951
rect 42182 182463 42472 182491
rect 42076 179353 42104 181900
rect 42062 179344 42118 179353
rect 42062 179279 42118 179288
rect 43456 44198 43484 212506
rect 44192 212129 44220 254759
rect 44560 254425 44588 297055
rect 44546 254416 44602 254425
rect 44546 254351 44602 254360
rect 44546 251152 44602 251161
rect 44546 251087 44602 251096
rect 44362 249112 44418 249121
rect 44362 249047 44418 249056
rect 44376 231849 44404 249047
rect 44362 231840 44418 231849
rect 44362 231775 44418 231784
rect 44560 226681 44588 251087
rect 44546 226672 44602 226681
rect 44546 226607 44602 226616
rect 44178 212120 44234 212129
rect 44178 212055 44234 212064
rect 44362 208448 44418 208457
rect 44362 208383 44418 208392
rect 43810 207768 43866 207777
rect 43810 207703 43866 207712
rect 43626 203688 43682 203697
rect 43626 203623 43682 203632
rect 43640 44334 43668 203623
rect 43824 183025 43852 207703
rect 44178 207224 44234 207233
rect 44178 207159 44234 207168
rect 43994 204096 44050 204105
rect 43994 204031 44050 204040
rect 44008 191593 44036 204031
rect 43994 191584 44050 191593
rect 43994 191519 44050 191528
rect 44192 186833 44220 207159
rect 44376 197305 44404 208383
rect 44546 205592 44602 205601
rect 44546 205527 44602 205536
rect 44362 197296 44418 197305
rect 44362 197231 44418 197240
rect 44560 190505 44588 205527
rect 44546 190496 44602 190505
rect 44546 190431 44602 190440
rect 44178 186824 44234 186833
rect 44178 186759 44234 186768
rect 43810 183016 43866 183025
rect 43810 182951 43866 182960
rect 44836 74534 44864 334047
rect 45480 314673 45508 336767
rect 45664 319161 45692 338399
rect 45650 319152 45706 319161
rect 45650 319087 45706 319096
rect 45466 314664 45522 314673
rect 45466 314599 45522 314608
rect 45006 298888 45062 298897
rect 45006 298823 45062 298832
rect 45020 256057 45048 298823
rect 45190 293584 45246 293593
rect 45190 293519 45246 293528
rect 45204 273057 45232 293519
rect 45190 273048 45246 273057
rect 45190 272983 45246 272992
rect 46216 264246 46244 611623
rect 46938 579184 46994 579193
rect 46938 579119 46994 579128
rect 46952 574054 46980 579119
rect 46940 574048 46992 574054
rect 46940 573990 46992 573996
rect 47582 558512 47638 558521
rect 47582 558447 47638 558456
rect 46386 547496 46442 547505
rect 46386 547431 46442 547440
rect 46400 399498 46428 547431
rect 47596 527134 47624 558447
rect 47584 527128 47636 527134
rect 47584 527070 47636 527076
rect 47766 430536 47822 430545
rect 47766 430471 47822 430480
rect 47582 419928 47638 419937
rect 47582 419863 47638 419872
rect 46388 399492 46440 399498
rect 46388 399434 46440 399440
rect 46386 376136 46442 376145
rect 46386 376071 46442 376080
rect 46400 309126 46428 376071
rect 46938 339280 46994 339289
rect 46938 339215 46994 339224
rect 46952 310185 46980 339215
rect 47122 338056 47178 338065
rect 47122 337991 47178 338000
rect 47136 324329 47164 337991
rect 47122 324320 47178 324329
rect 47122 324255 47178 324264
rect 46938 310176 46994 310185
rect 46938 310111 46994 310120
rect 46388 309120 46440 309126
rect 46388 309062 46440 309068
rect 47596 292194 47624 419863
rect 47780 398818 47808 430471
rect 47768 398812 47820 398818
rect 47768 398754 47820 398760
rect 47766 387696 47822 387705
rect 47766 387631 47822 387640
rect 47780 356046 47808 387631
rect 47768 356040 47820 356046
rect 47768 355982 47820 355988
rect 47952 353456 48004 353462
rect 47952 353398 48004 353404
rect 47768 309120 47820 309126
rect 47768 309062 47820 309068
rect 47584 292188 47636 292194
rect 47584 292130 47636 292136
rect 47780 292058 47808 309062
rect 47768 292052 47820 292058
rect 47768 291994 47820 292000
rect 47582 290728 47638 290737
rect 47582 290663 47638 290672
rect 46388 285728 46440 285734
rect 46388 285670 46440 285676
rect 46204 264240 46256 264246
rect 46204 264182 46256 264188
rect 46400 258097 46428 285670
rect 46386 258088 46442 258097
rect 46386 258023 46442 258032
rect 45006 256048 45062 256057
rect 45006 255983 45062 255992
rect 45650 255640 45706 255649
rect 45650 255575 45706 255584
rect 45006 248704 45062 248713
rect 45006 248639 45062 248648
rect 45020 234569 45048 248639
rect 45006 234560 45062 234569
rect 45006 234495 45062 234504
rect 45664 212945 45692 255575
rect 46202 254008 46258 254017
rect 46202 253943 46258 253952
rect 45926 252784 45982 252793
rect 45926 252719 45982 252728
rect 45940 225729 45968 252719
rect 45926 225720 45982 225729
rect 45926 225655 45982 225664
rect 45650 212936 45706 212945
rect 45650 212871 45706 212880
rect 46216 211313 46244 253943
rect 46938 251968 46994 251977
rect 46938 251903 46994 251912
rect 46386 248296 46442 248305
rect 46386 248231 46442 248240
rect 46400 235929 46428 248231
rect 46386 235920 46442 235929
rect 46386 235855 46442 235864
rect 46952 232257 46980 251903
rect 47122 251560 47178 251569
rect 47122 251495 47178 251504
rect 47136 240145 47164 251495
rect 47122 240136 47178 240145
rect 47122 240071 47178 240080
rect 46938 232248 46994 232257
rect 46938 232183 46994 232192
rect 46202 211304 46258 211313
rect 46202 211239 46258 211248
rect 46938 208856 46994 208865
rect 46938 208791 46994 208800
rect 46202 204368 46258 204377
rect 46202 204303 46258 204312
rect 44836 74506 45508 74534
rect 45480 49026 45508 74506
rect 46216 50386 46244 204303
rect 46952 187649 46980 208791
rect 46938 187640 46994 187649
rect 46938 187575 46994 187584
rect 47596 52018 47624 290663
rect 47768 282940 47820 282946
rect 47768 282882 47820 282888
rect 47780 179353 47808 282882
rect 47964 278186 47992 353398
rect 47952 278180 48004 278186
rect 47952 278122 48004 278128
rect 47766 179344 47822 179353
rect 47766 179279 47822 179288
rect 48976 53106 49004 761874
rect 50160 611312 50212 611318
rect 50160 611254 50212 611260
rect 50172 610162 50200 611254
rect 50160 610156 50212 610162
rect 50160 610098 50212 610104
rect 49146 291000 49202 291009
rect 49146 290935 49202 290944
rect 48964 53100 49016 53106
rect 48964 53042 49016 53048
rect 47584 52012 47636 52018
rect 47584 51954 47636 51960
rect 46204 50380 46256 50386
rect 46204 50322 46256 50328
rect 49160 49162 49188 290935
rect 50356 51882 50384 806074
rect 53104 799060 53156 799066
rect 53104 799002 53156 799008
rect 53116 790770 53144 799002
rect 57244 797700 57296 797706
rect 57244 797642 57296 797648
rect 53104 790764 53156 790770
rect 53104 790706 53156 790712
rect 57256 789206 57284 797642
rect 57244 789200 57296 789206
rect 57244 789142 57296 789148
rect 61396 786185 61424 816954
rect 62948 807968 63000 807974
rect 62948 807910 63000 807916
rect 62672 805996 62724 806002
rect 62672 805938 62724 805944
rect 62212 790764 62264 790770
rect 62212 790706 62264 790712
rect 62224 790537 62252 790706
rect 62210 790528 62266 790537
rect 62210 790463 62266 790472
rect 62120 789200 62172 789206
rect 62118 789168 62120 789177
rect 62172 789168 62174 789177
rect 62118 789103 62174 789112
rect 62118 787400 62174 787409
rect 62118 787335 62174 787344
rect 62132 786690 62160 787335
rect 62120 786684 62172 786690
rect 62120 786626 62172 786632
rect 61382 786176 61438 786185
rect 61382 786111 61438 786120
rect 62120 785188 62172 785194
rect 62120 785130 62172 785136
rect 62132 784961 62160 785130
rect 62118 784952 62174 784961
rect 62118 784887 62174 784896
rect 60004 774240 60056 774246
rect 60004 774182 60056 774188
rect 53104 763224 53156 763230
rect 53104 763166 53156 763172
rect 51724 712156 51776 712162
rect 51724 712098 51776 712104
rect 51736 705158 51764 712098
rect 51724 705152 51776 705158
rect 51724 705094 51776 705100
rect 51722 538248 51778 538257
rect 51722 538183 51778 538192
rect 51736 531282 51764 538183
rect 51724 531276 51776 531282
rect 51724 531218 51776 531224
rect 51446 404968 51502 404977
rect 51446 404903 51502 404912
rect 51460 402966 51488 404903
rect 51448 402960 51500 402966
rect 51448 402902 51500 402908
rect 51080 400240 51132 400246
rect 51080 400182 51132 400188
rect 51092 395729 51120 400182
rect 51078 395720 51134 395729
rect 51078 395655 51134 395664
rect 51078 362264 51134 362273
rect 51078 362199 51134 362208
rect 51092 360194 51120 362199
rect 51080 360188 51132 360194
rect 51080 360130 51132 360136
rect 51722 354376 51778 354385
rect 51722 354311 51778 354320
rect 51080 314764 51132 314770
rect 51080 314706 51132 314712
rect 51092 310457 51120 314706
rect 51078 310448 51134 310457
rect 51078 310383 51134 310392
rect 50528 295384 50580 295390
rect 50528 295326 50580 295332
rect 50540 278769 50568 295326
rect 50526 278760 50582 278769
rect 50526 278695 50582 278704
rect 51736 278322 51764 354311
rect 51908 292596 51960 292602
rect 51908 292538 51960 292544
rect 51724 278316 51776 278322
rect 51724 278258 51776 278264
rect 51920 266257 51948 292538
rect 53116 276729 53144 763166
rect 60016 742422 60044 774182
rect 61384 772880 61436 772886
rect 61384 772822 61436 772828
rect 61396 747318 61424 772822
rect 61384 747312 61436 747318
rect 61384 747254 61436 747260
rect 62120 746564 62172 746570
rect 62120 746506 62172 746512
rect 62132 746201 62160 746506
rect 62118 746192 62174 746201
rect 62118 746127 62174 746136
rect 62118 744152 62174 744161
rect 62118 744087 62174 744096
rect 62132 743918 62160 744087
rect 62120 743912 62172 743918
rect 62120 743854 62172 743860
rect 62120 743776 62172 743782
rect 62118 743744 62120 743753
rect 62172 743744 62174 743753
rect 62118 743679 62174 743688
rect 60004 742416 60056 742422
rect 62120 742416 62172 742422
rect 60004 742358 60056 742364
rect 62118 742384 62120 742393
rect 62172 742384 62174 742393
rect 62118 742319 62174 742328
rect 61384 730312 61436 730318
rect 61384 730254 61436 730260
rect 55864 719024 55916 719030
rect 55864 718966 55916 718972
rect 53286 301336 53342 301345
rect 53286 301271 53342 301280
rect 53300 291174 53328 301271
rect 53472 292188 53524 292194
rect 53472 292130 53524 292136
rect 53288 291168 53340 291174
rect 53288 291110 53340 291116
rect 53288 281580 53340 281586
rect 53288 281522 53340 281528
rect 53102 276720 53158 276729
rect 53102 276655 53158 276664
rect 51906 266248 51962 266257
rect 51906 266183 51962 266192
rect 51724 254584 51776 254590
rect 51724 254526 51776 254532
rect 50526 247480 50582 247489
rect 50526 247415 50582 247424
rect 50540 53242 50568 247415
rect 51736 223553 51764 254526
rect 51722 223544 51778 223553
rect 51722 223479 51778 223488
rect 53300 215121 53328 281522
rect 53484 277914 53512 292130
rect 53656 292052 53708 292058
rect 53656 291994 53708 292000
rect 53668 284986 53696 291994
rect 53656 284980 53708 284986
rect 53656 284922 53708 284928
rect 53472 277908 53524 277914
rect 53472 277850 53524 277856
rect 55876 264217 55904 718966
rect 61396 699689 61424 730254
rect 62120 705152 62172 705158
rect 62120 705094 62172 705100
rect 62132 704449 62160 705094
rect 62118 704440 62174 704449
rect 62118 704375 62174 704384
rect 62120 703792 62172 703798
rect 62120 703734 62172 703740
rect 62132 703361 62160 703734
rect 62118 703352 62174 703361
rect 62118 703287 62174 703296
rect 61382 699680 61438 699689
rect 61382 699615 61438 699624
rect 62212 698284 62264 698290
rect 62212 698226 62264 698232
rect 62224 698057 62252 698226
rect 62210 698048 62266 698057
rect 62210 697983 62266 697992
rect 61384 687540 61436 687546
rect 61384 687482 61436 687488
rect 60004 676252 60056 676258
rect 60004 676194 60056 676200
rect 57244 669384 57296 669390
rect 57244 669326 57296 669332
rect 57256 660958 57284 669326
rect 58624 667956 58676 667962
rect 58624 667898 58676 667904
rect 57244 660952 57296 660958
rect 57244 660894 57296 660900
rect 58636 659598 58664 667898
rect 58624 659592 58676 659598
rect 58624 659534 58676 659540
rect 58624 610156 58676 610162
rect 58624 610098 58676 610104
rect 56048 399492 56100 399498
rect 56048 399434 56100 399440
rect 56060 278458 56088 399434
rect 57244 294092 57296 294098
rect 57244 294034 57296 294040
rect 56324 284980 56376 284986
rect 56324 284922 56376 284928
rect 56048 278452 56100 278458
rect 56048 278394 56100 278400
rect 56336 277778 56364 284922
rect 56324 277772 56376 277778
rect 56324 277714 56376 277720
rect 57256 275913 57284 294034
rect 57242 275904 57298 275913
rect 57242 275839 57298 275848
rect 58636 264382 58664 610098
rect 58808 280220 58860 280226
rect 58808 280162 58860 280168
rect 58624 264376 58676 264382
rect 58624 264318 58676 264324
rect 55862 264208 55918 264217
rect 55862 264143 55918 264152
rect 57244 228404 57296 228410
rect 57244 228346 57296 228352
rect 56508 227044 56560 227050
rect 56508 226986 56560 226992
rect 56520 218210 56548 226986
rect 55680 218204 55732 218210
rect 55680 218146 55732 218152
rect 56508 218204 56560 218210
rect 56508 218146 56560 218152
rect 55692 217138 55720 218146
rect 57256 218074 57284 228346
rect 57428 218204 57480 218210
rect 57428 218146 57480 218152
rect 56508 218068 56560 218074
rect 56508 218010 56560 218016
rect 57244 218068 57296 218074
rect 57244 218010 57296 218016
rect 56520 217138 56548 218010
rect 57440 217274 57468 218146
rect 58164 218068 58216 218074
rect 58164 218010 58216 218016
rect 55646 217110 55720 217138
rect 56474 217110 56548 217138
rect 57302 217246 57468 217274
rect 55646 216988 55674 217110
rect 56474 216988 56502 217110
rect 57302 216988 57330 217246
rect 58176 217138 58204 218010
rect 58820 217977 58848 280162
rect 60016 278089 60044 676194
rect 61396 656577 61424 687482
rect 62120 660952 62172 660958
rect 62118 660920 62120 660929
rect 62172 660920 62174 660929
rect 62118 660855 62174 660864
rect 62120 659592 62172 659598
rect 62118 659560 62120 659569
rect 62172 659560 62174 659569
rect 62118 659495 62174 659504
rect 62118 658336 62174 658345
rect 62118 658271 62174 658280
rect 62132 657558 62160 658271
rect 62120 657552 62172 657558
rect 62120 657494 62172 657500
rect 61382 656568 61438 656577
rect 61382 656503 61438 656512
rect 62120 655512 62172 655518
rect 62120 655454 62172 655460
rect 62132 655353 62160 655454
rect 62118 655344 62174 655353
rect 62118 655279 62174 655288
rect 61384 643136 61436 643142
rect 61384 643078 61436 643084
rect 60188 633480 60240 633486
rect 60188 633422 60240 633428
rect 60200 278769 60228 633422
rect 61396 613873 61424 643078
rect 62120 616820 62172 616826
rect 62120 616762 62172 616768
rect 62132 616593 62160 616762
rect 62118 616584 62174 616593
rect 62118 616519 62174 616528
rect 62118 614680 62174 614689
rect 62118 614615 62174 614624
rect 62132 614174 62160 614615
rect 62120 614168 62172 614174
rect 62120 614110 62172 614116
rect 61382 613864 61438 613873
rect 61382 613799 61438 613808
rect 62120 613420 62172 613426
rect 62120 613362 62172 613368
rect 62132 612649 62160 613362
rect 62118 612640 62174 612649
rect 62118 612575 62174 612584
rect 61384 610020 61436 610026
rect 61384 609962 61436 609968
rect 60370 319424 60426 319433
rect 60370 319359 60426 319368
rect 60384 315994 60412 319359
rect 60372 315988 60424 315994
rect 60372 315930 60424 315936
rect 60372 284436 60424 284442
rect 60372 284378 60424 284384
rect 60186 278760 60242 278769
rect 60186 278695 60242 278704
rect 60002 278080 60058 278089
rect 60002 278015 60058 278024
rect 60384 256737 60412 284378
rect 60370 256728 60426 256737
rect 60370 256663 60426 256672
rect 61396 231334 61424 609962
rect 62486 594144 62542 594153
rect 62486 594079 62542 594088
rect 62302 590064 62358 590073
rect 62302 589999 62358 590008
rect 62120 575476 62172 575482
rect 62120 575418 62172 575424
rect 62132 574841 62160 575418
rect 62118 574832 62174 574841
rect 62118 574767 62174 574776
rect 62120 574048 62172 574054
rect 62120 573990 62172 573996
rect 62132 573617 62160 573990
rect 62118 573608 62174 573617
rect 62118 573543 62174 573552
rect 62316 569945 62344 589999
rect 62302 569936 62358 569945
rect 62302 569871 62358 569880
rect 62500 568585 62528 594079
rect 62486 568576 62542 568585
rect 62486 568511 62542 568520
rect 62486 550216 62542 550225
rect 62486 550151 62542 550160
rect 62120 532024 62172 532030
rect 62120 531966 62172 531972
rect 62132 531185 62160 531966
rect 62304 531276 62356 531282
rect 62304 531218 62356 531224
rect 62118 531176 62174 531185
rect 62118 531111 62174 531120
rect 62316 530641 62344 531218
rect 62302 530632 62358 530641
rect 62302 530567 62358 530576
rect 62120 528624 62172 528630
rect 62118 528592 62120 528601
rect 62172 528592 62174 528601
rect 62118 528527 62174 528536
rect 62120 527128 62172 527134
rect 62118 527096 62120 527105
rect 62172 527096 62174 527105
rect 62118 527031 62174 527040
rect 62500 525745 62528 550151
rect 62486 525736 62542 525745
rect 62486 525671 62542 525680
rect 62120 404320 62172 404326
rect 62120 404262 62172 404268
rect 62132 404161 62160 404262
rect 62118 404152 62174 404161
rect 62118 404087 62174 404096
rect 62120 402960 62172 402966
rect 62120 402902 62172 402908
rect 62132 402665 62160 402902
rect 62118 402656 62174 402665
rect 62118 402591 62174 402600
rect 62118 400752 62174 400761
rect 62118 400687 62174 400696
rect 62132 400246 62160 400687
rect 62120 400240 62172 400246
rect 62120 400182 62172 400188
rect 62120 400104 62172 400110
rect 62120 400046 62172 400052
rect 62132 399401 62160 400046
rect 62118 399392 62174 399401
rect 62118 399327 62174 399336
rect 62120 398812 62172 398818
rect 62120 398754 62172 398760
rect 62132 398313 62160 398754
rect 62118 398304 62174 398313
rect 62118 398239 62174 398248
rect 62486 381576 62542 381585
rect 62486 381511 62542 381520
rect 62120 361548 62172 361554
rect 62120 361490 62172 361496
rect 62132 360913 62160 361490
rect 62118 360904 62174 360913
rect 62118 360839 62174 360848
rect 62120 360188 62172 360194
rect 62120 360130 62172 360136
rect 62132 359825 62160 360130
rect 62118 359816 62174 359825
rect 62118 359751 62174 359760
rect 62118 357776 62174 357785
rect 62118 357711 62174 357720
rect 62132 357474 62160 357711
rect 62120 357468 62172 357474
rect 62120 357410 62172 357416
rect 62120 356040 62172 356046
rect 62118 356008 62120 356017
rect 62172 356008 62174 356017
rect 62118 355943 62174 355952
rect 62500 354521 62528 381511
rect 62486 354512 62542 354521
rect 62486 354447 62542 354456
rect 62394 341728 62450 341737
rect 62394 341663 62450 341672
rect 62212 341420 62264 341426
rect 62212 341362 62264 341368
rect 62224 325694 62252 341362
rect 62408 335354 62436 341663
rect 62316 335326 62436 335354
rect 62316 330562 62344 335326
rect 62486 332616 62542 332625
rect 62486 332551 62542 332560
rect 62316 330534 62436 330562
rect 62224 325666 62344 325694
rect 62026 320784 62082 320793
rect 62026 320719 62082 320728
rect 62040 317393 62068 320719
rect 62026 317384 62082 317393
rect 62026 317319 62082 317328
rect 62118 316024 62174 316033
rect 62118 315959 62120 315968
rect 62172 315959 62174 315968
rect 62120 315930 62172 315936
rect 62118 314800 62174 314809
rect 62118 314735 62120 314744
rect 62172 314735 62174 314744
rect 62120 314706 62172 314712
rect 62316 314129 62344 325666
rect 62408 316034 62436 330534
rect 62500 325694 62528 332551
rect 62500 325666 62620 325694
rect 62408 316006 62528 316034
rect 62302 314120 62358 314129
rect 62302 314055 62358 314064
rect 62500 313562 62528 316006
rect 62408 313534 62528 313562
rect 62408 313041 62436 313534
rect 62394 313032 62450 313041
rect 62394 312967 62450 312976
rect 62394 297392 62450 297401
rect 62394 297327 62450 297336
rect 62118 295760 62174 295769
rect 62118 295695 62174 295704
rect 62132 295390 62160 295695
rect 62120 295384 62172 295390
rect 62120 295326 62172 295332
rect 62118 294128 62174 294137
rect 62118 294063 62120 294072
rect 62172 294063 62174 294072
rect 62120 294034 62172 294040
rect 62118 292768 62174 292777
rect 62118 292703 62174 292712
rect 62132 292602 62160 292703
rect 62120 292596 62172 292602
rect 62120 292538 62172 292544
rect 62408 292505 62436 297327
rect 62394 292496 62450 292505
rect 62394 292431 62450 292440
rect 62120 291168 62172 291174
rect 62120 291110 62172 291116
rect 62132 291009 62160 291110
rect 62118 291000 62174 291009
rect 62118 290935 62174 290944
rect 62394 288552 62450 288561
rect 62394 288487 62450 288496
rect 62408 287424 62436 288487
rect 62408 287396 62528 287424
rect 62302 287192 62358 287201
rect 62302 287127 62358 287136
rect 62118 284472 62174 284481
rect 62118 284407 62120 284416
rect 62172 284407 62174 284416
rect 62120 284378 62172 284384
rect 62118 283248 62174 283257
rect 62118 283183 62174 283192
rect 62132 282946 62160 283183
rect 62120 282940 62172 282946
rect 62120 282882 62172 282888
rect 62118 282160 62174 282169
rect 62118 282095 62174 282104
rect 62132 281586 62160 282095
rect 62120 281580 62172 281586
rect 62120 281522 62172 281528
rect 62118 280392 62174 280401
rect 62118 280327 62174 280336
rect 62132 280226 62160 280327
rect 62120 280220 62172 280226
rect 62120 280162 62172 280168
rect 62316 277394 62344 287127
rect 62500 287054 62528 287396
rect 62224 277366 62344 277394
rect 62408 287026 62528 287054
rect 62224 273873 62252 277366
rect 62210 273864 62266 273873
rect 62210 273799 62266 273808
rect 62408 254590 62436 287026
rect 62592 278730 62620 325666
rect 62684 287054 62712 805938
rect 62960 787137 62988 807910
rect 653404 790832 653456 790838
rect 653404 790774 653456 790780
rect 62946 787128 63002 787137
rect 62946 787063 63002 787072
rect 651470 778424 651526 778433
rect 651470 778359 651526 778368
rect 651484 777646 651512 778359
rect 651472 777640 651524 777646
rect 651472 777582 651524 777588
rect 652022 777064 652078 777073
rect 652022 776999 652078 777008
rect 651470 776112 651526 776121
rect 651470 776047 651526 776056
rect 651484 775606 651512 776047
rect 651472 775600 651524 775606
rect 651472 775542 651524 775548
rect 651380 775328 651432 775334
rect 651378 775296 651380 775305
rect 651432 775296 651434 775305
rect 651378 775231 651434 775240
rect 651470 774208 651526 774217
rect 651470 774143 651472 774152
rect 651524 774143 651526 774152
rect 651472 774114 651524 774120
rect 651472 773832 651524 773838
rect 651472 773774 651524 773780
rect 651484 773401 651512 773774
rect 651470 773392 651526 773401
rect 651470 773327 651526 773336
rect 62948 755540 63000 755546
rect 62948 755482 63000 755488
rect 62960 747697 62988 755482
rect 62946 747688 63002 747697
rect 62946 747623 63002 747632
rect 63040 747312 63092 747318
rect 63040 747254 63092 747260
rect 63052 741849 63080 747254
rect 63038 741840 63094 741849
rect 63038 741775 63094 741784
rect 652036 736914 652064 776999
rect 653416 775334 653444 790774
rect 670608 784304 670660 784310
rect 670608 784246 670660 784252
rect 669228 784168 669280 784174
rect 669228 784110 669280 784116
rect 669044 782536 669096 782542
rect 669044 782478 669096 782484
rect 655520 781108 655572 781114
rect 655520 781050 655572 781056
rect 655060 778388 655112 778394
rect 655060 778330 655112 778336
rect 653404 775328 653456 775334
rect 653404 775270 653456 775276
rect 655072 773838 655100 778330
rect 655532 774178 655560 781050
rect 660304 777640 660356 777646
rect 660304 777582 660356 777588
rect 655520 774172 655572 774178
rect 655520 774114 655572 774120
rect 655060 773832 655112 773838
rect 655060 773774 655112 773780
rect 653404 746632 653456 746638
rect 653404 746574 653456 746580
rect 652024 736908 652076 736914
rect 652024 736850 652076 736856
rect 651470 734224 651526 734233
rect 651470 734159 651526 734168
rect 651484 733446 651512 734159
rect 651472 733440 651524 733446
rect 651472 733382 651524 733388
rect 652666 732864 652722 732873
rect 652666 732799 652722 732808
rect 651470 731776 651526 731785
rect 651470 731711 651526 731720
rect 651484 731474 651512 731711
rect 651472 731468 651524 731474
rect 651472 731410 651524 731416
rect 651380 731128 651432 731134
rect 651378 731096 651380 731105
rect 651432 731096 651434 731105
rect 651378 731031 651434 731040
rect 652680 730726 652708 732799
rect 653416 731134 653444 746574
rect 656164 736908 656216 736914
rect 656164 736850 656216 736856
rect 654784 734188 654836 734194
rect 654784 734130 654836 734136
rect 653404 731128 653456 731134
rect 653404 731070 653456 731076
rect 652668 730720 652720 730726
rect 652668 730662 652720 730668
rect 651472 730040 651524 730046
rect 651472 729982 651524 729988
rect 651484 729881 651512 729982
rect 651470 729872 651526 729881
rect 651470 729807 651526 729816
rect 62948 729360 63000 729366
rect 62948 729302 63000 729308
rect 62960 712094 62988 729302
rect 654796 728550 654824 734130
rect 651472 728544 651524 728550
rect 651470 728512 651472 728521
rect 654784 728544 654836 728550
rect 651524 728512 651526 728521
rect 654784 728486 654836 728492
rect 651470 728447 651526 728456
rect 656176 716310 656204 736850
rect 657544 735616 657596 735622
rect 657544 735558 657596 735564
rect 657556 730046 657584 735558
rect 658924 731468 658976 731474
rect 658924 731410 658976 731416
rect 657544 730040 657596 730046
rect 657544 729982 657596 729988
rect 656164 716304 656216 716310
rect 656164 716246 656216 716252
rect 62960 712066 63172 712094
rect 62946 701312 63002 701321
rect 62946 701247 63002 701256
rect 62960 701078 62988 701247
rect 62948 701072 63000 701078
rect 62948 701014 63000 701020
rect 63144 700913 63172 712066
rect 654784 701208 654836 701214
rect 654784 701150 654836 701156
rect 63130 700904 63186 700913
rect 63130 700839 63186 700848
rect 651470 689480 651526 689489
rect 651470 689415 651526 689424
rect 651484 688702 651512 689415
rect 652760 688832 652812 688838
rect 651654 688800 651710 688809
rect 652760 688774 652812 688780
rect 651654 688735 651710 688744
rect 651472 688696 651524 688702
rect 651472 688638 651524 688644
rect 651470 687440 651526 687449
rect 651470 687375 651526 687384
rect 651484 687274 651512 687375
rect 651472 687268 651524 687274
rect 651472 687210 651524 687216
rect 651472 687064 651524 687070
rect 651472 687006 651524 687012
rect 651484 686769 651512 687006
rect 651470 686760 651526 686769
rect 651470 686695 651526 686704
rect 651668 686526 651696 688735
rect 62948 686520 63000 686526
rect 62948 686462 63000 686468
rect 651656 686520 651708 686526
rect 651656 686462 651708 686468
rect 62960 657665 62988 686462
rect 651472 685568 651524 685574
rect 651472 685510 651524 685516
rect 651484 685273 651512 685510
rect 651470 685264 651526 685273
rect 651470 685199 651526 685208
rect 652574 684448 652630 684457
rect 652772 684434 652800 688774
rect 654796 687070 654824 701150
rect 656532 690260 656584 690266
rect 656532 690202 656584 690208
rect 654784 687064 654836 687070
rect 654784 687006 654836 687012
rect 656544 685574 656572 690202
rect 657544 688696 657596 688702
rect 657544 688638 657596 688644
rect 656532 685568 656584 685574
rect 656532 685510 656584 685516
rect 652630 684406 652800 684434
rect 652574 684383 652630 684392
rect 62946 657656 63002 657665
rect 62946 657591 63002 657600
rect 653404 655580 653456 655586
rect 653404 655522 653456 655528
rect 651470 643240 651526 643249
rect 651470 643175 651526 643184
rect 651484 642394 651512 643175
rect 62948 642388 63000 642394
rect 62948 642330 63000 642336
rect 651472 642388 651524 642394
rect 651472 642330 651524 642336
rect 62960 612105 62988 642330
rect 652022 641880 652078 641889
rect 652022 641815 652078 641824
rect 651470 640792 651526 640801
rect 651470 640727 651526 640736
rect 651484 640354 651512 640727
rect 651472 640348 651524 640354
rect 651472 640290 651524 640296
rect 651380 640144 651432 640150
rect 651378 640112 651380 640121
rect 651432 640112 651434 640121
rect 651378 640047 651434 640056
rect 651656 638920 651708 638926
rect 651656 638862 651708 638868
rect 651472 638784 651524 638790
rect 651472 638726 651524 638732
rect 651484 638625 651512 638726
rect 651470 638616 651526 638625
rect 651470 638551 651526 638560
rect 651668 638217 651696 638862
rect 651654 638208 651710 638217
rect 651654 638143 651710 638152
rect 652036 634098 652064 641815
rect 653416 640150 653444 655522
rect 655520 645924 655572 645930
rect 655520 645866 655572 645872
rect 655336 643136 655388 643142
rect 655336 643078 655388 643084
rect 653404 640144 653456 640150
rect 653404 640086 653456 640092
rect 655348 638926 655376 643078
rect 655336 638920 655388 638926
rect 655336 638862 655388 638868
rect 655532 638790 655560 645866
rect 655520 638784 655572 638790
rect 655520 638726 655572 638732
rect 652024 634092 652076 634098
rect 652024 634034 652076 634040
rect 63132 625864 63184 625870
rect 63132 625806 63184 625812
rect 63144 618089 63172 625806
rect 657556 625190 657584 688638
rect 658936 669526 658964 731410
rect 660316 715018 660344 777582
rect 668584 733440 668636 733446
rect 668584 733382 668636 733388
rect 661684 730720 661736 730726
rect 661684 730662 661736 730668
rect 660304 715012 660356 715018
rect 660304 714954 660356 714960
rect 661696 670750 661724 730662
rect 667848 705220 667900 705226
rect 667848 705162 667900 705168
rect 667020 703860 667072 703866
rect 667020 703802 667072 703808
rect 661684 670744 661736 670750
rect 661684 670686 661736 670692
rect 658924 669520 658976 669526
rect 658924 669462 658976 669468
rect 658924 642388 658976 642394
rect 658924 642330 658976 642336
rect 657544 625184 657596 625190
rect 657544 625126 657596 625132
rect 63130 618080 63186 618089
rect 63130 618015 63186 618024
rect 62946 612096 63002 612105
rect 62946 612031 63002 612040
rect 64142 611416 64198 611425
rect 64142 611351 64198 611360
rect 653404 611380 653456 611386
rect 63406 595776 63462 595785
rect 63406 595711 63462 595720
rect 63038 590744 63094 590753
rect 63038 590679 63094 590688
rect 62854 585712 62910 585721
rect 62854 585647 62910 585656
rect 62684 287026 62804 287054
rect 62580 278724 62632 278730
rect 62580 278666 62632 278672
rect 62776 277394 62804 287026
rect 62684 277366 62804 277394
rect 62396 254584 62448 254590
rect 62396 254526 62448 254532
rect 61384 231328 61436 231334
rect 61384 231270 61436 231276
rect 61384 228540 61436 228546
rect 61384 228482 61436 228488
rect 60648 227588 60700 227594
rect 60648 227530 60700 227536
rect 59360 221604 59412 221610
rect 59360 221546 59412 221552
rect 58992 218748 59044 218754
rect 58992 218690 59044 218696
rect 58806 217968 58862 217977
rect 58806 217903 58862 217912
rect 59004 217138 59032 218690
rect 59372 218074 59400 221546
rect 59820 218884 59872 218890
rect 59820 218826 59872 218832
rect 59360 218068 59412 218074
rect 59360 218010 59412 218016
rect 59832 217138 59860 218826
rect 60660 217274 60688 227530
rect 61396 218210 61424 228482
rect 62684 224233 62712 277366
rect 62670 224224 62726 224233
rect 62670 224159 62726 224168
rect 62868 223553 62896 585647
rect 63052 287054 63080 590679
rect 63420 571169 63448 595711
rect 63406 571160 63462 571169
rect 63406 571095 63462 571104
rect 63222 556744 63278 556753
rect 63222 556679 63278 556688
rect 63236 528057 63264 556679
rect 63222 528048 63278 528057
rect 63222 527983 63278 527992
rect 63314 427136 63370 427145
rect 63314 427071 63370 427080
rect 63328 400217 63356 427071
rect 63314 400208 63370 400217
rect 63314 400143 63370 400152
rect 63222 385928 63278 385937
rect 63222 385863 63278 385872
rect 63236 357377 63264 385863
rect 63222 357368 63278 357377
rect 63222 357303 63278 357312
rect 63314 341456 63370 341465
rect 63314 341391 63370 341400
rect 63328 311817 63356 341391
rect 63314 311808 63370 311817
rect 63314 311743 63370 311752
rect 63314 299568 63370 299577
rect 63314 299503 63370 299512
rect 63328 289785 63356 299503
rect 63314 289776 63370 289785
rect 63314 289711 63370 289720
rect 63052 287026 63448 287054
rect 63038 285968 63094 285977
rect 63038 285903 63094 285912
rect 63052 285734 63080 285903
rect 63040 285728 63092 285734
rect 63040 285670 63092 285676
rect 63222 280936 63278 280945
rect 63222 280871 63278 280880
rect 63040 227180 63092 227186
rect 63040 227122 63092 227128
rect 62854 223544 62910 223553
rect 62854 223479 62910 223488
rect 62764 222896 62816 222902
rect 62764 222838 62816 222844
rect 62304 219020 62356 219026
rect 62304 218962 62356 218968
rect 61384 218204 61436 218210
rect 61384 218146 61436 218152
rect 61476 218068 61528 218074
rect 61476 218010 61528 218016
rect 58130 217110 58204 217138
rect 58958 217110 59032 217138
rect 59786 217110 59860 217138
rect 60614 217246 60688 217274
rect 58130 216988 58158 217110
rect 58958 216988 58986 217110
rect 59786 216988 59814 217110
rect 60614 216988 60642 217246
rect 61488 217138 61516 218010
rect 62316 217138 62344 218962
rect 62776 218074 62804 222838
rect 63052 219434 63080 227122
rect 63236 224505 63264 280871
rect 63420 278594 63448 287026
rect 63408 278588 63460 278594
rect 63408 278530 63460 278536
rect 64156 278050 64184 611351
rect 653404 611322 653456 611328
rect 651470 597952 651526 597961
rect 651470 597887 651526 597896
rect 651484 597582 651512 597887
rect 651472 597576 651524 597582
rect 651472 597518 651524 597524
rect 651470 596728 651526 596737
rect 651470 596663 651526 596672
rect 651484 596222 651512 596663
rect 651472 596216 651524 596222
rect 651472 596158 651524 596164
rect 653416 595542 653444 611322
rect 657544 600500 657596 600506
rect 657544 600442 657596 600448
rect 654784 599004 654836 599010
rect 654784 598946 654836 598952
rect 651656 595536 651708 595542
rect 651656 595478 651708 595484
rect 653404 595536 653456 595542
rect 653404 595478 653456 595484
rect 651470 595368 651526 595377
rect 651470 595303 651526 595312
rect 651484 594862 651512 595303
rect 651668 595105 651696 595478
rect 651654 595096 651710 595105
rect 651654 595031 651710 595040
rect 651472 594856 651524 594862
rect 651472 594798 651524 594804
rect 651472 594720 651524 594726
rect 651472 594662 651524 594668
rect 651484 594153 651512 594662
rect 651470 594144 651526 594153
rect 651470 594079 651526 594088
rect 654796 593298 654824 598946
rect 657556 594726 657584 600442
rect 657544 594720 657596 594726
rect 657544 594662 657596 594668
rect 651472 593292 651524 593298
rect 651472 593234 651524 593240
rect 654784 593292 654836 593298
rect 654784 593234 654836 593240
rect 651484 592929 651512 593234
rect 651470 592920 651526 592929
rect 651470 592855 651526 592864
rect 658936 579698 658964 642330
rect 660304 634092 660356 634098
rect 660304 634034 660356 634040
rect 660316 581058 660344 634034
rect 664444 596216 664496 596222
rect 664444 596158 664496 596164
rect 661684 594856 661736 594862
rect 661684 594798 661736 594804
rect 660304 581052 660356 581058
rect 660304 580994 660356 581000
rect 658924 579692 658976 579698
rect 658924 579634 658976 579640
rect 653404 565888 653456 565894
rect 653404 565830 653456 565836
rect 651470 553480 651526 553489
rect 651470 553415 651526 553424
rect 651484 552702 651512 553415
rect 651472 552696 651524 552702
rect 651472 552638 651524 552644
rect 651654 552120 651710 552129
rect 651654 552055 651710 552064
rect 651470 551168 651526 551177
rect 651470 551103 651526 551112
rect 651484 550662 651512 551103
rect 651472 550656 651524 550662
rect 651472 550598 651524 550604
rect 651380 550384 651432 550390
rect 651378 550352 651380 550361
rect 651432 550352 651434 550361
rect 651378 550287 651434 550296
rect 651668 549914 651696 552055
rect 653416 550390 653444 565830
rect 657820 554804 657872 554810
rect 657820 554746 657872 554752
rect 655152 553444 655204 553450
rect 655152 553386 655204 553392
rect 653404 550384 653456 550390
rect 653404 550326 653456 550332
rect 651656 549908 651708 549914
rect 651656 549850 651708 549856
rect 651470 549264 651526 549273
rect 651470 549199 651472 549208
rect 651524 549199 651526 549208
rect 651472 549170 651524 549176
rect 655164 548826 655192 553386
rect 657832 549234 657860 554746
rect 660304 550656 660356 550662
rect 660304 550598 660356 550604
rect 657820 549228 657872 549234
rect 657820 549170 657872 549176
rect 651472 548820 651524 548826
rect 651472 548762 651524 548768
rect 655152 548820 655204 548826
rect 655152 548762 655204 548768
rect 651484 548457 651512 548762
rect 651470 548448 651526 548457
rect 651470 548383 651526 548392
rect 658464 518220 658516 518226
rect 658464 518162 658516 518168
rect 658476 509930 658504 518162
rect 650644 509924 650696 509930
rect 650644 509866 650696 509872
rect 658464 509924 658516 509930
rect 658464 509866 658516 509872
rect 64326 353424 64382 353433
rect 64326 353359 64382 353368
rect 64144 278044 64196 278050
rect 64144 277986 64196 277992
rect 64340 277642 64368 353359
rect 635004 278316 635056 278322
rect 635004 278258 635056 278264
rect 637592 278310 637974 278338
rect 64328 277636 64380 277642
rect 64328 277578 64380 277584
rect 65904 272542 65932 278052
rect 67100 274242 67128 278052
rect 67088 274236 67140 274242
rect 67088 274178 67140 274184
rect 65892 272536 65944 272542
rect 65892 272478 65944 272484
rect 68204 271182 68232 278052
rect 69400 273970 69428 278052
rect 69664 277908 69716 277914
rect 69664 277850 69716 277856
rect 69676 277506 69704 277850
rect 69664 277500 69716 277506
rect 69664 277442 69716 277448
rect 69388 273964 69440 273970
rect 69388 273906 69440 273912
rect 68192 271176 68244 271182
rect 68192 271118 68244 271124
rect 70596 269822 70624 278052
rect 71792 275330 71820 278052
rect 71780 275324 71832 275330
rect 71780 275266 71832 275272
rect 72988 272678 73016 278052
rect 74184 274718 74212 278052
rect 74172 274712 74224 274718
rect 74172 274654 74224 274660
rect 72976 272672 73028 272678
rect 72976 272614 73028 272620
rect 75380 271454 75408 278052
rect 76484 275602 76512 278052
rect 76472 275596 76524 275602
rect 76472 275538 76524 275544
rect 76840 274712 76892 274718
rect 76840 274654 76892 274660
rect 75368 271448 75420 271454
rect 75368 271390 75420 271396
rect 76852 271318 76880 274654
rect 77680 274106 77708 278052
rect 77668 274100 77720 274106
rect 77668 274042 77720 274048
rect 76840 271312 76892 271318
rect 76840 271254 76892 271260
rect 78876 270366 78904 278052
rect 78864 270360 78916 270366
rect 78864 270302 78916 270308
rect 80072 269822 80100 278052
rect 81268 274990 81296 278052
rect 81256 274984 81308 274990
rect 81256 274926 81308 274932
rect 82464 272814 82492 278052
rect 83674 278038 84148 278066
rect 84778 278038 85528 278066
rect 82452 272808 82504 272814
rect 82452 272750 82504 272756
rect 84120 270502 84148 278038
rect 84108 270496 84160 270502
rect 84108 270438 84160 270444
rect 85500 269958 85528 278038
rect 85960 274718 85988 278052
rect 86224 275596 86276 275602
rect 86224 275538 86276 275544
rect 85948 274712 86000 274718
rect 85948 274654 86000 274660
rect 85488 269952 85540 269958
rect 85488 269894 85540 269900
rect 70584 269816 70636 269822
rect 70584 269758 70636 269764
rect 79324 269816 79376 269822
rect 79324 269758 79376 269764
rect 80060 269816 80112 269822
rect 80060 269758 80112 269764
rect 79336 267034 79364 269758
rect 86236 267442 86264 275538
rect 87156 271590 87184 278052
rect 88352 273834 88380 278052
rect 89562 278038 89668 278066
rect 88340 273828 88392 273834
rect 88340 273770 88392 273776
rect 87144 271584 87196 271590
rect 87144 271526 87196 271532
rect 89640 270094 89668 278038
rect 90744 275602 90772 278052
rect 91862 278038 92428 278066
rect 90732 275596 90784 275602
rect 90732 275538 90784 275544
rect 90364 274712 90416 274718
rect 90364 274654 90416 274660
rect 89628 270088 89680 270094
rect 89628 270030 89680 270036
rect 86224 267436 86276 267442
rect 86224 267378 86276 267384
rect 90376 267170 90404 274654
rect 92400 268394 92428 278038
rect 93044 275738 93072 278052
rect 93032 275732 93084 275738
rect 93032 275674 93084 275680
rect 94240 272950 94268 278052
rect 95436 274378 95464 278052
rect 96632 275194 96660 278052
rect 96620 275188 96672 275194
rect 96620 275130 96672 275136
rect 95424 274372 95476 274378
rect 95424 274314 95476 274320
rect 94228 272944 94280 272950
rect 94228 272886 94280 272892
rect 97828 271726 97856 278052
rect 99038 278038 99328 278066
rect 97816 271720 97868 271726
rect 97816 271662 97868 271668
rect 99300 268530 99328 278038
rect 100128 275466 100156 278052
rect 100116 275460 100168 275466
rect 100116 275402 100168 275408
rect 101324 274514 101352 278052
rect 101312 274508 101364 274514
rect 101312 274450 101364 274456
rect 102520 273086 102548 278052
rect 103716 274718 103744 278052
rect 104912 277394 104940 278052
rect 104912 277366 105032 277394
rect 103704 274712 103756 274718
rect 103704 274654 103756 274660
rect 104808 274712 104860 274718
rect 104808 274654 104860 274660
rect 102508 273080 102560 273086
rect 102508 273022 102560 273028
rect 99288 268524 99340 268530
rect 99288 268466 99340 268472
rect 92388 268388 92440 268394
rect 92388 268330 92440 268336
rect 104820 267306 104848 274654
rect 105004 268666 105032 277366
rect 106016 271862 106044 278052
rect 107212 276010 107240 278052
rect 107200 276004 107252 276010
rect 107200 275946 107252 275952
rect 108408 273222 108436 278052
rect 109618 278038 110368 278066
rect 108396 273216 108448 273222
rect 108396 273158 108448 273164
rect 106004 271856 106056 271862
rect 106004 271798 106056 271804
rect 110340 268802 110368 278038
rect 110800 274718 110828 278052
rect 110788 274712 110840 274718
rect 110788 274654 110840 274660
rect 111708 274712 111760 274718
rect 111708 274654 111760 274660
rect 110328 268796 110380 268802
rect 110328 268738 110380 268744
rect 104992 268660 105044 268666
rect 104992 268602 105044 268608
rect 111720 267578 111748 274654
rect 111996 270230 112024 278052
rect 113206 278038 113496 278066
rect 113468 271046 113496 278038
rect 114388 274650 114416 278052
rect 115506 278038 115888 278066
rect 114376 274644 114428 274650
rect 114376 274586 114428 274592
rect 113456 271040 113508 271046
rect 113456 270982 113508 270988
rect 111984 270224 112036 270230
rect 111984 270166 112036 270172
rect 115860 268938 115888 278038
rect 116688 272406 116716 278052
rect 117898 278038 118648 278066
rect 116676 272400 116728 272406
rect 116676 272342 116728 272348
rect 118620 269074 118648 278038
rect 119080 273698 119108 278052
rect 120276 273834 120304 278052
rect 119344 273828 119396 273834
rect 119344 273770 119396 273776
rect 120264 273828 120316 273834
rect 120264 273770 120316 273776
rect 119068 273692 119120 273698
rect 119068 273634 119120 273640
rect 118608 269068 118660 269074
rect 118608 269010 118660 269016
rect 115848 268932 115900 268938
rect 115848 268874 115900 268880
rect 119356 267714 119384 273770
rect 121472 270638 121500 278052
rect 122590 278038 122788 278066
rect 121460 270632 121512 270638
rect 121460 270574 121512 270580
rect 122760 269686 122788 278038
rect 123772 270910 123800 278052
rect 124968 271998 124996 278052
rect 126178 278038 126928 278066
rect 124956 271992 125008 271998
rect 124956 271934 125008 271940
rect 123760 270904 123812 270910
rect 123760 270846 123812 270852
rect 122748 269680 122800 269686
rect 122748 269622 122800 269628
rect 126900 269414 126928 278038
rect 127360 272270 127388 278052
rect 128556 274786 128584 278052
rect 128544 274780 128596 274786
rect 128544 274722 128596 274728
rect 127348 272264 127400 272270
rect 127348 272206 127400 272212
rect 129660 269550 129688 278052
rect 130856 274242 130884 278052
rect 130384 274236 130436 274242
rect 130384 274178 130436 274184
rect 130844 274236 130896 274242
rect 130844 274178 130896 274184
rect 129648 269544 129700 269550
rect 129648 269486 129700 269492
rect 126888 269408 126940 269414
rect 126888 269350 126940 269356
rect 119344 267708 119396 267714
rect 119344 267650 119396 267656
rect 111708 267572 111760 267578
rect 111708 267514 111760 267520
rect 104808 267300 104860 267306
rect 104808 267242 104860 267248
rect 90364 267164 90416 267170
rect 90364 267106 90416 267112
rect 79324 267028 79376 267034
rect 79324 266970 79376 266976
rect 130396 266626 130424 274178
rect 132052 273562 132080 278052
rect 133262 278038 133828 278066
rect 132040 273556 132092 273562
rect 132040 273498 132092 273504
rect 133800 270366 133828 278038
rect 134444 270774 134472 278052
rect 134432 270768 134484 270774
rect 134432 270710 134484 270716
rect 132500 270360 132552 270366
rect 132500 270302 132552 270308
rect 133788 270360 133840 270366
rect 133788 270302 133840 270308
rect 130384 266620 130436 266626
rect 130384 266562 130436 266568
rect 132512 266490 132540 270302
rect 135640 268258 135668 278052
rect 136836 275058 136864 278052
rect 136824 275052 136876 275058
rect 136824 274994 136876 275000
rect 137652 275052 137704 275058
rect 137652 274994 137704 275000
rect 136824 272536 136876 272542
rect 136824 272478 136876 272484
rect 135628 268252 135680 268258
rect 135628 268194 135680 268200
rect 132500 266484 132552 266490
rect 132500 266426 132552 266432
rect 136836 264330 136864 272478
rect 137664 270502 137692 274994
rect 137940 272542 137968 278052
rect 139136 275874 139164 278052
rect 140346 278038 140728 278066
rect 139124 275868 139176 275874
rect 139124 275810 139176 275816
rect 139400 273964 139452 273970
rect 139400 273906 139452 273912
rect 137928 272536 137980 272542
rect 137928 272478 137980 272484
rect 138480 271176 138532 271182
rect 138480 271118 138532 271124
rect 137468 270496 137520 270502
rect 137468 270438 137520 270444
rect 137652 270496 137704 270502
rect 137652 270438 137704 270444
rect 137480 266762 137508 270438
rect 137468 266756 137520 266762
rect 137468 266698 137520 266704
rect 138112 266620 138164 266626
rect 138112 266562 138164 266568
rect 136836 264302 137310 264330
rect 138124 264316 138152 266562
rect 138492 264330 138520 271118
rect 139412 264330 139440 273906
rect 140700 268258 140728 278038
rect 141056 275324 141108 275330
rect 141056 275266 141108 275272
rect 140136 268252 140188 268258
rect 140136 268194 140188 268200
rect 140688 268252 140740 268258
rect 140688 268194 140740 268200
rect 140148 267034 140176 268194
rect 140136 267028 140188 267034
rect 140136 266970 140188 266976
rect 140596 266892 140648 266898
rect 140596 266834 140648 266840
rect 138492 264302 138966 264330
rect 139412 264302 139794 264330
rect 140608 264316 140636 266834
rect 141068 264330 141096 275266
rect 141528 271182 141556 278052
rect 142724 272678 142752 278052
rect 142160 272672 142212 272678
rect 142160 272614 142212 272620
rect 142712 272672 142764 272678
rect 142712 272614 142764 272620
rect 141516 271176 141568 271182
rect 141516 271118 141568 271124
rect 142172 264330 142200 272614
rect 142712 271448 142764 271454
rect 142712 271390 142764 271396
rect 142724 264330 142752 271390
rect 143540 271312 143592 271318
rect 143540 271254 143592 271260
rect 143552 264330 143580 271254
rect 143920 269278 143948 278052
rect 144920 274100 144972 274106
rect 144920 274042 144972 274048
rect 143908 269272 143960 269278
rect 143908 269214 143960 269220
rect 144932 267734 144960 274042
rect 145116 272134 145144 278052
rect 146220 275058 146248 278052
rect 146208 275052 146260 275058
rect 146208 274994 146260 275000
rect 145288 274916 145340 274922
rect 145288 274858 145340 274864
rect 145300 273426 145328 274858
rect 145288 273420 145340 273426
rect 145288 273362 145340 273368
rect 147416 272678 147444 278052
rect 148612 273970 148640 278052
rect 149612 275188 149664 275194
rect 149612 275130 149664 275136
rect 148600 273964 148652 273970
rect 148600 273906 148652 273912
rect 147864 273420 147916 273426
rect 147864 273362 147916 273368
rect 145564 272672 145616 272678
rect 145564 272614 145616 272620
rect 147404 272672 147456 272678
rect 147404 272614 147456 272620
rect 145104 272128 145156 272134
rect 145104 272070 145156 272076
rect 144932 267706 145144 267734
rect 144736 267436 144788 267442
rect 144736 267378 144788 267384
rect 141068 264302 141450 264330
rect 142172 264302 142278 264330
rect 142724 264302 143106 264330
rect 143552 264302 143934 264330
rect 144748 264316 144776 267378
rect 145116 264330 145144 267706
rect 145576 267442 145604 272614
rect 146392 269816 146444 269822
rect 146392 269758 146444 269764
rect 145564 267436 145616 267442
rect 145564 267378 145616 267384
rect 145116 264302 145590 264330
rect 146404 264316 146432 269758
rect 147220 266484 147272 266490
rect 147220 266426 147272 266432
rect 147232 264316 147260 266426
rect 147876 264330 147904 273362
rect 148416 272808 148468 272814
rect 148416 272750 148468 272756
rect 148428 264330 148456 272750
rect 149428 269952 149480 269958
rect 149428 269894 149480 269900
rect 149440 264330 149468 269894
rect 149624 266626 149652 275130
rect 149808 274922 149836 278052
rect 151018 278038 151768 278066
rect 149796 274916 149848 274922
rect 149796 274858 149848 274864
rect 151084 271992 151136 271998
rect 151084 271934 151136 271940
rect 150532 266892 150584 266898
rect 150532 266834 150584 266840
rect 149612 266620 149664 266626
rect 149612 266562 149664 266568
rect 147876 264302 148074 264330
rect 148428 264302 148902 264330
rect 149440 264302 149730 264330
rect 150544 264316 150572 266834
rect 151096 266762 151124 271934
rect 151740 268122 151768 278038
rect 152004 271584 152056 271590
rect 152004 271526 152056 271532
rect 151728 268116 151780 268122
rect 151728 268058 151780 268064
rect 151360 267164 151412 267170
rect 151360 267106 151412 267112
rect 151084 266756 151136 266762
rect 151084 266698 151136 266704
rect 151372 264316 151400 267106
rect 152016 264330 152044 271526
rect 152200 271318 152228 278052
rect 152832 275732 152884 275738
rect 152832 275674 152884 275680
rect 152188 271312 152240 271318
rect 152188 271254 152240 271260
rect 152844 269958 152872 275674
rect 153396 275194 153424 278052
rect 153384 275188 153436 275194
rect 153384 275130 153436 275136
rect 154500 274106 154528 278052
rect 154764 275596 154816 275602
rect 154764 275538 154816 275544
rect 154488 274100 154540 274106
rect 154488 274042 154540 274048
rect 153844 273556 153896 273562
rect 153844 273498 153896 273504
rect 153016 270088 153068 270094
rect 153016 270030 153068 270036
rect 152832 269952 152884 269958
rect 152832 269894 152884 269900
rect 152016 264302 152214 264330
rect 153028 264316 153056 270030
rect 153856 267714 153884 273498
rect 154776 267734 154804 275538
rect 155696 272814 155724 278052
rect 156892 275466 156920 278052
rect 158102 278038 158668 278066
rect 156880 275460 156932 275466
rect 156880 275402 156932 275408
rect 157616 274372 157668 274378
rect 157616 274314 157668 274320
rect 155960 272944 156012 272950
rect 155960 272886 156012 272892
rect 155684 272808 155736 272814
rect 155684 272750 155736 272756
rect 155500 268388 155552 268394
rect 155500 268330 155552 268336
rect 153476 267708 153528 267714
rect 153476 267650 153528 267656
rect 153844 267708 153896 267714
rect 153844 267650 153896 267656
rect 154684 267706 154804 267734
rect 153488 264330 153516 267650
rect 153488 264302 153870 264330
rect 154684 264316 154712 267706
rect 155512 264316 155540 268330
rect 155972 264330 156000 272886
rect 157156 269952 157208 269958
rect 157156 269894 157208 269900
rect 155972 264302 156354 264330
rect 157168 264316 157196 269894
rect 157628 264330 157656 274314
rect 158640 269822 158668 278038
rect 159284 274378 159312 278052
rect 160480 275738 160508 278052
rect 160468 275732 160520 275738
rect 160468 275674 160520 275680
rect 159456 275324 159508 275330
rect 159456 275266 159508 275272
rect 159272 274372 159324 274378
rect 159272 274314 159324 274320
rect 158812 271720 158864 271726
rect 158812 271662 158864 271668
rect 158628 269816 158680 269822
rect 158628 269758 158680 269764
rect 157628 264302 158010 264330
rect 158824 264316 158852 271662
rect 159468 266898 159496 275266
rect 160928 274508 160980 274514
rect 160928 274450 160980 274456
rect 160468 268524 160520 268530
rect 160468 268466 160520 268472
rect 159456 266892 159508 266898
rect 159456 266834 159508 266840
rect 159640 266620 159692 266626
rect 159640 266562 159692 266568
rect 159652 264316 159680 266562
rect 160480 264316 160508 268466
rect 160940 264330 160968 274450
rect 161584 268394 161612 278052
rect 162780 277394 162808 278052
rect 162688 277366 162808 277394
rect 162688 271454 162716 277366
rect 163504 276004 163556 276010
rect 163504 275946 163556 275952
rect 162860 273080 162912 273086
rect 162860 273022 162912 273028
rect 162676 271448 162728 271454
rect 162676 271390 162728 271396
rect 161572 268388 161624 268394
rect 161572 268330 161624 268336
rect 162124 266892 162176 266898
rect 162124 266834 162176 266840
rect 160940 264302 161322 264330
rect 162136 264316 162164 266834
rect 162872 264330 162900 273022
rect 163516 266422 163544 275946
rect 163976 275466 164004 278052
rect 163964 275460 164016 275466
rect 163964 275402 164016 275408
rect 164976 271856 165028 271862
rect 164976 271798 165028 271804
rect 163780 268660 163832 268666
rect 163780 268602 163832 268608
rect 163504 266416 163556 266422
rect 163504 266358 163556 266364
rect 162872 264302 162978 264330
rect 163792 264316 163820 268602
rect 164608 267300 164660 267306
rect 164608 267242 164660 267248
rect 164620 264316 164648 267242
rect 164988 264330 165016 271798
rect 165172 271590 165200 278052
rect 165896 273216 165948 273222
rect 165896 273158 165948 273164
rect 165160 271584 165212 271590
rect 165160 271526 165212 271532
rect 165908 264330 165936 273158
rect 166368 272950 166396 278052
rect 167564 276010 167592 278052
rect 167552 276004 167604 276010
rect 167552 275946 167604 275952
rect 168288 274780 168340 274786
rect 168288 274722 168340 274728
rect 166356 272944 166408 272950
rect 166356 272886 166408 272892
rect 168104 270632 168156 270638
rect 168104 270574 168156 270580
rect 167920 268796 167972 268802
rect 167920 268738 167972 268744
rect 167092 266416 167144 266422
rect 167092 266358 167144 266364
rect 164988 264302 165462 264330
rect 165908 264302 166290 264330
rect 167104 264316 167132 266358
rect 167932 264316 167960 268738
rect 168116 267170 168144 270574
rect 168300 268802 168328 274722
rect 168760 274514 168788 278052
rect 169024 275188 169076 275194
rect 169024 275130 169076 275136
rect 168748 274508 168800 274514
rect 168748 274450 168800 274456
rect 168748 270224 168800 270230
rect 168748 270166 168800 270172
rect 168288 268796 168340 268802
rect 168288 268738 168340 268744
rect 168564 267572 168616 267578
rect 168564 267514 168616 267520
rect 168104 267164 168156 267170
rect 168104 267106 168156 267112
rect 168576 266422 168604 267514
rect 168564 266416 168616 266422
rect 168564 266358 168616 266364
rect 168760 264316 168788 270166
rect 169036 267578 169064 275130
rect 169864 271726 169892 278052
rect 171060 275602 171088 278052
rect 171048 275596 171100 275602
rect 171048 275538 171100 275544
rect 171600 274644 171652 274650
rect 171600 274586 171652 274592
rect 169852 271720 169904 271726
rect 169852 271662 169904 271668
rect 169944 271040 169996 271046
rect 169944 270982 169996 270988
rect 169024 267572 169076 267578
rect 169024 267514 169076 267520
rect 169576 266416 169628 266422
rect 169576 266358 169628 266364
rect 169588 264316 169616 266358
rect 169956 264330 169984 270982
rect 171232 268932 171284 268938
rect 171232 268874 171284 268880
rect 169956 264302 170430 264330
rect 171244 264316 171272 268874
rect 171612 264330 171640 274586
rect 172256 273086 172284 278052
rect 173466 278038 173848 278066
rect 174662 278038 175136 278066
rect 175858 278038 176608 278066
rect 173256 273692 173308 273698
rect 173256 273634 173308 273640
rect 172244 273080 172296 273086
rect 172244 273022 172296 273028
rect 172520 272400 172572 272406
rect 172520 272342 172572 272348
rect 172532 264330 172560 272342
rect 173268 264330 173296 273634
rect 173820 269958 173848 278038
rect 174268 275868 174320 275874
rect 174268 275810 174320 275816
rect 174280 271862 174308 275810
rect 174268 271856 174320 271862
rect 174268 271798 174320 271804
rect 173808 269952 173860 269958
rect 173808 269894 173860 269900
rect 175108 269074 175136 278038
rect 175280 273828 175332 273834
rect 175280 273770 175332 273776
rect 174544 269068 174596 269074
rect 174544 269010 174596 269016
rect 175096 269068 175148 269074
rect 175096 269010 175148 269016
rect 171612 264302 172086 264330
rect 172532 264302 172914 264330
rect 173268 264302 173742 264330
rect 174556 264316 174584 269010
rect 175292 264330 175320 273770
rect 176580 270094 176608 278038
rect 176568 270088 176620 270094
rect 176568 270030 176620 270036
rect 176200 269680 176252 269686
rect 176200 269622 176252 269628
rect 175292 264302 175398 264330
rect 176212 264316 176240 269622
rect 176948 268666 176976 278052
rect 178144 275874 178172 278052
rect 178868 276004 178920 276010
rect 178868 275946 178920 275952
rect 178132 275868 178184 275874
rect 178132 275810 178184 275816
rect 177488 270904 177540 270910
rect 177488 270846 177540 270852
rect 176936 268660 176988 268666
rect 176936 268602 176988 268608
rect 177028 267164 177080 267170
rect 177028 267106 177080 267112
rect 177040 264316 177068 267106
rect 177500 264330 177528 270846
rect 178684 269408 178736 269414
rect 178684 269350 178736 269356
rect 177672 269068 177724 269074
rect 177672 269010 177724 269016
rect 177684 267170 177712 269010
rect 177672 267164 177724 267170
rect 177672 267106 177724 267112
rect 177500 264302 177882 264330
rect 178696 264316 178724 269350
rect 178880 266898 178908 275946
rect 179340 274650 179368 278052
rect 180536 277394 180564 278052
rect 180536 277366 180656 277394
rect 179328 274644 179380 274650
rect 179328 274586 179380 274592
rect 179880 272264 179932 272270
rect 179880 272206 179932 272212
rect 178868 266892 178920 266898
rect 178868 266834 178920 266840
rect 179512 266756 179564 266762
rect 179512 266698 179564 266704
rect 179524 264316 179552 266698
rect 179892 264330 179920 272206
rect 180628 268530 180656 277366
rect 181732 272542 181760 278052
rect 182942 278038 183508 278066
rect 184138 278038 184888 278066
rect 182456 274236 182508 274242
rect 182456 274178 182508 274184
rect 181720 272536 181772 272542
rect 181720 272478 181772 272484
rect 181168 269544 181220 269550
rect 181168 269486 181220 269492
rect 180616 268524 180668 268530
rect 180616 268466 180668 268472
rect 179892 264302 180366 264330
rect 181180 264316 181208 269486
rect 181996 268796 182048 268802
rect 181996 268738 182048 268744
rect 182008 264316 182036 268738
rect 182468 264330 182496 274178
rect 183480 269686 183508 278038
rect 183652 270360 183704 270366
rect 183652 270302 183704 270308
rect 183468 269680 183520 269686
rect 183468 269622 183520 269628
rect 182468 264302 182850 264330
rect 183664 264316 183692 270302
rect 184860 270230 184888 278038
rect 185228 276010 185256 278052
rect 185216 276004 185268 276010
rect 185216 275946 185268 275952
rect 185308 275052 185360 275058
rect 185308 274994 185360 275000
rect 185124 270768 185176 270774
rect 185124 270710 185176 270716
rect 184848 270224 184900 270230
rect 184848 270166 184900 270172
rect 184480 267708 184532 267714
rect 184480 267650 184532 267656
rect 184492 264316 184520 267650
rect 185136 264330 185164 270710
rect 185320 270366 185348 274994
rect 186424 273222 186452 278052
rect 187436 278038 187634 278066
rect 186412 273216 186464 273222
rect 186412 273158 186464 273164
rect 186964 272536 187016 272542
rect 186964 272478 187016 272484
rect 186136 270496 186188 270502
rect 186136 270438 186188 270444
rect 185308 270360 185360 270366
rect 185308 270302 185360 270308
rect 185136 264302 185334 264330
rect 186148 264316 186176 270438
rect 186976 267306 187004 272478
rect 187436 271046 187464 278038
rect 188816 277394 188844 278052
rect 188816 277366 188936 277394
rect 187700 272400 187752 272406
rect 187700 272342 187752 272348
rect 187424 271040 187476 271046
rect 187424 270982 187476 270988
rect 186964 267300 187016 267306
rect 186964 267242 187016 267248
rect 186964 267028 187016 267034
rect 186964 266970 187016 266976
rect 186976 264316 187004 266970
rect 187712 264330 187740 272342
rect 188908 268802 188936 277366
rect 190012 275194 190040 278052
rect 190000 275188 190052 275194
rect 190000 275130 190052 275136
rect 189080 274916 189132 274922
rect 189080 274858 189132 274864
rect 189092 272270 189120 274858
rect 189080 272264 189132 272270
rect 189080 272206 189132 272212
rect 189264 271856 189316 271862
rect 189264 271798 189316 271804
rect 189080 271176 189132 271182
rect 189080 271118 189132 271124
rect 188896 268796 188948 268802
rect 188896 268738 188948 268744
rect 188620 268252 188672 268258
rect 188620 268194 188672 268200
rect 187712 264302 187818 264330
rect 188632 264316 188660 268194
rect 189092 265674 189120 271118
rect 189080 265668 189132 265674
rect 189080 265610 189132 265616
rect 189276 264330 189304 271798
rect 191208 271182 191236 278052
rect 192404 273834 192432 278052
rect 193508 274242 193536 278052
rect 194718 278038 195008 278066
rect 193496 274236 193548 274242
rect 193496 274178 193548 274184
rect 194784 273964 194836 273970
rect 194784 273906 194836 273912
rect 192392 273828 192444 273834
rect 192392 273770 192444 273776
rect 193220 272672 193272 272678
rect 193220 272614 193272 272620
rect 192392 272128 192444 272134
rect 192392 272070 192444 272076
rect 191196 271176 191248 271182
rect 191196 271118 191248 271124
rect 191104 269272 191156 269278
rect 191104 269214 191156 269220
rect 190460 268796 190512 268802
rect 190460 268738 190512 268744
rect 190472 267034 190500 268738
rect 190460 267028 190512 267034
rect 190460 266970 190512 266976
rect 189908 265668 189960 265674
rect 189908 265610 189960 265616
rect 189920 264330 189948 265610
rect 189276 264302 189474 264330
rect 189920 264302 190302 264330
rect 191116 264316 191144 269214
rect 191932 267436 191984 267442
rect 191932 267378 191984 267384
rect 191944 264316 191972 267378
rect 192404 264330 192432 272070
rect 193232 264330 193260 272614
rect 194416 270360 194468 270366
rect 194416 270302 194468 270308
rect 192404 264302 192786 264330
rect 193232 264302 193614 264330
rect 194428 264316 194456 270302
rect 194796 264330 194824 273906
rect 194980 272406 195008 278038
rect 195900 272542 195928 278052
rect 197096 272678 197124 278052
rect 198096 274100 198148 274106
rect 198096 274042 198148 274048
rect 197084 272672 197136 272678
rect 197084 272614 197136 272620
rect 195888 272536 195940 272542
rect 195888 272478 195940 272484
rect 194968 272400 195020 272406
rect 194968 272342 195020 272348
rect 196440 272264 196492 272270
rect 196440 272206 196492 272212
rect 196072 268116 196124 268122
rect 196072 268058 196124 268064
rect 194796 264302 195270 264330
rect 196084 264316 196112 268058
rect 196452 264330 196480 272206
rect 197360 271312 197412 271318
rect 197360 271254 197412 271260
rect 197372 264330 197400 271254
rect 198108 264330 198136 274042
rect 198292 271318 198320 278052
rect 199502 278038 199976 278066
rect 199568 275732 199620 275738
rect 199568 275674 199620 275680
rect 198280 271312 198332 271318
rect 198280 271254 198332 271260
rect 199384 267572 199436 267578
rect 199384 267514 199436 267520
rect 196452 264302 196926 264330
rect 197372 264302 197754 264330
rect 198108 264302 198582 264330
rect 199396 264316 199424 267514
rect 199580 267442 199608 275674
rect 199948 270366 199976 278038
rect 200120 272808 200172 272814
rect 200120 272750 200172 272756
rect 199936 270360 199988 270366
rect 199936 270302 199988 270308
rect 199568 267436 199620 267442
rect 199568 267378 199620 267384
rect 200132 264330 200160 272750
rect 200592 268802 200620 278052
rect 201788 277394 201816 278052
rect 201696 277366 201816 277394
rect 200764 275324 200816 275330
rect 200764 275266 200816 275272
rect 200776 270502 200804 275266
rect 200764 270496 200816 270502
rect 200764 270438 200816 270444
rect 201696 269822 201724 277366
rect 202328 274372 202380 274378
rect 202328 274314 202380 274320
rect 201868 270496 201920 270502
rect 201868 270438 201920 270444
rect 201040 269816 201092 269822
rect 201040 269758 201092 269764
rect 201684 269816 201736 269822
rect 201684 269758 201736 269764
rect 200580 268796 200632 268802
rect 200580 268738 200632 268744
rect 200132 264302 200238 264330
rect 201052 264316 201080 269758
rect 201880 264316 201908 270438
rect 202340 264330 202368 274314
rect 202984 271862 203012 278052
rect 202972 271856 203024 271862
rect 202972 271798 203024 271804
rect 204180 269550 204208 278052
rect 205376 272814 205404 278052
rect 206586 278038 206876 278066
rect 206376 275460 206428 275466
rect 206376 275402 206428 275408
rect 205364 272808 205416 272814
rect 205364 272750 205416 272756
rect 205640 271584 205692 271590
rect 205640 271526 205692 271532
rect 204720 271448 204772 271454
rect 204720 271390 204772 271396
rect 204168 269544 204220 269550
rect 204168 269486 204220 269492
rect 203524 268388 203576 268394
rect 203524 268330 203576 268336
rect 202340 264302 202722 264330
rect 203536 264316 203564 268330
rect 204352 267436 204404 267442
rect 204352 267378 204404 267384
rect 204364 264316 204392 267378
rect 204732 264330 204760 271390
rect 205456 269680 205508 269686
rect 205456 269622 205508 269628
rect 205468 267442 205496 269622
rect 205456 267436 205508 267442
rect 205456 267378 205508 267384
rect 205652 264330 205680 271526
rect 206388 264330 206416 275402
rect 206848 270502 206876 278038
rect 207768 274786 207796 278052
rect 207756 274780 207808 274786
rect 207756 274722 207808 274728
rect 208400 274508 208452 274514
rect 208400 274450 208452 274456
rect 207296 272944 207348 272950
rect 207296 272886 207348 272892
rect 206836 270496 206888 270502
rect 206836 270438 206888 270444
rect 207308 264330 207336 272886
rect 208412 264330 208440 274450
rect 208872 273970 208900 278052
rect 210068 274106 210096 278052
rect 210700 274780 210752 274786
rect 210700 274722 210752 274728
rect 210056 274100 210108 274106
rect 210056 274042 210108 274048
rect 208860 273964 208912 273970
rect 208860 273906 208912 273912
rect 209780 273080 209832 273086
rect 209780 273022 209832 273028
rect 209320 266892 209372 266898
rect 209320 266834 209372 266840
rect 204732 264302 205206 264330
rect 205652 264302 206034 264330
rect 206388 264302 206862 264330
rect 207308 264302 207690 264330
rect 208412 264302 208518 264330
rect 209332 264316 209360 266834
rect 209792 265674 209820 273022
rect 209964 271720 210016 271726
rect 209964 271662 210016 271668
rect 209780 265668 209832 265674
rect 209780 265610 209832 265616
rect 209976 264330 210004 271662
rect 210712 268394 210740 274722
rect 211264 272950 211292 278052
rect 211620 275596 211672 275602
rect 211620 275538 211672 275544
rect 211252 272944 211304 272950
rect 211252 272886 211304 272892
rect 211160 270088 211212 270094
rect 211160 270030 211212 270036
rect 210700 268388 210752 268394
rect 210700 268330 210752 268336
rect 211172 266422 211200 270030
rect 211160 266416 211212 266422
rect 211160 266358 211212 266364
rect 210700 265668 210752 265674
rect 210700 265610 210752 265616
rect 210712 264330 210740 265610
rect 211632 264330 211660 275538
rect 212460 270094 212488 278052
rect 213656 271454 213684 278052
rect 214852 275330 214880 278052
rect 214840 275324 214892 275330
rect 214840 275266 214892 275272
rect 214564 274644 214616 274650
rect 214564 274586 214616 274592
rect 213644 271448 213696 271454
rect 213644 271390 213696 271396
rect 212448 270088 212500 270094
rect 212448 270030 212500 270036
rect 212632 269952 212684 269958
rect 212632 269894 212684 269900
rect 209976 264302 210174 264330
rect 210712 264302 211002 264330
rect 211632 264302 211830 264330
rect 212644 264316 212672 269894
rect 214288 267164 214340 267170
rect 214288 267106 214340 267112
rect 213460 266416 213512 266422
rect 213460 266358 213512 266364
rect 213472 264316 213500 266358
rect 214300 264316 214328 267106
rect 214576 266422 214604 274586
rect 215956 271590 215984 278052
rect 216680 275868 216732 275874
rect 216680 275810 216732 275816
rect 215944 271584 215996 271590
rect 215944 271526 215996 271532
rect 215944 271040 215996 271046
rect 215944 270982 215996 270988
rect 215116 268660 215168 268666
rect 215116 268602 215168 268608
rect 214564 266416 214616 266422
rect 214564 266358 214616 266364
rect 215128 264316 215156 268602
rect 215956 267578 215984 270982
rect 215944 267572 215996 267578
rect 215944 267514 215996 267520
rect 215944 266416 215996 266422
rect 215944 266358 215996 266364
rect 215956 264316 215984 266358
rect 216692 264330 216720 275810
rect 217152 275738 217180 278052
rect 217140 275732 217192 275738
rect 217140 275674 217192 275680
rect 218348 275602 218376 278052
rect 218336 275596 218388 275602
rect 218336 275538 218388 275544
rect 218704 273216 218756 273222
rect 218704 273158 218756 273164
rect 217600 268524 217652 268530
rect 217600 268466 217652 268472
rect 216692 264302 216798 264330
rect 217612 264316 217640 268466
rect 218428 267436 218480 267442
rect 218428 267378 218480 267384
rect 218440 264316 218468 267378
rect 218716 266898 218744 273158
rect 219544 273086 219572 278052
rect 219532 273080 219584 273086
rect 219532 273022 219584 273028
rect 220740 272950 220768 278052
rect 221280 276004 221332 276010
rect 221280 275946 221332 275952
rect 220084 272944 220136 272950
rect 220084 272886 220136 272892
rect 220728 272944 220780 272950
rect 220728 272886 220780 272892
rect 219348 270224 219400 270230
rect 219348 270166 219400 270172
rect 219360 267458 219388 270166
rect 219360 267430 219664 267458
rect 219256 267300 219308 267306
rect 219256 267242 219308 267248
rect 218704 266892 218756 266898
rect 218704 266834 218756 266840
rect 219268 264316 219296 267242
rect 219636 264330 219664 267430
rect 220096 267170 220124 272886
rect 220084 267164 220136 267170
rect 220084 267106 220136 267112
rect 220912 266892 220964 266898
rect 220912 266834 220964 266840
rect 219636 264302 220110 264330
rect 220924 264316 220952 266834
rect 221292 264330 221320 275946
rect 221936 275466 221964 278052
rect 221924 275460 221976 275466
rect 221924 275402 221976 275408
rect 222936 275188 222988 275194
rect 222936 275130 222988 275136
rect 222568 267572 222620 267578
rect 222568 267514 222620 267520
rect 221292 264302 221766 264330
rect 222580 264316 222608 267514
rect 222948 264330 222976 275130
rect 223132 274378 223160 278052
rect 224236 275874 224264 278052
rect 224224 275868 224276 275874
rect 224224 275810 224276 275816
rect 224224 275732 224276 275738
rect 224224 275674 224276 275680
rect 223120 274372 223172 274378
rect 223120 274314 223172 274320
rect 223488 269544 223540 269550
rect 223488 269486 223540 269492
rect 223500 267306 223528 269486
rect 224236 268666 224264 275674
rect 224960 273828 225012 273834
rect 224960 273770 225012 273776
rect 224224 268660 224276 268666
rect 224224 268602 224276 268608
rect 223488 267300 223540 267306
rect 223488 267242 223540 267248
rect 224224 267028 224276 267034
rect 224224 266970 224276 266976
rect 222948 264302 223422 264330
rect 224236 264316 224264 266970
rect 224972 265674 225000 273770
rect 225432 271726 225460 278052
rect 226432 274236 226484 274242
rect 226432 274178 226484 274184
rect 225420 271720 225472 271726
rect 225420 271662 225472 271668
rect 225144 271176 225196 271182
rect 225144 271118 225196 271124
rect 224960 265668 225012 265674
rect 224960 265610 225012 265616
rect 225156 265554 225184 271118
rect 225604 265668 225656 265674
rect 225604 265610 225656 265616
rect 225064 265526 225184 265554
rect 225064 264316 225092 265526
rect 225616 264330 225644 265610
rect 226444 264330 226472 274178
rect 226628 269958 226656 278052
rect 227838 278038 228128 278066
rect 228100 272542 228128 278038
rect 229020 275738 229048 278052
rect 229008 275732 229060 275738
rect 229008 275674 229060 275680
rect 229100 272672 229152 272678
rect 229100 272614 229152 272620
rect 227904 272536 227956 272542
rect 227904 272478 227956 272484
rect 228088 272536 228140 272542
rect 228088 272478 228140 272484
rect 227168 272400 227220 272406
rect 227168 272342 227220 272348
rect 226616 269952 226668 269958
rect 226616 269894 226668 269900
rect 227180 264330 227208 272342
rect 227916 264330 227944 272478
rect 228364 271720 228416 271726
rect 228364 271662 228416 271668
rect 228376 267034 228404 271662
rect 228364 267028 228416 267034
rect 228364 266970 228416 266976
rect 229112 264330 229140 272614
rect 229560 271312 229612 271318
rect 229560 271254 229612 271260
rect 229572 264330 229600 271254
rect 230216 271182 230244 278052
rect 231334 278038 231716 278066
rect 230204 271176 230256 271182
rect 230204 271118 230256 271124
rect 230848 270360 230900 270366
rect 230848 270302 230900 270308
rect 225616 264302 225906 264330
rect 226444 264302 226734 264330
rect 227180 264302 227562 264330
rect 227916 264302 228390 264330
rect 229112 264302 229218 264330
rect 229572 264302 230046 264330
rect 230860 264316 230888 270302
rect 231308 268796 231360 268802
rect 231308 268738 231360 268744
rect 231320 264330 231348 268738
rect 231688 268530 231716 278038
rect 232516 276010 232544 278052
rect 232504 276004 232556 276010
rect 232504 275946 232556 275952
rect 232688 275868 232740 275874
rect 232688 275810 232740 275816
rect 232700 270366 232728 275810
rect 233712 272678 233740 278052
rect 234922 278038 235304 278066
rect 233884 275596 233936 275602
rect 233884 275538 233936 275544
rect 233700 272672 233752 272678
rect 233700 272614 233752 272620
rect 233240 271856 233292 271862
rect 233240 271798 233292 271804
rect 232688 270360 232740 270366
rect 232688 270302 232740 270308
rect 232504 269816 232556 269822
rect 232504 269758 232556 269764
rect 231676 268524 231728 268530
rect 231676 268466 231728 268472
rect 231320 264302 231702 264330
rect 232516 264316 232544 269758
rect 233252 264330 233280 271798
rect 233896 267442 233924 275538
rect 234804 272808 234856 272814
rect 234804 272750 234856 272756
rect 233884 267436 233936 267442
rect 233884 267378 233936 267384
rect 234160 267300 234212 267306
rect 234160 267242 234212 267248
rect 233252 264302 233358 264330
rect 234172 264316 234200 267242
rect 234816 264330 234844 272750
rect 235276 271318 235304 278038
rect 236104 275874 236132 278052
rect 236092 275868 236144 275874
rect 236092 275810 236144 275816
rect 235264 271312 235316 271318
rect 235264 271254 235316 271260
rect 235816 270496 235868 270502
rect 235816 270438 235868 270444
rect 234816 264302 235014 264330
rect 235828 264316 235856 270438
rect 237300 269822 237328 278052
rect 237840 274100 237892 274106
rect 237840 274042 237892 274048
rect 237472 273964 237524 273970
rect 237472 273906 237524 273912
rect 237288 269816 237340 269822
rect 237288 269758 237340 269764
rect 236644 268388 236696 268394
rect 236644 268330 236696 268336
rect 236656 264316 236684 268330
rect 237484 264316 237512 273906
rect 237852 264330 237880 274042
rect 238496 273970 238524 278052
rect 239220 276004 239272 276010
rect 239220 275946 239272 275952
rect 239232 274242 239260 275946
rect 239600 275602 239628 278052
rect 239588 275596 239640 275602
rect 239588 275538 239640 275544
rect 239404 275324 239456 275330
rect 239404 275266 239456 275272
rect 239220 274236 239272 274242
rect 239220 274178 239272 274184
rect 238484 273964 238536 273970
rect 238484 273906 238536 273912
rect 239128 267164 239180 267170
rect 239128 267106 239180 267112
rect 237852 264302 238326 264330
rect 239140 264316 239168 267106
rect 239416 266422 239444 275266
rect 240796 271454 240824 278052
rect 241992 277394 242020 278052
rect 241900 277366 242020 277394
rect 240416 271448 240468 271454
rect 240416 271390 240468 271396
rect 240784 271448 240836 271454
rect 240784 271390 240836 271396
rect 239956 270088 240008 270094
rect 239956 270030 240008 270036
rect 239404 266416 239456 266422
rect 239404 266358 239456 266364
rect 239968 264316 239996 270030
rect 240428 264330 240456 271390
rect 241900 270094 241928 277366
rect 243188 275330 243216 278052
rect 243544 275732 243596 275738
rect 243544 275674 243596 275680
rect 243176 275324 243228 275330
rect 243176 275266 243228 275272
rect 242072 271584 242124 271590
rect 242072 271526 242124 271532
rect 241888 270088 241940 270094
rect 241888 270030 241940 270036
rect 241612 266416 241664 266422
rect 241612 266358 241664 266364
rect 240428 264302 240810 264330
rect 241624 264316 241652 266358
rect 242084 264330 242112 271526
rect 243268 268660 243320 268666
rect 243268 268602 243320 268608
rect 242084 264302 242466 264330
rect 243280 264316 243308 268602
rect 243556 267442 243584 275674
rect 243728 275460 243780 275466
rect 243728 275402 243780 275408
rect 243544 267436 243596 267442
rect 243544 267378 243596 267384
rect 243740 266422 243768 275402
rect 244384 270230 244412 278052
rect 245396 278038 245502 278066
rect 246790 278038 246988 278066
rect 244556 273080 244608 273086
rect 244556 273022 244608 273028
rect 244372 270224 244424 270230
rect 244372 270166 244424 270172
rect 244096 267300 244148 267306
rect 244096 267242 244148 267248
rect 243728 266416 243780 266422
rect 243728 266358 243780 266364
rect 244108 264316 244136 267242
rect 244568 264330 244596 273022
rect 245396 272814 245424 278038
rect 245752 272944 245804 272950
rect 245752 272886 245804 272892
rect 245384 272808 245436 272814
rect 245384 272750 245436 272756
rect 244568 264302 244950 264330
rect 245764 264316 245792 272886
rect 246960 267170 246988 278038
rect 247224 274372 247276 274378
rect 247224 274314 247276 274320
rect 246948 267164 247000 267170
rect 246948 267106 247000 267112
rect 246580 266416 246632 266422
rect 246580 266358 246632 266364
rect 246592 264316 246620 266358
rect 247236 264330 247264 274314
rect 247880 272950 247908 278052
rect 249076 274106 249104 278052
rect 250272 275738 250300 278052
rect 250444 275868 250496 275874
rect 250444 275810 250496 275816
rect 250260 275732 250312 275738
rect 250260 275674 250312 275680
rect 249064 274100 249116 274106
rect 249064 274042 249116 274048
rect 247868 272944 247920 272950
rect 247868 272886 247920 272892
rect 249064 272536 249116 272542
rect 249064 272478 249116 272484
rect 248236 270360 248288 270366
rect 248236 270302 248288 270308
rect 247236 264302 247434 264330
rect 248248 264316 248276 270302
rect 249076 267034 249104 272478
rect 249892 269952 249944 269958
rect 249892 269894 249944 269900
rect 249064 267028 249116 267034
rect 249064 266970 249116 266976
rect 249064 266892 249116 266898
rect 249064 266834 249116 266840
rect 249076 264316 249104 266834
rect 249904 264316 249932 269894
rect 250456 266422 250484 275810
rect 251468 271046 251496 278052
rect 252008 271176 252060 271182
rect 252008 271118 252060 271124
rect 251456 271040 251508 271046
rect 251456 270982 251508 270988
rect 251548 267436 251600 267442
rect 251548 267378 251600 267384
rect 250720 267028 250772 267034
rect 250720 266970 250772 266976
rect 250444 266416 250496 266422
rect 250444 266358 250496 266364
rect 250732 264316 250760 266970
rect 251560 264316 251588 267378
rect 252020 264330 252048 271118
rect 252664 268394 252692 278052
rect 253860 274718 253888 278052
rect 253848 274712 253900 274718
rect 253848 274654 253900 274660
rect 253940 274236 253992 274242
rect 253940 274178 253992 274184
rect 253204 268524 253256 268530
rect 253204 268466 253256 268472
rect 252652 268388 252704 268394
rect 252652 268330 252704 268336
rect 252020 264302 252402 264330
rect 253216 264316 253244 268466
rect 253952 264330 253980 274178
rect 254400 272672 254452 272678
rect 254400 272614 254452 272620
rect 254412 264330 254440 272614
rect 254964 272542 254992 278052
rect 255964 275596 256016 275602
rect 255964 275538 256016 275544
rect 254952 272536 255004 272542
rect 254952 272478 255004 272484
rect 255320 271312 255372 271318
rect 255320 271254 255372 271260
rect 255332 264330 255360 271254
rect 255976 267034 256004 275538
rect 256160 275466 256188 278052
rect 257356 275602 257384 278052
rect 257344 275596 257396 275602
rect 257344 275538 257396 275544
rect 256148 275460 256200 275466
rect 256148 275402 256200 275408
rect 256700 275324 256752 275330
rect 256700 275266 256752 275272
rect 256712 271318 256740 275266
rect 256884 274712 256936 274718
rect 256884 274654 256936 274660
rect 256700 271312 256752 271318
rect 256700 271254 256752 271260
rect 256896 269958 256924 274654
rect 258080 273828 258132 273834
rect 258080 273770 258132 273776
rect 256884 269952 256936 269958
rect 256884 269894 256936 269900
rect 257344 269816 257396 269822
rect 257344 269758 257396 269764
rect 255964 267028 256016 267034
rect 255964 266970 256016 266976
rect 256516 266416 256568 266422
rect 256516 266358 256568 266364
rect 253952 264302 254058 264330
rect 254412 264302 254886 264330
rect 255332 264302 255714 264330
rect 256528 264316 256556 266358
rect 257356 264316 257384 269758
rect 258092 264330 258120 273770
rect 258552 269822 258580 278052
rect 259762 278038 260144 278066
rect 259368 275732 259420 275738
rect 259368 275674 259420 275680
rect 259380 273834 259408 275674
rect 259368 273828 259420 273834
rect 259368 273770 259420 273776
rect 260116 271454 260144 278038
rect 260944 275806 260972 278052
rect 260932 275800 260984 275806
rect 260932 275742 260984 275748
rect 259644 271448 259696 271454
rect 259644 271390 259696 271396
rect 260104 271448 260156 271454
rect 260104 271390 260156 271396
rect 258540 269816 258592 269822
rect 258540 269758 258592 269764
rect 259000 267028 259052 267034
rect 259000 266970 259052 266976
rect 258092 264302 258198 264330
rect 259012 264316 259040 266970
rect 259656 264330 259684 271390
rect 262048 271318 262076 278052
rect 262312 275596 262364 275602
rect 262312 275538 262364 275544
rect 262324 272814 262352 275538
rect 263244 275126 263272 278052
rect 263232 275120 263284 275126
rect 263232 275062 263284 275068
rect 264244 272944 264296 272950
rect 264244 272886 264296 272892
rect 262312 272808 262364 272814
rect 262312 272750 262364 272756
rect 262680 272672 262732 272678
rect 262680 272614 262732 272620
rect 261024 271312 261076 271318
rect 261024 271254 261076 271260
rect 262036 271312 262088 271318
rect 262036 271254 262088 271260
rect 260656 270088 260708 270094
rect 260656 270030 260708 270036
rect 259656 264302 259854 264330
rect 260668 264316 260696 270030
rect 261036 264330 261064 271254
rect 262312 270224 262364 270230
rect 262312 270166 262364 270172
rect 261036 264302 261510 264330
rect 262324 264316 262352 270166
rect 262692 264330 262720 272614
rect 264256 267734 264284 272886
rect 264440 272678 264468 278052
rect 265650 278038 266216 278066
rect 265256 274100 265308 274106
rect 265256 274042 265308 274048
rect 264428 272672 264480 272678
rect 264428 272614 264480 272620
rect 264256 267706 264376 267734
rect 263968 267164 264020 267170
rect 263968 267106 264020 267112
rect 262692 264302 263166 264330
rect 263980 264316 264008 267106
rect 264348 264330 264376 267706
rect 265268 264330 265296 274042
rect 266188 270094 266216 278038
rect 266360 275800 266412 275806
rect 266360 275742 266412 275748
rect 266372 274106 266400 275742
rect 266832 275602 266860 278052
rect 266820 275596 266872 275602
rect 266820 275538 266872 275544
rect 266360 274100 266412 274106
rect 266360 274042 266412 274048
rect 266360 273828 266412 273834
rect 266360 273770 266412 273776
rect 266176 270088 266228 270094
rect 266176 270030 266228 270036
rect 266372 264330 266400 273770
rect 268028 271182 268056 278052
rect 269224 275398 269252 278052
rect 269212 275392 269264 275398
rect 269212 275334 269264 275340
rect 270132 275256 270184 275262
rect 270132 275198 270184 275204
rect 269304 272536 269356 272542
rect 269304 272478 269356 272484
rect 268016 271176 268068 271182
rect 268016 271118 268068 271124
rect 266912 271040 266964 271046
rect 266912 270982 266964 270988
rect 266924 264330 266952 270982
rect 268936 269952 268988 269958
rect 268936 269894 268988 269900
rect 268108 268388 268160 268394
rect 268108 268330 268160 268336
rect 264348 264302 264822 264330
rect 265268 264302 265650 264330
rect 266372 264302 266478 264330
rect 266924 264302 267306 264330
rect 268120 264316 268148 268330
rect 268948 264316 268976 269894
rect 269316 264330 269344 272478
rect 270144 272354 270172 275198
rect 270328 272542 270356 278052
rect 271524 273970 271552 278052
rect 272734 278038 273116 278066
rect 273930 278038 274312 278066
rect 271512 273964 271564 273970
rect 271512 273906 271564 273912
rect 270960 272808 271012 272814
rect 270960 272750 271012 272756
rect 270316 272536 270368 272542
rect 270316 272478 270368 272484
rect 270144 272326 270540 272354
rect 270512 264330 270540 272326
rect 270972 264330 271000 272750
rect 272616 271448 272668 271454
rect 272616 271390 272668 271396
rect 272248 269816 272300 269822
rect 272248 269758 272300 269764
rect 269316 264302 269790 264330
rect 270512 264302 270618 264330
rect 270972 264302 271446 264330
rect 272260 264316 272288 269758
rect 272628 264330 272656 271390
rect 273088 269822 273116 278038
rect 273260 275120 273312 275126
rect 273260 275062 273312 275068
rect 273076 269816 273128 269822
rect 273076 269758 273128 269764
rect 273272 269074 273300 275062
rect 273536 274100 273588 274106
rect 273536 274042 273588 274048
rect 273260 269068 273312 269074
rect 273260 269010 273312 269016
rect 273548 264330 273576 274042
rect 274284 272814 274312 278038
rect 274640 275392 274692 275398
rect 274640 275334 274692 275340
rect 274272 272808 274324 272814
rect 274272 272750 274324 272756
rect 274652 271862 274680 275334
rect 275112 274718 275140 278052
rect 276308 275330 276336 278052
rect 276480 275596 276532 275602
rect 276480 275538 276532 275544
rect 276296 275324 276348 275330
rect 276296 275266 276348 275272
rect 275100 274712 275152 274718
rect 275100 274654 275152 274660
rect 276020 272672 276072 272678
rect 276020 272614 276072 272620
rect 274640 271856 274692 271862
rect 274640 271798 274692 271804
rect 274640 271312 274692 271318
rect 274640 271254 274692 271260
rect 274652 264330 274680 271254
rect 275560 269068 275612 269074
rect 275560 269010 275612 269016
rect 272628 264302 273102 264330
rect 273548 264302 273930 264330
rect 274652 264302 274758 264330
rect 275572 264316 275600 269010
rect 276032 264330 276060 272614
rect 276492 267782 276520 275538
rect 277504 275534 277532 278052
rect 277492 275528 277544 275534
rect 277492 275470 277544 275476
rect 278320 274712 278372 274718
rect 278320 274654 278372 274660
rect 278332 270502 278360 274654
rect 278608 274106 278636 278052
rect 278596 274100 278648 274106
rect 278596 274042 278648 274048
rect 279240 271856 279292 271862
rect 279240 271798 279292 271804
rect 278780 271176 278832 271182
rect 278780 271118 278832 271124
rect 278320 270496 278372 270502
rect 278320 270438 278372 270444
rect 277216 270088 277268 270094
rect 277216 270030 277268 270036
rect 276480 267776 276532 267782
rect 276480 267718 276532 267724
rect 276032 264302 276414 264330
rect 277228 264316 277256 270030
rect 278044 267776 278096 267782
rect 278044 267718 278096 267724
rect 278056 264316 278084 267718
rect 278792 264330 278820 271118
rect 279252 264330 279280 271798
rect 279804 271182 279832 278052
rect 280344 273964 280396 273970
rect 280344 273906 280396 273912
rect 279792 271176 279844 271182
rect 279792 271118 279844 271124
rect 280356 265674 280384 273906
rect 281000 273086 281028 278052
rect 282210 278038 282776 278066
rect 280988 273080 281040 273086
rect 280988 273022 281040 273028
rect 280528 272536 280580 272542
rect 280528 272478 280580 272484
rect 280344 265668 280396 265674
rect 280344 265610 280396 265616
rect 278792 264302 278898 264330
rect 279252 264302 279726 264330
rect 280540 264316 280568 272478
rect 282184 269816 282236 269822
rect 282184 269758 282236 269764
rect 280988 265668 281040 265674
rect 280988 265610 281040 265616
rect 281000 264330 281028 265610
rect 281000 264302 281382 264330
rect 282196 264316 282224 269758
rect 282748 269278 282776 278038
rect 283104 275324 283156 275330
rect 283104 275266 283156 275272
rect 282920 272808 282972 272814
rect 282920 272750 282972 272756
rect 282736 269272 282788 269278
rect 282736 269214 282788 269220
rect 282932 264330 282960 272750
rect 283116 270366 283144 275266
rect 283392 274718 283420 278052
rect 284588 275738 284616 278052
rect 284576 275732 284628 275738
rect 284576 275674 284628 275680
rect 285128 275528 285180 275534
rect 285128 275470 285180 275476
rect 283380 274712 283432 274718
rect 283380 274654 283432 274660
rect 283840 270496 283892 270502
rect 283840 270438 283892 270444
rect 283104 270360 283156 270366
rect 283104 270302 283156 270308
rect 282932 264302 283038 264330
rect 283852 264316 283880 270438
rect 284668 270360 284720 270366
rect 284668 270302 284720 270308
rect 284680 264316 284708 270302
rect 285140 264330 285168 275470
rect 285692 275330 285720 278052
rect 286888 275874 286916 278052
rect 286876 275868 286928 275874
rect 286876 275810 286928 275816
rect 285680 275324 285732 275330
rect 285680 275266 285732 275272
rect 288084 275058 288112 278052
rect 288072 275052 288124 275058
rect 288072 274994 288124 275000
rect 289280 274922 289308 278052
rect 290096 275732 290148 275738
rect 290096 275674 290148 275680
rect 289268 274916 289320 274922
rect 289268 274858 289320 274864
rect 289176 274712 289228 274718
rect 289176 274654 289228 274660
rect 285864 274100 285916 274106
rect 285864 274042 285916 274048
rect 285876 264330 285904 274042
rect 286324 273080 286376 273086
rect 286324 273022 286376 273028
rect 286336 267034 286364 273022
rect 287060 271176 287112 271182
rect 287060 271118 287112 271124
rect 286324 267028 286376 267034
rect 286324 266970 286376 266976
rect 287072 264330 287100 271118
rect 288808 269272 288860 269278
rect 288808 269214 288860 269220
rect 287980 267028 288032 267034
rect 287980 266970 288032 266976
rect 285140 264302 285522 264330
rect 285876 264302 286350 264330
rect 287072 264302 287178 264330
rect 287992 264316 288020 266970
rect 288820 264316 288848 269214
rect 289188 264330 289216 274654
rect 290108 264330 290136 275674
rect 290476 274718 290504 278052
rect 291672 275330 291700 278052
rect 291844 275868 291896 275874
rect 291844 275810 291896 275816
rect 291292 275324 291344 275330
rect 291292 275266 291344 275272
rect 291660 275324 291712 275330
rect 291660 275266 291712 275272
rect 290464 274712 290516 274718
rect 290464 274654 290516 274660
rect 289188 264302 289662 264330
rect 290108 264302 290490 264330
rect 291304 264316 291332 275266
rect 291856 264330 291884 275810
rect 292868 275194 292896 278052
rect 292856 275188 292908 275194
rect 292856 275130 292908 275136
rect 292856 275052 292908 275058
rect 292856 274994 292908 275000
rect 292672 274916 292724 274922
rect 292672 274858 292724 274864
rect 292684 265674 292712 274858
rect 292672 265668 292724 265674
rect 292672 265610 292724 265616
rect 292868 264330 292896 274994
rect 293972 274990 294000 278052
rect 293960 274984 294012 274990
rect 293960 274926 294012 274932
rect 295168 274718 295196 278052
rect 295340 275324 295392 275330
rect 295340 275266 295392 275272
rect 294144 274712 294196 274718
rect 294144 274654 294196 274660
rect 295156 274712 295208 274718
rect 295156 274654 295208 274660
rect 293500 265668 293552 265674
rect 293500 265610 293552 265616
rect 293512 264330 293540 265610
rect 294156 264330 294184 274654
rect 295352 264330 295380 275266
rect 295800 275188 295852 275194
rect 295800 275130 295852 275136
rect 295812 264330 295840 275130
rect 296364 274854 296392 278052
rect 297180 274984 297232 274990
rect 297180 274926 297232 274932
rect 296352 274848 296404 274854
rect 296352 274790 296404 274796
rect 296812 274712 296864 274718
rect 296812 274654 296864 274660
rect 296824 265674 296852 274654
rect 297192 267734 297220 274926
rect 297560 274718 297588 278052
rect 298756 275194 298784 278052
rect 299952 275330 299980 278052
rect 300964 278038 301070 278066
rect 302266 278038 302464 278066
rect 299940 275324 299992 275330
rect 299940 275266 299992 275272
rect 298744 275188 298796 275194
rect 298744 275130 298796 275136
rect 300032 275188 300084 275194
rect 300032 275130 300084 275136
rect 298376 274848 298428 274854
rect 298376 274790 298428 274796
rect 297548 274712 297600 274718
rect 297548 274654 297600 274660
rect 297100 267706 297220 267734
rect 296812 265668 296864 265674
rect 296812 265610 296864 265616
rect 291856 264302 292146 264330
rect 292868 264302 292974 264330
rect 293512 264302 293802 264330
rect 294156 264302 294630 264330
rect 295352 264302 295458 264330
rect 295812 264302 296286 264330
rect 297100 264316 297128 267706
rect 297548 265668 297600 265674
rect 297548 265610 297600 265616
rect 297560 264330 297588 265610
rect 298388 264330 298416 274790
rect 299480 274712 299532 274718
rect 299480 274654 299532 274660
rect 299492 264330 299520 274654
rect 300044 264330 300072 275130
rect 300964 266422 300992 278038
rect 301136 275324 301188 275330
rect 301136 275266 301188 275272
rect 300952 266416 301004 266422
rect 300952 266358 301004 266364
rect 301148 264330 301176 275266
rect 302056 266416 302108 266422
rect 302056 266358 302108 266364
rect 297560 264302 297942 264330
rect 298388 264302 298770 264330
rect 299492 264302 299598 264330
rect 300044 264302 300426 264330
rect 301148 264302 301254 264330
rect 302068 264316 302096 266358
rect 302436 264330 302464 278038
rect 303448 274718 303476 278052
rect 303724 278038 304658 278066
rect 305012 278038 305854 278066
rect 306392 278038 307050 278066
rect 307772 278038 308154 278066
rect 309152 278038 309350 278066
rect 303436 274712 303488 274718
rect 303436 274654 303488 274660
rect 303724 266422 303752 278038
rect 303988 274712 304040 274718
rect 303988 274654 304040 274660
rect 303712 266416 303764 266422
rect 303712 266358 303764 266364
rect 304000 264330 304028 274654
rect 304540 266416 304592 266422
rect 304540 266358 304592 266364
rect 302436 264302 302910 264330
rect 303738 264302 304028 264330
rect 304552 264316 304580 266358
rect 305012 264330 305040 278038
rect 306392 266370 306420 278038
rect 307772 267734 307800 278038
rect 306208 266342 306420 266370
rect 307496 267706 307800 267734
rect 305012 264302 305394 264330
rect 306208 264316 306236 266342
rect 307496 264330 307524 267706
rect 308680 266688 308732 266694
rect 308680 266630 308732 266636
rect 307852 266416 307904 266422
rect 307852 266358 307904 266364
rect 307050 264302 307524 264330
rect 307864 264316 307892 266358
rect 308692 264316 308720 266630
rect 309152 266422 309180 278038
rect 310532 266694 310560 278052
rect 310716 278038 311742 278066
rect 311912 278038 312938 278066
rect 313292 278038 314134 278066
rect 314672 278038 315238 278066
rect 316052 278038 316434 278066
rect 317432 278038 317630 278066
rect 318826 278038 319024 278066
rect 310520 266688 310572 266694
rect 310520 266630 310572 266636
rect 310336 266552 310388 266558
rect 310336 266494 310388 266500
rect 309140 266416 309192 266422
rect 309140 266358 309192 266364
rect 309508 266416 309560 266422
rect 309508 266358 309560 266364
rect 309520 264316 309548 266358
rect 310348 264316 310376 266494
rect 310716 266422 310744 278038
rect 311912 266558 311940 278038
rect 312820 267164 312872 267170
rect 312820 267106 312872 267112
rect 311900 266552 311952 266558
rect 311900 266494 311952 266500
rect 312268 266552 312320 266558
rect 312268 266494 312320 266500
rect 310704 266416 310756 266422
rect 310704 266358 310756 266364
rect 311164 266416 311216 266422
rect 311164 266358 311216 266364
rect 311176 264316 311204 266358
rect 312280 264330 312308 266494
rect 312018 264302 312308 264330
rect 312832 264316 312860 267106
rect 313292 266422 313320 278038
rect 314476 267028 314528 267034
rect 314476 266970 314528 266976
rect 313648 266688 313700 266694
rect 313648 266630 313700 266636
rect 313280 266416 313332 266422
rect 313280 266358 313332 266364
rect 313660 264316 313688 266630
rect 314488 264316 314516 266970
rect 314672 266558 314700 278038
rect 315304 267436 315356 267442
rect 315304 267378 315356 267384
rect 314660 266552 314712 266558
rect 314660 266494 314712 266500
rect 315316 264316 315344 267378
rect 316052 267170 316080 278038
rect 316040 267164 316092 267170
rect 316040 267106 316092 267112
rect 316960 266824 317012 266830
rect 316960 266766 317012 266772
rect 316132 266552 316184 266558
rect 316132 266494 316184 266500
rect 316144 264316 316172 266494
rect 316972 264316 317000 266766
rect 317432 266694 317460 278038
rect 318708 272400 318760 272406
rect 318708 272342 318760 272348
rect 318720 267734 318748 272342
rect 318628 267706 318748 267734
rect 317420 266688 317472 266694
rect 317420 266630 317472 266636
rect 317788 266688 317840 266694
rect 317788 266630 317840 266636
rect 317800 264316 317828 266630
rect 318628 264316 318656 267706
rect 318996 267034 319024 278038
rect 319180 278038 320022 278066
rect 320192 278038 321218 278066
rect 321572 278038 322414 278066
rect 322952 278038 323518 278066
rect 319180 267442 319208 278038
rect 319444 269136 319496 269142
rect 319444 269078 319496 269084
rect 319168 267436 319220 267442
rect 319168 267378 319220 267384
rect 318984 267028 319036 267034
rect 318984 266970 319036 266976
rect 319456 264316 319484 269078
rect 320192 266558 320220 278038
rect 321192 274712 321244 274718
rect 321192 274654 321244 274660
rect 321204 267734 321232 274654
rect 321376 270768 321428 270774
rect 321376 270710 321428 270716
rect 321112 267706 321232 267734
rect 320180 266552 320232 266558
rect 320180 266494 320232 266500
rect 320272 266416 320324 266422
rect 320272 266358 320324 266364
rect 320284 264316 320312 266358
rect 321112 264316 321140 267706
rect 321388 266422 321416 270710
rect 321572 266830 321600 278038
rect 322756 273964 322808 273970
rect 322756 273906 322808 273912
rect 321928 267300 321980 267306
rect 321928 267242 321980 267248
rect 321560 266824 321612 266830
rect 321560 266766 321612 266772
rect 321376 266416 321428 266422
rect 321376 266358 321428 266364
rect 321940 264316 321968 267242
rect 322768 264316 322796 273906
rect 322952 266694 322980 278038
rect 324044 272672 324096 272678
rect 324044 272614 324096 272620
rect 322940 266688 322992 266694
rect 322940 266630 322992 266636
rect 324056 264330 324084 272614
rect 324700 272406 324728 278052
rect 325712 278038 325910 278066
rect 325332 272808 325384 272814
rect 325332 272750 325384 272756
rect 324688 272400 324740 272406
rect 324688 272342 324740 272348
rect 325344 266422 325372 272750
rect 325516 271448 325568 271454
rect 325516 271390 325568 271396
rect 324412 266416 324464 266422
rect 324412 266358 324464 266364
rect 325332 266416 325384 266422
rect 325332 266358 325384 266364
rect 323610 264302 324084 264330
rect 324424 264316 324452 266358
rect 325528 264330 325556 271390
rect 325712 269142 325740 278038
rect 326436 275324 326488 275330
rect 326436 275266 326488 275272
rect 325700 269136 325752 269142
rect 325700 269078 325752 269084
rect 326448 264330 326476 275266
rect 327092 270774 327120 278052
rect 328288 274718 328316 278052
rect 328276 274712 328328 274718
rect 328276 274654 328328 274660
rect 329484 273290 329512 278052
rect 330588 273970 330616 278052
rect 331416 278038 331798 278066
rect 330576 273964 330628 273970
rect 330576 273906 330628 273912
rect 327724 273284 327776 273290
rect 327724 273226 327776 273232
rect 329472 273284 329524 273290
rect 329472 273226 329524 273232
rect 327080 270768 327132 270774
rect 327080 270710 327132 270716
rect 326896 269816 326948 269822
rect 326896 269758 326948 269764
rect 325266 264302 325556 264330
rect 326094 264302 326476 264330
rect 326908 264316 326936 269758
rect 327736 267306 327764 273226
rect 331416 272678 331444 278038
rect 331864 274304 331916 274310
rect 331864 274246 331916 274252
rect 331404 272672 331456 272678
rect 331404 272614 331456 272620
rect 329748 272536 329800 272542
rect 329748 272478 329800 272484
rect 329564 271312 329616 271318
rect 329564 271254 329616 271260
rect 327724 267300 327776 267306
rect 327724 267242 327776 267248
rect 327724 266552 327776 266558
rect 327724 266494 327776 266500
rect 327736 264316 327764 266494
rect 328552 266416 328604 266422
rect 328552 266358 328604 266364
rect 328564 264316 328592 266358
rect 329576 264330 329604 271254
rect 329760 266422 329788 272478
rect 331128 271176 331180 271182
rect 331128 271118 331180 271124
rect 330208 269952 330260 269958
rect 330208 269894 330260 269900
rect 329748 266416 329800 266422
rect 329748 266358 329800 266364
rect 329406 264302 329604 264330
rect 330220 264316 330248 269894
rect 331140 267734 331168 271118
rect 331048 267706 331168 267734
rect 331048 264316 331076 267706
rect 331876 266558 331904 274246
rect 332980 272814 333008 278052
rect 333796 272944 333848 272950
rect 333796 272886 333848 272892
rect 332968 272808 333020 272814
rect 332968 272750 333020 272756
rect 332324 272672 332376 272678
rect 332324 272614 332376 272620
rect 331864 266552 331916 266558
rect 331864 266494 331916 266500
rect 332336 264330 332364 272614
rect 332692 266892 332744 266898
rect 332692 266834 332744 266840
rect 331890 264302 332364 264330
rect 332704 264316 332732 266834
rect 333808 264330 333836 272886
rect 334176 271454 334204 278052
rect 335372 275330 335400 278052
rect 335556 278038 336582 278066
rect 335360 275324 335412 275330
rect 335360 275266 335412 275272
rect 335268 273964 335320 273970
rect 335268 273906 335320 273912
rect 334164 271448 334216 271454
rect 334164 271390 334216 271396
rect 334348 270224 334400 270230
rect 334348 270166 334400 270172
rect 333546 264302 333836 264330
rect 334360 264316 334388 270166
rect 335280 267734 335308 273906
rect 335556 269822 335584 278038
rect 337764 274310 337792 278052
rect 337752 274304 337804 274310
rect 337752 274246 337804 274252
rect 337752 274100 337804 274106
rect 337752 274042 337804 274048
rect 335544 269816 335596 269822
rect 335544 269758 335596 269764
rect 336004 269816 336056 269822
rect 336004 269758 336056 269764
rect 335188 267706 335308 267734
rect 335188 264316 335216 267706
rect 336016 264316 336044 269758
rect 337764 267734 337792 274042
rect 338868 272542 338896 278052
rect 338856 272536 338908 272542
rect 338856 272478 338908 272484
rect 339224 272536 339276 272542
rect 339224 272478 339276 272484
rect 337936 271584 337988 271590
rect 337936 271526 337988 271532
rect 337672 267706 337792 267734
rect 336832 266416 336884 266422
rect 336832 266358 336884 266364
rect 336844 264316 336872 266358
rect 337672 264316 337700 267706
rect 337948 266422 337976 271526
rect 338488 268524 338540 268530
rect 338488 268466 338540 268472
rect 337936 266416 337988 266422
rect 337936 266358 337988 266364
rect 338500 264316 338528 268466
rect 339236 264330 339264 272478
rect 340064 271318 340092 278052
rect 340892 278038 341274 278066
rect 340052 271312 340104 271318
rect 340052 271254 340104 271260
rect 340604 271312 340656 271318
rect 340604 271254 340656 271260
rect 340616 264330 340644 271254
rect 340892 269958 340920 278038
rect 342456 271182 342484 278052
rect 343652 272678 343680 278052
rect 343836 278038 344862 278066
rect 343640 272672 343692 272678
rect 343640 272614 343692 272620
rect 342444 271176 342496 271182
rect 342444 271118 342496 271124
rect 343548 271176 343600 271182
rect 343548 271118 343600 271124
rect 340880 269952 340932 269958
rect 340880 269894 340932 269900
rect 341800 269952 341852 269958
rect 341800 269894 341852 269900
rect 340972 267436 341024 267442
rect 340972 267378 341024 267384
rect 339236 264302 339342 264330
rect 340170 264302 340644 264330
rect 340984 264316 341012 267378
rect 341812 264316 341840 269894
rect 343560 267734 343588 271118
rect 343468 267706 343588 267734
rect 342628 266416 342680 266422
rect 342628 266358 342680 266364
rect 342640 264316 342668 266358
rect 343468 264316 343496 267706
rect 343836 266898 343864 278038
rect 345952 272950 345980 278052
rect 346412 278038 347162 278066
rect 345940 272944 345992 272950
rect 345940 272886 345992 272892
rect 344652 272808 344704 272814
rect 344652 272750 344704 272756
rect 343824 266892 343876 266898
rect 343824 266834 343876 266840
rect 344664 264330 344692 272750
rect 346216 272672 346268 272678
rect 346216 272614 346268 272620
rect 345296 270088 345348 270094
rect 345296 270030 345348 270036
rect 345112 266552 345164 266558
rect 345112 266494 345164 266500
rect 344310 264302 344692 264330
rect 345124 264316 345152 266494
rect 345308 266422 345336 270030
rect 345296 266416 345348 266422
rect 345296 266358 345348 266364
rect 346228 264330 346256 272614
rect 346412 270230 346440 278038
rect 348344 273970 348372 278052
rect 349172 278038 349554 278066
rect 348332 273964 348384 273970
rect 348332 273906 348384 273912
rect 348424 272944 348476 272950
rect 348424 272886 348476 272892
rect 347688 271448 347740 271454
rect 347688 271390 347740 271396
rect 346400 270224 346452 270230
rect 346400 270166 346452 270172
rect 347504 266688 347556 266694
rect 347504 266630 347556 266636
rect 346768 266416 346820 266422
rect 346768 266358 346820 266364
rect 345966 264302 346256 264330
rect 346780 264316 346808 266358
rect 347516 264330 347544 266630
rect 347700 266422 347728 271390
rect 348436 266558 348464 272886
rect 349172 269822 349200 278038
rect 350356 273964 350408 273970
rect 350356 273906 350408 273912
rect 349160 269816 349212 269822
rect 349160 269758 349212 269764
rect 348792 268388 348844 268394
rect 348792 268330 348844 268336
rect 348424 266552 348476 266558
rect 348424 266494 348476 266500
rect 347688 266416 347740 266422
rect 347688 266358 347740 266364
rect 348804 264330 348832 268330
rect 350080 266552 350132 266558
rect 350080 266494 350132 266500
rect 349252 266416 349304 266422
rect 349252 266358 349304 266364
rect 347516 264302 347622 264330
rect 348450 264302 348832 264330
rect 349264 264316 349292 266358
rect 350092 264316 350120 266494
rect 350368 266422 350396 273906
rect 350736 271590 350764 278052
rect 351932 274106 351960 278052
rect 352116 278038 353142 278066
rect 351920 274100 351972 274106
rect 351920 274042 351972 274048
rect 351184 271720 351236 271726
rect 351184 271662 351236 271668
rect 350724 271584 350776 271590
rect 350724 271526 350776 271532
rect 350908 267300 350960 267306
rect 350908 267242 350960 267248
rect 350356 266416 350408 266422
rect 350356 266358 350408 266364
rect 350920 264316 350948 267242
rect 351196 266694 351224 271662
rect 351736 269816 351788 269822
rect 351736 269758 351788 269764
rect 351184 266688 351236 266694
rect 351184 266630 351236 266636
rect 351748 264316 351776 269758
rect 352116 268530 352144 278038
rect 353944 274100 353996 274106
rect 353944 274042 353996 274048
rect 352564 268660 352616 268666
rect 352564 268602 352616 268608
rect 352104 268524 352156 268530
rect 352104 268466 352156 268472
rect 352576 264316 352604 268602
rect 353392 267028 353444 267034
rect 353392 266970 353444 266976
rect 353404 264316 353432 266970
rect 353956 266558 353984 274042
rect 354232 272542 354260 278052
rect 355152 278038 355442 278066
rect 354220 272536 354272 272542
rect 354220 272478 354272 272484
rect 354496 272536 354548 272542
rect 354496 272478 354548 272484
rect 353944 266552 353996 266558
rect 353944 266494 353996 266500
rect 354508 264330 354536 272478
rect 355152 271318 355180 278038
rect 356624 271862 356652 278052
rect 357452 278038 357834 278066
rect 358832 278038 359030 278066
rect 355324 271856 355376 271862
rect 355324 271798 355376 271804
rect 356612 271856 356664 271862
rect 356612 271798 356664 271804
rect 355140 271312 355192 271318
rect 355140 271254 355192 271260
rect 355048 270360 355100 270366
rect 355048 270302 355100 270308
rect 354246 264302 354536 264330
rect 355060 264316 355088 270302
rect 355336 267442 355364 271798
rect 357164 271312 357216 271318
rect 357164 271254 357216 271260
rect 355324 267436 355376 267442
rect 355324 267378 355376 267384
rect 355876 266552 355928 266558
rect 355876 266494 355928 266500
rect 355888 264316 355916 266494
rect 357176 264330 357204 271254
rect 357452 269958 357480 278038
rect 358636 275460 358688 275466
rect 358636 275402 358688 275408
rect 357440 269952 357492 269958
rect 357440 269894 357492 269900
rect 357532 266416 357584 266422
rect 357532 266358 357584 266364
rect 356730 264302 357204 264330
rect 357544 264316 357572 266358
rect 358648 264330 358676 275402
rect 358832 270094 358860 278038
rect 359464 274236 359516 274242
rect 359464 274178 359516 274184
rect 358820 270088 358872 270094
rect 358820 270030 358872 270036
rect 359188 269952 359240 269958
rect 359188 269894 359240 269900
rect 358386 264302 358676 264330
rect 359200 264316 359228 269894
rect 359476 266422 359504 274178
rect 360212 271182 360240 278052
rect 361212 273080 361264 273086
rect 361212 273022 361264 273028
rect 360844 271584 360896 271590
rect 360844 271526 360896 271532
rect 360200 271176 360252 271182
rect 360200 271118 360252 271124
rect 360016 267164 360068 267170
rect 360016 267106 360068 267112
rect 359464 266416 359516 266422
rect 359464 266358 359516 266364
rect 360028 264316 360056 267106
rect 360856 266558 360884 271526
rect 360844 266552 360896 266558
rect 360844 266494 360896 266500
rect 361224 264330 361252 273022
rect 361408 272814 361436 278052
rect 362512 272950 362540 278052
rect 362776 273216 362828 273222
rect 362776 273158 362828 273164
rect 362500 272944 362552 272950
rect 362500 272886 362552 272892
rect 361396 272808 361448 272814
rect 361396 272750 361448 272756
rect 362224 272808 362276 272814
rect 362224 272750 362276 272756
rect 362236 267306 362264 272750
rect 362500 267436 362552 267442
rect 362500 267378 362552 267384
rect 362224 267300 362276 267306
rect 362224 267242 362276 267248
rect 361672 266416 361724 266422
rect 361672 266358 361724 266364
rect 360870 264302 361252 264330
rect 361684 264316 361712 266358
rect 362512 264316 362540 267378
rect 362788 266422 362816 273158
rect 363708 272678 363736 278052
rect 363880 275596 363932 275602
rect 363880 275538 363932 275544
rect 363696 272672 363748 272678
rect 363696 272614 363748 272620
rect 363892 267734 363920 275538
rect 364904 271454 364932 278052
rect 365444 272944 365496 272950
rect 365444 272886 365496 272892
rect 364892 271448 364944 271454
rect 364892 271390 364944 271396
rect 364156 271176 364208 271182
rect 364156 271118 364208 271124
rect 363800 267706 363920 267734
rect 362776 266416 362828 266422
rect 362776 266358 362828 266364
rect 363800 264330 363828 267706
rect 363354 264302 363828 264330
rect 364168 264316 364196 271118
rect 365456 264330 365484 272886
rect 366100 271726 366128 278052
rect 367112 278038 367310 278066
rect 366088 271720 366140 271726
rect 366088 271662 366140 271668
rect 366364 271448 366416 271454
rect 366364 271390 366416 271396
rect 365812 267708 365864 267714
rect 365812 267650 365864 267656
rect 365010 264302 365484 264330
rect 365824 264316 365852 267650
rect 366376 267170 366404 271390
rect 366640 270088 366692 270094
rect 366640 270030 366692 270036
rect 366364 267164 366416 267170
rect 366364 267106 366416 267112
rect 366652 264316 366680 270030
rect 367112 268394 367140 278038
rect 368492 273970 368520 278052
rect 369124 274372 369176 274378
rect 369124 274314 369176 274320
rect 368480 273964 368532 273970
rect 368480 273906 368532 273912
rect 367468 268524 367520 268530
rect 367468 268466 367520 268472
rect 367100 268388 367152 268394
rect 367100 268330 367152 268336
rect 367480 264316 367508 268466
rect 369136 267442 369164 274314
rect 369596 274106 369624 278052
rect 370332 278038 370806 278066
rect 371252 278038 372002 278066
rect 372632 278038 373198 278066
rect 369584 274100 369636 274106
rect 369584 274042 369636 274048
rect 370332 272814 370360 278038
rect 371056 275324 371108 275330
rect 371056 275266 371108 275272
rect 370320 272808 370372 272814
rect 370320 272750 370372 272756
rect 370504 272808 370556 272814
rect 370504 272750 370556 272756
rect 369124 267436 369176 267442
rect 369124 267378 369176 267384
rect 368296 266892 368348 266898
rect 368296 266834 368348 266840
rect 368308 264316 368336 266834
rect 369952 266552 370004 266558
rect 369952 266494 370004 266500
rect 369124 266416 369176 266422
rect 369124 266358 369176 266364
rect 369136 264316 369164 266358
rect 369964 264316 369992 266494
rect 370516 266422 370544 272750
rect 370504 266416 370556 266422
rect 370504 266358 370556 266364
rect 371068 264330 371096 275266
rect 371252 269822 371280 278038
rect 372252 270224 372304 270230
rect 372252 270166 372304 270172
rect 371240 269816 371292 269822
rect 371240 269758 371292 269764
rect 371608 267572 371660 267578
rect 371608 267514 371660 267520
rect 370806 264302 371096 264330
rect 371620 264316 371648 267514
rect 372264 266558 372292 270166
rect 372632 268666 372660 278038
rect 374380 277394 374408 278052
rect 374380 277366 374500 277394
rect 373264 274100 373316 274106
rect 373264 274042 373316 274048
rect 372620 268660 372672 268666
rect 372620 268602 372672 268608
rect 372436 268388 372488 268394
rect 372436 268330 372488 268336
rect 372252 266552 372304 266558
rect 372252 266494 372304 266500
rect 372448 264316 372476 268330
rect 373276 267578 373304 274042
rect 373264 267572 373316 267578
rect 373264 267514 373316 267520
rect 374472 267442 374500 277366
rect 375576 272542 375604 278052
rect 376786 278038 376984 278066
rect 376116 272672 376168 272678
rect 376116 272614 376168 272620
rect 375564 272536 375616 272542
rect 375564 272478 375616 272484
rect 375288 271856 375340 271862
rect 375288 271798 375340 271804
rect 374460 267436 374512 267442
rect 374460 267378 374512 267384
rect 373264 267300 373316 267306
rect 373264 267242 373316 267248
rect 373276 264316 373304 267242
rect 374920 266552 374972 266558
rect 374920 266494 374972 266500
rect 374092 266416 374144 266422
rect 374092 266358 374144 266364
rect 374104 264316 374132 266358
rect 374932 264316 374960 266494
rect 375300 266422 375328 271798
rect 375288 266416 375340 266422
rect 375288 266358 375340 266364
rect 376128 264330 376156 272614
rect 376956 270366 376984 278038
rect 377600 278038 377890 278066
rect 377600 271590 377628 278038
rect 377772 273964 377824 273970
rect 377772 273906 377824 273912
rect 377588 271584 377640 271590
rect 377588 271526 377640 271532
rect 376944 270360 376996 270366
rect 376944 270302 376996 270308
rect 376576 269816 376628 269822
rect 376576 269758 376628 269764
rect 375774 264302 376156 264330
rect 376588 264316 376616 269758
rect 377784 264330 377812 273906
rect 379072 271318 379100 278052
rect 380268 274242 380296 278052
rect 381464 275466 381492 278052
rect 382292 278038 382674 278066
rect 381452 275460 381504 275466
rect 381452 275402 381504 275408
rect 381544 274508 381596 274514
rect 381544 274450 381596 274456
rect 380256 274236 380308 274242
rect 380256 274178 380308 274184
rect 379428 272536 379480 272542
rect 379428 272478 379480 272484
rect 379060 271312 379112 271318
rect 379060 271254 379112 271260
rect 378232 266892 378284 266898
rect 378232 266834 378284 266840
rect 377430 264302 377812 264330
rect 378244 264316 378272 266834
rect 379440 264330 379468 272478
rect 379704 270360 379756 270366
rect 379704 270302 379756 270308
rect 379716 266558 379744 270302
rect 381556 267714 381584 274450
rect 382004 271720 382056 271726
rect 382004 271662 382056 271668
rect 381544 267708 381596 267714
rect 381544 267650 381596 267656
rect 380716 267436 380768 267442
rect 380716 267378 380768 267384
rect 379704 266552 379756 266558
rect 379704 266494 379756 266500
rect 379888 266416 379940 266422
rect 379888 266358 379940 266364
rect 379086 264302 379468 264330
rect 379900 264316 379928 266358
rect 380728 264316 380756 267378
rect 382016 264330 382044 271662
rect 382292 269958 382320 278038
rect 383856 271454 383884 278052
rect 385052 274666 385080 278052
rect 384960 274638 385080 274666
rect 385880 278038 386170 278066
rect 384960 273086 384988 274638
rect 385880 273222 385908 278038
rect 386052 275460 386104 275466
rect 386052 275402 386104 275408
rect 385868 273216 385920 273222
rect 385868 273158 385920 273164
rect 384948 273080 385000 273086
rect 384948 273022 385000 273028
rect 385684 273080 385736 273086
rect 385684 273022 385736 273028
rect 384948 272128 385000 272134
rect 384948 272070 385000 272076
rect 383844 271448 383896 271454
rect 383844 271390 383896 271396
rect 384764 271448 384816 271454
rect 384764 271390 384816 271396
rect 382280 269952 382332 269958
rect 382280 269894 382332 269900
rect 383016 269952 383068 269958
rect 383016 269894 383068 269900
rect 382372 268932 382424 268938
rect 382372 268874 382424 268880
rect 381570 264302 382044 264330
rect 382384 264316 382412 268874
rect 383028 266422 383056 269894
rect 383200 267028 383252 267034
rect 383200 266970 383252 266976
rect 383016 266416 383068 266422
rect 383016 266358 383068 266364
rect 383212 264316 383240 266970
rect 384028 266416 384080 266422
rect 384028 266358 384080 266364
rect 384040 264316 384068 266358
rect 384776 264330 384804 271390
rect 384960 266422 384988 272070
rect 385696 267170 385724 273022
rect 385684 267164 385736 267170
rect 385684 267106 385736 267112
rect 384948 266416 385000 266422
rect 384948 266358 385000 266364
rect 386064 264330 386092 275402
rect 387352 274378 387380 278052
rect 388548 275602 388576 278052
rect 388536 275596 388588 275602
rect 388536 275538 388588 275544
rect 387340 274372 387392 274378
rect 387340 274314 387392 274320
rect 388996 274236 389048 274242
rect 388996 274178 389048 274184
rect 387708 271584 387760 271590
rect 387708 271526 387760 271532
rect 387340 268796 387392 268802
rect 387340 268738 387392 268744
rect 386512 266416 386564 266422
rect 386512 266358 386564 266364
rect 384776 264302 384882 264330
rect 385710 264302 386092 264330
rect 386524 264316 386552 266358
rect 387352 264316 387380 268738
rect 387720 266422 387748 271526
rect 388168 267708 388220 267714
rect 388168 267650 388220 267656
rect 387708 266416 387760 266422
rect 387708 266358 387760 266364
rect 388180 264316 388208 267650
rect 389008 264316 389036 274178
rect 389744 271182 389772 278052
rect 390940 272950 390968 278052
rect 392136 274514 392164 278052
rect 392124 274508 392176 274514
rect 392124 274450 392176 274456
rect 390928 272944 390980 272950
rect 390928 272886 390980 272892
rect 391848 272264 391900 272270
rect 391848 272206 391900 272212
rect 390284 271312 390336 271318
rect 390284 271254 390336 271260
rect 389732 271176 389784 271182
rect 389732 271118 389784 271124
rect 390296 264330 390324 271254
rect 390652 267572 390704 267578
rect 390652 267514 390704 267520
rect 389850 264302 390324 264330
rect 390664 264316 390692 267514
rect 391860 264330 391888 272206
rect 393332 270094 393360 278052
rect 393516 278038 394450 278066
rect 393320 270088 393372 270094
rect 393320 270030 393372 270036
rect 392032 269680 392084 269686
rect 392032 269622 392084 269628
rect 392044 267306 392072 269622
rect 393516 268530 393544 278038
rect 395632 273086 395660 278052
rect 395620 273080 395672 273086
rect 395620 273022 395672 273028
rect 396828 272814 396856 278052
rect 397472 278038 398038 278066
rect 397000 273828 397052 273834
rect 397000 273770 397052 273776
rect 396816 272808 396868 272814
rect 396816 272750 396868 272756
rect 395988 272400 396040 272406
rect 395988 272342 396040 272348
rect 394332 271176 394384 271182
rect 394332 271118 394384 271124
rect 393688 268660 393740 268666
rect 393688 268602 393740 268608
rect 393504 268524 393556 268530
rect 393504 268466 393556 268472
rect 392032 267300 392084 267306
rect 392032 267242 392084 267248
rect 393136 267164 393188 267170
rect 393136 267106 393188 267112
rect 392308 266416 392360 266422
rect 392308 266358 392360 266364
rect 391506 264302 391888 264330
rect 392320 264316 392348 266358
rect 393148 264316 393176 267106
rect 393700 266422 393728 268602
rect 393688 266416 393740 266422
rect 393688 266358 393740 266364
rect 394344 264330 394372 271118
rect 394700 270088 394752 270094
rect 394700 270030 394752 270036
rect 394712 266898 394740 270030
rect 394700 266892 394752 266898
rect 394700 266834 394752 266840
rect 394792 266756 394844 266762
rect 394792 266698 394844 266704
rect 393990 264302 394372 264330
rect 394804 264316 394832 266698
rect 396000 264330 396028 272342
rect 397012 267734 397040 273770
rect 397472 270230 397500 278038
rect 399220 275330 399248 278052
rect 399208 275324 399260 275330
rect 399208 275266 399260 275272
rect 400324 274106 400352 278052
rect 400508 278038 401534 278066
rect 401704 278038 402730 278066
rect 400312 274100 400364 274106
rect 400312 274042 400364 274048
rect 400036 273216 400088 273222
rect 400036 273158 400088 273164
rect 397460 270224 397512 270230
rect 397460 270166 397512 270172
rect 398748 269544 398800 269550
rect 398748 269486 398800 269492
rect 397276 268524 397328 268530
rect 397276 268466 397328 268472
rect 396920 267706 397040 267734
rect 396920 264330 396948 267706
rect 395646 264302 396028 264330
rect 396474 264302 396948 264330
rect 397288 264316 397316 268466
rect 398760 267442 398788 269486
rect 398748 267436 398800 267442
rect 398748 267378 398800 267384
rect 398104 267300 398156 267306
rect 398104 267242 398156 267248
rect 398116 264316 398144 267242
rect 399760 266620 399812 266626
rect 399760 266562 399812 266568
rect 398932 266416 398984 266422
rect 398932 266358 398984 266364
rect 398944 264316 398972 266358
rect 399772 264316 399800 266562
rect 400048 266422 400076 273158
rect 400508 268394 400536 278038
rect 401508 274100 401560 274106
rect 401508 274042 401560 274048
rect 400864 270496 400916 270502
rect 400864 270438 400916 270444
rect 400496 268388 400548 268394
rect 400496 268330 400548 268336
rect 400036 266416 400088 266422
rect 400036 266358 400088 266364
rect 400876 264330 400904 270438
rect 401520 267734 401548 274042
rect 401704 269686 401732 278038
rect 403912 271862 403940 278052
rect 404372 278038 405122 278066
rect 404176 273080 404228 273086
rect 404176 273022 404228 273028
rect 403900 271856 403952 271862
rect 403900 271798 403952 271804
rect 403624 270632 403676 270638
rect 403624 270574 403676 270580
rect 401692 269680 401744 269686
rect 401692 269622 401744 269628
rect 401692 269272 401744 269278
rect 401692 269214 401744 269220
rect 400614 264302 400904 264330
rect 401428 267706 401548 267734
rect 401428 264316 401456 267706
rect 401704 267034 401732 269214
rect 402244 268388 402296 268394
rect 402244 268330 402296 268336
rect 401692 267028 401744 267034
rect 401692 266970 401744 266976
rect 402256 264316 402284 268330
rect 403072 267436 403124 267442
rect 403072 267378 403124 267384
rect 403084 264316 403112 267378
rect 403636 266762 403664 270574
rect 403624 266756 403676 266762
rect 403624 266698 403676 266704
rect 404188 264330 404216 273022
rect 404372 270366 404400 278038
rect 405556 272944 405608 272950
rect 405556 272886 405608 272892
rect 404360 270360 404412 270366
rect 404360 270302 404412 270308
rect 404360 269680 404412 269686
rect 404360 269622 404412 269628
rect 404372 267714 404400 269622
rect 404360 267708 404412 267714
rect 404360 267650 404412 267656
rect 404728 266892 404780 266898
rect 404728 266834 404780 266840
rect 403926 264302 404216 264330
rect 404740 264316 404768 266834
rect 405568 264316 405596 272886
rect 406304 272678 406332 278052
rect 407132 278038 407514 278066
rect 406844 272808 406896 272814
rect 406844 272750 406896 272756
rect 406292 272672 406344 272678
rect 406292 272614 406344 272620
rect 406856 264330 406884 272750
rect 407132 269822 407160 278038
rect 408604 273970 408632 278052
rect 408788 278038 409814 278066
rect 408592 273964 408644 273970
rect 408592 273906 408644 273912
rect 407764 270904 407816 270910
rect 407764 270846 407816 270852
rect 407120 269816 407172 269822
rect 407120 269758 407172 269764
rect 407212 266756 407264 266762
rect 407212 266698 407264 266704
rect 406410 264302 406884 264330
rect 407224 264316 407252 266698
rect 407776 266626 407804 270846
rect 408788 270094 408816 278038
rect 410800 276004 410852 276010
rect 410800 275946 410852 275952
rect 409788 274644 409840 274650
rect 409788 274586 409840 274592
rect 409604 270224 409656 270230
rect 409604 270166 409656 270172
rect 408776 270088 408828 270094
rect 408776 270030 408828 270036
rect 408408 269408 408460 269414
rect 408408 269350 408460 269356
rect 408040 267708 408092 267714
rect 408040 267650 408092 267656
rect 407764 266620 407816 266626
rect 407764 266562 407816 266568
rect 408052 264316 408080 267650
rect 408420 267578 408448 269350
rect 408408 267572 408460 267578
rect 408408 267514 408460 267520
rect 408868 266416 408920 266422
rect 408868 266358 408920 266364
rect 408880 264316 408908 266358
rect 409616 264330 409644 270166
rect 409800 266422 409828 274586
rect 409788 266416 409840 266422
rect 409788 266358 409840 266364
rect 410812 264330 410840 275946
rect 410996 272542 411024 278052
rect 411272 278038 412206 278066
rect 412652 278038 413402 278066
rect 410984 272536 411036 272542
rect 410984 272478 411036 272484
rect 411272 269958 411300 278038
rect 412272 272672 412324 272678
rect 412272 272614 412324 272620
rect 411260 269952 411312 269958
rect 411260 269894 411312 269900
rect 412284 266422 412312 272614
rect 412456 270088 412508 270094
rect 412456 270030 412508 270036
rect 411352 266416 411404 266422
rect 411352 266358 411404 266364
rect 412272 266416 412324 266422
rect 412272 266358 412324 266364
rect 409616 264302 409722 264330
rect 410550 264302 410840 264330
rect 411364 264316 411392 266358
rect 412468 264330 412496 270030
rect 412652 269550 412680 278038
rect 413836 274508 413888 274514
rect 413836 274450 413888 274456
rect 412640 269544 412692 269550
rect 412640 269486 412692 269492
rect 413008 267028 413060 267034
rect 413008 266970 413060 266976
rect 412206 264302 412496 264330
rect 413020 264316 413048 266970
rect 413848 264316 413876 274450
rect 414584 271726 414612 278052
rect 415412 278038 415794 278066
rect 416792 278038 416898 278066
rect 414572 271720 414624 271726
rect 414572 271662 414624 271668
rect 414664 270768 414716 270774
rect 414664 270710 414716 270716
rect 414676 266762 414704 270710
rect 415032 270360 415084 270366
rect 415032 270302 415084 270308
rect 414664 266756 414716 266762
rect 414664 266698 414716 266704
rect 415044 264330 415072 270302
rect 415412 268938 415440 278038
rect 416412 275732 416464 275738
rect 416412 275674 416464 275680
rect 415400 268932 415452 268938
rect 415400 268874 415452 268880
rect 416228 268252 416280 268258
rect 416228 268194 416280 268200
rect 416240 266898 416268 268194
rect 416228 266892 416280 266898
rect 416228 266834 416280 266840
rect 416424 266422 416452 275674
rect 416596 272536 416648 272542
rect 416596 272478 416648 272484
rect 415492 266416 415544 266422
rect 415492 266358 415544 266364
rect 416412 266416 416464 266422
rect 416412 266358 416464 266364
rect 414690 264302 415072 264330
rect 415504 264316 415532 266358
rect 416608 264330 416636 272478
rect 416792 269278 416820 278038
rect 418080 272134 418108 278052
rect 418804 275324 418856 275330
rect 418804 275266 418856 275272
rect 418068 272128 418120 272134
rect 418068 272070 418120 272076
rect 417424 271040 417476 271046
rect 417424 270982 417476 270988
rect 417148 269816 417200 269822
rect 417148 269758 417200 269764
rect 416780 269272 416832 269278
rect 416780 269214 416832 269220
rect 416346 264302 416636 264330
rect 417160 264316 417188 269758
rect 417436 267306 417464 270982
rect 417424 267300 417476 267306
rect 417424 267242 417476 267248
rect 418816 266422 418844 275266
rect 419080 274372 419132 274378
rect 419080 274314 419132 274320
rect 417976 266416 418028 266422
rect 417976 266358 418028 266364
rect 418804 266416 418856 266422
rect 418804 266358 418856 266364
rect 417988 264316 418016 266358
rect 419092 264330 419120 274314
rect 419276 271454 419304 278052
rect 420472 275466 420500 278052
rect 420460 275460 420512 275466
rect 420460 275402 420512 275408
rect 420552 275052 420604 275058
rect 420552 274994 420604 275000
rect 419264 271448 419316 271454
rect 419264 271390 419316 271396
rect 420184 271448 420236 271454
rect 420184 271390 420236 271396
rect 419632 269952 419684 269958
rect 419632 269894 419684 269900
rect 418830 264302 419120 264330
rect 419644 264316 419672 269894
rect 420196 267170 420224 271390
rect 420564 267734 420592 274994
rect 421668 271590 421696 278052
rect 422312 278038 422878 278066
rect 423692 278038 423982 278066
rect 422116 273964 422168 273970
rect 422116 273906 422168 273912
rect 421656 271584 421708 271590
rect 421656 271526 421708 271532
rect 420472 267706 420592 267734
rect 420184 267164 420236 267170
rect 420184 267106 420236 267112
rect 420472 264316 420500 267706
rect 421288 267572 421340 267578
rect 421288 267514 421340 267520
rect 421300 264316 421328 267514
rect 422128 264316 422156 273906
rect 422312 268802 422340 278038
rect 423692 269686 423720 278038
rect 425164 274242 425192 278052
rect 425152 274236 425204 274242
rect 425152 274178 425204 274184
rect 425704 274236 425756 274242
rect 425704 274178 425756 274184
rect 423680 269680 423732 269686
rect 423680 269622 423732 269628
rect 423864 269680 423916 269686
rect 423864 269622 423916 269628
rect 422300 268796 422352 268802
rect 422300 268738 422352 268744
rect 422300 268116 422352 268122
rect 422300 268058 422352 268064
rect 422312 267442 422340 268058
rect 423876 267714 423904 269622
rect 424600 269544 424652 269550
rect 424600 269486 424652 269492
rect 423864 267708 423916 267714
rect 423864 267650 423916 267656
rect 422300 267436 422352 267442
rect 422300 267378 422352 267384
rect 422944 266892 422996 266898
rect 422944 266834 422996 266840
rect 422956 264316 422984 266834
rect 423772 266552 423824 266558
rect 423772 266494 423824 266500
rect 423784 264316 423812 266494
rect 424612 264316 424640 269486
rect 425716 266558 425744 274178
rect 426360 271318 426388 278052
rect 426544 278038 427570 278066
rect 426348 271312 426400 271318
rect 426348 271254 426400 271260
rect 426544 269414 426572 278038
rect 427084 275188 427136 275194
rect 427084 275130 427136 275136
rect 426532 269408 426584 269414
rect 426532 269350 426584 269356
rect 425704 266552 425756 266558
rect 425704 266494 425756 266500
rect 426256 266552 426308 266558
rect 426256 266494 426308 266500
rect 425428 266416 425480 266422
rect 425428 266358 425480 266364
rect 425440 264316 425468 266358
rect 426268 264316 426296 266494
rect 427096 266422 427124 275130
rect 428752 272270 428780 278052
rect 429212 278038 429962 278066
rect 428740 272264 428792 272270
rect 428740 272206 428792 272212
rect 428464 272128 428516 272134
rect 428464 272070 428516 272076
rect 427452 271040 427504 271046
rect 427452 270982 427504 270988
rect 427084 266416 427136 266422
rect 427084 266358 427136 266364
rect 427464 264330 427492 270982
rect 427912 266688 427964 266694
rect 427912 266630 427964 266636
rect 427110 264302 427492 264330
rect 427924 264316 427952 266630
rect 428476 266558 428504 272070
rect 429212 268666 429240 278038
rect 430212 275868 430264 275874
rect 430212 275810 430264 275816
rect 429200 268660 429252 268666
rect 429200 268602 429252 268608
rect 428740 267436 428792 267442
rect 428740 267378 428792 267384
rect 428464 266552 428516 266558
rect 428464 266494 428516 266500
rect 428752 264316 428780 267378
rect 429568 266416 429620 266422
rect 429568 266358 429620 266364
rect 429580 264316 429608 266358
rect 430224 264330 430252 275810
rect 430396 271720 430448 271726
rect 430396 271662 430448 271668
rect 430408 266422 430436 271662
rect 431144 271454 431172 278052
rect 431684 271992 431736 271998
rect 431684 271934 431736 271940
rect 431132 271448 431184 271454
rect 431132 271390 431184 271396
rect 430396 266416 430448 266422
rect 430396 266358 430448 266364
rect 431696 264330 431724 271934
rect 432248 271318 432276 278052
rect 433156 271856 433208 271862
rect 433156 271798 433208 271804
rect 432236 271312 432288 271318
rect 432236 271254 432288 271260
rect 432880 267164 432932 267170
rect 432880 267106 432932 267112
rect 432052 266416 432104 266422
rect 432052 266358 432104 266364
rect 430224 264302 430422 264330
rect 431250 264302 431724 264330
rect 432064 264316 432092 266358
rect 432892 264316 432920 267106
rect 433168 266422 433196 271798
rect 433444 270638 433472 278052
rect 434640 272406 434668 278052
rect 435640 275460 435692 275466
rect 435640 275402 435692 275408
rect 434628 272400 434680 272406
rect 434628 272342 434680 272348
rect 433432 270632 433484 270638
rect 433432 270574 433484 270580
rect 433708 269068 433760 269074
rect 433708 269010 433760 269016
rect 433156 266416 433208 266422
rect 433156 266358 433208 266364
rect 433720 264316 433748 269010
rect 434536 266552 434588 266558
rect 434536 266494 434588 266500
rect 434548 264316 434576 266494
rect 435652 264330 435680 275402
rect 435836 273834 435864 278052
rect 436112 278038 437046 278066
rect 437952 278038 438242 278066
rect 435824 273828 435876 273834
rect 435824 273770 435876 273776
rect 436112 268530 436140 278038
rect 437204 271584 437256 271590
rect 437204 271526 437256 271532
rect 436560 268932 436612 268938
rect 436560 268874 436612 268880
rect 436100 268524 436152 268530
rect 436100 268466 436152 268472
rect 436572 264330 436600 268874
rect 436744 267300 436796 267306
rect 436744 267242 436796 267248
rect 436756 266694 436784 267242
rect 436744 266688 436796 266694
rect 436744 266630 436796 266636
rect 437216 264330 437244 271526
rect 437952 271182 437980 278038
rect 438124 273828 438176 273834
rect 438124 273770 438176 273776
rect 437940 271176 437992 271182
rect 437940 271118 437992 271124
rect 438136 266898 438164 273770
rect 439332 273222 439360 278052
rect 439320 273216 439372 273222
rect 439320 273158 439372 273164
rect 439964 271448 440016 271454
rect 439964 271390 440016 271396
rect 438676 268796 438728 268802
rect 438676 268738 438728 268744
rect 438124 266892 438176 266898
rect 438124 266834 438176 266840
rect 437848 266552 437900 266558
rect 437848 266494 437900 266500
rect 435390 264302 435680 264330
rect 436218 264302 436600 264330
rect 437046 264302 437244 264330
rect 437860 264316 437888 266494
rect 438688 264316 438716 268738
rect 439976 264330 440004 271390
rect 440528 270910 440556 278052
rect 441724 277394 441752 278052
rect 441632 277366 441752 277394
rect 440884 273556 440936 273562
rect 440884 273498 440936 273504
rect 440516 270904 440568 270910
rect 440516 270846 440568 270852
rect 440896 267578 440924 273498
rect 441344 271176 441396 271182
rect 441344 271118 441396 271124
rect 441160 268660 441212 268666
rect 441160 268602 441212 268608
rect 440884 267572 440936 267578
rect 440884 267514 440936 267520
rect 440332 266416 440384 266422
rect 440332 266358 440384 266364
rect 439530 264302 440004 264330
rect 440344 264316 440372 266358
rect 441172 264316 441200 268602
rect 441356 266422 441384 271118
rect 441632 270502 441660 277366
rect 442920 274106 442948 278052
rect 443104 278038 444130 278066
rect 444392 278038 445326 278066
rect 442908 274100 442960 274106
rect 442908 274042 442960 274048
rect 442908 271312 442960 271318
rect 442908 271254 442960 271260
rect 441620 270496 441672 270502
rect 441620 270438 441672 270444
rect 441620 269408 441672 269414
rect 441620 269350 441672 269356
rect 441632 266898 441660 269350
rect 441620 266892 441672 266898
rect 441620 266834 441672 266840
rect 442724 266892 442776 266898
rect 442724 266834 442776 266840
rect 441344 266416 441396 266422
rect 441344 266358 441396 266364
rect 441988 266416 442040 266422
rect 441988 266358 442040 266364
rect 442000 264316 442028 266358
rect 442736 264330 442764 266834
rect 442920 266422 442948 271254
rect 443104 268394 443132 278038
rect 444012 273216 444064 273222
rect 444012 273158 444064 273164
rect 443092 268388 443144 268394
rect 443092 268330 443144 268336
rect 442908 266416 442960 266422
rect 442908 266358 442960 266364
rect 444024 264330 444052 273158
rect 444392 268122 444420 278038
rect 445024 275596 445076 275602
rect 445024 275538 445076 275544
rect 445036 271182 445064 275538
rect 446508 273086 446536 278052
rect 447152 278038 447626 278066
rect 446496 273080 446548 273086
rect 446496 273022 446548 273028
rect 446864 273080 446916 273086
rect 446864 273022 446916 273028
rect 445024 271176 445076 271182
rect 445024 271118 445076 271124
rect 445668 271176 445720 271182
rect 445668 271118 445720 271124
rect 444380 268116 444432 268122
rect 444380 268058 444432 268064
rect 445300 267708 445352 267714
rect 445300 267650 445352 267656
rect 444472 266416 444524 266422
rect 444472 266358 444524 266364
rect 442736 264302 442842 264330
rect 443670 264302 444052 264330
rect 444484 264316 444512 266358
rect 445312 264316 445340 267650
rect 445680 266422 445708 271118
rect 446128 268524 446180 268530
rect 446128 268466 446180 268472
rect 445668 266416 445720 266422
rect 445668 266358 445720 266364
rect 446140 264316 446168 268466
rect 446876 264330 446904 273022
rect 447152 268258 447180 278038
rect 447600 273692 447652 273698
rect 447600 273634 447652 273640
rect 447140 268252 447192 268258
rect 447140 268194 447192 268200
rect 447612 267442 447640 273634
rect 448808 272950 448836 278052
rect 448796 272944 448848 272950
rect 448796 272886 448848 272892
rect 450004 272814 450032 278052
rect 450832 278038 451214 278066
rect 451384 278038 452410 278066
rect 449992 272808 450044 272814
rect 449992 272750 450044 272756
rect 449716 272400 449768 272406
rect 449716 272342 449768 272348
rect 449164 270904 449216 270910
rect 449164 270846 449216 270852
rect 448428 268252 448480 268258
rect 448428 268194 448480 268200
rect 447784 267572 447836 267578
rect 447784 267514 447836 267520
rect 447600 267436 447652 267442
rect 447600 267378 447652 267384
rect 446876 264302 446982 264330
rect 447796 264316 447824 267514
rect 448440 266558 448468 268194
rect 449176 266762 449204 270846
rect 449164 266756 449216 266762
rect 449164 266698 449216 266704
rect 448428 266552 448480 266558
rect 448428 266494 448480 266500
rect 448612 266416 448664 266422
rect 448612 266358 448664 266364
rect 448624 264316 448652 266358
rect 449728 264330 449756 272342
rect 450544 272264 450596 272270
rect 450544 272206 450596 272212
rect 450268 267436 450320 267442
rect 450268 267378 450320 267384
rect 449466 264302 449756 264330
rect 450280 264316 450308 267378
rect 450556 266422 450584 272206
rect 450832 270774 450860 278038
rect 451188 274100 451240 274106
rect 451188 274042 451240 274048
rect 450820 270768 450872 270774
rect 450820 270710 450872 270716
rect 451200 267734 451228 274042
rect 451384 269686 451412 278038
rect 453592 274650 453620 278052
rect 454052 278038 454710 278066
rect 453580 274644 453632 274650
rect 453580 274586 453632 274592
rect 452292 272808 452344 272814
rect 452292 272750 452344 272756
rect 451372 269680 451424 269686
rect 451372 269622 451424 269628
rect 451108 267706 451228 267734
rect 450544 266416 450596 266422
rect 450544 266358 450596 266364
rect 451108 264316 451136 267706
rect 452304 264330 452332 272750
rect 453304 270632 453356 270638
rect 453304 270574 453356 270580
rect 453316 267170 453344 270574
rect 454052 270230 454080 278038
rect 455892 276010 455920 278052
rect 456812 278038 457102 278066
rect 455880 276004 455932 276010
rect 455880 275946 455932 275952
rect 456064 276004 456116 276010
rect 456064 275946 456116 275952
rect 455328 272944 455380 272950
rect 455328 272886 455380 272892
rect 454040 270224 454092 270230
rect 454040 270166 454092 270172
rect 453580 269680 453632 269686
rect 453580 269622 453632 269628
rect 453304 267164 453356 267170
rect 453304 267106 453356 267112
rect 452752 266620 452804 266626
rect 452752 266562 452804 266568
rect 451950 264302 452332 264330
rect 452764 264316 452792 266562
rect 453592 264316 453620 269622
rect 455144 267164 455196 267170
rect 455144 267106 455196 267112
rect 454408 266416 454460 266422
rect 454408 266358 454460 266364
rect 454420 264316 454448 266358
rect 455156 264330 455184 267106
rect 455340 266422 455368 272886
rect 456076 267578 456104 275946
rect 456812 272678 456840 278038
rect 458284 277394 458312 278052
rect 458192 277366 458312 277394
rect 458468 278038 459494 278066
rect 457444 274644 457496 274650
rect 457444 274586 457496 274592
rect 456800 272672 456852 272678
rect 456800 272614 456852 272620
rect 457168 272672 457220 272678
rect 457168 272614 457220 272620
rect 456432 270496 456484 270502
rect 456432 270438 456484 270444
rect 456064 267572 456116 267578
rect 456064 267514 456116 267520
rect 455328 266416 455380 266422
rect 455328 266358 455380 266364
rect 456444 264330 456472 270438
rect 457180 264330 457208 272614
rect 457456 267306 457484 274586
rect 458192 270094 458220 277366
rect 458180 270088 458232 270094
rect 458180 270030 458232 270036
rect 458468 269414 458496 278038
rect 460676 274514 460704 278052
rect 461228 278038 461886 278066
rect 460664 274508 460716 274514
rect 460664 274450 460716 274456
rect 461030 272912 461086 272921
rect 461030 272847 461086 272856
rect 461044 272678 461072 272847
rect 461032 272672 461084 272678
rect 460846 272640 460902 272649
rect 461032 272614 461084 272620
rect 460846 272575 460902 272584
rect 458824 270224 458876 270230
rect 458824 270166 458876 270172
rect 458456 269408 458508 269414
rect 458456 269350 458508 269356
rect 457444 267300 457496 267306
rect 457444 267242 457496 267248
rect 457720 266756 457772 266762
rect 457720 266698 457772 266704
rect 455156 264302 455262 264330
rect 456090 264302 456472 264330
rect 456918 264302 457208 264330
rect 457732 264316 457760 266698
rect 458836 264330 458864 270166
rect 460204 267572 460256 267578
rect 460204 267514 460256 267520
rect 459376 267300 459428 267306
rect 459376 267242 459428 267248
rect 458574 264302 458864 264330
rect 459388 264316 459416 267242
rect 460216 264316 460244 267514
rect 460860 267306 460888 272575
rect 461228 270366 461256 278038
rect 462976 275738 463004 278052
rect 463712 278038 464186 278066
rect 465092 278038 465382 278066
rect 462964 275732 463016 275738
rect 462964 275674 463016 275680
rect 463148 275732 463200 275738
rect 463148 275674 463200 275680
rect 463160 274666 463188 275674
rect 462976 274638 463188 274666
rect 461400 272944 461452 272950
rect 461400 272886 461452 272892
rect 461412 272678 461440 272886
rect 461400 272672 461452 272678
rect 461860 272672 461912 272678
rect 461400 272614 461452 272620
rect 461858 272640 461860 272649
rect 461912 272640 461914 272649
rect 461858 272575 461914 272584
rect 461216 270360 461268 270366
rect 461216 270302 461268 270308
rect 461400 270360 461452 270366
rect 461400 270302 461452 270308
rect 460848 267300 460900 267306
rect 460848 267242 460900 267248
rect 461412 264330 461440 270302
rect 461860 268388 461912 268394
rect 461860 268330 461912 268336
rect 461058 264302 461440 264330
rect 461872 264316 461900 268330
rect 462976 266626 463004 274638
rect 463240 274508 463292 274514
rect 463240 274450 463292 274456
rect 463252 273254 463280 274450
rect 463160 273226 463280 273254
rect 462964 266620 463016 266626
rect 462964 266562 463016 266568
rect 463160 264330 463188 273226
rect 463712 272542 463740 278038
rect 463700 272536 463752 272542
rect 463700 272478 463752 272484
rect 464710 272504 464766 272513
rect 464710 272439 464766 272448
rect 463516 270088 463568 270094
rect 463516 270030 463568 270036
rect 462714 264302 463188 264330
rect 463528 264316 463556 270030
rect 464724 264330 464752 272439
rect 465092 269822 465120 278038
rect 466564 275330 466592 278052
rect 466552 275324 466604 275330
rect 466552 275266 466604 275272
rect 467564 275324 467616 275330
rect 467564 275266 467616 275272
rect 466274 272912 466330 272921
rect 466274 272847 466330 272856
rect 466288 272626 466316 272847
rect 466414 272672 466466 272678
rect 466288 272620 466414 272626
rect 466288 272614 466466 272620
rect 466288 272598 466454 272614
rect 465080 269816 465132 269822
rect 465080 269758 465132 269764
rect 466000 269816 466052 269822
rect 466000 269758 466052 269764
rect 465172 267300 465224 267306
rect 465172 267242 465224 267248
rect 464370 264302 464752 264330
rect 465184 264316 465212 267242
rect 466012 264316 466040 269758
rect 466828 265124 466880 265130
rect 466828 265066 466880 265072
rect 466840 264316 466868 265066
rect 467576 264330 467604 275266
rect 467760 274378 467788 278052
rect 467944 278038 468970 278066
rect 467748 274372 467800 274378
rect 467748 274314 467800 274320
rect 467944 269958 467972 278038
rect 470152 275058 470180 278052
rect 470140 275052 470192 275058
rect 470140 274994 470192 275000
rect 471256 273562 471284 278052
rect 471612 276276 471664 276282
rect 471612 276218 471664 276224
rect 471244 273556 471296 273562
rect 471244 273498 471296 273504
rect 470554 272536 470606 272542
rect 470692 272536 470744 272542
rect 470554 272478 470606 272484
rect 470690 272504 470692 272513
rect 470744 272504 470746 272513
rect 470566 272354 470594 272478
rect 470690 272439 470746 272448
rect 470566 272326 470640 272354
rect 470612 272218 470640 272326
rect 470612 272190 470824 272218
rect 470796 272134 470824 272190
rect 470554 272128 470606 272134
rect 470784 272128 470836 272134
rect 470606 272076 470640 272082
rect 470554 272070 470640 272076
rect 470784 272070 470836 272076
rect 470566 272054 470640 272070
rect 470612 271969 470640 272054
rect 470598 271960 470654 271969
rect 470598 271895 470654 271904
rect 467932 269952 467984 269958
rect 467932 269894 467984 269900
rect 468484 269952 468536 269958
rect 468484 269894 468536 269900
rect 467576 264302 467682 264330
rect 468496 264316 468524 269894
rect 470968 269408 471020 269414
rect 470968 269350 471020 269356
rect 470140 267028 470192 267034
rect 470140 266970 470192 266976
rect 469312 265260 469364 265266
rect 469312 265202 469364 265208
rect 469324 264316 469352 265202
rect 470152 264316 470180 266970
rect 470980 264316 471008 269350
rect 471624 264330 471652 276218
rect 472452 273970 472480 278052
rect 473084 274916 473136 274922
rect 473084 274858 473136 274864
rect 472440 273964 472492 273970
rect 472440 273906 472492 273912
rect 473096 264330 473124 274858
rect 473648 273834 473676 278052
rect 474844 274242 474872 278052
rect 475028 278038 476054 278066
rect 474832 274236 474884 274242
rect 474832 274178 474884 274184
rect 474648 273964 474700 273970
rect 474648 273906 474700 273912
rect 473636 273828 473688 273834
rect 473636 273770 473688 273776
rect 474280 269272 474332 269278
rect 474280 269214 474332 269220
rect 473452 266416 473504 266422
rect 473452 266358 473504 266364
rect 471624 264302 471822 264330
rect 472650 264302 473124 264330
rect 473464 264316 473492 266358
rect 474292 264316 474320 269214
rect 474660 266422 474688 273906
rect 475028 269550 475056 278038
rect 477040 276412 477092 276418
rect 477040 276354 477092 276360
rect 476764 274780 476816 274786
rect 476764 274722 476816 274728
rect 476028 273556 476080 273562
rect 476028 273498 476080 273504
rect 475016 269544 475068 269550
rect 475016 269486 475068 269492
rect 476040 267734 476068 273498
rect 475948 267706 476068 267734
rect 474648 266416 474700 266422
rect 474648 266358 474700 266364
rect 475108 266416 475160 266422
rect 475108 266358 475160 266364
rect 475120 264316 475148 266358
rect 475948 264316 475976 267706
rect 476776 266762 476804 274722
rect 476764 266756 476816 266762
rect 476764 266698 476816 266704
rect 477052 264330 477080 276354
rect 477236 275194 477264 278052
rect 478064 278038 478354 278066
rect 479168 278038 479550 278066
rect 477224 275188 477276 275194
rect 477224 275130 477276 275136
rect 478064 271969 478092 278038
rect 478696 273420 478748 273426
rect 478696 273362 478748 273368
rect 478050 271960 478106 271969
rect 478050 271895 478106 271904
rect 477592 265396 477644 265402
rect 477592 265338 477644 265344
rect 476790 264302 477080 264330
rect 477604 264316 477632 265338
rect 478708 264330 478736 273362
rect 479168 271046 479196 278038
rect 479984 276548 480036 276554
rect 479984 276490 480036 276496
rect 479522 272096 479578 272105
rect 479522 272031 479578 272040
rect 479156 271040 479208 271046
rect 479156 270982 479208 270988
rect 479536 266422 479564 272031
rect 479524 266416 479576 266422
rect 479524 266358 479576 266364
rect 479248 265532 479300 265538
rect 479248 265474 479300 265480
rect 478446 264302 478736 264330
rect 479260 264316 479288 265474
rect 479996 264330 480024 276490
rect 480732 274650 480760 278052
rect 480720 274644 480772 274650
rect 480720 274586 480772 274592
rect 481364 273828 481416 273834
rect 481364 273770 481416 273776
rect 480536 272128 480588 272134
rect 480534 272096 480536 272105
rect 480588 272096 480590 272105
rect 480534 272031 480590 272040
rect 480168 271992 480220 271998
rect 480220 271940 480484 271946
rect 480168 271934 480484 271940
rect 480180 271918 480484 271934
rect 480456 271862 480484 271918
rect 480168 271856 480220 271862
rect 480444 271856 480496 271862
rect 480220 271804 480300 271810
rect 480168 271798 480300 271804
rect 480444 271798 480496 271804
rect 480180 271782 480300 271798
rect 480272 271046 480300 271782
rect 480260 271040 480312 271046
rect 480260 270982 480312 270988
rect 481376 264330 481404 273770
rect 481928 273698 481956 278052
rect 483138 278038 483612 278066
rect 482836 277364 482888 277370
rect 482836 277306 482888 277312
rect 481916 273692 481968 273698
rect 481916 273634 481968 273640
rect 482848 266422 482876 277306
rect 483584 271726 483612 278038
rect 484320 275874 484348 278052
rect 484872 278038 485530 278066
rect 484308 275868 484360 275874
rect 484308 275810 484360 275816
rect 484308 275052 484360 275058
rect 484308 274994 484360 275000
rect 484320 274514 484348 274994
rect 484308 274508 484360 274514
rect 484308 274450 484360 274456
rect 484216 273692 484268 273698
rect 484216 273634 484268 273640
rect 483572 271720 483624 271726
rect 483572 271662 483624 271668
rect 484228 266422 484256 273634
rect 484872 271862 484900 278038
rect 485044 275460 485096 275466
rect 485044 275402 485096 275408
rect 485228 275460 485280 275466
rect 485228 275402 485280 275408
rect 485056 275194 485084 275402
rect 485044 275188 485096 275194
rect 485044 275130 485096 275136
rect 485240 275058 485268 275402
rect 485228 275052 485280 275058
rect 485228 274994 485280 275000
rect 484860 271856 484912 271862
rect 484860 271798 484912 271804
rect 485044 271720 485096 271726
rect 485044 271662 485096 271668
rect 485056 266898 485084 271662
rect 486620 271046 486648 278052
rect 486792 274644 486844 274650
rect 486792 274586 486844 274592
rect 486608 271040 486660 271046
rect 486608 270982 486660 270988
rect 485044 266892 485096 266898
rect 485044 266834 485096 266840
rect 485044 266756 485096 266762
rect 485044 266698 485096 266704
rect 481732 266416 481784 266422
rect 481732 266358 481784 266364
rect 482836 266416 482888 266422
rect 482836 266358 482888 266364
rect 483388 266416 483440 266422
rect 483388 266358 483440 266364
rect 484216 266416 484268 266422
rect 484216 266358 484268 266364
rect 479996 264302 480102 264330
rect 480930 264302 481404 264330
rect 481744 264316 481772 266358
rect 482560 266076 482612 266082
rect 482560 266018 482612 266024
rect 482572 264316 482600 266018
rect 483400 264316 483428 266358
rect 484216 266212 484268 266218
rect 484216 266154 484268 266160
rect 484228 264316 484256 266154
rect 485056 264316 485084 266698
rect 486804 266422 486832 274586
rect 486976 270768 487028 270774
rect 486976 270710 487028 270716
rect 485872 266416 485924 266422
rect 485872 266358 485924 266364
rect 486792 266416 486844 266422
rect 486792 266358 486844 266364
rect 485884 264316 485912 266358
rect 486988 264330 487016 270710
rect 487816 270638 487844 278052
rect 488552 278038 489026 278066
rect 487988 277228 488040 277234
rect 487988 277170 488040 277176
rect 487804 270632 487856 270638
rect 487804 270574 487856 270580
rect 487160 266348 487212 266354
rect 487160 266290 487212 266296
rect 487172 266082 487200 266290
rect 487160 266076 487212 266082
rect 487160 266018 487212 266024
rect 488000 264330 488028 277170
rect 488356 274508 488408 274514
rect 488356 274450 488408 274456
rect 486726 264302 487016 264330
rect 487554 264302 488028 264330
rect 488368 264316 488396 274450
rect 488552 269074 488580 278038
rect 490208 270910 490236 278052
rect 490564 275868 490616 275874
rect 490564 275810 490616 275816
rect 490196 270904 490248 270910
rect 490196 270846 490248 270852
rect 489644 270632 489696 270638
rect 489644 270574 489696 270580
rect 488540 269068 488592 269074
rect 488540 269010 488592 269016
rect 489656 264330 489684 270574
rect 490576 267714 490604 275810
rect 491404 275194 491432 278052
rect 491680 278038 492614 278066
rect 491392 275188 491444 275194
rect 491392 275130 491444 275136
rect 491680 268938 491708 278038
rect 493704 271590 493732 278052
rect 494072 278038 494914 278066
rect 495452 278038 496110 278066
rect 493692 271584 493744 271590
rect 493692 271526 493744 271532
rect 492588 270904 492640 270910
rect 492588 270846 492640 270852
rect 491668 268932 491720 268938
rect 491668 268874 491720 268880
rect 490840 267980 490892 267986
rect 490840 267922 490892 267928
rect 490564 267708 490616 267714
rect 490564 267650 490616 267656
rect 490012 266756 490064 266762
rect 490012 266698 490064 266704
rect 489210 264302 489684 264330
rect 490024 264316 490052 266698
rect 490852 264316 490880 267922
rect 492600 266490 492628 270846
rect 493324 269068 493376 269074
rect 493324 269010 493376 269016
rect 491668 266484 491720 266490
rect 491668 266426 491720 266432
rect 492588 266484 492640 266490
rect 492588 266426 492640 266432
rect 491680 264316 491708 266426
rect 492496 266076 492548 266082
rect 492496 266018 492548 266024
rect 492508 264316 492536 266018
rect 493336 264316 493364 269010
rect 494072 268258 494100 278038
rect 495072 271040 495124 271046
rect 495072 270982 495124 270988
rect 494060 268252 494112 268258
rect 494060 268194 494112 268200
rect 495084 266490 495112 270982
rect 495256 269544 495308 269550
rect 495256 269486 495308 269492
rect 494152 266484 494204 266490
rect 494152 266426 494204 266432
rect 495072 266484 495124 266490
rect 495072 266426 495124 266432
rect 494164 264316 494192 266426
rect 495268 264330 495296 269486
rect 495452 268802 495480 278038
rect 496544 271720 496596 271726
rect 496544 271662 496596 271668
rect 495440 268796 495492 268802
rect 495440 268738 495492 268744
rect 495808 268252 495860 268258
rect 495808 268194 495860 268200
rect 495006 264302 495296 264330
rect 495820 264316 495848 268194
rect 496556 264330 496584 271662
rect 497292 271454 497320 278052
rect 497924 277092 497976 277098
rect 497924 277034 497976 277040
rect 497280 271448 497332 271454
rect 497280 271390 497332 271396
rect 497936 264330 497964 277034
rect 498488 275602 498516 278052
rect 499684 277394 499712 278052
rect 499592 277366 499712 277394
rect 498476 275596 498528 275602
rect 498476 275538 498528 275544
rect 498844 275596 498896 275602
rect 498844 275538 498896 275544
rect 498292 268932 498344 268938
rect 498292 268874 498344 268880
rect 496556 264302 496662 264330
rect 497490 264302 497964 264330
rect 498304 264316 498332 268874
rect 498856 267442 498884 275538
rect 499304 271584 499356 271590
rect 499304 271526 499356 271532
rect 498844 267436 498896 267442
rect 498844 267378 498896 267384
rect 499316 264330 499344 271526
rect 499592 268666 499620 277366
rect 500880 271318 500908 278052
rect 501432 278038 501998 278066
rect 501432 271862 501460 278038
rect 503180 273222 503208 278052
rect 504008 278038 504390 278066
rect 503444 275052 503496 275058
rect 503444 274994 503496 275000
rect 503168 273216 503220 273222
rect 503168 273158 503220 273164
rect 501602 271960 501658 271969
rect 501602 271895 501658 271904
rect 501420 271856 501472 271862
rect 501420 271798 501472 271804
rect 500868 271312 500920 271318
rect 500868 271254 500920 271260
rect 500776 268796 500828 268802
rect 500776 268738 500828 268744
rect 499580 268660 499632 268666
rect 499580 268602 499632 268608
rect 499948 266892 500000 266898
rect 499948 266834 500000 266840
rect 499146 264302 499344 264330
rect 499960 264316 499988 266834
rect 500788 264316 500816 268738
rect 501616 266626 501644 271895
rect 501972 271448 502024 271454
rect 501972 271390 502024 271396
rect 501604 266620 501656 266626
rect 501604 266562 501656 266568
rect 501984 264330 502012 271390
rect 503260 268660 503312 268666
rect 503260 268602 503312 268608
rect 502432 266484 502484 266490
rect 502432 266426 502484 266432
rect 501630 264302 502012 264330
rect 502444 264316 502472 266426
rect 503272 264316 503300 268602
rect 503456 266490 503484 274994
rect 504008 271182 504036 278038
rect 505572 275874 505600 278052
rect 506492 278038 506782 278066
rect 505560 275868 505612 275874
rect 505560 275810 505612 275816
rect 506204 274372 506256 274378
rect 506204 274314 506256 274320
rect 504180 273216 504232 273222
rect 504180 273158 504232 273164
rect 504192 272406 504220 273158
rect 504180 272400 504232 272406
rect 504180 272342 504232 272348
rect 504364 272400 504416 272406
rect 504364 272342 504416 272348
rect 504376 271998 504404 272342
rect 504364 271992 504416 271998
rect 504548 271992 504600 271998
rect 504364 271934 504416 271940
rect 504546 271960 504548 271969
rect 504600 271960 504602 271969
rect 504546 271895 504602 271904
rect 504548 271720 504600 271726
rect 504548 271662 504600 271668
rect 504560 271454 504588 271662
rect 504548 271448 504600 271454
rect 504548 271390 504600 271396
rect 505008 271448 505060 271454
rect 505008 271390 505060 271396
rect 503996 271176 504048 271182
rect 503996 271118 504048 271124
rect 504824 266620 504876 266626
rect 504824 266562 504876 266568
rect 503444 266484 503496 266490
rect 503444 266426 503496 266432
rect 504088 266484 504140 266490
rect 504088 266426 504140 266432
rect 504100 264316 504128 266426
rect 504836 264330 504864 266562
rect 505020 266490 505048 271390
rect 505008 266484 505060 266490
rect 505008 266426 505060 266432
rect 506216 264330 506244 274314
rect 506492 268530 506520 278038
rect 507492 275188 507544 275194
rect 507492 275130 507544 275136
rect 506480 268524 506532 268530
rect 506480 268466 506532 268472
rect 507504 267734 507532 275130
rect 507964 273086 507992 278052
rect 509068 276010 509096 278052
rect 509056 276004 509108 276010
rect 509056 275946 509108 275952
rect 507952 273080 508004 273086
rect 507952 273022 508004 273028
rect 509700 273080 509752 273086
rect 509700 273022 509752 273028
rect 507676 271312 507728 271318
rect 507676 271254 507728 271260
rect 507412 267706 507532 267734
rect 506572 266484 506624 266490
rect 506572 266426 506624 266432
rect 504836 264302 504942 264330
rect 505770 264302 506244 264330
rect 506584 264316 506612 266426
rect 507412 264316 507440 267706
rect 507688 266490 507716 271254
rect 509238 269920 509294 269929
rect 509238 269855 509294 269864
rect 509252 269686 509280 269855
rect 509240 269680 509292 269686
rect 509240 269622 509292 269628
rect 509146 269512 509202 269521
rect 509146 269447 509202 269456
rect 508228 268524 508280 268530
rect 508228 268466 508280 268472
rect 507860 266892 507912 266898
rect 507860 266834 507912 266840
rect 507872 266490 507900 266834
rect 507676 266484 507728 266490
rect 507676 266426 507728 266432
rect 507860 266484 507912 266490
rect 507860 266426 507912 266432
rect 508240 264316 508268 268466
rect 509160 267734 509188 269447
rect 509068 267706 509188 267734
rect 509068 264316 509096 267706
rect 509712 266762 509740 273022
rect 510264 272270 510292 278052
rect 511460 273222 511488 278052
rect 511632 276956 511684 276962
rect 511632 276898 511684 276904
rect 511448 273216 511500 273222
rect 511448 273158 511500 273164
rect 510252 272264 510304 272270
rect 510252 272206 510304 272212
rect 509884 269544 509936 269550
rect 509882 269512 509884 269521
rect 509936 269512 509938 269521
rect 509882 269447 509938 269456
rect 511644 267734 511672 276898
rect 512656 275602 512684 278052
rect 513196 276004 513248 276010
rect 513196 275946 513248 275952
rect 512644 275596 512696 275602
rect 512644 275538 512696 275544
rect 511816 274236 511868 274242
rect 511816 274178 511868 274184
rect 509884 267708 509936 267714
rect 509884 267650 509936 267656
rect 511552 267706 511672 267734
rect 509700 266756 509752 266762
rect 509700 266698 509752 266704
rect 509896 264316 509924 267650
rect 510712 266756 510764 266762
rect 510712 266698 510764 266704
rect 510724 264316 510752 266698
rect 511552 264316 511580 267706
rect 511828 266762 511856 274178
rect 513208 266762 513236 275946
rect 513852 274106 513880 278052
rect 514484 276820 514536 276826
rect 514484 276762 514536 276768
rect 513840 274100 513892 274106
rect 513840 274042 513892 274048
rect 513840 273080 513892 273086
rect 513840 273022 513892 273028
rect 513852 272814 513880 273022
rect 513840 272808 513892 272814
rect 513840 272750 513892 272756
rect 514024 272808 514076 272814
rect 514024 272750 514076 272756
rect 514036 272406 514064 272750
rect 514024 272400 514076 272406
rect 514024 272342 514076 272348
rect 511816 266756 511868 266762
rect 511816 266698 511868 266704
rect 512368 266756 512420 266762
rect 512368 266698 512420 266704
rect 513196 266756 513248 266762
rect 513196 266698 513248 266704
rect 512380 264316 512408 266698
rect 513196 265940 513248 265946
rect 513196 265882 513248 265888
rect 513208 264316 513236 265882
rect 514496 264330 514524 276762
rect 515048 272950 515076 278052
rect 516244 275738 516272 278052
rect 516612 278038 517362 278066
rect 516232 275732 516284 275738
rect 516232 275674 516284 275680
rect 515220 273216 515272 273222
rect 515220 273158 515272 273164
rect 515404 273216 515456 273222
rect 515404 273158 515456 273164
rect 515232 272950 515260 273158
rect 515036 272944 515088 272950
rect 515036 272886 515088 272892
rect 515220 272944 515272 272950
rect 515220 272886 515272 272892
rect 514852 267436 514904 267442
rect 514852 267378 514904 267384
rect 514050 264302 514524 264330
rect 514864 264316 514892 267378
rect 515416 267170 515444 273158
rect 516612 269929 516640 278038
rect 516784 275596 516836 275602
rect 516784 275538 516836 275544
rect 516598 269920 516654 269929
rect 516598 269855 516654 269864
rect 516796 267578 516824 275538
rect 518544 273086 518572 278052
rect 518716 276684 518768 276690
rect 518716 276626 518768 276632
rect 518532 273080 518584 273086
rect 518532 273022 518584 273028
rect 517428 272400 517480 272406
rect 517428 272342 517480 272348
rect 516784 267572 516836 267578
rect 516784 267514 516836 267520
rect 515404 267164 515456 267170
rect 515404 267106 515456 267112
rect 517244 267164 517296 267170
rect 517244 267106 517296 267112
rect 516508 266756 516560 266762
rect 516508 266698 516560 266704
rect 515680 265804 515732 265810
rect 515680 265746 515732 265752
rect 515692 264316 515720 265746
rect 516520 264316 516548 266698
rect 517256 264330 517284 267106
rect 517440 266762 517468 272342
rect 518728 267734 518756 276626
rect 519740 273222 519768 278052
rect 520292 278038 520950 278066
rect 519728 273216 519780 273222
rect 519728 273158 519780 273164
rect 520096 272264 520148 272270
rect 520096 272206 520148 272212
rect 518544 267706 518756 267734
rect 517428 266756 517480 266762
rect 517428 266698 517480 266704
rect 518544 264330 518572 267706
rect 519820 267572 519872 267578
rect 519820 267514 519872 267520
rect 518992 266756 519044 266762
rect 518992 266698 519044 266704
rect 517256 264302 517362 264330
rect 518190 264302 518572 264330
rect 519004 264316 519032 266698
rect 519832 264316 519860 267514
rect 520108 266762 520136 272206
rect 520292 270502 520320 278038
rect 521476 273216 521528 273222
rect 521476 273158 521528 273164
rect 520280 270496 520332 270502
rect 520280 270438 520332 270444
rect 520096 266756 520148 266762
rect 520096 266698 520148 266704
rect 520648 265668 520700 265674
rect 520648 265610 520700 265616
rect 520660 264316 520688 265610
rect 521488 264316 521516 273158
rect 522132 272678 522160 278052
rect 522764 275868 522816 275874
rect 522764 275810 522816 275816
rect 522120 272672 522172 272678
rect 522120 272614 522172 272620
rect 522776 264330 522804 275810
rect 523328 274786 523356 278052
rect 524432 278038 524538 278066
rect 523316 274780 523368 274786
rect 523316 274722 523368 274728
rect 523684 274780 523736 274786
rect 523684 274722 523736 274728
rect 523132 270496 523184 270502
rect 523132 270438 523184 270444
rect 522330 264302 522804 264330
rect 523144 264316 523172 270438
rect 523696 267306 523724 274722
rect 524052 271176 524104 271182
rect 524052 271118 524104 271124
rect 524064 267734 524092 271118
rect 524432 270230 524460 278038
rect 525628 272814 525656 278052
rect 526824 275602 526852 278052
rect 527192 278038 528034 278066
rect 528572 278038 529230 278066
rect 526812 275596 526864 275602
rect 526812 275538 526864 275544
rect 525616 272808 525668 272814
rect 525616 272750 525668 272756
rect 526812 272672 526864 272678
rect 526812 272614 526864 272620
rect 525616 270360 525668 270366
rect 525616 270302 525668 270308
rect 524420 270224 524472 270230
rect 524420 270166 524472 270172
rect 523972 267706 524092 267734
rect 523684 267300 523736 267306
rect 523684 267242 523736 267248
rect 523972 264316 524000 267706
rect 524788 267300 524840 267306
rect 524788 267242 524840 267248
rect 524800 264316 524828 267242
rect 525628 264316 525656 270302
rect 526824 264330 526852 272614
rect 527192 270230 527220 278038
rect 528192 275732 528244 275738
rect 528192 275674 528244 275680
rect 527180 270224 527232 270230
rect 527180 270166 527232 270172
rect 527180 268116 527232 268122
rect 527180 268058 527232 268064
rect 527192 267170 527220 268058
rect 527180 267164 527232 267170
rect 527180 267106 527232 267112
rect 528204 266762 528232 275674
rect 528376 270224 528428 270230
rect 528376 270166 528428 270172
rect 527272 266756 527324 266762
rect 527272 266698 527324 266704
rect 528192 266756 528244 266762
rect 528192 266698 528244 266704
rect 526470 264302 526852 264330
rect 527284 264316 527312 266698
rect 528388 264330 528416 270166
rect 528572 268394 528600 278038
rect 530412 275466 530440 278052
rect 531332 278038 531622 278066
rect 530400 275460 530452 275466
rect 530400 275402 530452 275408
rect 529848 272808 529900 272814
rect 529848 272750 529900 272756
rect 528560 268388 528612 268394
rect 528560 268330 528612 268336
rect 529664 267164 529716 267170
rect 529664 267106 529716 267112
rect 528928 266756 528980 266762
rect 528928 266698 528980 266704
rect 528126 264302 528416 264330
rect 528940 264316 528968 266698
rect 529676 264330 529704 267106
rect 529860 266762 529888 272750
rect 530398 270192 530454 270201
rect 531332 270178 531360 278038
rect 532332 275596 532384 275602
rect 532332 275538 532384 275544
rect 530398 270127 530454 270136
rect 530780 270150 531360 270178
rect 530412 269822 530440 270127
rect 530780 270094 530808 270150
rect 530768 270088 530820 270094
rect 530768 270030 530820 270036
rect 530952 270088 531004 270094
rect 530952 270030 531004 270036
rect 530400 269816 530452 269822
rect 530400 269758 530452 269764
rect 529848 266756 529900 266762
rect 529848 266698 529900 266704
rect 530964 264330 530992 270030
rect 532344 267734 532372 275538
rect 532516 272944 532568 272950
rect 532516 272886 532568 272892
rect 532252 267706 532372 267734
rect 531412 266756 531464 266762
rect 531412 266698 531464 266704
rect 529676 264302 529782 264330
rect 530610 264302 530992 264330
rect 531424 264316 531452 266698
rect 532252 264316 532280 267706
rect 532528 266762 532556 272886
rect 532712 272542 532740 278052
rect 533908 274786 533936 278052
rect 534092 278038 535118 278066
rect 535748 278038 536314 278066
rect 533896 274780 533948 274786
rect 533896 274722 533948 274728
rect 532884 272808 532936 272814
rect 532884 272750 532936 272756
rect 533712 272808 533764 272814
rect 533712 272750 533764 272756
rect 532896 272542 532924 272750
rect 532700 272536 532752 272542
rect 532700 272478 532752 272484
rect 532884 272536 532936 272542
rect 532884 272478 532936 272484
rect 532884 270496 532936 270502
rect 532884 270438 532936 270444
rect 532896 269686 532924 270438
rect 533528 270360 533580 270366
rect 533172 270308 533528 270314
rect 533172 270302 533580 270308
rect 533172 270286 533568 270302
rect 533172 270094 533200 270286
rect 533160 270088 533212 270094
rect 533160 270030 533212 270036
rect 532884 269680 532936 269686
rect 532884 269622 532936 269628
rect 532516 266756 532568 266762
rect 532516 266698 532568 266704
rect 533068 266756 533120 266762
rect 533068 266698 533120 266704
rect 533080 264316 533108 266698
rect 533724 264330 533752 272750
rect 534092 270201 534120 278038
rect 534724 274780 534776 274786
rect 534724 274722 534776 274728
rect 534078 270192 534134 270201
rect 534078 270127 534134 270136
rect 533988 269952 534040 269958
rect 533988 269894 534040 269900
rect 534000 266762 534028 269894
rect 534736 267034 534764 274722
rect 534724 267028 534776 267034
rect 534724 266970 534776 266976
rect 535552 267028 535604 267034
rect 535552 266970 535604 266976
rect 534724 266892 534776 266898
rect 534724 266834 534776 266840
rect 533988 266756 534040 266762
rect 533988 266698 534040 266704
rect 533724 264302 533922 264330
rect 534736 264316 534764 266834
rect 535564 264316 535592 266970
rect 535748 265130 535776 278038
rect 537496 275330 537524 278052
rect 538508 278038 538706 278066
rect 537668 275460 537720 275466
rect 537668 275402 537720 275408
rect 537484 275324 537536 275330
rect 537484 275266 537536 275272
rect 536748 274100 536800 274106
rect 536748 274042 536800 274048
rect 536562 272504 536618 272513
rect 536562 272439 536618 272448
rect 535736 265124 535788 265130
rect 535736 265066 535788 265072
rect 536576 264330 536604 272439
rect 536760 267034 536788 274042
rect 536748 267028 536800 267034
rect 536748 266970 536800 266976
rect 537680 264330 537708 275402
rect 538508 273254 538536 278038
rect 539888 277394 539916 278052
rect 539888 277366 540008 277394
rect 539322 274000 539378 274009
rect 539322 273935 539378 273944
rect 538324 273226 538536 273254
rect 538324 270094 538352 273226
rect 539048 272944 539100 272950
rect 538508 272892 539048 272898
rect 538508 272886 539100 272892
rect 538508 272870 539088 272886
rect 538508 272542 538536 272870
rect 538680 272808 538732 272814
rect 538680 272750 538732 272756
rect 538692 272542 538720 272750
rect 538496 272536 538548 272542
rect 538496 272478 538548 272484
rect 538680 272536 538732 272542
rect 538680 272478 538732 272484
rect 538312 270088 538364 270094
rect 538312 270030 538364 270036
rect 538324 269878 538720 269906
rect 538034 269784 538090 269793
rect 538034 269719 538090 269728
rect 536406 264302 536604 264330
rect 537234 264302 537708 264330
rect 538048 264316 538076 269719
rect 538324 269414 538352 269878
rect 538692 269822 538720 269878
rect 538496 269816 538548 269822
rect 538496 269758 538548 269764
rect 538680 269816 538732 269822
rect 538680 269758 538732 269764
rect 538508 269414 538536 269758
rect 538312 269408 538364 269414
rect 538312 269350 538364 269356
rect 538496 269408 538548 269414
rect 538496 269350 538548 269356
rect 539336 264330 539364 273935
rect 539692 267028 539744 267034
rect 539692 266970 539744 266976
rect 538890 264302 539364 264330
rect 539704 264316 539732 266970
rect 539980 265266 540008 277366
rect 540992 274786 541020 278052
rect 541176 278038 542202 278066
rect 540980 274780 541032 274786
rect 540980 274722 541032 274728
rect 540520 269952 540572 269958
rect 540520 269894 540572 269900
rect 539968 265260 540020 265266
rect 539968 265202 540020 265208
rect 540532 264316 540560 269894
rect 541176 269822 541204 278038
rect 543384 276282 543412 278052
rect 543372 276276 543424 276282
rect 543372 276218 543424 276224
rect 542268 275324 542320 275330
rect 542268 275266 542320 275272
rect 542280 273254 542308 275266
rect 544580 274922 544608 278052
rect 544568 274916 544620 274922
rect 544568 274858 544620 274864
rect 545776 273970 545804 278052
rect 546512 278038 546986 278066
rect 547892 278038 548090 278066
rect 545946 274000 546002 274009
rect 545764 273964 545816 273970
rect 545946 273935 545948 273944
rect 545764 273906 545816 273912
rect 546000 273935 546002 273944
rect 545948 273906 546000 273912
rect 542188 273226 542308 273254
rect 541164 269816 541216 269822
rect 541348 269816 541400 269822
rect 541164 269758 541216 269764
rect 541346 269784 541348 269793
rect 541400 269784 541402 269793
rect 541346 269719 541402 269728
rect 541348 268388 541400 268394
rect 541348 268330 541400 268336
rect 541360 264316 541388 268330
rect 542188 264316 542216 273226
rect 546512 269210 546540 278038
rect 547694 272504 547750 272513
rect 547694 272439 547750 272448
rect 547708 272134 547736 272439
rect 547512 272128 547564 272134
rect 547510 272096 547512 272105
rect 547696 272128 547748 272134
rect 547564 272096 547566 272105
rect 547892 272105 547920 278038
rect 549272 273562 549300 278052
rect 550468 276418 550496 278052
rect 550652 278038 551678 278066
rect 550456 276412 550508 276418
rect 550456 276354 550508 276360
rect 549260 273556 549312 273562
rect 549260 273498 549312 273504
rect 549904 273556 549956 273562
rect 549904 273498 549956 273504
rect 547696 272070 547748 272076
rect 547878 272096 547934 272105
rect 547510 272031 547566 272040
rect 547878 272031 547934 272040
rect 546500 269204 546552 269210
rect 546500 269146 546552 269152
rect 543004 266756 543056 266762
rect 543004 266698 543056 266704
rect 543016 264316 543044 266698
rect 549916 266490 549944 273498
rect 549904 266484 549956 266490
rect 549904 266426 549956 266432
rect 550652 265402 550680 278038
rect 552860 273426 552888 278052
rect 553412 278038 554070 278066
rect 552848 273420 552900 273426
rect 552848 273362 552900 273368
rect 553412 265538 553440 278038
rect 555252 276554 555280 278052
rect 555240 276548 555292 276554
rect 555240 276490 555292 276496
rect 556356 273834 556384 278052
rect 557552 277370 557580 278052
rect 557736 278038 558762 278066
rect 557540 277364 557592 277370
rect 557540 277306 557592 277312
rect 556344 273828 556396 273834
rect 556344 273770 556396 273776
rect 556804 273828 556856 273834
rect 556804 273770 556856 273776
rect 556816 266626 556844 273770
rect 556804 266620 556856 266626
rect 556804 266562 556856 266568
rect 557736 266354 557764 278038
rect 559944 273698 559972 278052
rect 560312 278038 561154 278066
rect 559932 273692 559984 273698
rect 559932 273634 559984 273640
rect 557724 266348 557776 266354
rect 557724 266290 557776 266296
rect 560312 266218 560340 278038
rect 562336 271998 562364 278052
rect 563440 274650 563468 278052
rect 563428 274644 563480 274650
rect 563428 274586 563480 274592
rect 562324 271992 562376 271998
rect 562324 271934 562376 271940
rect 564636 270774 564664 278052
rect 565832 277234 565860 278052
rect 565820 277228 565872 277234
rect 565820 277170 565872 277176
rect 567028 274514 567056 278052
rect 567016 274508 567068 274514
rect 567016 274450 567068 274456
rect 564624 270768 564676 270774
rect 564624 270710 564676 270716
rect 567844 270768 567896 270774
rect 567844 270710 567896 270716
rect 567856 267714 567884 270710
rect 568224 270638 568252 278052
rect 569420 273086 569448 278052
rect 569972 278038 570630 278066
rect 569408 273080 569460 273086
rect 569408 273022 569460 273028
rect 568212 270632 568264 270638
rect 568212 270574 568264 270580
rect 569972 267986 570000 278038
rect 571720 270910 571748 278052
rect 572732 278038 572930 278066
rect 571708 270904 571760 270910
rect 571708 270846 571760 270852
rect 569960 267980 570012 267986
rect 569960 267922 570012 267928
rect 567844 267708 567896 267714
rect 567844 267650 567896 267656
rect 560300 266212 560352 266218
rect 560300 266154 560352 266160
rect 572732 266082 572760 278038
rect 574112 269074 574140 278052
rect 575308 271046 575336 278052
rect 575492 278038 576518 278066
rect 576872 278038 577714 278066
rect 578528 278038 578910 278066
rect 575296 271040 575348 271046
rect 575296 270982 575348 270988
rect 575492 269414 575520 278038
rect 575480 269408 575532 269414
rect 575480 269350 575532 269356
rect 574100 269068 574152 269074
rect 574100 269010 574152 269016
rect 576872 268258 576900 278038
rect 578528 271862 578556 278038
rect 580000 277098 580028 278052
rect 581012 278038 581210 278066
rect 579988 277092 580040 277098
rect 579988 277034 580040 277040
rect 578516 271856 578568 271862
rect 578516 271798 578568 271804
rect 578884 271856 578936 271862
rect 578884 271798 578936 271804
rect 576860 268252 576912 268258
rect 576860 268194 576912 268200
rect 578896 267442 578924 271798
rect 581012 268938 581040 278038
rect 582392 271590 582420 278052
rect 583588 273562 583616 278052
rect 583772 278038 584798 278066
rect 583576 273556 583628 273562
rect 583576 273498 583628 273504
rect 582380 271584 582432 271590
rect 582380 271526 582432 271532
rect 583024 271584 583076 271590
rect 583024 271526 583076 271532
rect 581000 268932 581052 268938
rect 581000 268874 581052 268880
rect 583036 267578 583064 271526
rect 583772 268802 583800 278038
rect 585980 271726 586008 278052
rect 587084 275058 587112 278052
rect 587912 278038 588294 278066
rect 587072 275052 587124 275058
rect 587072 274994 587124 275000
rect 585968 271720 586020 271726
rect 585968 271662 586020 271668
rect 583760 268796 583812 268802
rect 583760 268738 583812 268744
rect 587912 268666 587940 278038
rect 589476 271454 589504 278052
rect 590672 273834 590700 278052
rect 591868 274378 591896 278052
rect 591856 274372 591908 274378
rect 591856 274314 591908 274320
rect 590660 273828 590712 273834
rect 590660 273770 590712 273776
rect 589464 271448 589516 271454
rect 589464 271390 589516 271396
rect 589924 271448 589976 271454
rect 589924 271390 589976 271396
rect 587900 268660 587952 268666
rect 587900 268602 587952 268608
rect 583024 267572 583076 267578
rect 583024 267514 583076 267520
rect 578884 267436 578936 267442
rect 578884 267378 578936 267384
rect 589936 266898 589964 271390
rect 593064 271318 593092 278052
rect 594260 275194 594288 278052
rect 594812 278038 595378 278066
rect 596192 278038 596574 278066
rect 594248 275188 594300 275194
rect 594248 275130 594300 275136
rect 593052 271312 593104 271318
rect 593052 271254 593104 271260
rect 594812 268530 594840 278038
rect 596192 269550 596220 278038
rect 597756 270774 597784 278052
rect 598952 274242 598980 278052
rect 600148 276962 600176 278052
rect 600136 276956 600188 276962
rect 600136 276898 600188 276904
rect 601344 276010 601372 278052
rect 601712 278038 602462 278066
rect 601332 276004 601384 276010
rect 601332 275946 601384 275952
rect 598940 274236 598992 274242
rect 598940 274178 598992 274184
rect 600964 272400 601016 272406
rect 600964 272342 601016 272348
rect 601148 272400 601200 272406
rect 601148 272342 601200 272348
rect 600976 272134 601004 272342
rect 600964 272128 601016 272134
rect 600964 272070 601016 272076
rect 601160 271998 601188 272342
rect 601148 271992 601200 271998
rect 601148 271934 601200 271940
rect 598204 271312 598256 271318
rect 598204 271254 598256 271260
rect 597744 270768 597796 270774
rect 597744 270710 597796 270716
rect 596180 269544 596232 269550
rect 596180 269486 596232 269492
rect 594800 268524 594852 268530
rect 594800 268466 594852 268472
rect 589924 266892 589976 266898
rect 589924 266834 589976 266840
rect 598216 266762 598244 271254
rect 598204 266756 598256 266762
rect 598204 266698 598256 266704
rect 572720 266076 572772 266082
rect 572720 266018 572772 266024
rect 601712 265946 601740 278038
rect 603644 276826 603672 278052
rect 603632 276820 603684 276826
rect 603632 276762 603684 276768
rect 604840 271862 604868 278052
rect 605852 278038 606050 278066
rect 604828 271856 604880 271862
rect 604828 271798 604880 271804
rect 601700 265940 601752 265946
rect 601700 265882 601752 265888
rect 605852 265810 605880 278038
rect 607232 272134 607260 278052
rect 607416 278038 608442 278066
rect 607220 272128 607272 272134
rect 607220 272070 607272 272076
rect 607416 268122 607444 278038
rect 609624 276690 609652 278052
rect 609612 276684 609664 276690
rect 609612 276626 609664 276632
rect 610728 272270 610756 278052
rect 611648 278038 611938 278066
rect 612752 278038 613134 278066
rect 610716 272264 610768 272270
rect 610716 272206 610768 272212
rect 611648 271590 611676 278038
rect 611636 271584 611688 271590
rect 611636 271526 611688 271532
rect 612004 271584 612056 271590
rect 612004 271526 612056 271532
rect 607404 268116 607456 268122
rect 607404 268058 607456 268064
rect 612016 267306 612044 271526
rect 612004 267300 612056 267306
rect 612004 267242 612056 267248
rect 605840 265804 605892 265810
rect 605840 265746 605892 265752
rect 612752 265674 612780 278038
rect 614316 273222 614344 278052
rect 615512 275874 615540 278052
rect 616432 278038 616722 278066
rect 617352 278038 617826 278066
rect 615500 275868 615552 275874
rect 615500 275810 615552 275816
rect 614304 273216 614356 273222
rect 614304 273158 614356 273164
rect 616432 269686 616460 278038
rect 617352 271182 617380 278038
rect 619008 271590 619036 278052
rect 619652 278038 620218 278066
rect 618996 271584 619048 271590
rect 618996 271526 619048 271532
rect 617340 271176 617392 271182
rect 617340 271118 617392 271124
rect 617524 271176 617576 271182
rect 617524 271118 617576 271124
rect 616420 269680 616472 269686
rect 616420 269622 616472 269628
rect 617536 267170 617564 271118
rect 619652 270502 619680 278038
rect 621400 272678 621428 278052
rect 622596 275738 622624 278052
rect 623806 278038 624004 278066
rect 622584 275732 622636 275738
rect 622584 275674 622636 275680
rect 621388 272672 621440 272678
rect 621388 272614 621440 272620
rect 619640 270496 619692 270502
rect 619640 270438 619692 270444
rect 623976 270230 624004 278038
rect 624988 272950 625016 278052
rect 624976 272944 625028 272950
rect 624976 272886 625028 272892
rect 626092 271182 626120 278052
rect 626552 278038 627302 278066
rect 626080 271176 626132 271182
rect 626080 271118 626132 271124
rect 626552 270366 626580 278038
rect 628484 272814 628512 278052
rect 629484 277908 629536 277914
rect 629484 277850 629536 277856
rect 629496 277506 629524 277850
rect 629484 277500 629536 277506
rect 629484 277442 629536 277448
rect 629680 275602 629708 278052
rect 630692 278038 630890 278066
rect 629668 275596 629720 275602
rect 629668 275538 629720 275544
rect 628472 272808 628524 272814
rect 628472 272750 628524 272756
rect 626540 270360 626592 270366
rect 626540 270302 626592 270308
rect 623964 270224 624016 270230
rect 623964 270166 624016 270172
rect 630692 270094 630720 278038
rect 632072 272950 632100 278052
rect 632060 272944 632112 272950
rect 632060 272886 632112 272892
rect 633268 271454 633296 278052
rect 634372 274106 634400 278052
rect 634360 274100 634412 274106
rect 634360 274042 634412 274048
rect 634084 272672 634136 272678
rect 634084 272614 634136 272620
rect 633256 271448 633308 271454
rect 633256 271390 633308 271396
rect 630680 270088 630732 270094
rect 630680 270030 630732 270036
rect 617524 267164 617576 267170
rect 617524 267106 617576 267112
rect 634096 267034 634124 272614
rect 634084 267028 634136 267034
rect 634084 266970 634136 266976
rect 612740 265668 612792 265674
rect 612740 265610 612792 265616
rect 553400 265532 553452 265538
rect 553400 265474 553452 265480
rect 550640 265396 550692 265402
rect 550640 265338 550692 265344
rect 554410 262168 554466 262177
rect 554410 262103 554466 262112
rect 554424 260914 554452 262103
rect 570604 261520 570656 261526
rect 570604 261462 570656 261468
rect 554412 260908 554464 260914
rect 554412 260850 554464 260856
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 554318 259992 554374 260001
rect 554318 259927 554374 259936
rect 554332 259486 554360 259927
rect 554320 259480 554372 259486
rect 554320 259422 554372 259428
rect 563704 259480 563756 259486
rect 563704 259422 563756 259428
rect 553950 257816 554006 257825
rect 553950 257751 554006 257760
rect 553964 256766 553992 257751
rect 553952 256760 554004 256766
rect 553952 256702 554004 256708
rect 560944 256760 560996 256766
rect 560944 256702 560996 256708
rect 554502 255640 554558 255649
rect 554502 255575 554504 255584
rect 554556 255575 554558 255584
rect 558184 255604 558236 255610
rect 554504 255546 554556 255552
rect 558184 255546 558236 255552
rect 554410 253464 554466 253473
rect 554410 253399 554466 253408
rect 554424 252618 554452 253399
rect 554412 252612 554464 252618
rect 554412 252554 554464 252560
rect 554134 251288 554190 251297
rect 554134 251223 554136 251232
rect 554188 251223 554190 251232
rect 556804 251252 556856 251258
rect 554136 251194 554188 251200
rect 556804 251194 556856 251200
rect 554042 249112 554098 249121
rect 554042 249047 554098 249056
rect 553858 246936 553914 246945
rect 553858 246871 553914 246880
rect 553872 245682 553900 246871
rect 553860 245676 553912 245682
rect 553860 245618 553912 245624
rect 553490 244760 553546 244769
rect 553490 244695 553546 244704
rect 553504 244322 553532 244695
rect 553492 244316 553544 244322
rect 553492 244258 553544 244264
rect 553674 242584 553730 242593
rect 553674 242519 553730 242528
rect 553688 241534 553716 242519
rect 553676 241528 553728 241534
rect 553676 241470 553728 241476
rect 553768 236836 553820 236842
rect 553768 236778 553820 236784
rect 553780 236065 553808 236778
rect 553766 236056 553822 236065
rect 553766 235991 553822 236000
rect 134984 231464 135036 231470
rect 134984 231406 135036 231412
rect 137652 231464 137704 231470
rect 137652 231406 137704 231412
rect 92388 231192 92440 231198
rect 92388 231134 92440 231140
rect 82084 230036 82136 230042
rect 82084 229978 82136 229984
rect 86224 230036 86276 230042
rect 86224 229978 86276 229984
rect 68284 229764 68336 229770
rect 68284 229706 68336 229712
rect 67548 228676 67600 228682
rect 67548 228618 67600 228624
rect 64788 227724 64840 227730
rect 64788 227666 64840 227672
rect 63222 224496 63278 224505
rect 63222 224431 63278 224440
rect 63052 219406 63172 219434
rect 62764 218068 62816 218074
rect 62764 218010 62816 218016
rect 63144 217274 63172 219406
rect 64604 219156 64656 219162
rect 64604 219098 64656 219104
rect 63960 218068 64012 218074
rect 63960 218010 64012 218016
rect 61442 217110 61516 217138
rect 62270 217110 62344 217138
rect 63098 217246 63172 217274
rect 61442 216988 61470 217110
rect 62270 216988 62298 217110
rect 63098 216988 63126 217246
rect 63972 217138 64000 218010
rect 64616 217274 64644 219098
rect 64800 218074 64828 227666
rect 66168 225616 66220 225622
rect 66168 225558 66220 225564
rect 66180 218074 66208 225558
rect 66904 223304 66956 223310
rect 66904 223246 66956 223252
rect 66916 219162 66944 223246
rect 66904 219156 66956 219162
rect 66904 219098 66956 219104
rect 67560 218210 67588 228618
rect 66444 218204 66496 218210
rect 66444 218146 66496 218152
rect 67548 218204 67600 218210
rect 67548 218146 67600 218152
rect 68100 218204 68152 218210
rect 68100 218146 68152 218152
rect 64788 218068 64840 218074
rect 64788 218010 64840 218016
rect 65616 218068 65668 218074
rect 65616 218010 65668 218016
rect 66168 218068 66220 218074
rect 66168 218010 66220 218016
rect 64616 217246 64782 217274
rect 63926 217110 64000 217138
rect 63926 216988 63954 217110
rect 64754 216988 64782 217246
rect 65628 217138 65656 218010
rect 66456 217138 66484 218146
rect 67272 218068 67324 218074
rect 67272 218010 67324 218016
rect 67284 217138 67312 218010
rect 68112 217138 68140 218146
rect 68296 218074 68324 229706
rect 72424 226024 72476 226030
rect 72424 225966 72476 225972
rect 68928 224120 68980 224126
rect 68928 224062 68980 224068
rect 68284 218068 68336 218074
rect 68284 218010 68336 218016
rect 68940 217274 68968 224062
rect 69572 223168 69624 223174
rect 69572 223110 69624 223116
rect 69584 218210 69612 223110
rect 71412 223032 71464 223038
rect 71412 222974 71464 222980
rect 69756 220516 69808 220522
rect 69756 220458 69808 220464
rect 69572 218204 69624 218210
rect 69572 218146 69624 218152
rect 69768 217274 69796 220458
rect 70584 219428 70636 219434
rect 70584 219370 70636 219376
rect 65582 217110 65656 217138
rect 66410 217110 66484 217138
rect 67238 217110 67312 217138
rect 68066 217110 68140 217138
rect 68894 217246 68968 217274
rect 69722 217246 69796 217274
rect 65582 216988 65610 217110
rect 66410 216988 66438 217110
rect 67238 216988 67266 217110
rect 68066 216988 68094 217110
rect 68894 216988 68922 217246
rect 69722 216988 69750 217246
rect 70596 217138 70624 219370
rect 71424 217274 71452 222974
rect 72436 219026 72464 225966
rect 76564 225752 76616 225758
rect 76564 225694 76616 225700
rect 73712 224392 73764 224398
rect 73712 224334 73764 224340
rect 73068 220380 73120 220386
rect 73068 220322 73120 220328
rect 72424 219020 72476 219026
rect 72424 218962 72476 218968
rect 72240 218068 72292 218074
rect 72240 218010 72292 218016
rect 70550 217110 70624 217138
rect 71378 217246 71452 217274
rect 70550 216988 70578 217110
rect 71378 216988 71406 217246
rect 72252 217138 72280 218010
rect 73080 217274 73108 220322
rect 73724 218074 73752 224334
rect 75828 223440 75880 223446
rect 75828 223382 75880 223388
rect 73896 221468 73948 221474
rect 73896 221410 73948 221416
rect 73712 218068 73764 218074
rect 73712 218010 73764 218016
rect 73908 217274 73936 221410
rect 75552 218204 75604 218210
rect 75552 218146 75604 218152
rect 74724 218068 74776 218074
rect 74724 218010 74776 218016
rect 72206 217110 72280 217138
rect 73034 217246 73108 217274
rect 73862 217246 73936 217274
rect 72206 216988 72234 217110
rect 73034 216988 73062 217246
rect 73862 216988 73890 217246
rect 74736 217138 74764 218010
rect 75564 217138 75592 218146
rect 75840 218074 75868 223382
rect 76380 220108 76432 220114
rect 76380 220050 76432 220056
rect 75828 218068 75880 218074
rect 75828 218010 75880 218016
rect 76392 217274 76420 220050
rect 76576 218210 76604 225694
rect 79968 224664 80020 224670
rect 79968 224606 80020 224612
rect 78588 223576 78640 223582
rect 78588 223518 78640 223524
rect 77208 219020 77260 219026
rect 77208 218962 77260 218968
rect 76564 218204 76616 218210
rect 76564 218146 76616 218152
rect 74690 217110 74764 217138
rect 75518 217110 75592 217138
rect 76346 217246 76420 217274
rect 74690 216988 74718 217110
rect 75518 216988 75546 217110
rect 76346 216988 76374 217246
rect 77220 217138 77248 218962
rect 78600 218074 78628 223518
rect 79692 220244 79744 220250
rect 79692 220186 79744 220192
rect 78036 218068 78088 218074
rect 78036 218010 78088 218016
rect 78588 218068 78640 218074
rect 78588 218010 78640 218016
rect 78864 218068 78916 218074
rect 78864 218010 78916 218016
rect 78048 217138 78076 218010
rect 78876 217138 78904 218010
rect 79704 217274 79732 220186
rect 79980 218074 80008 224606
rect 81348 222760 81400 222766
rect 81348 222702 81400 222708
rect 80520 221740 80572 221746
rect 80520 221682 80572 221688
rect 79968 218068 80020 218074
rect 79968 218010 80020 218016
rect 80532 217274 80560 221682
rect 81360 217274 81388 222702
rect 82096 221474 82124 229978
rect 83464 225888 83516 225894
rect 83464 225830 83516 225836
rect 82084 221468 82136 221474
rect 82084 221410 82136 221416
rect 83004 220924 83056 220930
rect 83004 220866 83056 220872
rect 82176 218068 82228 218074
rect 82176 218010 82228 218016
rect 77174 217110 77248 217138
rect 78002 217110 78076 217138
rect 78830 217110 78904 217138
rect 79658 217246 79732 217274
rect 80486 217246 80560 217274
rect 81314 217246 81388 217274
rect 77174 216988 77202 217110
rect 78002 216988 78030 217110
rect 78830 216988 78858 217110
rect 79658 216988 79686 217246
rect 80486 216988 80514 217246
rect 81314 216988 81342 217246
rect 82188 217138 82216 218010
rect 83016 217274 83044 220866
rect 83476 218074 83504 225830
rect 85488 224528 85540 224534
rect 85488 224470 85540 224476
rect 85304 222352 85356 222358
rect 85304 222294 85356 222300
rect 83832 219156 83884 219162
rect 83832 219098 83884 219104
rect 83464 218068 83516 218074
rect 83464 218010 83516 218016
rect 82142 217110 82216 217138
rect 82970 217246 83044 217274
rect 82142 216988 82170 217110
rect 82970 216988 82998 217246
rect 83844 217138 83872 219098
rect 85316 218074 85344 222294
rect 84660 218068 84712 218074
rect 84660 218010 84712 218016
rect 85304 218068 85356 218074
rect 85304 218010 85356 218016
rect 84672 217138 84700 218010
rect 85500 217274 85528 224470
rect 86236 221746 86264 229978
rect 88248 227860 88300 227866
rect 88248 227802 88300 227808
rect 87972 222488 88024 222494
rect 87972 222430 88024 222436
rect 86224 221740 86276 221746
rect 86224 221682 86276 221688
rect 86316 221468 86368 221474
rect 86316 221410 86368 221416
rect 86328 217274 86356 221410
rect 87144 218068 87196 218074
rect 87144 218010 87196 218016
rect 83798 217110 83872 217138
rect 84626 217110 84700 217138
rect 85454 217246 85528 217274
rect 86282 217246 86356 217274
rect 83798 216988 83826 217110
rect 84626 216988 84654 217110
rect 85454 216988 85482 217246
rect 86282 216988 86310 217246
rect 87156 217138 87184 218010
rect 87984 217274 88012 222430
rect 88260 218074 88288 227802
rect 89628 227316 89680 227322
rect 89628 227258 89680 227264
rect 88984 224392 89036 224398
rect 88984 224334 89036 224340
rect 89444 224392 89496 224398
rect 89444 224334 89496 224340
rect 88996 224126 89024 224334
rect 88984 224120 89036 224126
rect 88984 224062 89036 224068
rect 89456 218074 89484 224334
rect 88248 218068 88300 218074
rect 88248 218010 88300 218016
rect 88800 218068 88852 218074
rect 88800 218010 88852 218016
rect 89444 218068 89496 218074
rect 89444 218010 89496 218016
rect 87110 217110 87184 217138
rect 87938 217246 88012 217274
rect 87110 216988 87138 217110
rect 87938 216988 87966 217246
rect 88812 217138 88840 218010
rect 89640 217274 89668 227258
rect 91284 221332 91336 221338
rect 91284 221274 91336 221280
rect 91296 217274 91324 221274
rect 92400 219434 92428 231134
rect 128268 231056 128320 231062
rect 128268 230998 128320 231004
rect 104808 230920 104860 230926
rect 104808 230862 104860 230868
rect 94504 230648 94556 230654
rect 94504 230590 94556 230596
rect 93584 228812 93636 228818
rect 93584 228754 93636 228760
rect 92124 219406 92428 219434
rect 92124 217274 92152 219406
rect 93596 218074 93624 228754
rect 94516 219434 94544 230590
rect 95240 230172 95292 230178
rect 95240 230114 95292 230120
rect 95252 227866 95280 230114
rect 102140 229492 102192 229498
rect 102140 229434 102192 229440
rect 100668 229084 100720 229090
rect 100668 229026 100720 229032
rect 95240 227860 95292 227866
rect 95240 227802 95292 227808
rect 96436 227452 96488 227458
rect 96436 227394 96488 227400
rect 96252 224936 96304 224942
rect 96252 224878 96304 224884
rect 94688 221740 94740 221746
rect 94688 221682 94740 221688
rect 94700 219434 94728 221682
rect 94424 219406 94544 219434
rect 94608 219406 94728 219434
rect 94424 219298 94452 219406
rect 93768 219292 93820 219298
rect 93768 219234 93820 219240
rect 94412 219292 94464 219298
rect 94412 219234 94464 219240
rect 92940 218068 92992 218074
rect 92940 218010 92992 218016
rect 93584 218068 93636 218074
rect 93584 218010 93636 218016
rect 88766 217110 88840 217138
rect 89594 217246 89668 217274
rect 90410 217252 90462 217258
rect 88766 216988 88794 217110
rect 89594 216988 89622 217246
rect 90410 217194 90462 217200
rect 91250 217246 91324 217274
rect 92078 217246 92152 217274
rect 90422 216988 90450 217194
rect 91250 216988 91278 217246
rect 92078 216988 92106 217246
rect 92952 217138 92980 218010
rect 93780 217138 93808 219234
rect 94608 217274 94636 219406
rect 96264 218074 96292 224878
rect 95424 218068 95476 218074
rect 95424 218010 95476 218016
rect 96252 218068 96304 218074
rect 96252 218010 96304 218016
rect 92906 217110 92980 217138
rect 93734 217110 93808 217138
rect 94562 217246 94636 217274
rect 92906 216988 92934 217110
rect 93734 216988 93762 217110
rect 94562 216988 94590 217246
rect 95436 217138 95464 218010
rect 96448 217274 96476 227394
rect 99288 222624 99340 222630
rect 99288 222566 99340 222572
rect 97908 222012 97960 222018
rect 97908 221954 97960 221960
rect 97080 218204 97132 218210
rect 97080 218146 97132 218152
rect 95390 217110 95464 217138
rect 96218 217246 96476 217274
rect 95390 216988 95418 217110
rect 96218 216988 96246 217246
rect 97092 217138 97120 218146
rect 97920 217274 97948 221954
rect 99300 218074 99328 222566
rect 100392 218340 100444 218346
rect 100392 218282 100444 218288
rect 98736 218068 98788 218074
rect 98736 218010 98788 218016
rect 99288 218068 99340 218074
rect 99288 218010 99340 218016
rect 99564 218068 99616 218074
rect 99564 218010 99616 218016
rect 97046 217110 97120 217138
rect 97874 217246 97948 217274
rect 97046 216988 97074 217110
rect 97874 216988 97902 217246
rect 98748 217138 98776 218010
rect 99576 217138 99604 218010
rect 100404 217138 100432 218282
rect 100680 218074 100708 229026
rect 102152 227594 102180 229434
rect 102140 227588 102192 227594
rect 102140 227530 102192 227536
rect 103428 227588 103480 227594
rect 103428 227530 103480 227536
rect 102048 224800 102100 224806
rect 102048 224742 102100 224748
rect 101220 220652 101272 220658
rect 101220 220594 101272 220600
rect 100668 218068 100720 218074
rect 100668 218010 100720 218016
rect 101232 217274 101260 220594
rect 102060 217274 102088 224742
rect 103440 218142 103468 227530
rect 104532 221876 104584 221882
rect 104532 221818 104584 221824
rect 102876 218136 102928 218142
rect 102876 218078 102928 218084
rect 103428 218136 103480 218142
rect 103428 218078 103480 218084
rect 98702 217110 98776 217138
rect 99530 217110 99604 217138
rect 100358 217110 100432 217138
rect 101186 217246 101260 217274
rect 102014 217246 102088 217274
rect 98702 216988 98730 217110
rect 99530 216988 99558 217110
rect 100358 216988 100386 217110
rect 101186 216988 101214 217246
rect 102014 216988 102042 217246
rect 102888 217138 102916 218078
rect 103704 218068 103756 218074
rect 103704 218010 103756 218016
rect 103716 217138 103744 218010
rect 104544 217274 104572 221818
rect 104820 218074 104848 230862
rect 118608 230784 118660 230790
rect 118608 230726 118660 230732
rect 110328 229356 110380 229362
rect 110328 229298 110380 229304
rect 106188 228948 106240 228954
rect 106188 228890 106240 228896
rect 106004 223984 106056 223990
rect 106004 223926 106056 223932
rect 106016 218074 106044 223926
rect 104808 218068 104860 218074
rect 104808 218010 104860 218016
rect 105360 218068 105412 218074
rect 105360 218010 105412 218016
rect 106004 218068 106056 218074
rect 106004 218010 106056 218016
rect 102842 217110 102916 217138
rect 103670 217110 103744 217138
rect 104498 217246 104572 217274
rect 102842 216988 102870 217110
rect 103670 216988 103698 217110
rect 104498 216988 104526 217246
rect 105372 217138 105400 218010
rect 106200 217274 106228 228890
rect 110340 227730 110368 229298
rect 112996 228268 113048 228274
rect 112996 228210 113048 228216
rect 110328 227724 110380 227730
rect 110328 227666 110380 227672
rect 110512 227724 110564 227730
rect 110512 227666 110564 227672
rect 110524 227610 110552 227666
rect 110340 227582 110552 227610
rect 110144 225480 110196 225486
rect 110144 225422 110196 225428
rect 108672 223848 108724 223854
rect 108672 223790 108724 223796
rect 107844 219972 107896 219978
rect 107844 219914 107896 219920
rect 107016 218612 107068 218618
rect 107016 218554 107068 218560
rect 105326 217110 105400 217138
rect 106154 217246 106228 217274
rect 105326 216988 105354 217110
rect 106154 216988 106182 217246
rect 107028 217138 107056 218554
rect 107856 217274 107884 219914
rect 108684 217274 108712 223790
rect 110156 219434 110184 225422
rect 110156 219406 110276 219434
rect 109500 218068 109552 218074
rect 109500 218010 109552 218016
rect 106982 217110 107056 217138
rect 107810 217246 107884 217274
rect 108638 217246 108712 217274
rect 106982 216988 107010 217110
rect 107810 216988 107838 217246
rect 108638 216988 108666 217246
rect 109512 217138 109540 218010
rect 110248 217274 110276 219406
rect 110340 218090 110368 227582
rect 112812 223712 112864 223718
rect 112812 223654 112864 223660
rect 111156 221060 111208 221066
rect 111156 221002 111208 221008
rect 110340 218074 110460 218090
rect 110340 218068 110472 218074
rect 110340 218062 110420 218068
rect 110420 218010 110472 218016
rect 111168 217274 111196 221002
rect 112824 218074 112852 223654
rect 111984 218068 112036 218074
rect 111984 218010 112036 218016
rect 112812 218068 112864 218074
rect 112812 218010 112864 218016
rect 110248 217246 110322 217274
rect 109466 217110 109540 217138
rect 109466 216988 109494 217110
rect 110294 216988 110322 217246
rect 111122 217246 111196 217274
rect 111122 216988 111150 217246
rect 111996 217138 112024 218010
rect 113008 217274 113036 228210
rect 117228 226772 117280 226778
rect 117228 226714 117280 226720
rect 114284 220788 114336 220794
rect 114284 220730 114336 220736
rect 114296 219978 114324 220730
rect 114284 219972 114336 219978
rect 114284 219914 114336 219920
rect 114468 219972 114520 219978
rect 114468 219914 114520 219920
rect 113640 218340 113692 218346
rect 113640 218282 113692 218288
rect 111950 217110 112024 217138
rect 112778 217246 113036 217274
rect 111950 216988 111978 217110
rect 112778 216988 112806 217246
rect 113652 217138 113680 218282
rect 114480 217274 114508 219914
rect 117240 218074 117268 226714
rect 118424 222216 118476 222222
rect 118424 222158 118476 222164
rect 118148 221332 118200 221338
rect 118148 221274 118200 221280
rect 118160 221066 118188 221274
rect 118148 221060 118200 221066
rect 118148 221002 118200 221008
rect 118436 219434 118464 222158
rect 118620 219434 118648 230726
rect 126888 230308 126940 230314
rect 126888 230250 126940 230256
rect 123484 229220 123536 229226
rect 123484 229162 123536 229168
rect 119988 228132 120040 228138
rect 119988 228074 120040 228080
rect 117596 219428 117648 219434
rect 117596 219370 117648 219376
rect 117780 219428 117832 219434
rect 118436 219406 118556 219434
rect 118620 219428 118752 219434
rect 118620 219406 118700 219428
rect 117780 219370 117832 219376
rect 117608 218210 117636 219370
rect 117596 218204 117648 218210
rect 117596 218146 117648 218152
rect 116124 218068 116176 218074
rect 116124 218010 116176 218016
rect 117228 218068 117280 218074
rect 117228 218010 117280 218016
rect 115296 217456 115348 217462
rect 115296 217398 115348 217404
rect 113606 217110 113680 217138
rect 114434 217246 114508 217274
rect 113606 216988 113634 217110
rect 114434 216988 114462 217246
rect 115308 217138 115336 217398
rect 116136 217138 116164 218010
rect 116952 217592 117004 217598
rect 116952 217534 117004 217540
rect 116964 217138 116992 217534
rect 117792 217138 117820 219370
rect 117964 219292 118016 219298
rect 117964 219234 118016 219240
rect 117976 218618 118004 219234
rect 117964 218612 118016 218618
rect 117964 218554 118016 218560
rect 118148 218612 118200 218618
rect 118148 218554 118200 218560
rect 118160 218346 118188 218554
rect 118148 218340 118200 218346
rect 118148 218282 118200 218288
rect 118528 217274 118556 219406
rect 118700 219370 118752 219376
rect 118712 219339 118740 219370
rect 120000 218074 120028 228074
rect 122748 226908 122800 226914
rect 122748 226850 122800 226856
rect 122564 226296 122616 226302
rect 122564 226238 122616 226244
rect 121092 219836 121144 219842
rect 121092 219778 121144 219784
rect 120264 218340 120316 218346
rect 120264 218282 120316 218288
rect 119436 218068 119488 218074
rect 119436 218010 119488 218016
rect 119988 218068 120040 218074
rect 119988 218010 120040 218016
rect 118528 217246 118602 217274
rect 115262 217110 115336 217138
rect 116090 217110 116164 217138
rect 116918 217110 116992 217138
rect 117746 217110 117820 217138
rect 115262 216988 115290 217110
rect 116090 216988 116118 217110
rect 116918 216988 116946 217110
rect 117746 216988 117774 217110
rect 118574 216988 118602 217246
rect 119448 217138 119476 218010
rect 120276 217138 120304 218282
rect 121104 217274 121132 219778
rect 122576 218074 122604 226238
rect 121920 218068 121972 218074
rect 121920 218010 121972 218016
rect 122564 218068 122616 218074
rect 122564 218010 122616 218016
rect 119402 217110 119476 217138
rect 120230 217110 120304 217138
rect 121058 217246 121132 217274
rect 119402 216988 119430 217110
rect 120230 216988 120258 217110
rect 121058 216988 121086 217246
rect 121932 217138 121960 218010
rect 122760 217274 122788 226850
rect 123496 219434 123524 229162
rect 126704 227996 126756 228002
rect 126704 227938 126756 227944
rect 125232 225344 125284 225350
rect 125232 225286 125284 225292
rect 124404 221060 124456 221066
rect 124404 221002 124456 221008
rect 123404 219406 123524 219434
rect 123404 218210 123432 219406
rect 123392 218204 123444 218210
rect 123392 218146 123444 218152
rect 123576 218204 123628 218210
rect 123576 218146 123628 218152
rect 121886 217110 121960 217138
rect 122714 217246 122788 217274
rect 121886 216988 121914 217110
rect 122714 216988 122742 217246
rect 123588 217138 123616 218146
rect 124416 217274 124444 221002
rect 125244 217274 125272 225286
rect 126716 218074 126744 227938
rect 126060 218068 126112 218074
rect 126060 218010 126112 218016
rect 126704 218068 126756 218074
rect 126704 218010 126756 218016
rect 123542 217110 123616 217138
rect 124370 217246 124444 217274
rect 125198 217246 125272 217274
rect 123542 216988 123570 217110
rect 124370 216988 124398 217246
rect 125198 216988 125226 217246
rect 126072 217138 126100 218010
rect 126900 217274 126928 230250
rect 127624 226160 127676 226166
rect 127624 226102 127676 226108
rect 127636 225486 127664 226102
rect 127624 225480 127676 225486
rect 127624 225422 127676 225428
rect 127440 221332 127492 221338
rect 127440 221274 127492 221280
rect 127452 221066 127480 221274
rect 127256 221060 127308 221066
rect 127256 221002 127308 221008
rect 127440 221060 127492 221066
rect 127440 221002 127492 221008
rect 127900 221060 127952 221066
rect 127900 221002 127952 221008
rect 127268 220946 127296 221002
rect 127912 220946 127940 221002
rect 127268 220918 127940 220946
rect 127624 219972 127676 219978
rect 127624 219914 127676 219920
rect 127636 219706 127664 219914
rect 127624 219700 127676 219706
rect 127624 219642 127676 219648
rect 128280 218074 128308 230998
rect 133788 230444 133840 230450
rect 133788 230386 133840 230392
rect 133512 227860 133564 227866
rect 133512 227802 133564 227808
rect 129556 226636 129608 226642
rect 129556 226578 129608 226584
rect 129372 225344 129424 225350
rect 129372 225286 129424 225292
rect 129384 218074 129412 225286
rect 127716 218068 127768 218074
rect 127716 218010 127768 218016
rect 128268 218068 128320 218074
rect 128268 218010 128320 218016
rect 128544 218068 128596 218074
rect 128544 218010 128596 218016
rect 129372 218068 129424 218074
rect 129372 218010 129424 218016
rect 126026 217110 126100 217138
rect 126854 217246 126928 217274
rect 126026 216988 126054 217110
rect 126854 216988 126882 217246
rect 127728 217138 127756 218010
rect 128556 217138 128584 218010
rect 129568 217274 129596 226578
rect 132408 225072 132460 225078
rect 132408 225014 132460 225020
rect 131028 219700 131080 219706
rect 131028 219642 131080 219648
rect 130200 218068 130252 218074
rect 130200 218010 130252 218016
rect 127682 217110 127756 217138
rect 128510 217110 128584 217138
rect 129338 217246 129596 217274
rect 127682 216988 127710 217110
rect 128510 216988 128538 217110
rect 129338 216988 129366 217246
rect 130212 217138 130240 218010
rect 131040 217274 131068 219642
rect 132420 219434 132448 225014
rect 131856 219428 131908 219434
rect 131856 219370 131908 219376
rect 132408 219428 132460 219434
rect 132408 219370 132460 219376
rect 132592 219428 132644 219434
rect 132592 219370 132644 219376
rect 130166 217110 130240 217138
rect 130994 217246 131068 217274
rect 130166 216988 130194 217110
rect 130994 216988 131022 217246
rect 131868 217138 131896 219370
rect 132604 218226 132632 219370
rect 132512 218198 132632 218226
rect 132512 218074 132540 218198
rect 133524 218074 133552 227802
rect 133800 219434 133828 230386
rect 134996 219434 135024 231406
rect 137664 230518 137692 231406
rect 137652 230512 137704 230518
rect 137652 230454 137704 230460
rect 137468 230444 137520 230450
rect 137468 230386 137520 230392
rect 137480 230042 137508 230386
rect 137284 230036 137336 230042
rect 137284 229978 137336 229984
rect 137468 230036 137520 230042
rect 137468 229978 137520 229984
rect 137296 229634 137324 229978
rect 137284 229628 137336 229634
rect 137284 229570 137336 229576
rect 140042 229120 140098 229129
rect 140042 229055 140098 229064
rect 137376 228540 137428 228546
rect 137376 228482 137428 228488
rect 136824 228404 136876 228410
rect 136824 228346 136876 228352
rect 136638 227896 136694 227905
rect 136836 227866 136864 228346
rect 137388 228290 137416 228482
rect 139308 228404 139360 228410
rect 139308 228346 139360 228352
rect 137204 228274 137416 228290
rect 137192 228268 137416 228274
rect 137244 228262 137416 228268
rect 137192 228210 137244 228216
rect 136638 227831 136640 227840
rect 136692 227831 136694 227840
rect 136824 227860 136876 227866
rect 136640 227802 136692 227808
rect 136824 227802 136876 227808
rect 136548 226500 136600 226506
rect 136548 226442 136600 226448
rect 135168 225208 135220 225214
rect 135168 225150 135220 225156
rect 135180 219434 135208 225150
rect 133708 219406 133828 219434
rect 134352 219406 135024 219434
rect 135088 219406 135208 219434
rect 132500 218068 132552 218074
rect 132500 218010 132552 218016
rect 132684 218068 132736 218074
rect 132684 218010 132736 218016
rect 133512 218068 133564 218074
rect 133512 218010 133564 218016
rect 132696 217138 132724 218010
rect 133708 217274 133736 219406
rect 134352 217274 134380 219406
rect 131822 217110 131896 217138
rect 132650 217110 132724 217138
rect 133478 217246 133736 217274
rect 134306 217246 134380 217274
rect 135088 217274 135116 219406
rect 136560 218074 136588 226442
rect 137282 223952 137338 223961
rect 137282 223887 137338 223896
rect 136916 220516 136968 220522
rect 136916 220458 136968 220464
rect 137100 220516 137152 220522
rect 137100 220458 137152 220464
rect 136928 219570 136956 220458
rect 137112 219842 137140 220458
rect 137100 219836 137152 219842
rect 137100 219778 137152 219784
rect 136916 219564 136968 219570
rect 136916 219506 136968 219512
rect 136916 218204 136968 218210
rect 136916 218146 136968 218152
rect 135996 218068 136048 218074
rect 135996 218010 136048 218016
rect 136548 218068 136600 218074
rect 136548 218010 136600 218016
rect 135088 217246 135162 217274
rect 131822 216988 131850 217110
rect 132650 216988 132678 217110
rect 133478 216988 133506 217246
rect 134306 216988 134334 217246
rect 135134 216988 135162 217246
rect 136008 217138 136036 218010
rect 136928 217274 136956 218146
rect 137296 218074 137324 223887
rect 138294 221640 138350 221649
rect 138294 221575 138296 221584
rect 138348 221575 138350 221584
rect 138480 221604 138532 221610
rect 138296 221546 138348 221552
rect 138480 221546 138532 221552
rect 137652 219564 137704 219570
rect 137652 219506 137704 219512
rect 137284 218068 137336 218074
rect 137284 218010 137336 218016
rect 137664 217274 137692 219506
rect 138492 217274 138520 221546
rect 139320 217274 139348 228346
rect 140056 219434 140084 229055
rect 141160 227866 141188 231676
rect 141344 231662 141818 231690
rect 141148 227860 141200 227866
rect 141148 227802 141200 227808
rect 140778 222048 140834 222057
rect 140778 221983 140834 221992
rect 140792 221610 140820 221983
rect 141344 221649 141372 231662
rect 141514 227896 141570 227905
rect 141514 227831 141516 227840
rect 141568 227831 141570 227840
rect 141516 227802 141568 227808
rect 142448 227050 142476 231676
rect 143092 228274 143120 231676
rect 143552 231662 143750 231690
rect 144012 231662 144394 231690
rect 143552 229129 143580 231662
rect 143538 229120 143594 229129
rect 143538 229055 143594 229064
rect 143080 228268 143132 228274
rect 143080 228210 143132 228216
rect 143448 228268 143500 228274
rect 143448 228210 143500 228216
rect 142436 227044 142488 227050
rect 142436 226986 142488 226992
rect 143264 227044 143316 227050
rect 143264 226986 143316 226992
rect 141606 226536 141662 226545
rect 141606 226471 141608 226480
rect 141660 226471 141662 226480
rect 142250 226536 142306 226545
rect 142250 226471 142252 226480
rect 141608 226442 141660 226448
rect 142304 226471 142306 226480
rect 142252 226442 142304 226448
rect 141792 226432 141844 226438
rect 141792 226374 141844 226380
rect 142114 226432 142166 226438
rect 142166 226380 142292 226386
rect 142114 226374 142292 226380
rect 141330 221640 141386 221649
rect 140780 221604 140832 221610
rect 140780 221546 140832 221552
rect 140964 221604 141016 221610
rect 141330 221575 141386 221584
rect 140964 221546 141016 221552
rect 139964 219406 140084 219434
rect 139964 218890 139992 219406
rect 139952 218884 140004 218890
rect 139952 218826 140004 218832
rect 140136 218068 140188 218074
rect 140136 218010 140188 218016
rect 135962 217110 136036 217138
rect 136790 217246 136956 217274
rect 137618 217246 137692 217274
rect 138446 217246 138520 217274
rect 139274 217246 139348 217274
rect 135962 216988 135990 217110
rect 136790 216988 136818 217246
rect 137618 216988 137646 217246
rect 138446 216988 138474 217246
rect 139274 216988 139302 217246
rect 140148 217138 140176 218010
rect 140976 217274 141004 221546
rect 141804 217274 141832 226374
rect 142126 226358 142292 226374
rect 142264 226166 142292 226358
rect 142114 226160 142166 226166
rect 142114 226102 142166 226108
rect 142252 226160 142304 226166
rect 142252 226102 142304 226108
rect 142126 226012 142154 226102
rect 142126 225984 142292 226012
rect 142264 225622 142292 225984
rect 142114 225616 142166 225622
rect 142112 225584 142114 225593
rect 142252 225616 142304 225622
rect 142166 225584 142168 225593
rect 142252 225558 142304 225564
rect 142112 225519 142168 225528
rect 142126 224182 142476 224210
rect 142126 224126 142154 224182
rect 142114 224120 142166 224126
rect 142114 224062 142166 224068
rect 142252 224120 142304 224126
rect 142252 224062 142304 224068
rect 142264 223961 142292 224062
rect 142448 223961 142476 224182
rect 142250 223952 142306 223961
rect 142250 223887 142306 223896
rect 142434 223952 142490 223961
rect 142434 223887 142490 223896
rect 141976 222896 142028 222902
rect 141974 222864 141976 222873
rect 142160 222896 142212 222902
rect 142028 222864 142030 222873
rect 141974 222799 142030 222808
rect 142158 222864 142160 222873
rect 142212 222864 142214 222873
rect 142158 222799 142214 222808
rect 141988 222686 142200 222714
rect 141988 222222 142016 222686
rect 142172 222222 142200 222686
rect 141976 222216 142028 222222
rect 141976 222158 142028 222164
rect 142160 222216 142212 222222
rect 142160 222158 142212 222164
rect 141974 222048 142030 222057
rect 142030 222006 142292 222034
rect 141974 221983 142030 221992
rect 142112 220960 142168 220969
rect 142264 220930 142292 222006
rect 142112 220895 142114 220904
rect 142166 220895 142168 220904
rect 142252 220924 142304 220930
rect 142114 220866 142166 220872
rect 142252 220866 142304 220872
rect 142252 218884 142304 218890
rect 142252 218826 142304 218832
rect 142264 218482 142292 218826
rect 142252 218476 142304 218482
rect 142252 218418 142304 218424
rect 142436 218476 142488 218482
rect 142436 218418 142488 218424
rect 142448 218074 142476 218418
rect 143276 218074 143304 226986
rect 142436 218068 142488 218074
rect 142436 218010 142488 218016
rect 142620 218068 142672 218074
rect 142620 218010 142672 218016
rect 143264 218068 143316 218074
rect 143264 218010 143316 218016
rect 140102 217110 140176 217138
rect 140930 217246 141004 217274
rect 141758 217246 141832 217274
rect 140102 216988 140130 217110
rect 140930 216988 140958 217246
rect 141758 216988 141786 217246
rect 142632 217138 142660 218010
rect 143460 217274 143488 228210
rect 144012 222902 144040 231662
rect 144642 230480 144698 230489
rect 144642 230415 144698 230424
rect 144458 229800 144514 229809
rect 144458 229735 144460 229744
rect 144512 229735 144514 229744
rect 144460 229706 144512 229712
rect 144000 222896 144052 222902
rect 144000 222838 144052 222844
rect 144656 219706 144684 230415
rect 144828 229764 144880 229770
rect 144828 229706 144880 229712
rect 144840 227186 144868 229706
rect 145024 229094 145052 231676
rect 145668 229498 145696 231676
rect 146312 229770 146340 231676
rect 146680 231662 146970 231690
rect 146300 229764 146352 229770
rect 146300 229706 146352 229712
rect 145656 229492 145708 229498
rect 145656 229434 145708 229440
rect 146024 229424 146076 229430
rect 145838 229392 145894 229401
rect 146024 229366 146076 229372
rect 145838 229327 145840 229336
rect 145892 229327 145894 229336
rect 145840 229298 145892 229304
rect 145024 229066 145144 229094
rect 144828 227180 144880 227186
rect 144828 227122 144880 227128
rect 144644 219700 144696 219706
rect 144644 219642 144696 219648
rect 144828 219700 144880 219706
rect 144828 219642 144880 219648
rect 144840 218074 144868 219642
rect 145116 218754 145144 229066
rect 146036 228274 146064 229366
rect 146208 228676 146260 228682
rect 146208 228618 146260 228624
rect 146220 228274 146248 228618
rect 146024 228268 146076 228274
rect 146024 228210 146076 228216
rect 146208 228268 146260 228274
rect 146208 228210 146260 228216
rect 146206 228032 146262 228041
rect 146206 227967 146262 227976
rect 146024 222896 146076 222902
rect 146024 222838 146076 222844
rect 145562 221232 145618 221241
rect 145562 221167 145618 221176
rect 145576 220930 145604 221167
rect 145564 220924 145616 220930
rect 145564 220866 145616 220872
rect 145840 220788 145892 220794
rect 145840 220730 145892 220736
rect 145654 220416 145710 220425
rect 145852 220386 145880 220730
rect 145654 220351 145656 220360
rect 145708 220351 145710 220360
rect 145840 220380 145892 220386
rect 145656 220322 145708 220328
rect 145840 220322 145892 220328
rect 146036 219434 146064 222838
rect 146220 219434 146248 227967
rect 146680 223310 146708 231662
rect 147128 228540 147180 228546
rect 147128 228482 147180 228488
rect 147140 228041 147168 228482
rect 147126 228032 147182 228041
rect 147126 227967 147182 227976
rect 147600 226030 147628 231676
rect 147968 231662 148258 231690
rect 147968 229401 147996 231662
rect 148324 229424 148376 229430
rect 147954 229392 148010 229401
rect 148324 229366 148376 229372
rect 147954 229327 148010 229336
rect 147588 226024 147640 226030
rect 147588 225966 147640 225972
rect 147772 226024 147824 226030
rect 147772 225966 147824 225972
rect 147784 225593 147812 225966
rect 147770 225584 147826 225593
rect 147770 225519 147826 225528
rect 146668 223304 146720 223310
rect 146668 223246 146720 223252
rect 147312 223304 147364 223310
rect 147312 223246 147364 223252
rect 146390 221232 146446 221241
rect 146390 221167 146446 221176
rect 146404 221066 146432 221167
rect 146392 221060 146444 221066
rect 146392 221002 146444 221008
rect 146944 220788 146996 220794
rect 146944 220730 146996 220736
rect 146956 220522 146984 220730
rect 146944 220516 146996 220522
rect 146944 220458 146996 220464
rect 147128 220516 147180 220522
rect 147128 220458 147180 220464
rect 147140 219722 147168 220458
rect 146772 219706 147168 219722
rect 146760 219700 147168 219706
rect 146812 219694 147168 219700
rect 146760 219642 146812 219648
rect 147324 219434 147352 223246
rect 148336 220425 148364 229366
rect 148888 228274 148916 231676
rect 148876 228268 148928 228274
rect 148876 228210 148928 228216
rect 148874 225992 148930 226001
rect 148874 225927 148930 225936
rect 148322 220416 148378 220425
rect 148322 220351 148378 220360
rect 147588 219564 147640 219570
rect 147588 219506 147640 219512
rect 145944 219406 146064 219434
rect 146128 219406 146248 219434
rect 146956 219406 147352 219434
rect 145104 218748 145156 218754
rect 145104 218690 145156 218696
rect 145944 218074 145972 219406
rect 144276 218068 144328 218074
rect 144276 218010 144328 218016
rect 144828 218068 144880 218074
rect 144828 218010 144880 218016
rect 145104 218068 145156 218074
rect 145104 218010 145156 218016
rect 145932 218068 145984 218074
rect 145932 218010 145984 218016
rect 142586 217110 142660 217138
rect 143414 217246 143488 217274
rect 142586 216988 142614 217110
rect 143414 216988 143442 217246
rect 144288 217138 144316 218010
rect 145116 217138 145144 218010
rect 146128 217274 146156 219406
rect 146956 218890 146984 219406
rect 146944 218884 146996 218890
rect 146944 218826 146996 218832
rect 146760 218748 146812 218754
rect 146760 218690 146812 218696
rect 146772 217274 146800 218690
rect 147600 217274 147628 219506
rect 148888 218074 148916 225927
rect 149532 223174 149560 231676
rect 149808 231662 150190 231690
rect 150544 231662 150834 231690
rect 151096 231662 151478 231690
rect 149808 226030 149836 231662
rect 150346 230208 150402 230217
rect 150346 230143 150402 230152
rect 150072 227180 150124 227186
rect 150072 227122 150124 227128
rect 149796 226024 149848 226030
rect 149796 225966 149848 225972
rect 149520 223168 149572 223174
rect 149520 223110 149572 223116
rect 150084 218074 150112 227122
rect 150360 219434 150388 230143
rect 150544 229809 150572 231662
rect 151096 230489 151124 231662
rect 151082 230480 151138 230489
rect 151082 230415 151138 230424
rect 151910 230208 151966 230217
rect 151910 230143 151966 230152
rect 151924 229906 151952 230143
rect 151728 229900 151780 229906
rect 151728 229842 151780 229848
rect 151912 229900 151964 229906
rect 151912 229842 151964 229848
rect 150530 229800 150586 229809
rect 150530 229735 150586 229744
rect 151004 229758 151400 229786
rect 151004 229566 151032 229758
rect 151176 229628 151228 229634
rect 151176 229570 151228 229576
rect 150992 229560 151044 229566
rect 150992 229502 151044 229508
rect 151188 220969 151216 229570
rect 151372 229514 151400 229758
rect 151740 229616 151768 229842
rect 151740 229588 151952 229616
rect 151372 229498 151814 229514
rect 151372 229492 151826 229498
rect 151372 229486 151774 229492
rect 151774 229434 151826 229440
rect 151636 229424 151688 229430
rect 151636 229366 151688 229372
rect 151648 229265 151676 229366
rect 151634 229256 151690 229265
rect 151924 229226 151952 229588
rect 151634 229191 151690 229200
rect 151912 229220 151964 229226
rect 151912 229162 151964 229168
rect 151912 226024 151964 226030
rect 151910 225992 151912 226001
rect 151964 225992 151966 226001
rect 151910 225927 151966 225936
rect 151464 225814 151952 225842
rect 151174 220960 151230 220969
rect 151174 220895 151230 220904
rect 150268 219406 150388 219434
rect 151464 219434 151492 225814
rect 151924 225758 151952 225814
rect 151728 225752 151780 225758
rect 151726 225720 151728 225729
rect 151912 225752 151964 225758
rect 151780 225720 151782 225729
rect 151912 225694 151964 225700
rect 151726 225655 151782 225664
rect 151634 224496 151690 224505
rect 151634 224431 151690 224440
rect 151648 224262 151676 224431
rect 151636 224256 151688 224262
rect 151636 224198 151688 224204
rect 151774 224256 151826 224262
rect 151774 224198 151826 224204
rect 151786 224074 151814 224198
rect 151648 224046 151814 224074
rect 151648 223961 151676 224046
rect 151634 223952 151690 223961
rect 151634 223887 151690 223896
rect 152108 223174 152136 231676
rect 152384 231662 152766 231690
rect 152384 224505 152412 231662
rect 153396 229362 153424 231676
rect 153672 231662 154054 231690
rect 154698 231662 154988 231690
rect 153384 229356 153436 229362
rect 153384 229298 153436 229304
rect 153672 229265 153700 231662
rect 154026 229800 154082 229809
rect 154026 229735 154028 229744
rect 154080 229735 154082 229744
rect 154212 229764 154264 229770
rect 154028 229706 154080 229712
rect 154212 229706 154264 229712
rect 153844 229356 153896 229362
rect 153844 229298 153896 229304
rect 153658 229256 153714 229265
rect 153658 229191 153714 229200
rect 153106 228440 153162 228449
rect 153106 228375 153162 228384
rect 153476 228404 153528 228410
rect 152370 224496 152426 224505
rect 152370 224431 152426 224440
rect 152096 223168 152148 223174
rect 152096 223110 152148 223116
rect 151464 219406 151676 219434
rect 148416 218068 148468 218074
rect 148416 218010 148468 218016
rect 148876 218068 148928 218074
rect 148876 218010 148928 218016
rect 149244 218068 149296 218074
rect 149244 218010 149296 218016
rect 150072 218068 150124 218074
rect 150072 218010 150124 218016
rect 144242 217110 144316 217138
rect 145070 217110 145144 217138
rect 145898 217246 146156 217274
rect 146726 217246 146800 217274
rect 147554 217246 147628 217274
rect 144242 216988 144270 217110
rect 145070 216988 145098 217110
rect 145898 216988 145926 217246
rect 146726 216988 146754 217246
rect 147554 216988 147582 217246
rect 148428 217138 148456 218010
rect 149256 217138 149284 218010
rect 150268 217274 150296 219406
rect 150624 219020 150676 219026
rect 150624 218962 150676 218968
rect 150636 218482 150664 218962
rect 150900 218884 150952 218890
rect 150900 218826 150952 218832
rect 150440 218476 150492 218482
rect 150440 218418 150492 218424
rect 150624 218476 150676 218482
rect 150624 218418 150676 218424
rect 150452 218210 150480 218418
rect 150440 218204 150492 218210
rect 150440 218146 150492 218152
rect 148382 217110 148456 217138
rect 149210 217110 149284 217138
rect 150038 217246 150296 217274
rect 148382 216988 148410 217110
rect 149210 216988 149238 217110
rect 150038 216988 150066 217246
rect 150912 217138 150940 218826
rect 151648 217274 151676 219406
rect 152372 219020 152424 219026
rect 152372 218962 152424 218968
rect 152384 218482 152412 218962
rect 153120 218482 153148 228375
rect 153476 228346 153528 228352
rect 153488 220386 153516 228346
rect 153660 223032 153712 223038
rect 153660 222974 153712 222980
rect 153672 222766 153700 222974
rect 153660 222760 153712 222766
rect 153660 222702 153712 222708
rect 153476 220380 153528 220386
rect 153476 220322 153528 220328
rect 153856 219026 153884 229298
rect 154224 228410 154252 229706
rect 154394 228440 154450 228449
rect 154212 228404 154264 228410
rect 154394 228375 154396 228384
rect 154212 228346 154264 228352
rect 154448 228375 154450 228384
rect 154396 228346 154448 228352
rect 154304 225752 154356 225758
rect 154356 225700 154712 225706
rect 154304 225694 154712 225700
rect 154316 225678 154712 225694
rect 154684 225622 154712 225678
rect 154672 225616 154724 225622
rect 154672 225558 154724 225564
rect 154028 223576 154080 223582
rect 154028 223518 154080 223524
rect 154212 223576 154264 223582
rect 154212 223518 154264 223524
rect 154040 222766 154068 223518
rect 154028 222760 154080 222766
rect 154028 222702 154080 222708
rect 154224 222358 154252 223518
rect 154960 223446 154988 231662
rect 155328 224262 155356 231676
rect 155972 229226 156000 231676
rect 156156 231662 156630 231690
rect 156984 231662 157274 231690
rect 157536 231662 157918 231690
rect 158088 231662 158562 231690
rect 158916 231662 159206 231690
rect 155960 229220 156012 229226
rect 155960 229162 156012 229168
rect 155866 227080 155922 227089
rect 155866 227015 155922 227024
rect 155316 224256 155368 224262
rect 155316 224198 155368 224204
rect 154948 223440 155000 223446
rect 154948 223382 155000 223388
rect 155500 223440 155552 223446
rect 155500 223382 155552 223388
rect 154396 223168 154448 223174
rect 154396 223110 154448 223116
rect 154212 222352 154264 222358
rect 154212 222294 154264 222300
rect 154408 221354 154436 223110
rect 155512 223038 155540 223382
rect 155500 223032 155552 223038
rect 155500 222974 155552 222980
rect 155684 223032 155736 223038
rect 155684 222974 155736 222980
rect 154224 221326 154436 221354
rect 153844 219020 153896 219026
rect 153844 218962 153896 218968
rect 154028 219020 154080 219026
rect 154028 218962 154080 218968
rect 154040 218482 154068 218962
rect 152372 218476 152424 218482
rect 152372 218418 152424 218424
rect 152556 218476 152608 218482
rect 152556 218418 152608 218424
rect 153108 218476 153160 218482
rect 153108 218418 153160 218424
rect 153384 218476 153436 218482
rect 153384 218418 153436 218424
rect 154028 218476 154080 218482
rect 154028 218418 154080 218424
rect 151648 217246 151722 217274
rect 150866 217110 150940 217138
rect 150866 216988 150894 217110
rect 151694 216988 151722 217246
rect 152568 217138 152596 218418
rect 153396 217138 153424 218418
rect 154224 217274 154252 221326
rect 154396 220380 154448 220386
rect 154396 220322 154448 220328
rect 154408 218890 154436 220322
rect 154396 218884 154448 218890
rect 154396 218826 154448 218832
rect 155696 218482 155724 222974
rect 155040 218476 155092 218482
rect 155040 218418 155092 218424
rect 155684 218476 155736 218482
rect 155684 218418 155736 218424
rect 152522 217110 152596 217138
rect 153350 217110 153424 217138
rect 154178 217246 154252 217274
rect 152522 216988 152550 217110
rect 153350 216988 153378 217110
rect 154178 216988 154206 217246
rect 155052 217138 155080 218418
rect 155880 217274 155908 227015
rect 156156 220114 156184 231662
rect 156984 222766 157012 231662
rect 157248 229220 157300 229226
rect 157248 229162 157300 229168
rect 156972 222760 157024 222766
rect 156972 222702 157024 222708
rect 156144 220108 156196 220114
rect 156144 220050 156196 220056
rect 157260 218482 157288 229162
rect 157536 225729 157564 231662
rect 158088 229514 158116 231662
rect 157812 229486 158116 229514
rect 157812 229362 157840 229486
rect 157800 229356 157852 229362
rect 157800 229298 157852 229304
rect 157984 229356 158036 229362
rect 157984 229298 158036 229304
rect 157522 225720 157578 225729
rect 157522 225655 157578 225664
rect 157524 220108 157576 220114
rect 157524 220050 157576 220056
rect 156696 218476 156748 218482
rect 156696 218418 156748 218424
rect 157248 218476 157300 218482
rect 157248 218418 157300 218424
rect 155006 217110 155080 217138
rect 155834 217246 155908 217274
rect 155006 216988 155034 217110
rect 155834 216988 155862 217246
rect 156708 217138 156736 218418
rect 157536 217274 157564 220050
rect 157996 219162 158024 229298
rect 158350 220960 158406 220969
rect 158350 220895 158406 220904
rect 157984 219156 158036 219162
rect 157984 219098 158036 219104
rect 158364 217274 158392 220895
rect 158916 220250 158944 231662
rect 159836 229094 159864 231676
rect 159192 229066 159864 229094
rect 159192 223446 159220 229066
rect 160006 228440 160062 228449
rect 160006 228375 160062 228384
rect 159180 223440 159232 223446
rect 159180 223382 159232 223388
rect 159364 223440 159416 223446
rect 159364 223382 159416 223388
rect 158904 220244 158956 220250
rect 158904 220186 158956 220192
rect 159376 219298 159404 223382
rect 159364 219292 159416 219298
rect 159364 219234 159416 219240
rect 159824 218884 159876 218890
rect 159824 218826 159876 218832
rect 159180 218476 159232 218482
rect 159180 218418 159232 218424
rect 156662 217110 156736 217138
rect 157490 217246 157564 217274
rect 158318 217246 158392 217274
rect 156662 216988 156690 217110
rect 157490 216988 157518 217246
rect 158318 216988 158346 217246
rect 159192 217138 159220 218418
rect 159836 217274 159864 218826
rect 160020 218482 160048 228375
rect 160480 224670 160508 231676
rect 160848 231662 161138 231690
rect 160848 229809 160876 231662
rect 160834 229800 160890 229809
rect 161768 229770 161796 231676
rect 162136 231662 162426 231690
rect 160834 229735 160890 229744
rect 161388 229764 161440 229770
rect 161388 229706 161440 229712
rect 161756 229764 161808 229770
rect 161756 229706 161808 229712
rect 161400 229514 161428 229706
rect 161756 229628 161808 229634
rect 161756 229570 161808 229576
rect 161400 229486 161474 229514
rect 161294 229392 161350 229401
rect 161294 229327 161350 229336
rect 161308 229226 161336 229327
rect 161446 229242 161474 229486
rect 161768 229401 161796 229570
rect 161754 229392 161810 229401
rect 161754 229327 161810 229336
rect 161446 229226 161520 229242
rect 161296 229220 161348 229226
rect 161446 229220 161532 229226
rect 161446 229214 161480 229220
rect 161296 229162 161348 229168
rect 161480 229162 161532 229168
rect 162136 229094 162164 231662
rect 161952 229066 162164 229094
rect 161432 228848 161488 228857
rect 161432 228783 161434 228792
rect 161486 228783 161488 228792
rect 161572 228812 161624 228818
rect 161434 228754 161486 228760
rect 161572 228754 161624 228760
rect 161584 228449 161612 228754
rect 161570 228440 161626 228449
rect 161570 228375 161626 228384
rect 161432 227352 161488 227361
rect 161432 227287 161434 227296
rect 161486 227287 161488 227296
rect 161572 227316 161624 227322
rect 161434 227258 161486 227264
rect 161572 227258 161624 227264
rect 161584 227089 161612 227258
rect 161570 227080 161626 227089
rect 161570 227015 161626 227024
rect 160468 224664 160520 224670
rect 160468 224606 160520 224612
rect 161952 223582 161980 229066
rect 163056 225894 163084 231676
rect 163700 229362 163728 231676
rect 164344 230194 164372 231676
rect 164344 230166 164464 230194
rect 163964 229764 164016 229770
rect 163964 229706 164016 229712
rect 163688 229356 163740 229362
rect 163688 229298 163740 229304
rect 163044 225888 163096 225894
rect 163044 225830 163096 225836
rect 162768 224664 162820 224670
rect 162768 224606 162820 224612
rect 161940 223576 161992 223582
rect 161940 223518 161992 223524
rect 162124 223576 162176 223582
rect 162124 223518 162176 223524
rect 160836 222148 160888 222154
rect 160836 222090 160888 222096
rect 160192 219020 160244 219026
rect 160192 218962 160244 218968
rect 160204 218482 160232 218962
rect 160008 218476 160060 218482
rect 160008 218418 160060 218424
rect 160192 218476 160244 218482
rect 160192 218418 160244 218424
rect 160848 217274 160876 222090
rect 161432 221776 161488 221785
rect 161432 221711 161434 221720
rect 161486 221711 161488 221720
rect 161572 221740 161624 221746
rect 161434 221682 161486 221688
rect 161572 221682 161624 221688
rect 161584 221626 161612 221682
rect 161446 221598 161612 221626
rect 161446 221338 161474 221598
rect 161756 221468 161808 221474
rect 161756 221410 161808 221416
rect 161434 221332 161486 221338
rect 161434 221274 161486 221280
rect 161768 221082 161796 221410
rect 161446 221054 161796 221082
rect 161446 220930 161474 221054
rect 161570 220960 161626 220969
rect 161434 220924 161486 220930
rect 161570 220895 161572 220904
rect 161434 220866 161486 220872
rect 161624 220895 161626 220904
rect 161572 220866 161624 220872
rect 161480 219020 161532 219026
rect 161480 218962 161532 218968
rect 161492 218346 161520 218962
rect 162136 218618 162164 223518
rect 162492 219292 162544 219298
rect 162492 219234 162544 219240
rect 162124 218612 162176 218618
rect 162124 218554 162176 218560
rect 161480 218340 161532 218346
rect 161480 218282 161532 218288
rect 161664 218340 161716 218346
rect 161664 218282 161716 218288
rect 159836 217246 160002 217274
rect 159146 217110 159220 217138
rect 159146 216988 159174 217110
rect 159974 216988 160002 217246
rect 160802 217246 160876 217274
rect 160802 216988 160830 217246
rect 161676 217138 161704 218282
rect 162504 217138 162532 219234
rect 162780 218346 162808 224606
rect 163976 218346 164004 229706
rect 164240 229356 164292 229362
rect 164240 229298 164292 229304
rect 164252 228857 164280 229298
rect 164238 228848 164294 228857
rect 164238 228783 164294 228792
rect 164436 221338 164464 230166
rect 164988 222494 165016 231676
rect 165632 224534 165660 231676
rect 166000 231662 166290 231690
rect 166000 230178 166028 231662
rect 165988 230172 166040 230178
rect 165988 230114 166040 230120
rect 166264 230172 166316 230178
rect 166264 230114 166316 230120
rect 166276 229906 166304 230114
rect 166264 229900 166316 229906
rect 166264 229842 166316 229848
rect 166540 228812 166592 228818
rect 166540 228754 166592 228760
rect 166552 228698 166580 228754
rect 166000 228682 166580 228698
rect 165988 228676 166580 228682
rect 166040 228670 166580 228676
rect 165988 228618 166040 228624
rect 166920 227361 166948 231676
rect 167196 231662 167578 231690
rect 167840 231662 168222 231690
rect 168576 231662 168866 231690
rect 169128 231662 169510 231690
rect 169772 231662 170154 231690
rect 166906 227352 166962 227361
rect 166906 227287 166962 227296
rect 165620 224528 165672 224534
rect 165620 224470 165672 224476
rect 165528 224256 165580 224262
rect 165528 224198 165580 224204
rect 164976 222488 165028 222494
rect 164976 222430 165028 222436
rect 164424 221332 164476 221338
rect 164424 221274 164476 221280
rect 164148 220244 164200 220250
rect 164148 220186 164200 220192
rect 162768 218340 162820 218346
rect 162768 218282 162820 218288
rect 163320 218340 163372 218346
rect 163320 218282 163372 218288
rect 163964 218340 164016 218346
rect 163964 218282 164016 218288
rect 163332 217138 163360 218282
rect 164160 217274 164188 220186
rect 165540 218346 165568 224198
rect 166264 222760 166316 222766
rect 166264 222702 166316 222708
rect 166080 222148 166132 222154
rect 166080 222090 166132 222096
rect 166092 221202 166120 222090
rect 166080 221196 166132 221202
rect 166080 221138 166132 221144
rect 165804 219156 165856 219162
rect 165804 219098 165856 219104
rect 164976 218340 165028 218346
rect 164976 218282 165028 218288
rect 165528 218340 165580 218346
rect 165528 218282 165580 218288
rect 161630 217110 161704 217138
rect 162458 217110 162532 217138
rect 163286 217110 163360 217138
rect 164114 217246 164188 217274
rect 161630 216988 161658 217110
rect 162458 216988 162486 217110
rect 163286 216988 163314 217110
rect 164114 216988 164142 217246
rect 164988 217138 165016 218282
rect 165816 217138 165844 219098
rect 166276 219026 166304 222702
rect 167000 222012 167052 222018
rect 167000 221954 167052 221960
rect 167012 221785 167040 221954
rect 166998 221776 167054 221785
rect 167196 221746 167224 231662
rect 167840 224398 167868 231662
rect 167828 224392 167880 224398
rect 167828 224334 167880 224340
rect 168288 224392 168340 224398
rect 168288 224334 168340 224340
rect 166998 221711 167054 221720
rect 167184 221740 167236 221746
rect 167184 221682 167236 221688
rect 167460 221740 167512 221746
rect 167460 221682 167512 221688
rect 166264 219020 166316 219026
rect 166264 218962 166316 218968
rect 166632 218612 166684 218618
rect 166632 218554 166684 218560
rect 166644 217138 166672 218554
rect 167472 217138 167500 221682
rect 168300 217138 168328 224334
rect 168576 217326 168604 231662
rect 169128 229362 169156 231662
rect 169116 229356 169168 229362
rect 169116 229298 169168 229304
rect 169574 227216 169630 227225
rect 169574 227151 169630 227160
rect 168930 219464 168986 219473
rect 169588 219434 169616 227151
rect 169772 222018 169800 231662
rect 170784 231198 170812 231676
rect 170772 231192 170824 231198
rect 170772 231134 170824 231140
rect 171428 230654 171456 231676
rect 171704 231662 172086 231690
rect 171416 230648 171468 230654
rect 171416 230590 171468 230596
rect 170956 229356 171008 229362
rect 170956 229298 171008 229304
rect 170770 227488 170826 227497
rect 170770 227423 170772 227432
rect 170824 227423 170826 227432
rect 170772 227394 170824 227400
rect 169760 222012 169812 222018
rect 169760 221954 169812 221960
rect 169758 219464 169814 219473
rect 168930 219399 168932 219408
rect 168984 219399 168986 219408
rect 169116 219428 169168 219434
rect 168932 219370 168984 219376
rect 169116 219370 169168 219376
rect 169576 219428 169628 219434
rect 169758 219399 169760 219408
rect 169576 219370 169628 219376
rect 169812 219399 169814 219408
rect 169760 219370 169812 219376
rect 168564 217320 168616 217326
rect 168564 217262 168616 217268
rect 169128 217138 169156 219370
rect 169760 219020 169812 219026
rect 169760 218962 169812 218968
rect 169772 218618 169800 218962
rect 170968 218618 170996 229298
rect 171704 227497 171732 231662
rect 171690 227488 171746 227497
rect 171094 227452 171146 227458
rect 171690 227423 171746 227432
rect 171094 227394 171146 227400
rect 171106 227225 171134 227394
rect 171092 227216 171148 227225
rect 171092 227151 171148 227160
rect 172152 222420 172204 222426
rect 172152 222362 172204 222368
rect 171784 222012 171836 222018
rect 171784 221954 171836 221960
rect 171416 221740 171468 221746
rect 171416 221682 171468 221688
rect 171600 221740 171652 221746
rect 171600 221682 171652 221688
rect 171428 221513 171456 221682
rect 171414 221504 171470 221513
rect 171414 221439 171470 221448
rect 171612 221338 171640 221682
rect 171600 221332 171652 221338
rect 171600 221274 171652 221280
rect 171600 219292 171652 219298
rect 171600 219234 171652 219240
rect 171612 218618 171640 219234
rect 169760 218612 169812 218618
rect 169760 218554 169812 218560
rect 169944 218612 169996 218618
rect 169944 218554 169996 218560
rect 170956 218612 171008 218618
rect 170956 218554 171008 218560
rect 171600 218612 171652 218618
rect 171600 218554 171652 218560
rect 169956 217138 169984 218554
rect 171796 218498 171824 221954
rect 171966 221504 172022 221513
rect 171966 221439 171968 221448
rect 172020 221439 172022 221448
rect 171968 221410 172020 221416
rect 172164 219434 172192 222362
rect 172716 222154 172744 231676
rect 173162 228848 173218 228857
rect 173162 228783 173218 228792
rect 172704 222148 172756 222154
rect 172704 222090 172756 222096
rect 173176 219434 173204 228783
rect 173360 224942 173388 231676
rect 174018 231662 174216 231690
rect 173716 229764 173768 229770
rect 173716 229706 173768 229712
rect 173728 229226 173756 229706
rect 173716 229220 173768 229226
rect 173716 229162 173768 229168
rect 173900 229220 173952 229226
rect 173900 229162 173952 229168
rect 173912 228954 173940 229162
rect 173900 228948 173952 228954
rect 173900 228890 173952 228896
rect 174188 224954 174216 231662
rect 174648 229090 174676 231676
rect 175306 231662 175596 231690
rect 174820 229220 174872 229226
rect 174820 229162 174872 229168
rect 174832 229090 174860 229162
rect 174636 229084 174688 229090
rect 174636 229026 174688 229032
rect 174820 229084 174872 229090
rect 174820 229026 174872 229032
rect 175370 227624 175426 227633
rect 175370 227559 175372 227568
rect 175424 227559 175426 227568
rect 175372 227530 175424 227536
rect 175568 224954 175596 231662
rect 173348 224936 173400 224942
rect 174188 224926 174308 224954
rect 173348 224878 173400 224884
rect 174084 222148 174136 222154
rect 174084 222090 174136 222096
rect 172152 219428 172204 219434
rect 172152 219370 172204 219376
rect 172428 219428 172480 219434
rect 172428 219370 172480 219376
rect 173164 219428 173216 219434
rect 173164 219370 173216 219376
rect 171968 219156 172020 219162
rect 171968 219098 172020 219104
rect 171612 218470 171824 218498
rect 171414 218376 171470 218385
rect 170772 218340 170824 218346
rect 171414 218311 171470 218320
rect 170772 218282 170824 218288
rect 170784 217138 170812 218282
rect 171428 218210 171456 218311
rect 171416 218204 171468 218210
rect 171416 218146 171468 218152
rect 171612 217274 171640 218470
rect 171980 218385 172008 219098
rect 171966 218376 172022 218385
rect 171966 218311 172022 218320
rect 164942 217110 165016 217138
rect 165770 217110 165844 217138
rect 166598 217110 166672 217138
rect 167426 217110 167500 217138
rect 168254 217110 168328 217138
rect 169082 217110 169156 217138
rect 169910 217110 169984 217138
rect 170738 217110 170812 217138
rect 171566 217246 171640 217274
rect 164942 216988 164970 217110
rect 165770 216988 165798 217110
rect 166598 216988 166626 217110
rect 167426 216988 167454 217110
rect 168254 216988 168282 217110
rect 169082 216988 169110 217110
rect 169910 216988 169938 217110
rect 170738 216988 170766 217110
rect 171566 216988 171594 217246
rect 172440 217138 172468 219370
rect 173256 218068 173308 218074
rect 173256 218010 173308 218016
rect 173268 217138 173296 218010
rect 174096 217138 174124 222090
rect 174280 217938 174308 224926
rect 174912 224936 174964 224942
rect 174912 224878 174964 224884
rect 175292 224926 175596 224954
rect 175752 231662 175950 231690
rect 174268 217932 174320 217938
rect 174268 217874 174320 217880
rect 174924 217138 174952 224878
rect 175292 220810 175320 224926
rect 175752 222630 175780 231662
rect 175924 229764 175976 229770
rect 175924 229706 175976 229712
rect 176384 229764 176436 229770
rect 176384 229706 176436 229712
rect 175936 229226 175964 229706
rect 175924 229220 175976 229226
rect 175924 229162 175976 229168
rect 176106 228848 176162 228857
rect 176106 228783 176108 228792
rect 176160 228783 176162 228792
rect 176108 228754 176160 228760
rect 175924 227520 175976 227526
rect 175924 227462 175976 227468
rect 175936 227361 175964 227462
rect 175922 227352 175978 227361
rect 175922 227287 175978 227296
rect 176396 224954 176424 229706
rect 176396 224926 176516 224954
rect 175740 222624 175792 222630
rect 175740 222566 175792 222572
rect 175924 222556 175976 222562
rect 175924 222498 175976 222504
rect 175108 220782 175320 220810
rect 175108 220658 175136 220782
rect 175096 220652 175148 220658
rect 175096 220594 175148 220600
rect 175280 220652 175332 220658
rect 175280 220594 175332 220600
rect 175292 218346 175320 220594
rect 175936 219162 175964 222498
rect 176290 221912 176346 221921
rect 176290 221847 176292 221856
rect 176344 221847 176346 221856
rect 176292 221818 176344 221824
rect 175924 219156 175976 219162
rect 175924 219098 175976 219104
rect 175280 218340 175332 218346
rect 175280 218282 175332 218288
rect 175740 218340 175792 218346
rect 175740 218282 175792 218288
rect 175752 217138 175780 218282
rect 176488 217274 176516 224926
rect 176580 223394 176608 231676
rect 177224 227633 177252 231676
rect 177408 231662 177882 231690
rect 177210 227624 177266 227633
rect 177210 227559 177266 227568
rect 176750 227352 176806 227361
rect 176750 227287 176752 227296
rect 176804 227287 176806 227296
rect 176752 227258 176804 227264
rect 176580 223366 176700 223394
rect 176672 223310 176700 223366
rect 176660 223304 176712 223310
rect 176660 223246 176712 223252
rect 177408 221921 177436 231662
rect 178512 224806 178540 231676
rect 179156 230926 179184 231676
rect 179144 230920 179196 230926
rect 179144 230862 179196 230868
rect 179800 229090 179828 231676
rect 180444 229226 180472 231676
rect 180432 229220 180484 229226
rect 180432 229162 180484 229168
rect 179788 229084 179840 229090
rect 179788 229026 179840 229032
rect 180064 229084 180116 229090
rect 180064 229026 180116 229032
rect 179326 224904 179382 224913
rect 179326 224839 179382 224848
rect 178500 224800 178552 224806
rect 178500 224742 178552 224748
rect 178776 224800 178828 224806
rect 178776 224742 178828 224748
rect 177394 221912 177450 221921
rect 177394 221847 177450 221856
rect 177210 220824 177266 220833
rect 177210 220759 177212 220768
rect 177264 220759 177266 220768
rect 177396 220788 177448 220794
rect 177212 220730 177264 220736
rect 177396 220730 177448 220736
rect 176488 217246 176562 217274
rect 172394 217110 172468 217138
rect 173222 217110 173296 217138
rect 174050 217110 174124 217138
rect 174878 217110 174952 217138
rect 175706 217110 175780 217138
rect 172394 216988 172422 217110
rect 173222 216988 173250 217110
rect 174050 216988 174078 217110
rect 174878 216988 174906 217110
rect 175706 216988 175734 217110
rect 176534 216988 176562 217246
rect 177408 217138 177436 220730
rect 178788 219434 178816 224742
rect 178960 222012 179012 222018
rect 178960 221954 179012 221960
rect 178972 221746 179000 221954
rect 178960 221740 179012 221746
rect 178960 221682 179012 221688
rect 178224 219428 178276 219434
rect 178224 219370 178276 219376
rect 178776 219428 178828 219434
rect 178776 219370 178828 219376
rect 178236 217138 178264 219370
rect 179052 219020 179104 219026
rect 179052 218962 179104 218968
rect 179064 217138 179092 218962
rect 179340 218210 179368 224839
rect 180076 219298 180104 229026
rect 181088 223990 181116 231676
rect 181732 229094 181760 231676
rect 181732 229066 181852 229094
rect 181444 228676 181496 228682
rect 181444 228618 181496 228624
rect 181628 228676 181680 228682
rect 181628 228618 181680 228624
rect 181456 228138 181484 228618
rect 181260 228132 181312 228138
rect 181260 228074 181312 228080
rect 181444 228132 181496 228138
rect 181444 228074 181496 228080
rect 181272 228018 181300 228074
rect 181640 228018 181668 228618
rect 181272 227990 181668 228018
rect 181536 227588 181588 227594
rect 181536 227530 181588 227536
rect 181352 224936 181404 224942
rect 181352 224878 181404 224884
rect 181364 224534 181392 224878
rect 181352 224528 181404 224534
rect 181352 224470 181404 224476
rect 181076 223984 181128 223990
rect 181076 223926 181128 223932
rect 181548 220946 181576 227530
rect 181824 223446 181852 229066
rect 182376 227730 182404 231676
rect 182652 231662 183034 231690
rect 183678 231662 183876 231690
rect 182364 227724 182416 227730
rect 182364 227666 182416 227672
rect 181996 224936 182048 224942
rect 181994 224904 181996 224913
rect 182048 224904 182050 224913
rect 181994 224839 182050 224848
rect 181812 223440 181864 223446
rect 181812 223382 181864 223388
rect 182652 221882 182680 231662
rect 183376 229220 183428 229226
rect 183376 229162 183428 229168
rect 183388 224954 183416 229162
rect 183204 224926 183416 224954
rect 182640 221876 182692 221882
rect 182640 221818 182692 221824
rect 182824 221876 182876 221882
rect 182824 221818 182876 221824
rect 182836 221762 182864 221818
rect 181088 220918 181576 220946
rect 182100 221734 182864 221762
rect 180064 219292 180116 219298
rect 180064 219234 180116 219240
rect 180522 218784 180578 218793
rect 180522 218719 180524 218728
rect 180576 218719 180578 218728
rect 180708 218748 180760 218754
rect 180524 218690 180576 218696
rect 180708 218690 180760 218696
rect 179328 218204 179380 218210
rect 179328 218146 179380 218152
rect 179880 218204 179932 218210
rect 179880 218146 179932 218152
rect 179892 217138 179920 218146
rect 180720 217138 180748 218690
rect 181088 218618 181116 220918
rect 181260 220788 181312 220794
rect 181260 220730 181312 220736
rect 181444 220788 181496 220794
rect 181444 220730 181496 220736
rect 181272 219858 181300 220730
rect 181456 219978 181484 220730
rect 181444 219972 181496 219978
rect 181444 219914 181496 219920
rect 181628 219972 181680 219978
rect 181628 219914 181680 219920
rect 181640 219858 181668 219914
rect 181272 219830 181668 219858
rect 182100 219434 182128 221734
rect 181628 219428 181680 219434
rect 181628 219370 181680 219376
rect 182088 219428 182140 219434
rect 182088 219370 182140 219376
rect 182272 219428 182324 219434
rect 182272 219370 182324 219376
rect 181444 219292 181496 219298
rect 181444 219234 181496 219240
rect 181076 218612 181128 218618
rect 181076 218554 181128 218560
rect 181456 218346 181484 219234
rect 181444 218340 181496 218346
rect 181444 218282 181496 218288
rect 181640 217274 181668 219370
rect 182284 218793 182312 219370
rect 182270 218784 182326 218793
rect 182270 218719 182326 218728
rect 182364 218612 182416 218618
rect 182364 218554 182416 218560
rect 177362 217110 177436 217138
rect 178190 217110 178264 217138
rect 179018 217110 179092 217138
rect 179846 217110 179920 217138
rect 180674 217110 180748 217138
rect 181502 217246 181668 217274
rect 177362 216988 177390 217110
rect 178190 216988 178218 217110
rect 179018 216988 179046 217110
rect 179846 216988 179874 217110
rect 180674 216988 180702 217110
rect 181502 216988 181530 217246
rect 182376 217138 182404 218554
rect 183204 217274 183232 224926
rect 183848 223854 183876 231662
rect 184308 225758 184336 231676
rect 184952 228954 184980 231676
rect 185136 231662 185610 231690
rect 185872 231662 186254 231690
rect 186608 231662 186898 231690
rect 184940 228948 184992 228954
rect 184940 228890 184992 228896
rect 184296 225752 184348 225758
rect 184296 225694 184348 225700
rect 184480 225752 184532 225758
rect 184480 225694 184532 225700
rect 183836 223848 183888 223854
rect 183836 223790 183888 223796
rect 184020 223440 184072 223446
rect 184020 223382 184072 223388
rect 182330 217110 182404 217138
rect 183158 217246 183232 217274
rect 182330 216988 182358 217110
rect 183158 216988 183186 217246
rect 184032 217138 184060 223382
rect 184492 219434 184520 225694
rect 184848 223848 184900 223854
rect 184848 223790 184900 223796
rect 184480 219428 184532 219434
rect 184480 219370 184532 219376
rect 184860 217138 184888 223790
rect 185136 220833 185164 231662
rect 185584 230172 185636 230178
rect 185584 230114 185636 230120
rect 185398 229936 185454 229945
rect 185398 229871 185454 229880
rect 185412 229770 185440 229871
rect 185596 229770 185624 230114
rect 185400 229764 185452 229770
rect 185400 229706 185452 229712
rect 185584 229764 185636 229770
rect 185584 229706 185636 229712
rect 185872 229094 185900 231662
rect 186044 230172 186096 230178
rect 186044 230114 186096 230120
rect 186056 229945 186084 230114
rect 186042 229936 186098 229945
rect 186042 229871 186098 229880
rect 185584 229084 185636 229090
rect 185872 229066 185992 229094
rect 185584 229026 185636 229032
rect 185400 228948 185452 228954
rect 185400 228890 185452 228896
rect 185412 228682 185440 228890
rect 185596 228682 185624 229026
rect 185400 228676 185452 228682
rect 185400 228618 185452 228624
rect 185584 228676 185636 228682
rect 185584 228618 185636 228624
rect 185400 227724 185452 227730
rect 185400 227666 185452 227672
rect 185412 226914 185440 227666
rect 185584 227452 185636 227458
rect 185584 227394 185636 227400
rect 185596 226914 185624 227394
rect 185400 226908 185452 226914
rect 185400 226850 185452 226856
rect 185584 226908 185636 226914
rect 185584 226850 185636 226856
rect 185412 224998 185808 225026
rect 185412 224806 185440 224998
rect 185780 224942 185808 224998
rect 185768 224936 185820 224942
rect 185768 224878 185820 224884
rect 185400 224800 185452 224806
rect 185400 224742 185452 224748
rect 185964 223718 185992 229066
rect 186136 227588 186188 227594
rect 186136 227530 186188 227536
rect 185952 223712 186004 223718
rect 185952 223654 186004 223660
rect 185122 220824 185178 220833
rect 185122 220759 185178 220768
rect 185950 220824 186006 220833
rect 185950 220759 186006 220768
rect 185676 219428 185728 219434
rect 185676 219370 185728 219376
rect 185688 217138 185716 219370
rect 185964 218754 185992 220759
rect 186148 219434 186176 227530
rect 186608 223582 186636 231662
rect 187528 226778 187556 231676
rect 188172 230790 188200 231676
rect 188356 231662 188830 231690
rect 189092 231662 189474 231690
rect 188160 230784 188212 230790
rect 188160 230726 188212 230732
rect 187516 226772 187568 226778
rect 187516 226714 187568 226720
rect 186964 223848 187016 223854
rect 186964 223790 187016 223796
rect 186596 223576 186648 223582
rect 186596 223518 186648 223524
rect 186136 219428 186188 219434
rect 186136 219370 186188 219376
rect 186274 219428 186326 219434
rect 186274 219370 186326 219376
rect 186286 219314 186314 219370
rect 186240 219286 186314 219314
rect 185952 218748 186004 218754
rect 185952 218690 186004 218696
rect 186240 218074 186268 219286
rect 186504 218748 186556 218754
rect 186504 218690 186556 218696
rect 186228 218068 186280 218074
rect 186228 218010 186280 218016
rect 186516 217138 186544 218690
rect 186976 218482 187004 223790
rect 187332 223576 187384 223582
rect 187332 223518 187384 223524
rect 186964 218476 187016 218482
rect 186964 218418 187016 218424
rect 187344 217274 187372 223518
rect 188356 219434 188384 231662
rect 189092 229094 189120 231662
rect 189092 229066 189212 229094
rect 188896 223304 188948 223310
rect 188896 223246 188948 223252
rect 187988 219406 188384 219434
rect 187988 217462 188016 219406
rect 188908 218074 188936 223246
rect 188160 218068 188212 218074
rect 188160 218010 188212 218016
rect 188896 218068 188948 218074
rect 188896 218010 188948 218016
rect 187976 217456 188028 217462
rect 187976 217398 188028 217404
rect 183986 217110 184060 217138
rect 184814 217110 184888 217138
rect 185642 217110 185716 217138
rect 186470 217110 186544 217138
rect 187298 217246 187372 217274
rect 183986 216988 184014 217110
rect 184814 216988 184842 217110
rect 185642 216988 185670 217110
rect 186470 216988 186498 217110
rect 187298 216988 187326 217246
rect 188172 217138 188200 218010
rect 188896 217932 188948 217938
rect 188896 217874 188948 217880
rect 188126 217110 188200 217138
rect 188908 217138 188936 217874
rect 189184 217598 189212 229066
rect 189724 229084 189776 229090
rect 189724 229026 189776 229032
rect 189736 218618 189764 229026
rect 190104 228954 190132 231676
rect 190656 231662 190762 231690
rect 191024 231662 191406 231690
rect 190656 229094 190684 231662
rect 190472 229066 190684 229094
rect 190092 228948 190144 228954
rect 190092 228890 190144 228896
rect 190000 226772 190052 226778
rect 190000 226714 190052 226720
rect 190012 219298 190040 226714
rect 190472 220946 190500 229066
rect 191024 222222 191052 231662
rect 192036 222766 192064 231676
rect 192680 227730 192708 231676
rect 192852 229084 192904 229090
rect 192852 229026 192904 229032
rect 192864 228002 192892 229026
rect 193034 228984 193090 228993
rect 193034 228919 193090 228928
rect 192852 227996 192904 228002
rect 192852 227938 192904 227944
rect 192668 227724 192720 227730
rect 192668 227666 192720 227672
rect 192024 222760 192076 222766
rect 192024 222702 192076 222708
rect 191012 222216 191064 222222
rect 191012 222158 191064 222164
rect 191472 222148 191524 222154
rect 191472 222090 191524 222096
rect 190380 220918 190500 220946
rect 190380 220794 190408 220918
rect 190550 220824 190606 220833
rect 190368 220788 190420 220794
rect 190550 220759 190552 220768
rect 190368 220730 190420 220736
rect 190604 220759 190606 220768
rect 190552 220730 190604 220736
rect 190000 219292 190052 219298
rect 190000 219234 190052 219240
rect 190644 219292 190696 219298
rect 190644 219234 190696 219240
rect 189724 218612 189776 218618
rect 189724 218554 189776 218560
rect 189816 218476 189868 218482
rect 189816 218418 189868 218424
rect 189172 217592 189224 217598
rect 189172 217534 189224 217540
rect 189828 217138 189856 218418
rect 190656 217138 190684 219234
rect 191484 217274 191512 222090
rect 192852 218612 192904 218618
rect 192852 218554 192904 218560
rect 192024 218340 192076 218346
rect 192024 218282 192076 218288
rect 192036 218074 192064 218282
rect 192024 218068 192076 218074
rect 192024 218010 192076 218016
rect 192300 218068 192352 218074
rect 192300 218010 192352 218016
rect 188908 217110 188982 217138
rect 188126 216988 188154 217110
rect 188954 216988 188982 217110
rect 189782 217110 189856 217138
rect 190610 217110 190684 217138
rect 191438 217246 191512 217274
rect 189782 216988 189810 217110
rect 190610 216988 190638 217110
rect 191438 216988 191466 217246
rect 192312 217138 192340 218010
rect 192864 217274 192892 218554
rect 193048 218074 193076 228919
rect 193324 221338 193352 231676
rect 193968 226302 193996 231676
rect 194416 230648 194468 230654
rect 194416 230590 194468 230596
rect 194428 230314 194456 230590
rect 194416 230308 194468 230314
rect 194416 230250 194468 230256
rect 193956 226296 194008 226302
rect 193956 226238 194008 226244
rect 194140 226296 194192 226302
rect 194140 226238 194192 226244
rect 194152 225894 194180 226238
rect 193588 225888 193640 225894
rect 193588 225830 193640 225836
rect 194140 225888 194192 225894
rect 194140 225830 194192 225836
rect 193312 221332 193364 221338
rect 193312 221274 193364 221280
rect 193600 218346 193628 225830
rect 194612 224126 194640 231676
rect 194876 230308 194928 230314
rect 194876 230250 194928 230256
rect 194888 229770 194916 230250
rect 195060 230036 195112 230042
rect 195060 229978 195112 229984
rect 195072 229770 195100 229978
rect 194876 229764 194928 229770
rect 194876 229706 194928 229712
rect 195060 229764 195112 229770
rect 195060 229706 195112 229712
rect 195256 229090 195284 231676
rect 195900 231062 195928 231676
rect 196176 231662 196558 231690
rect 196912 231662 197202 231690
rect 197372 231662 197846 231690
rect 198016 231662 198490 231690
rect 195888 231056 195940 231062
rect 195888 230998 195940 231004
rect 195428 230308 195480 230314
rect 195428 230250 195480 230256
rect 195612 230308 195664 230314
rect 195612 230250 195664 230256
rect 195440 230042 195468 230250
rect 195428 230036 195480 230042
rect 195428 229978 195480 229984
rect 195244 229084 195296 229090
rect 195244 229026 195296 229032
rect 195426 228984 195482 228993
rect 195244 228948 195296 228954
rect 195426 228919 195428 228928
rect 195244 228890 195296 228896
rect 195480 228919 195482 228928
rect 195428 228890 195480 228896
rect 195256 228138 195284 228890
rect 195244 228132 195296 228138
rect 195244 228074 195296 228080
rect 195244 224936 195296 224942
rect 195244 224878 195296 224884
rect 195428 224936 195480 224942
rect 195428 224878 195480 224884
rect 195256 224126 195284 224878
rect 194600 224120 194652 224126
rect 194600 224062 194652 224068
rect 195244 224120 195296 224126
rect 195244 224062 195296 224068
rect 195440 223718 195468 224878
rect 195428 223712 195480 223718
rect 195428 223654 195480 223660
rect 194508 222760 194560 222766
rect 194508 222702 194560 222708
rect 193588 218340 193640 218346
rect 193588 218282 193640 218288
rect 194520 218074 194548 222702
rect 195624 219434 195652 230250
rect 196176 225486 196204 231662
rect 196912 230654 196940 231662
rect 196900 230648 196952 230654
rect 196900 230590 196952 230596
rect 197372 226642 197400 231662
rect 198016 229094 198044 231662
rect 197648 229066 198044 229094
rect 197360 226636 197412 226642
rect 197360 226578 197412 226584
rect 196164 225480 196216 225486
rect 196164 225422 196216 225428
rect 196348 225480 196400 225486
rect 196348 225422 196400 225428
rect 195888 223712 195940 223718
rect 195888 223654 195940 223660
rect 195256 219406 195652 219434
rect 194874 219328 194930 219337
rect 194874 219263 194876 219272
rect 194928 219263 194930 219272
rect 195060 219292 195112 219298
rect 194876 219234 194928 219240
rect 195060 219234 195112 219240
rect 195072 218754 195100 219234
rect 195060 218748 195112 218754
rect 195060 218690 195112 218696
rect 195256 218482 195284 219406
rect 195612 218748 195664 218754
rect 195612 218690 195664 218696
rect 195244 218476 195296 218482
rect 195244 218418 195296 218424
rect 193036 218068 193088 218074
rect 193036 218010 193088 218016
rect 193956 218068 194008 218074
rect 193956 218010 194008 218016
rect 194508 218068 194560 218074
rect 194508 218010 194560 218016
rect 194784 218068 194836 218074
rect 194784 218010 194836 218016
rect 192864 217246 193122 217274
rect 192266 217110 192340 217138
rect 192266 216988 192294 217110
rect 193094 216988 193122 217246
rect 193968 217138 193996 218010
rect 194796 217138 194824 218010
rect 195624 217138 195652 218690
rect 195900 218074 195928 223654
rect 196360 219434 196388 225422
rect 197176 222624 197228 222630
rect 197176 222566 197228 222572
rect 196268 219406 196388 219434
rect 196268 219026 196296 219406
rect 196256 219020 196308 219026
rect 196256 218962 196308 218968
rect 196440 218340 196492 218346
rect 196440 218282 196492 218288
rect 195888 218068 195940 218074
rect 195888 218010 195940 218016
rect 196452 217138 196480 218282
rect 197188 217274 197216 222566
rect 197648 219842 197676 229066
rect 198004 225888 198056 225894
rect 198004 225830 198056 225836
rect 197636 219836 197688 219842
rect 197636 219778 197688 219784
rect 197820 219836 197872 219842
rect 197820 219778 197872 219784
rect 197832 219337 197860 219778
rect 197818 219328 197874 219337
rect 197818 219263 197874 219272
rect 198016 218754 198044 225830
rect 199120 225350 199148 231676
rect 199108 225344 199160 225350
rect 199108 225286 199160 225292
rect 199764 222358 199792 231676
rect 200408 229094 200436 231676
rect 201052 230518 201080 231676
rect 201040 230512 201092 230518
rect 201040 230454 201092 230460
rect 200408 229066 200528 229094
rect 200120 228540 200172 228546
rect 200120 228482 200172 228488
rect 200304 228540 200356 228546
rect 200304 228482 200356 228488
rect 200132 227746 200160 228482
rect 200316 228002 200344 228482
rect 200304 227996 200356 228002
rect 200304 227938 200356 227944
rect 200500 227866 200528 229066
rect 201408 229084 201460 229090
rect 201408 229026 201460 229032
rect 200488 227860 200540 227866
rect 200488 227802 200540 227808
rect 200672 227860 200724 227866
rect 200672 227802 200724 227808
rect 200684 227746 200712 227802
rect 200132 227718 200712 227746
rect 200040 227594 200252 227610
rect 200040 227588 200264 227594
rect 200040 227582 200212 227588
rect 199752 222352 199804 222358
rect 199752 222294 199804 222300
rect 198004 218748 198056 218754
rect 198004 218690 198056 218696
rect 198280 218748 198332 218754
rect 198280 218690 198332 218696
rect 198096 218612 198148 218618
rect 198096 218554 198148 218560
rect 197188 217246 197262 217274
rect 193922 217110 193996 217138
rect 194750 217110 194824 217138
rect 195578 217110 195652 217138
rect 196406 217110 196480 217138
rect 193922 216988 193950 217110
rect 194750 216988 194778 217110
rect 195578 216988 195606 217110
rect 196406 216988 196434 217110
rect 197234 216988 197262 217246
rect 198108 217138 198136 218554
rect 198292 218482 198320 218690
rect 198280 218476 198332 218482
rect 198280 218418 198332 218424
rect 199752 218476 199804 218482
rect 199752 218418 199804 218424
rect 198924 218068 198976 218074
rect 198924 218010 198976 218016
rect 198936 217138 198964 218010
rect 199764 217138 199792 218418
rect 200040 218074 200068 227582
rect 200212 227530 200264 227536
rect 201224 223984 201276 223990
rect 201224 223926 201276 223932
rect 201236 219434 201264 223926
rect 201236 219406 201356 219434
rect 200212 219020 200264 219026
rect 200212 218962 200264 218968
rect 200224 218618 200252 218962
rect 200212 218612 200264 218618
rect 200212 218554 200264 218560
rect 200396 218612 200448 218618
rect 200396 218554 200448 218560
rect 200408 218210 200436 218554
rect 200396 218204 200448 218210
rect 200396 218146 200448 218152
rect 200580 218204 200632 218210
rect 200580 218146 200632 218152
rect 200028 218068 200080 218074
rect 200028 218010 200080 218016
rect 200592 217138 200620 218146
rect 201328 217274 201356 219406
rect 201420 218226 201448 229026
rect 201696 225078 201724 231676
rect 202340 229770 202368 231676
rect 202328 229764 202380 229770
rect 202328 229706 202380 229712
rect 202984 226506 203012 231676
rect 203168 231662 203642 231690
rect 202972 226500 203024 226506
rect 202972 226442 203024 226448
rect 201684 225072 201736 225078
rect 201684 225014 201736 225020
rect 202236 225072 202288 225078
rect 202236 225014 202288 225020
rect 201420 218210 201540 218226
rect 201420 218204 201552 218210
rect 201420 218198 201500 218204
rect 201500 218146 201552 218152
rect 202248 217274 202276 225014
rect 203168 219706 203196 231662
rect 203524 226636 203576 226642
rect 203524 226578 203576 226584
rect 203156 219700 203208 219706
rect 203156 219642 203208 219648
rect 203536 218890 203564 226578
rect 203708 226160 203760 226166
rect 203708 226102 203760 226108
rect 203892 226160 203944 226166
rect 203892 226102 203944 226108
rect 203720 225350 203748 226102
rect 203904 225894 203932 226102
rect 203892 225888 203944 225894
rect 203892 225830 203944 225836
rect 203708 225344 203760 225350
rect 203708 225286 203760 225292
rect 204272 225214 204300 231676
rect 204640 231662 204930 231690
rect 204640 229094 204668 231662
rect 204904 230308 204956 230314
rect 204904 230250 204956 230256
rect 204916 229770 204944 230250
rect 204904 229764 204956 229770
rect 204904 229706 204956 229712
rect 204548 229066 204668 229094
rect 204260 225208 204312 225214
rect 204260 225150 204312 225156
rect 204548 224806 204576 229066
rect 205560 228274 205588 231676
rect 205928 231662 206218 231690
rect 206480 231662 206862 231690
rect 205548 228268 205600 228274
rect 205548 228210 205600 228216
rect 205732 228268 205784 228274
rect 205732 228210 205784 228216
rect 205744 228154 205772 228210
rect 205468 228126 205772 228154
rect 204904 225888 204956 225894
rect 204904 225830 204956 225836
rect 204916 225486 204944 225830
rect 204904 225480 204956 225486
rect 204904 225422 204956 225428
rect 204536 224800 204588 224806
rect 204536 224742 204588 224748
rect 204720 224800 204772 224806
rect 204720 224742 204772 224748
rect 204732 224126 204760 224742
rect 204720 224120 204772 224126
rect 204720 224062 204772 224068
rect 204904 224120 204956 224126
rect 204904 224062 204956 224068
rect 204916 223718 204944 224062
rect 204904 223712 204956 223718
rect 204904 223654 204956 223660
rect 204168 221332 204220 221338
rect 204168 221274 204220 221280
rect 203892 219700 203944 219706
rect 203892 219642 203944 219648
rect 203524 218884 203576 218890
rect 203524 218826 203576 218832
rect 203064 218068 203116 218074
rect 203064 218010 203116 218016
rect 201328 217246 201402 217274
rect 198062 217110 198136 217138
rect 198890 217110 198964 217138
rect 199718 217110 199792 217138
rect 200546 217110 200620 217138
rect 198062 216988 198090 217110
rect 198890 216988 198918 217110
rect 199718 216988 199746 217110
rect 200546 216988 200574 217110
rect 201374 216988 201402 217246
rect 202202 217246 202276 217274
rect 202202 216988 202230 217246
rect 203076 217138 203104 218010
rect 203904 217274 203932 219642
rect 204180 219026 204208 221274
rect 204168 219020 204220 219026
rect 204168 218962 204220 218968
rect 204720 219020 204772 219026
rect 204720 218962 204772 218968
rect 204732 218482 204760 218962
rect 204720 218476 204772 218482
rect 204720 218418 204772 218424
rect 204720 218204 204772 218210
rect 204720 218146 204772 218152
rect 203030 217110 203104 217138
rect 203858 217246 203932 217274
rect 203030 216988 203058 217110
rect 203858 216988 203886 217246
rect 204732 217138 204760 218146
rect 205468 217274 205496 228126
rect 205928 221610 205956 231662
rect 206284 230308 206336 230314
rect 206284 230250 206336 230256
rect 205916 221604 205968 221610
rect 205916 221546 205968 221552
rect 206296 218074 206324 230250
rect 206480 221066 206508 231662
rect 207492 222494 207520 231676
rect 208136 227050 208164 231676
rect 208596 231662 208794 231690
rect 208124 227044 208176 227050
rect 208124 226986 208176 226992
rect 208124 225480 208176 225486
rect 208124 225422 208176 225428
rect 207480 222488 207532 222494
rect 207480 222430 207532 222436
rect 207664 222488 207716 222494
rect 207664 222430 207716 222436
rect 206468 221060 206520 221066
rect 206468 221002 206520 221008
rect 206468 218884 206520 218890
rect 206468 218826 206520 218832
rect 206284 218068 206336 218074
rect 206284 218010 206336 218016
rect 206480 217274 206508 218826
rect 207676 218210 207704 222430
rect 207848 219156 207900 219162
rect 207848 219098 207900 219104
rect 207860 218210 207888 219098
rect 207664 218204 207716 218210
rect 207664 218146 207716 218152
rect 207848 218204 207900 218210
rect 207848 218146 207900 218152
rect 208136 218074 208164 225422
rect 208400 221604 208452 221610
rect 208400 221546 208452 221552
rect 208412 219434 208440 221546
rect 208596 220522 208624 231662
rect 209424 225350 209452 231676
rect 210068 229498 210096 231676
rect 210252 231662 210726 231690
rect 210056 229492 210108 229498
rect 210056 229434 210108 229440
rect 210252 227866 210280 231662
rect 210424 227996 210476 228002
rect 210424 227938 210476 227944
rect 210240 227860 210292 227866
rect 210240 227802 210292 227808
rect 209412 225344 209464 225350
rect 209412 225286 209464 225292
rect 209688 225344 209740 225350
rect 209688 225286 209740 225292
rect 208584 220516 208636 220522
rect 208584 220458 208636 220464
rect 208320 219406 208440 219434
rect 207204 218068 207256 218074
rect 207204 218010 207256 218016
rect 208124 218068 208176 218074
rect 208124 218010 208176 218016
rect 205468 217246 205542 217274
rect 204686 217110 204760 217138
rect 204686 216988 204714 217110
rect 205514 216988 205542 217246
rect 206342 217246 206508 217274
rect 206342 216988 206370 217246
rect 207216 217138 207244 218010
rect 208320 217274 208348 219406
rect 209700 219162 209728 225286
rect 210436 220674 210464 227938
rect 210344 220646 210464 220674
rect 208860 219156 208912 219162
rect 208860 219098 208912 219104
rect 209688 219156 209740 219162
rect 209688 219098 209740 219104
rect 207170 217110 207244 217138
rect 207998 217246 208348 217274
rect 207170 216988 207198 217110
rect 207998 216988 208026 217246
rect 208872 217138 208900 219098
rect 210344 218618 210372 220646
rect 210516 220516 210568 220522
rect 210516 220458 210568 220464
rect 210332 218612 210384 218618
rect 210332 218554 210384 218560
rect 209688 218340 209740 218346
rect 209688 218282 209740 218288
rect 209700 217138 209728 218282
rect 210528 217274 210556 220458
rect 211356 219570 211384 231676
rect 212000 222902 212028 231676
rect 212552 231662 212658 231690
rect 212172 226500 212224 226506
rect 212172 226442 212224 226448
rect 211988 222896 212040 222902
rect 211988 222838 212040 222844
rect 211804 222352 211856 222358
rect 211804 222294 211856 222300
rect 211344 219564 211396 219570
rect 211344 219506 211396 219512
rect 211344 219156 211396 219162
rect 211344 219098 211396 219104
rect 208826 217110 208900 217138
rect 209654 217110 209728 217138
rect 210482 217246 210556 217274
rect 208826 216988 208854 217110
rect 209654 216988 209682 217110
rect 210482 216988 210510 217246
rect 211356 217138 211384 219098
rect 211816 218210 211844 222294
rect 211804 218204 211856 218210
rect 211804 218146 211856 218152
rect 212184 217274 212212 226442
rect 212552 225758 212580 231662
rect 213092 230444 213144 230450
rect 213092 230386 213144 230392
rect 213104 229094 213132 230386
rect 213288 229094 213316 231676
rect 213946 231662 214144 231690
rect 213104 229066 213224 229094
rect 213288 229066 213408 229094
rect 212540 225752 212592 225758
rect 212540 225694 212592 225700
rect 213000 218612 213052 218618
rect 213000 218554 213052 218560
rect 211310 217110 211384 217138
rect 212138 217246 212212 217274
rect 211310 216988 211338 217110
rect 212138 216988 212166 217246
rect 213012 217138 213040 218554
rect 213196 218346 213224 229066
rect 213380 227186 213408 229066
rect 213368 227180 213420 227186
rect 213368 227122 213420 227128
rect 213828 226908 213880 226914
rect 213828 226850 213880 226856
rect 213184 218340 213236 218346
rect 213184 218282 213236 218288
rect 213840 217274 213868 226850
rect 214116 220386 214144 231662
rect 214380 227724 214432 227730
rect 214380 227666 214432 227672
rect 214392 227186 214420 227666
rect 214380 227180 214432 227186
rect 214380 227122 214432 227128
rect 214576 226114 214604 231676
rect 215220 230042 215248 231676
rect 215208 230036 215260 230042
rect 215208 229978 215260 229984
rect 215864 228410 215892 231676
rect 216232 231662 216522 231690
rect 215852 228404 215904 228410
rect 215852 228346 215904 228352
rect 214748 227724 214800 227730
rect 214748 227666 214800 227672
rect 214760 226506 214788 227666
rect 214748 226500 214800 226506
rect 214748 226442 214800 226448
rect 214392 226086 214604 226114
rect 214748 226160 214800 226166
rect 214748 226102 214800 226108
rect 214392 226030 214420 226086
rect 214380 226024 214432 226030
rect 214380 225966 214432 225972
rect 214760 225350 214788 226102
rect 215208 225752 215260 225758
rect 215208 225694 215260 225700
rect 214748 225344 214800 225350
rect 214748 225286 214800 225292
rect 214104 220380 214156 220386
rect 214104 220322 214156 220328
rect 214288 220380 214340 220386
rect 214288 220322 214340 220328
rect 214104 220108 214156 220114
rect 214104 220050 214156 220056
rect 214116 219570 214144 220050
rect 214300 219978 214328 220322
rect 214288 219972 214340 219978
rect 214288 219914 214340 219920
rect 214104 219564 214156 219570
rect 214104 219506 214156 219512
rect 215220 218074 215248 225694
rect 216232 223174 216260 231662
rect 216404 228404 216456 228410
rect 216404 228346 216456 228352
rect 216220 223168 216272 223174
rect 216220 223110 216272 223116
rect 215944 222896 215996 222902
rect 215944 222838 215996 222844
rect 215956 219434 215984 222838
rect 216416 219434 216444 228346
rect 217152 225622 217180 231676
rect 217140 225616 217192 225622
rect 217140 225558 217192 225564
rect 217796 223854 217824 231676
rect 218440 227050 218468 231676
rect 218716 231662 219098 231690
rect 219544 231662 219742 231690
rect 218428 227044 218480 227050
rect 218428 226986 218480 226992
rect 217784 223848 217836 223854
rect 217784 223790 217836 223796
rect 217140 219836 217192 219842
rect 217140 219778 217192 219784
rect 215944 219428 215996 219434
rect 215944 219370 215996 219376
rect 216140 219406 216444 219434
rect 216140 218074 216168 219406
rect 216312 218476 216364 218482
rect 216312 218418 216364 218424
rect 214656 218068 214708 218074
rect 214656 218010 214708 218016
rect 215208 218068 215260 218074
rect 215208 218010 215260 218016
rect 215484 218068 215536 218074
rect 215484 218010 215536 218016
rect 216128 218068 216180 218074
rect 216128 218010 216180 218016
rect 212966 217110 213040 217138
rect 213794 217246 213868 217274
rect 212966 216988 212994 217110
rect 213794 216988 213822 217246
rect 214668 217138 214696 218010
rect 215496 217138 215524 218010
rect 216324 217138 216352 218418
rect 217152 217274 217180 219778
rect 218716 219570 218744 231662
rect 219348 226636 219400 226642
rect 219348 226578 219400 226584
rect 218704 219564 218756 219570
rect 218704 219506 218756 219512
rect 219360 219162 219388 226578
rect 219544 223038 219572 231662
rect 220372 229634 220400 231676
rect 220360 229628 220412 229634
rect 220360 229570 220412 229576
rect 220452 229492 220504 229498
rect 220452 229434 220504 229440
rect 219900 227452 219952 227458
rect 219900 227394 219952 227400
rect 220084 227452 220136 227458
rect 220084 227394 220136 227400
rect 219912 227066 219940 227394
rect 220096 227186 220124 227394
rect 220084 227180 220136 227186
rect 220084 227122 220136 227128
rect 220268 227180 220320 227186
rect 220268 227122 220320 227128
rect 220280 227066 220308 227122
rect 219912 227038 220308 227066
rect 220268 226908 220320 226914
rect 220268 226850 220320 226856
rect 220280 226642 220308 226850
rect 220268 226636 220320 226642
rect 220268 226578 220320 226584
rect 220084 226024 220136 226030
rect 220084 225966 220136 225972
rect 220268 226024 220320 226030
rect 220268 225966 220320 225972
rect 220096 225758 220124 225966
rect 220084 225752 220136 225758
rect 220084 225694 220136 225700
rect 220280 225622 220308 225966
rect 220268 225616 220320 225622
rect 220268 225558 220320 225564
rect 220464 224954 220492 229434
rect 221016 228546 221044 231676
rect 221292 231662 221674 231690
rect 221004 228540 221056 228546
rect 221004 228482 221056 228488
rect 220096 224926 220492 224954
rect 219532 223032 219584 223038
rect 219532 222974 219584 222980
rect 219808 221060 219860 221066
rect 219808 221002 219860 221008
rect 219624 219428 219676 219434
rect 219624 219370 219676 219376
rect 217324 219156 217376 219162
rect 217324 219098 217376 219104
rect 218796 219156 218848 219162
rect 218796 219098 218848 219104
rect 219348 219156 219400 219162
rect 219348 219098 219400 219104
rect 217336 218482 217364 219098
rect 217324 218476 217376 218482
rect 217324 218418 217376 218424
rect 217968 218204 218020 218210
rect 217968 218146 218020 218152
rect 214622 217110 214696 217138
rect 215450 217110 215524 217138
rect 216278 217110 216352 217138
rect 217106 217246 217180 217274
rect 214622 216988 214650 217110
rect 215450 216988 215478 217110
rect 216278 216988 216306 217110
rect 217106 216988 217134 217246
rect 217980 217138 218008 218146
rect 218808 217138 218836 219098
rect 219636 217138 219664 219370
rect 219820 218482 219848 221002
rect 219808 218476 219860 218482
rect 219808 218418 219860 218424
rect 220096 218074 220124 224926
rect 221292 221202 221320 231662
rect 221832 226500 221884 226506
rect 221832 226442 221884 226448
rect 221280 221196 221332 221202
rect 221280 221138 221332 221144
rect 220452 219700 220504 219706
rect 220452 219642 220504 219648
rect 220084 218068 220136 218074
rect 220084 218010 220136 218016
rect 220464 217274 220492 219642
rect 221844 218074 221872 226442
rect 222016 225616 222068 225622
rect 222016 225558 222068 225564
rect 221280 218068 221332 218074
rect 221280 218010 221332 218016
rect 221832 218068 221884 218074
rect 221832 218010 221884 218016
rect 217934 217110 218008 217138
rect 218762 217110 218836 217138
rect 219590 217110 219664 217138
rect 220418 217246 220492 217274
rect 217934 216988 217962 217110
rect 218762 216988 218790 217110
rect 219590 216988 219618 217110
rect 220418 216988 220446 217246
rect 221292 217138 221320 218010
rect 222028 217274 222056 225558
rect 222304 220930 222332 231676
rect 222948 226642 222976 231676
rect 223592 227186 223620 231676
rect 223776 231662 224250 231690
rect 224512 231662 224894 231690
rect 223580 227180 223632 227186
rect 223580 227122 223632 227128
rect 222936 226636 222988 226642
rect 222936 226578 222988 226584
rect 223776 224754 223804 231662
rect 224512 224954 224540 231662
rect 225524 229906 225552 231676
rect 225512 229900 225564 229906
rect 225512 229842 225564 229848
rect 225696 229900 225748 229906
rect 225696 229842 225748 229848
rect 224776 228404 224828 228410
rect 224776 228346 224828 228352
rect 223684 224726 223804 224754
rect 223868 224926 224540 224954
rect 222752 221196 222804 221202
rect 222752 221138 222804 221144
rect 222292 220924 222344 220930
rect 222292 220866 222344 220872
rect 222764 218210 222792 221138
rect 223684 220250 223712 224726
rect 223868 224670 223896 224926
rect 224224 224800 224276 224806
rect 224224 224742 224276 224748
rect 223856 224664 223908 224670
rect 223856 224606 223908 224612
rect 224236 224398 224264 224742
rect 224408 224664 224460 224670
rect 224408 224606 224460 224612
rect 224592 224664 224644 224670
rect 224592 224606 224644 224612
rect 224420 224398 224448 224606
rect 224224 224392 224276 224398
rect 224224 224334 224276 224340
rect 224408 224392 224460 224398
rect 224408 224334 224460 224340
rect 224224 220652 224276 220658
rect 224224 220594 224276 220600
rect 223672 220244 223724 220250
rect 223672 220186 223724 220192
rect 224236 219570 224264 220594
rect 224408 220380 224460 220386
rect 224408 220322 224460 220328
rect 224420 219706 224448 220322
rect 224408 219700 224460 219706
rect 224408 219642 224460 219648
rect 224224 219564 224276 219570
rect 224224 219506 224276 219512
rect 224040 219292 224092 219298
rect 224040 219234 224092 219240
rect 224052 218482 224080 219234
rect 224224 219156 224276 219162
rect 224224 219098 224276 219104
rect 224236 218618 224264 219098
rect 224224 218612 224276 218618
rect 224224 218554 224276 218560
rect 224040 218476 224092 218482
rect 224040 218418 224092 218424
rect 222752 218204 222804 218210
rect 222752 218146 222804 218152
rect 222936 218204 222988 218210
rect 222936 218146 222988 218152
rect 222028 217246 222102 217274
rect 221246 217110 221320 217138
rect 221246 216988 221274 217110
rect 222074 216988 222102 217246
rect 222948 217138 222976 218146
rect 224604 218074 224632 224606
rect 223764 218068 223816 218074
rect 223764 218010 223816 218016
rect 224592 218068 224644 218074
rect 224592 218010 224644 218016
rect 223776 217138 223804 218010
rect 224788 217274 224816 228346
rect 225708 219434 225736 229842
rect 226168 228682 226196 231676
rect 226536 231662 226826 231690
rect 226156 228676 226208 228682
rect 226156 228618 226208 228624
rect 226340 228676 226392 228682
rect 226340 228618 226392 228624
rect 226352 228562 226380 228618
rect 225616 219406 225736 219434
rect 226168 228534 226380 228562
rect 225616 218210 225644 219406
rect 225972 218612 226024 218618
rect 225972 218554 226024 218560
rect 225604 218204 225656 218210
rect 225604 218146 225656 218152
rect 225420 218068 225472 218074
rect 225420 218010 225472 218016
rect 222902 217110 222976 217138
rect 223730 217110 223804 217138
rect 224558 217246 224816 217274
rect 222902 216988 222930 217110
rect 223730 216988 223758 217110
rect 224558 216988 224586 217246
rect 225432 217138 225460 218010
rect 225984 217274 226012 218554
rect 226168 218074 226196 228534
rect 226536 221474 226564 231662
rect 227456 224262 227484 231676
rect 227444 224256 227496 224262
rect 227444 224198 227496 224204
rect 228100 222358 228128 231676
rect 228744 227322 228772 231676
rect 229296 231662 229402 231690
rect 228732 227316 228784 227322
rect 228732 227258 228784 227264
rect 228916 227044 228968 227050
rect 228916 226986 228968 226992
rect 228928 226506 228956 226986
rect 228916 226500 228968 226506
rect 228916 226442 228968 226448
rect 228732 223848 228784 223854
rect 228732 223790 228784 223796
rect 228088 222352 228140 222358
rect 228088 222294 228140 222300
rect 226524 221468 226576 221474
rect 226524 221410 226576 221416
rect 227904 221468 227956 221474
rect 227904 221410 227956 221416
rect 227076 219700 227128 219706
rect 227076 219642 227128 219648
rect 226156 218068 226208 218074
rect 226156 218010 226208 218016
rect 227088 217274 227116 219642
rect 227916 217274 227944 221410
rect 228744 217274 228772 223790
rect 229296 219570 229324 231662
rect 230032 224806 230060 231676
rect 230480 230036 230532 230042
rect 230480 229978 230532 229984
rect 230020 224800 230072 224806
rect 230020 224742 230072 224748
rect 230492 224210 230520 229978
rect 230676 229362 230704 231676
rect 230664 229356 230716 229362
rect 230664 229298 230716 229304
rect 231320 228818 231348 231676
rect 231872 231662 231978 231690
rect 232240 231662 232622 231690
rect 231308 228812 231360 228818
rect 231308 228754 231360 228760
rect 231032 226636 231084 226642
rect 231032 226578 231084 226584
rect 230400 224182 230520 224210
rect 230204 223032 230256 223038
rect 230204 222974 230256 222980
rect 229284 219564 229336 219570
rect 229284 219506 229336 219512
rect 230216 219434 230244 222974
rect 230216 219406 230336 219434
rect 229560 218068 229612 218074
rect 229560 218010 229612 218016
rect 225984 217246 226242 217274
rect 225386 217110 225460 217138
rect 225386 216988 225414 217110
rect 226214 216988 226242 217246
rect 227042 217246 227116 217274
rect 227870 217246 227944 217274
rect 228698 217246 228772 217274
rect 227042 216988 227070 217246
rect 227870 216988 227898 217246
rect 228698 216988 228726 217246
rect 229572 217138 229600 218010
rect 230308 217274 230336 219406
rect 230400 218090 230428 224182
rect 231044 218482 231072 226578
rect 231492 225888 231544 225894
rect 231492 225830 231544 225836
rect 231504 225350 231532 225830
rect 231492 225344 231544 225350
rect 231492 225286 231544 225292
rect 231676 224256 231728 224262
rect 231676 224198 231728 224204
rect 231032 218476 231084 218482
rect 231032 218418 231084 218424
rect 230400 218074 230520 218090
rect 231688 218074 231716 224198
rect 231872 222018 231900 231662
rect 231860 222012 231912 222018
rect 231860 221954 231912 221960
rect 232240 221746 232268 231662
rect 233252 229094 233280 231676
rect 233252 229066 233372 229094
rect 232964 224800 233016 224806
rect 232964 224742 233016 224748
rect 232976 224398 233004 224742
rect 232964 224392 233016 224398
rect 232964 224334 233016 224340
rect 233148 224392 233200 224398
rect 233148 224334 233200 224340
rect 232228 221740 232280 221746
rect 232228 221682 232280 221688
rect 232872 218340 232924 218346
rect 232872 218282 232924 218288
rect 230400 218068 230532 218074
rect 230400 218062 230480 218068
rect 230480 218010 230532 218016
rect 231216 218068 231268 218074
rect 231216 218010 231268 218016
rect 231676 218068 231728 218074
rect 231676 218010 231728 218016
rect 232044 218068 232096 218074
rect 232044 218010 232096 218016
rect 230308 217246 230382 217274
rect 229526 217110 229600 217138
rect 229526 216988 229554 217110
rect 230354 216988 230382 217246
rect 231228 217138 231256 218010
rect 232056 217138 232084 218010
rect 232884 217274 232912 218282
rect 233160 218074 233188 224334
rect 233344 222902 233372 229066
rect 233896 226778 233924 231676
rect 234172 231662 234554 231690
rect 233884 226772 233936 226778
rect 233884 226714 233936 226720
rect 233332 222896 233384 222902
rect 233332 222838 233384 222844
rect 233700 222012 233752 222018
rect 233700 221954 233752 221960
rect 233148 218068 233200 218074
rect 233148 218010 233200 218016
rect 233712 217274 233740 221954
rect 234172 220250 234200 231662
rect 235184 224534 235212 231676
rect 235828 230178 235856 231676
rect 235816 230172 235868 230178
rect 235816 230114 235868 230120
rect 235816 227316 235868 227322
rect 235816 227258 235868 227264
rect 235172 224528 235224 224534
rect 235172 224470 235224 224476
rect 234528 222896 234580 222902
rect 234528 222838 234580 222844
rect 234160 220244 234212 220250
rect 234160 220186 234212 220192
rect 234540 217274 234568 222838
rect 235828 218074 235856 227258
rect 236472 225350 236500 231676
rect 236656 231662 237130 231690
rect 236460 225344 236512 225350
rect 236460 225286 236512 225292
rect 236656 220794 236684 231662
rect 237288 225752 237340 225758
rect 237288 225694 237340 225700
rect 236644 220788 236696 220794
rect 236644 220730 236696 220736
rect 237012 220244 237064 220250
rect 237012 220186 237064 220192
rect 235356 218068 235408 218074
rect 235356 218010 235408 218016
rect 235816 218068 235868 218074
rect 235816 218010 235868 218016
rect 236184 218068 236236 218074
rect 236184 218010 236236 218016
rect 231182 217110 231256 217138
rect 232010 217110 232084 217138
rect 232838 217246 232912 217274
rect 233666 217246 233740 217274
rect 234494 217246 234568 217274
rect 231182 216988 231210 217110
rect 232010 216988 232038 217110
rect 232838 216988 232866 217246
rect 233666 216988 233694 217246
rect 234494 216988 234522 217246
rect 235368 217138 235396 218010
rect 236196 217138 236224 218010
rect 237024 217274 237052 220186
rect 237300 218074 237328 225694
rect 237760 224806 237788 231676
rect 238404 228002 238432 231676
rect 238576 228812 238628 228818
rect 238576 228754 238628 228760
rect 238392 227996 238444 228002
rect 238392 227938 238444 227944
rect 237748 224800 237800 224806
rect 237748 224742 237800 224748
rect 238024 223712 238076 223718
rect 238024 223654 238076 223660
rect 237840 219292 237892 219298
rect 237840 219234 237892 219240
rect 237288 218068 237340 218074
rect 237288 218010 237340 218016
rect 235322 217110 235396 217138
rect 236150 217110 236224 217138
rect 236978 217246 237052 217274
rect 235322 216988 235350 217110
rect 236150 216988 236178 217110
rect 236978 216988 237006 217246
rect 237852 217138 237880 219234
rect 238036 218482 238064 223654
rect 238024 218476 238076 218482
rect 238024 218418 238076 218424
rect 238588 217274 238616 228754
rect 239048 228138 239076 231676
rect 239036 228132 239088 228138
rect 239036 228074 239088 228080
rect 239692 223446 239720 231676
rect 240152 231662 240350 231690
rect 239680 223440 239732 223446
rect 239680 223382 239732 223388
rect 240152 221882 240180 231662
rect 240324 230172 240376 230178
rect 240324 230114 240376 230120
rect 240336 225758 240364 230114
rect 240980 229226 241008 231676
rect 240968 229220 241020 229226
rect 240968 229162 241020 229168
rect 241624 227458 241652 231676
rect 241612 227452 241664 227458
rect 241612 227394 241664 227400
rect 240324 225752 240376 225758
rect 240324 225694 240376 225700
rect 241152 225344 241204 225350
rect 241152 225286 241204 225292
rect 240140 221876 240192 221882
rect 240140 221818 240192 221824
rect 239220 221740 239272 221746
rect 239220 221682 239272 221688
rect 239232 219298 239260 221682
rect 239220 219292 239272 219298
rect 239220 219234 239272 219240
rect 239496 219292 239548 219298
rect 239496 219234 239548 219240
rect 238588 217246 238662 217274
rect 237806 217110 237880 217138
rect 237806 216988 237834 217110
rect 238634 216988 238662 217246
rect 239508 217138 239536 219234
rect 240324 218068 240376 218074
rect 240324 218010 240376 218016
rect 240336 217138 240364 218010
rect 241164 217274 241192 225286
rect 242268 223582 242296 231676
rect 242716 225208 242768 225214
rect 242716 225150 242768 225156
rect 242256 223576 242308 223582
rect 242256 223518 242308 223524
rect 241336 223168 241388 223174
rect 241336 223110 241388 223116
rect 241348 218074 241376 223110
rect 242728 220946 242756 225150
rect 242912 224942 242940 231676
rect 243280 231662 243570 231690
rect 243280 226642 243308 231662
rect 243452 226704 243504 226710
rect 243452 226646 243504 226652
rect 243268 226636 243320 226642
rect 243268 226578 243320 226584
rect 242900 224936 242952 224942
rect 242900 224878 242952 224884
rect 242728 220918 242848 220946
rect 242624 220788 242676 220794
rect 242624 220730 242676 220736
rect 242636 219434 242664 220730
rect 242636 219406 242756 219434
rect 241980 218204 242032 218210
rect 241980 218146 242032 218152
rect 241336 218068 241388 218074
rect 241336 218010 241388 218016
rect 239462 217110 239536 217138
rect 240290 217110 240364 217138
rect 241118 217246 241192 217274
rect 239462 216988 239490 217110
rect 240290 216988 240318 217110
rect 241118 216988 241146 217246
rect 241992 217138 242020 218146
rect 242728 217274 242756 219406
rect 242820 218226 242848 220918
rect 243464 218754 243492 226646
rect 244200 226302 244228 231676
rect 244476 231662 244858 231690
rect 245120 231662 245502 231690
rect 244476 229094 244504 231662
rect 244384 229066 244504 229094
rect 244188 226296 244240 226302
rect 244188 226238 244240 226244
rect 244096 223440 244148 223446
rect 244096 223382 244148 223388
rect 243452 218748 243504 218754
rect 243452 218690 243504 218696
rect 242820 218210 242940 218226
rect 242820 218204 242952 218210
rect 242820 218198 242900 218204
rect 242900 218146 242952 218152
rect 244108 218074 244136 223382
rect 244384 220266 244412 229066
rect 245120 223310 245148 231662
rect 246132 229770 246160 231676
rect 246120 229764 246172 229770
rect 246120 229706 246172 229712
rect 246488 229764 246540 229770
rect 246488 229706 246540 229712
rect 246304 228132 246356 228138
rect 246304 228074 246356 228080
rect 245292 224800 245344 224806
rect 245292 224742 245344 224748
rect 245108 223304 245160 223310
rect 245108 223246 245160 223252
rect 244292 220238 244412 220266
rect 244292 220114 244320 220238
rect 244280 220108 244332 220114
rect 244280 220050 244332 220056
rect 244464 220108 244516 220114
rect 244464 220050 244516 220056
rect 243636 218068 243688 218074
rect 243636 218010 243688 218016
rect 244096 218068 244148 218074
rect 244096 218010 244148 218016
rect 242728 217246 242802 217274
rect 241946 217110 242020 217138
rect 241946 216988 241974 217110
rect 242774 216988 242802 217246
rect 243648 217138 243676 218010
rect 244476 217274 244504 220050
rect 245304 217274 245332 224742
rect 246316 219026 246344 228074
rect 246500 220794 246528 229706
rect 246776 228954 246804 231676
rect 246764 228948 246816 228954
rect 246764 228890 246816 228896
rect 246856 223304 246908 223310
rect 246856 223246 246908 223252
rect 246488 220788 246540 220794
rect 246488 220730 246540 220736
rect 246304 219020 246356 219026
rect 246304 218962 246356 218968
rect 246120 218340 246172 218346
rect 246120 218282 246172 218288
rect 243602 217110 243676 217138
rect 244430 217246 244504 217274
rect 245258 217246 245332 217274
rect 243602 216988 243630 217110
rect 244430 216988 244458 217246
rect 245258 216988 245286 217246
rect 246132 217138 246160 218282
rect 246868 217274 246896 223246
rect 247420 222766 247448 231676
rect 247604 231662 248078 231690
rect 247408 222760 247460 222766
rect 247408 222702 247460 222708
rect 247604 222154 247632 231662
rect 248236 228948 248288 228954
rect 248236 228890 248288 228896
rect 247592 222148 247644 222154
rect 247592 222090 247644 222096
rect 248248 218074 248276 228890
rect 248708 226710 248736 231676
rect 248696 226704 248748 226710
rect 248696 226646 248748 226652
rect 249352 225894 249380 231676
rect 249616 226772 249668 226778
rect 249616 226714 249668 226720
rect 249340 225888 249392 225894
rect 249340 225830 249392 225836
rect 249432 218204 249484 218210
rect 249432 218146 249484 218152
rect 247776 218068 247828 218074
rect 247776 218010 247828 218016
rect 248236 218068 248288 218074
rect 248236 218010 248288 218016
rect 248604 218068 248656 218074
rect 248604 218010 248656 218016
rect 246868 217246 246942 217274
rect 246086 217110 246160 217138
rect 246086 216988 246114 217110
rect 246914 216988 246942 217246
rect 247788 217138 247816 218010
rect 248616 217138 248644 218010
rect 249444 217138 249472 218146
rect 249628 218074 249656 226714
rect 249996 222630 250024 231676
rect 250640 224126 250668 231676
rect 251284 229634 251312 231676
rect 251272 229628 251324 229634
rect 251272 229570 251324 229576
rect 251732 229628 251784 229634
rect 251732 229570 251784 229576
rect 251088 224528 251140 224534
rect 251088 224470 251140 224476
rect 250628 224120 250680 224126
rect 250628 224062 250680 224068
rect 250904 223576 250956 223582
rect 250904 223518 250956 223524
rect 249984 222624 250036 222630
rect 249984 222566 250036 222572
rect 250916 218074 250944 223518
rect 249616 218068 249668 218074
rect 249616 218010 249668 218016
rect 250260 218068 250312 218074
rect 250260 218010 250312 218016
rect 250904 218068 250956 218074
rect 250904 218010 250956 218016
rect 250272 217138 250300 218010
rect 251100 217274 251128 224470
rect 251744 218210 251772 229570
rect 251928 227594 251956 231676
rect 252572 229090 252600 231676
rect 252756 231662 253230 231690
rect 252560 229084 252612 229090
rect 252560 229026 252612 229032
rect 251916 227588 251968 227594
rect 251916 227530 251968 227536
rect 252468 225888 252520 225894
rect 252468 225830 252520 225836
rect 251732 218204 251784 218210
rect 251732 218146 251784 218152
rect 252480 218074 252508 225830
rect 252756 221338 252784 231662
rect 253860 228138 253888 231676
rect 253848 228132 253900 228138
rect 253848 228074 253900 228080
rect 254504 225078 254532 231676
rect 254780 231662 255162 231690
rect 254492 225072 254544 225078
rect 254492 225014 254544 225020
rect 252744 221332 252796 221338
rect 252744 221274 252796 221280
rect 253848 220856 253900 220862
rect 253848 220798 253900 220804
rect 253572 220652 253624 220658
rect 253572 220594 253624 220600
rect 253388 219156 253440 219162
rect 253388 219098 253440 219104
rect 252744 219020 252796 219026
rect 252744 218962 252796 218968
rect 251916 218068 251968 218074
rect 251916 218010 251968 218016
rect 252468 218068 252520 218074
rect 252468 218010 252520 218016
rect 247742 217110 247816 217138
rect 248570 217110 248644 217138
rect 249398 217110 249472 217138
rect 250226 217110 250300 217138
rect 251054 217246 251128 217274
rect 247742 216988 247770 217110
rect 248570 216988 248598 217110
rect 249398 216988 249426 217110
rect 250226 216988 250254 217110
rect 251054 216988 251082 217246
rect 251928 217138 251956 218010
rect 252756 217138 252784 218962
rect 253204 218748 253256 218754
rect 253204 218690 253256 218696
rect 253216 218346 253244 218690
rect 253400 218346 253428 219098
rect 253204 218340 253256 218346
rect 253204 218282 253256 218288
rect 253388 218340 253440 218346
rect 253388 218282 253440 218288
rect 253584 217274 253612 220594
rect 253860 218890 253888 220798
rect 254780 219978 254808 231662
rect 255228 229084 255280 229090
rect 255228 229026 255280 229032
rect 255044 225752 255096 225758
rect 255044 225694 255096 225700
rect 254768 219972 254820 219978
rect 254768 219914 254820 219920
rect 253848 218884 253900 218890
rect 253848 218826 253900 218832
rect 255056 218074 255084 225694
rect 254400 218068 254452 218074
rect 254400 218010 254452 218016
rect 255044 218068 255096 218074
rect 255044 218010 255096 218016
rect 251882 217110 251956 217138
rect 252710 217110 252784 217138
rect 253538 217246 253612 217274
rect 251882 216988 251910 217110
rect 252710 216988 252738 217110
rect 253538 216988 253566 217246
rect 254412 217138 254440 218010
rect 255240 217274 255268 229026
rect 255792 223990 255820 231676
rect 256436 230314 256464 231676
rect 256424 230308 256476 230314
rect 256424 230250 256476 230256
rect 256608 230308 256660 230314
rect 256608 230250 256660 230256
rect 255780 223984 255832 223990
rect 255780 223926 255832 223932
rect 256620 219434 256648 230250
rect 257080 228274 257108 231676
rect 257448 231662 257738 231690
rect 257068 228268 257120 228274
rect 257068 228210 257120 228216
rect 257448 225486 257476 231662
rect 257620 228268 257672 228274
rect 257620 228210 257672 228216
rect 257436 225480 257488 225486
rect 257436 225422 257488 225428
rect 257632 219434 257660 228210
rect 257804 227452 257856 227458
rect 257804 227394 257856 227400
rect 257816 219434 257844 227394
rect 258368 222494 258396 231676
rect 258644 231662 259026 231690
rect 258356 222488 258408 222494
rect 258356 222430 258408 222436
rect 258080 222148 258132 222154
rect 258080 222090 258132 222096
rect 256528 219406 256648 219434
rect 257540 219406 257660 219434
rect 257724 219406 257844 219434
rect 256528 218074 256556 219406
rect 257540 218074 257568 219406
rect 256056 218068 256108 218074
rect 256056 218010 256108 218016
rect 256516 218068 256568 218074
rect 256516 218010 256568 218016
rect 256884 218068 256936 218074
rect 256884 218010 256936 218016
rect 257528 218068 257580 218074
rect 257528 218010 257580 218016
rect 254366 217110 254440 217138
rect 255194 217246 255268 217274
rect 254366 216988 254394 217110
rect 255194 216988 255222 217246
rect 256068 217138 256096 218010
rect 256896 217138 256924 218010
rect 257724 217274 257752 219406
rect 258092 218346 258120 222090
rect 258644 220862 258672 231662
rect 259276 227588 259328 227594
rect 259276 227530 259328 227536
rect 258632 220856 258684 220862
rect 258632 220798 258684 220804
rect 259092 218884 259144 218890
rect 259092 218826 259144 218832
rect 258080 218340 258132 218346
rect 258080 218282 258132 218288
rect 258540 218068 258592 218074
rect 258540 218010 258592 218016
rect 256022 217110 256096 217138
rect 256850 217110 256924 217138
rect 257678 217246 257752 217274
rect 256022 216988 256050 217110
rect 256850 216988 256878 217110
rect 257678 216988 257706 217246
rect 258552 217138 258580 218010
rect 259104 217274 259132 218826
rect 259288 218074 259316 227530
rect 259656 226166 259684 231676
rect 259932 231662 260314 231690
rect 260852 231662 260958 231690
rect 259644 226160 259696 226166
rect 259644 226102 259696 226108
rect 259932 220522 259960 231662
rect 260852 221610 260880 231662
rect 261588 230450 261616 231676
rect 261576 230444 261628 230450
rect 261576 230386 261628 230392
rect 262232 227730 262260 231676
rect 262220 227724 262272 227730
rect 262220 227666 262272 227672
rect 262876 227186 262904 231676
rect 263060 231662 263534 231690
rect 263704 231662 264178 231690
rect 262864 227180 262916 227186
rect 262864 227122 262916 227128
rect 261852 226160 261904 226166
rect 261852 226102 261904 226108
rect 260840 221604 260892 221610
rect 260840 221546 260892 221552
rect 261024 221604 261076 221610
rect 261024 221546 261076 221552
rect 260196 220788 260248 220794
rect 260196 220730 260248 220736
rect 259920 220516 259972 220522
rect 259920 220458 259972 220464
rect 259276 218068 259328 218074
rect 259276 218010 259328 218016
rect 260208 217274 260236 220730
rect 261036 217274 261064 221546
rect 261208 219428 261260 219434
rect 261208 219370 261260 219376
rect 261220 219162 261248 219370
rect 261208 219156 261260 219162
rect 261208 219098 261260 219104
rect 261864 217274 261892 226102
rect 263060 221066 263088 231662
rect 263508 227180 263560 227186
rect 263508 227122 263560 227128
rect 263324 221876 263376 221882
rect 263324 221818 263376 221824
rect 263048 221060 263100 221066
rect 263048 221002 263100 221008
rect 263336 219434 263364 221818
rect 263520 219434 263548 227122
rect 263704 222154 263732 231662
rect 264808 228546 264836 231676
rect 265176 231662 265466 231690
rect 264796 228540 264848 228546
rect 264796 228482 264848 228488
rect 264244 226568 264296 226574
rect 264244 226510 264296 226516
rect 263692 222148 263744 222154
rect 263692 222090 263744 222096
rect 262680 219428 262732 219434
rect 263336 219406 263456 219434
rect 263520 219428 263652 219434
rect 263520 219406 263600 219428
rect 262680 219370 262732 219376
rect 259104 217246 259362 217274
rect 258506 217110 258580 217138
rect 258506 216988 258534 217110
rect 259334 216988 259362 217246
rect 260162 217246 260236 217274
rect 260990 217246 261064 217274
rect 261818 217246 261892 217274
rect 260162 216988 260190 217246
rect 260990 216988 261018 217246
rect 261818 216988 261846 217246
rect 262692 217138 262720 219370
rect 263428 217274 263456 219406
rect 263600 219370 263652 219376
rect 264256 219162 264284 226510
rect 264796 222760 264848 222766
rect 264796 222702 264848 222708
rect 264244 219156 264296 219162
rect 264244 219098 264296 219104
rect 264428 219156 264480 219162
rect 264428 219098 264480 219104
rect 264440 218618 264468 219098
rect 264428 218612 264480 218618
rect 264428 218554 264480 218560
rect 264808 218074 264836 222702
rect 265176 219842 265204 231662
rect 266096 226030 266124 231676
rect 266084 226024 266136 226030
rect 266084 225966 266136 225972
rect 266176 224936 266228 224942
rect 266176 224878 266228 224884
rect 265164 219836 265216 219842
rect 265164 219778 265216 219784
rect 265992 218612 266044 218618
rect 265992 218554 266044 218560
rect 264336 218068 264388 218074
rect 264336 218010 264388 218016
rect 264796 218068 264848 218074
rect 264796 218010 264848 218016
rect 265164 218068 265216 218074
rect 265164 218010 265216 218016
rect 263428 217246 263502 217274
rect 262646 217110 262720 217138
rect 262646 216988 262674 217110
rect 263474 216988 263502 217246
rect 264348 217138 264376 218010
rect 265176 217138 265204 218010
rect 266004 217138 266032 218554
rect 266188 218074 266216 224878
rect 266740 223718 266768 231676
rect 267384 226914 267412 231676
rect 267936 231662 268042 231690
rect 268304 231662 268686 231690
rect 267372 226908 267424 226914
rect 267372 226850 267424 226856
rect 267004 226024 267056 226030
rect 267004 225966 267056 225972
rect 266728 223712 266780 223718
rect 266728 223654 266780 223660
rect 266820 221332 266872 221338
rect 266820 221274 266872 221280
rect 266176 218068 266228 218074
rect 266176 218010 266228 218016
rect 266832 217274 266860 221274
rect 267016 219162 267044 225966
rect 267648 220516 267700 220522
rect 267648 220458 267700 220464
rect 267004 219156 267056 219162
rect 267004 219098 267056 219104
rect 267660 217274 267688 220458
rect 267936 220386 267964 231662
rect 268304 221202 268332 231662
rect 268936 228132 268988 228138
rect 268936 228074 268988 228080
rect 268292 221196 268344 221202
rect 268292 221138 268344 221144
rect 267924 220380 267976 220386
rect 267924 220322 267976 220328
rect 268948 218074 268976 228074
rect 269316 226574 269344 231676
rect 269304 226568 269356 226574
rect 269304 226510 269356 226516
rect 269960 225622 269988 231676
rect 269948 225616 270000 225622
rect 269948 225558 270000 225564
rect 270224 225616 270276 225622
rect 270224 225558 270276 225564
rect 270040 222148 270092 222154
rect 270040 222090 270092 222096
rect 268476 218068 268528 218074
rect 268476 218010 268528 218016
rect 268936 218068 268988 218074
rect 268936 218010 268988 218016
rect 269304 218068 269356 218074
rect 269304 218010 269356 218016
rect 264302 217110 264376 217138
rect 265130 217110 265204 217138
rect 265958 217110 266032 217138
rect 266786 217246 266860 217274
rect 267614 217246 267688 217274
rect 264302 216988 264330 217110
rect 265130 216988 265158 217110
rect 265958 216988 265986 217110
rect 266786 216988 266814 217246
rect 267614 216988 267642 217246
rect 268488 217138 268516 218010
rect 269316 217138 269344 218010
rect 270052 217274 270080 222090
rect 270236 218074 270264 225558
rect 270604 224670 270632 231676
rect 271248 227050 271276 231676
rect 271892 229906 271920 231676
rect 271880 229900 271932 229906
rect 271880 229842 271932 229848
rect 272536 228682 272564 231676
rect 272720 231662 273194 231690
rect 272524 228676 272576 228682
rect 272524 228618 272576 228624
rect 272524 228540 272576 228546
rect 272524 228482 272576 228488
rect 271236 227044 271288 227050
rect 271236 226986 271288 226992
rect 271788 227044 271840 227050
rect 271788 226986 271840 226992
rect 271144 226432 271196 226438
rect 271144 226374 271196 226380
rect 270592 224664 270644 224670
rect 270592 224606 270644 224612
rect 271156 218482 271184 226374
rect 271144 218476 271196 218482
rect 271144 218418 271196 218424
rect 270224 218068 270276 218074
rect 270224 218010 270276 218016
rect 270960 218068 271012 218074
rect 270960 218010 271012 218016
rect 270052 217246 270126 217274
rect 268442 217110 268516 217138
rect 269270 217110 269344 217138
rect 268442 216988 268470 217110
rect 269270 216988 269298 217110
rect 270098 216988 270126 217246
rect 270972 217138 271000 218010
rect 271800 217274 271828 226986
rect 272340 219428 272392 219434
rect 272340 219370 272392 219376
rect 270926 217110 271000 217138
rect 271754 217246 271828 217274
rect 272352 217274 272380 219370
rect 272536 218074 272564 228482
rect 272720 219706 272748 231662
rect 273824 228410 273852 231676
rect 273812 228404 273864 228410
rect 273812 228346 273864 228352
rect 274468 226030 274496 231676
rect 275112 229094 275140 231676
rect 274928 229066 275140 229094
rect 275480 231662 275770 231690
rect 276124 231662 276414 231690
rect 274456 226024 274508 226030
rect 274456 225966 274508 225972
rect 274272 224664 274324 224670
rect 274272 224606 274324 224612
rect 273444 220380 273496 220386
rect 273444 220322 273496 220328
rect 272708 219700 272760 219706
rect 272708 219642 272760 219648
rect 272892 219292 272944 219298
rect 272892 219234 272944 219240
rect 272708 219156 272760 219162
rect 272708 219098 272760 219104
rect 272720 218618 272748 219098
rect 272904 218618 272932 219234
rect 272708 218612 272760 218618
rect 272708 218554 272760 218560
rect 272892 218612 272944 218618
rect 272892 218554 272944 218560
rect 272524 218068 272576 218074
rect 272524 218010 272576 218016
rect 273456 217274 273484 220322
rect 274284 217274 274312 224606
rect 274928 223854 274956 229066
rect 275100 224120 275152 224126
rect 275100 224062 275152 224068
rect 274916 223848 274968 223854
rect 274916 223790 274968 223796
rect 275112 217274 275140 224062
rect 275480 223038 275508 231662
rect 275652 229900 275704 229906
rect 275652 229842 275704 229848
rect 275664 229094 275692 229842
rect 275664 229066 275876 229094
rect 275468 223032 275520 223038
rect 275468 222974 275520 222980
rect 272352 217246 272610 217274
rect 270926 216988 270954 217110
rect 271754 216988 271782 217246
rect 272582 216988 272610 217246
rect 273410 217246 273484 217274
rect 274238 217246 274312 217274
rect 275066 217246 275140 217274
rect 275848 217274 275876 229066
rect 276124 221474 276152 231662
rect 277044 230042 277072 231676
rect 277032 230036 277084 230042
rect 277032 229978 277084 229984
rect 277216 230036 277268 230042
rect 277216 229978 277268 229984
rect 277032 227724 277084 227730
rect 277032 227666 277084 227672
rect 276112 221468 276164 221474
rect 276112 221410 276164 221416
rect 277044 219434 277072 227666
rect 277228 227186 277256 229978
rect 277216 227180 277268 227186
rect 277216 227122 277268 227128
rect 277688 224398 277716 231676
rect 277964 231662 278346 231690
rect 277676 224392 277728 224398
rect 277676 224334 277728 224340
rect 277964 222018 277992 231662
rect 278412 226024 278464 226030
rect 278412 225966 278464 225972
rect 277952 222012 278004 222018
rect 277952 221954 278004 221960
rect 277044 219406 277256 219434
rect 277228 218074 277256 219406
rect 276756 218068 276808 218074
rect 276756 218010 276808 218016
rect 277216 218068 277268 218074
rect 277216 218010 277268 218016
rect 277584 218068 277636 218074
rect 277584 218010 277636 218016
rect 275848 217246 275922 217274
rect 273410 216988 273438 217246
rect 274238 216988 274266 217246
rect 275066 216988 275094 217246
rect 275894 216988 275922 217246
rect 276768 217138 276796 218010
rect 277596 217138 277624 218010
rect 278424 217274 278452 225966
rect 278976 224262 279004 231676
rect 279620 226438 279648 231676
rect 280264 227322 280292 231676
rect 280448 231662 280922 231690
rect 280252 227316 280304 227322
rect 280252 227258 280304 227264
rect 279608 226432 279660 226438
rect 279608 226374 279660 226380
rect 278964 224256 279016 224262
rect 278964 224198 279016 224204
rect 279424 223916 279476 223922
rect 279424 223858 279476 223864
rect 278596 223032 278648 223038
rect 278596 222974 278648 222980
rect 278608 218074 278636 222974
rect 279436 218618 279464 223858
rect 280068 222012 280120 222018
rect 280068 221954 280120 221960
rect 279424 218612 279476 218618
rect 279424 218554 279476 218560
rect 279240 218476 279292 218482
rect 279240 218418 279292 218424
rect 278596 218068 278648 218074
rect 278596 218010 278648 218016
rect 276722 217110 276796 217138
rect 277550 217110 277624 217138
rect 278378 217246 278452 217274
rect 276722 216988 276750 217110
rect 277550 216988 277578 217110
rect 278378 216988 278406 217246
rect 279252 217138 279280 218418
rect 280080 217274 280108 221954
rect 280448 220250 280476 231662
rect 281356 227180 281408 227186
rect 281356 227122 281408 227128
rect 280436 220244 280488 220250
rect 280436 220186 280488 220192
rect 281368 219434 281396 227122
rect 281552 222902 281580 231676
rect 282196 230178 282224 231676
rect 282184 230172 282236 230178
rect 282184 230114 282236 230120
rect 282644 230172 282696 230178
rect 282644 230114 282696 230120
rect 282656 225622 282684 230114
rect 282840 228818 282868 231676
rect 282828 228812 282880 228818
rect 282828 228754 282880 228760
rect 282644 225616 282696 225622
rect 282644 225558 282696 225564
rect 283484 223174 283512 231676
rect 283668 231662 284142 231690
rect 283472 223168 283524 223174
rect 283472 223110 283524 223116
rect 281540 222896 281592 222902
rect 281540 222838 281592 222844
rect 282460 222896 282512 222902
rect 282460 222838 282512 222844
rect 281368 219406 281488 219434
rect 281460 218074 281488 219406
rect 282184 219020 282236 219026
rect 282184 218962 282236 218968
rect 282196 218482 282224 218962
rect 282184 218476 282236 218482
rect 282184 218418 282236 218424
rect 282472 218074 282500 222838
rect 283668 221746 283696 231662
rect 284116 225616 284168 225622
rect 284116 225558 284168 225564
rect 283656 221740 283708 221746
rect 283656 221682 283708 221688
rect 282644 220924 282696 220930
rect 282644 220866 282696 220872
rect 280896 218068 280948 218074
rect 280896 218010 280948 218016
rect 281448 218068 281500 218074
rect 281448 218010 281500 218016
rect 281724 218068 281776 218074
rect 281724 218010 281776 218016
rect 282460 218068 282512 218074
rect 282460 218010 282512 218016
rect 279206 217110 279280 217138
rect 280034 217246 280108 217274
rect 279206 216988 279234 217110
rect 280034 216988 280062 217246
rect 280908 217138 280936 218010
rect 281736 217138 281764 218010
rect 282656 217274 282684 220866
rect 283380 220244 283432 220250
rect 283380 220186 283432 220192
rect 283392 217274 283420 220186
rect 280862 217110 280936 217138
rect 281690 217110 281764 217138
rect 282518 217246 282684 217274
rect 283346 217246 283420 217274
rect 284128 217274 284156 225558
rect 284772 223922 284800 231676
rect 285416 225214 285444 231676
rect 285588 228404 285640 228410
rect 285588 228346 285640 228352
rect 285404 225208 285456 225214
rect 285404 225150 285456 225156
rect 284760 223916 284812 223922
rect 284760 223858 284812 223864
rect 285600 219434 285628 228346
rect 286060 223446 286088 231676
rect 286324 226296 286376 226302
rect 286324 226238 286376 226244
rect 286048 223440 286100 223446
rect 286048 223382 286100 223388
rect 285508 219406 285628 219434
rect 285508 218074 285536 219406
rect 285864 219292 285916 219298
rect 285864 219234 285916 219240
rect 285036 218068 285088 218074
rect 285036 218010 285088 218016
rect 285496 218068 285548 218074
rect 285496 218010 285548 218016
rect 284128 217246 284202 217274
rect 280862 216988 280890 217110
rect 281690 216988 281718 217110
rect 282518 216988 282546 217246
rect 283346 216988 283374 217246
rect 284174 216988 284202 217246
rect 285048 217138 285076 218010
rect 285876 217138 285904 219234
rect 286336 218754 286364 226238
rect 286704 225350 286732 231676
rect 287348 229770 287376 231676
rect 287336 229764 287388 229770
rect 287336 229706 287388 229712
rect 287704 229764 287756 229770
rect 287704 229706 287756 229712
rect 286692 225344 286744 225350
rect 286692 225286 286744 225292
rect 286692 223984 286744 223990
rect 286692 223926 286744 223932
rect 286324 218748 286376 218754
rect 286324 218690 286376 218696
rect 286704 217274 286732 223926
rect 287716 220930 287744 229706
rect 287992 224806 288020 231676
rect 287980 224800 288032 224806
rect 287980 224742 288032 224748
rect 288636 223310 288664 231676
rect 288820 231662 289294 231690
rect 288624 223304 288676 223310
rect 288624 223246 288676 223252
rect 288256 223168 288308 223174
rect 288256 223110 288308 223116
rect 287888 222352 287940 222358
rect 287888 222294 287940 222300
rect 287704 220924 287756 220930
rect 287704 220866 287756 220872
rect 287900 218482 287928 222294
rect 287888 218476 287940 218482
rect 287888 218418 287940 218424
rect 287520 218068 287572 218074
rect 287520 218010 287572 218016
rect 285002 217110 285076 217138
rect 285830 217110 285904 217138
rect 286658 217246 286732 217274
rect 285002 216988 285030 217110
rect 285830 216988 285858 217110
rect 286658 216988 286686 217246
rect 287532 217138 287560 218010
rect 288268 217274 288296 223110
rect 288820 222194 288848 231662
rect 289924 226302 289952 231676
rect 290568 226778 290596 231676
rect 290556 226772 290608 226778
rect 290556 226714 290608 226720
rect 289912 226296 289964 226302
rect 289912 226238 289964 226244
rect 291016 226296 291068 226302
rect 291016 226238 291068 226244
rect 290832 224256 290884 224262
rect 290832 224198 290884 224204
rect 289728 223304 289780 223310
rect 289728 223246 289780 223252
rect 288544 222166 288848 222194
rect 288544 220114 288572 222166
rect 288532 220108 288584 220114
rect 288532 220050 288584 220056
rect 288716 220108 288768 220114
rect 288716 220050 288768 220056
rect 288728 218074 288756 220050
rect 289740 218074 289768 223246
rect 288716 218068 288768 218074
rect 288716 218010 288768 218016
rect 289176 218068 289228 218074
rect 289176 218010 289228 218016
rect 289728 218068 289780 218074
rect 289728 218010 289780 218016
rect 290004 218068 290056 218074
rect 290004 218010 290056 218016
rect 288268 217246 288342 217274
rect 287486 217110 287560 217138
rect 287486 216988 287514 217110
rect 288314 216988 288342 217246
rect 289188 217138 289216 218010
rect 290016 217138 290044 218010
rect 290844 217274 290872 224198
rect 291028 219434 291056 226238
rect 291212 223582 291240 231676
rect 291856 228954 291884 231676
rect 292500 229634 292528 231676
rect 292488 229628 292540 229634
rect 292488 229570 292540 229576
rect 291844 228948 291896 228954
rect 291844 228890 291896 228896
rect 291844 228812 291896 228818
rect 291844 228754 291896 228760
rect 291200 223576 291252 223582
rect 291200 223518 291252 223524
rect 291028 219406 291148 219434
rect 291120 218074 291148 219406
rect 291660 218884 291712 218890
rect 291660 218826 291712 218832
rect 291108 218068 291160 218074
rect 291108 218010 291160 218016
rect 289142 217110 289216 217138
rect 289970 217110 290044 217138
rect 290798 217246 290872 217274
rect 289142 216988 289170 217110
rect 289970 216988 289998 217110
rect 290798 216988 290826 217246
rect 291672 217138 291700 218826
rect 291856 218754 291884 228754
rect 293144 225894 293172 231676
rect 293328 231662 293802 231690
rect 293132 225888 293184 225894
rect 293132 225830 293184 225836
rect 292488 221468 292540 221474
rect 292488 221410 292540 221416
rect 291844 218748 291896 218754
rect 291844 218690 291896 218696
rect 292500 217274 292528 221410
rect 293328 220658 293356 231662
rect 293776 226908 293828 226914
rect 293776 226850 293828 226856
rect 293316 220652 293368 220658
rect 293316 220594 293368 220600
rect 293788 218074 293816 226850
rect 294432 224534 294460 231676
rect 294420 224528 294472 224534
rect 294420 224470 294472 224476
rect 295076 222358 295104 231676
rect 295720 229090 295748 231676
rect 295708 229084 295760 229090
rect 295708 229026 295760 229032
rect 296364 228274 296392 231676
rect 296628 228676 296680 228682
rect 296628 228618 296680 228624
rect 296352 228268 296404 228274
rect 296352 228210 296404 228216
rect 296444 225888 296496 225894
rect 296444 225830 296496 225836
rect 295064 222352 295116 222358
rect 295064 222294 295116 222300
rect 294972 220652 295024 220658
rect 294972 220594 295024 220600
rect 294144 218476 294196 218482
rect 294144 218418 294196 218424
rect 293316 218068 293368 218074
rect 293316 218010 293368 218016
rect 293776 218068 293828 218074
rect 293776 218010 293828 218016
rect 291626 217110 291700 217138
rect 292454 217246 292528 217274
rect 291626 216988 291654 217110
rect 292454 216988 292482 217246
rect 293328 217138 293356 218010
rect 294156 217138 294184 218418
rect 294984 217274 295012 220594
rect 296456 219434 296484 225830
rect 296456 219406 296576 219434
rect 295800 219156 295852 219162
rect 295800 219098 295852 219104
rect 293282 217110 293356 217138
rect 294110 217110 294184 217138
rect 294938 217246 295012 217274
rect 293282 216988 293310 217110
rect 294110 216988 294138 217110
rect 294938 216988 294966 217246
rect 295812 217138 295840 219098
rect 296548 217274 296576 219406
rect 296640 219178 296668 228618
rect 297008 225758 297036 231676
rect 297652 230314 297680 231676
rect 297640 230308 297692 230314
rect 297640 230250 297692 230256
rect 297824 230308 297876 230314
rect 297824 230250 297876 230256
rect 297836 229094 297864 230250
rect 297744 229066 297864 229094
rect 296996 225752 297048 225758
rect 296996 225694 297048 225700
rect 297272 225004 297324 225010
rect 297272 224946 297324 224952
rect 296640 219162 296760 219178
rect 296640 219156 296772 219162
rect 296640 219150 296720 219156
rect 296720 219098 296772 219104
rect 297284 219026 297312 224946
rect 297744 223310 297772 229066
rect 298296 227594 298324 231676
rect 298572 231662 298954 231690
rect 298284 227588 298336 227594
rect 298284 227530 298336 227536
rect 297916 223576 297968 223582
rect 297916 223518 297968 223524
rect 297732 223304 297784 223310
rect 297732 223246 297784 223252
rect 297272 219020 297324 219026
rect 297272 218962 297324 218968
rect 297928 218074 297956 223518
rect 298572 220794 298600 231662
rect 299584 227458 299612 231676
rect 300228 228818 300256 231676
rect 300216 228812 300268 228818
rect 300216 228754 300268 228760
rect 300676 228812 300728 228818
rect 300676 228754 300728 228760
rect 299572 227452 299624 227458
rect 299572 227394 299624 227400
rect 299296 224392 299348 224398
rect 299296 224334 299348 224340
rect 299112 223304 299164 223310
rect 299112 223246 299164 223252
rect 298560 220788 298612 220794
rect 298560 220730 298612 220736
rect 299124 218074 299152 223246
rect 297456 218068 297508 218074
rect 297456 218010 297508 218016
rect 297916 218068 297968 218074
rect 297916 218010 297968 218016
rect 298284 218068 298336 218074
rect 298284 218010 298336 218016
rect 299112 218068 299164 218074
rect 299112 218010 299164 218016
rect 296548 217246 296622 217274
rect 295766 217110 295840 217138
rect 295766 216988 295794 217110
rect 296594 216988 296622 217246
rect 297468 217138 297496 218010
rect 298296 217138 298324 218010
rect 299308 217274 299336 224334
rect 300492 218884 300544 218890
rect 300492 218826 300544 218832
rect 299940 218068 299992 218074
rect 299940 218010 299992 218016
rect 297422 217110 297496 217138
rect 298250 217110 298324 217138
rect 299078 217246 299336 217274
rect 297422 216988 297450 217110
rect 298250 216988 298278 217110
rect 299078 216988 299106 217246
rect 299952 217138 299980 218010
rect 300504 217274 300532 218826
rect 300688 218074 300716 228754
rect 300872 226166 300900 231676
rect 301240 231662 301530 231690
rect 301792 231662 302174 231690
rect 300860 226160 300912 226166
rect 300860 226102 300912 226108
rect 301240 221882 301268 231662
rect 301504 227588 301556 227594
rect 301504 227530 301556 227536
rect 301516 227050 301544 227530
rect 301504 227044 301556 227050
rect 301504 226986 301556 226992
rect 301228 221876 301280 221882
rect 301228 221818 301280 221824
rect 301412 221876 301464 221882
rect 301412 221818 301464 221824
rect 301424 219434 301452 221818
rect 301792 221610 301820 231662
rect 302804 230042 302832 231676
rect 302792 230036 302844 230042
rect 302792 229978 302844 229984
rect 303252 230036 303304 230042
rect 303252 229978 303304 229984
rect 302148 228948 302200 228954
rect 302148 228890 302200 228896
rect 301780 221604 301832 221610
rect 301780 221546 301832 221552
rect 301412 219428 301464 219434
rect 301412 219370 301464 219376
rect 302160 218074 302188 228890
rect 303264 223582 303292 229978
rect 303448 224874 303476 231676
rect 303816 231662 304106 231690
rect 304368 231662 304750 231690
rect 303436 224868 303488 224874
rect 303436 224810 303488 224816
rect 303252 223576 303304 223582
rect 303252 223518 303304 223524
rect 303252 221740 303304 221746
rect 303252 221682 303304 221688
rect 302424 220788 302476 220794
rect 302424 220730 302476 220736
rect 300676 218068 300728 218074
rect 300676 218010 300728 218016
rect 301596 218068 301648 218074
rect 301596 218010 301648 218016
rect 302148 218068 302200 218074
rect 302148 218010 302200 218016
rect 300504 217246 300762 217274
rect 299906 217110 299980 217138
rect 299906 216988 299934 217110
rect 300734 216988 300762 217246
rect 301608 217138 301636 218010
rect 302436 217274 302464 220730
rect 303264 217274 303292 221682
rect 303816 221338 303844 231662
rect 304368 222766 304396 231662
rect 304908 227452 304960 227458
rect 304908 227394 304960 227400
rect 304724 223440 304776 223446
rect 304724 223382 304776 223388
rect 304356 222760 304408 222766
rect 304356 222702 304408 222708
rect 303804 221332 303856 221338
rect 303804 221274 303856 221280
rect 304736 218074 304764 223382
rect 304080 218068 304132 218074
rect 304080 218010 304132 218016
rect 304724 218068 304776 218074
rect 304724 218010 304776 218016
rect 301562 217110 301636 217138
rect 302390 217246 302464 217274
rect 303218 217246 303292 217274
rect 301562 216988 301590 217110
rect 302390 216988 302418 217246
rect 303218 216988 303246 217246
rect 304092 217138 304120 218010
rect 304920 217274 304948 227394
rect 305380 225010 305408 231676
rect 305552 229084 305604 229090
rect 305552 229026 305604 229032
rect 305368 225004 305420 225010
rect 305368 224946 305420 224952
rect 305564 218618 305592 229026
rect 306024 228138 306052 231676
rect 306392 231662 306682 231690
rect 306852 231662 307326 231690
rect 306012 228132 306064 228138
rect 306012 228074 306064 228080
rect 306196 227316 306248 227322
rect 306196 227258 306248 227264
rect 305552 218612 305604 218618
rect 305552 218554 305604 218560
rect 306208 218074 306236 227258
rect 306392 222154 306420 231662
rect 306380 222148 306432 222154
rect 306380 222090 306432 222096
rect 306852 220522 306880 231662
rect 307956 230178 307984 231676
rect 307944 230172 307996 230178
rect 307944 230114 307996 230120
rect 308128 230172 308180 230178
rect 308128 230114 308180 230120
rect 307668 223576 307720 223582
rect 307668 223518 307720 223524
rect 306840 220516 306892 220522
rect 306840 220458 306892 220464
rect 307392 219020 307444 219026
rect 307392 218962 307444 218968
rect 305736 218068 305788 218074
rect 305736 218010 305788 218016
rect 306196 218068 306248 218074
rect 306196 218010 306248 218016
rect 306564 218068 306616 218074
rect 306564 218010 306616 218016
rect 304046 217110 304120 217138
rect 304874 217246 304948 217274
rect 304046 216988 304074 217110
rect 304874 216988 304902 217246
rect 305748 217138 305776 218010
rect 306576 217138 306604 218010
rect 307404 217138 307432 218962
rect 307680 218074 307708 223518
rect 308140 223446 308168 230114
rect 308600 227594 308628 231676
rect 308588 227588 308640 227594
rect 308588 227530 308640 227536
rect 309048 226160 309100 226166
rect 309048 226102 309100 226108
rect 308128 223440 308180 223446
rect 308128 223382 308180 223388
rect 308864 221604 308916 221610
rect 308864 221546 308916 221552
rect 308876 219434 308904 221546
rect 309060 219434 309088 226102
rect 309244 220386 309272 231676
rect 309888 228546 309916 231676
rect 310546 231662 310744 231690
rect 310716 229094 310744 231662
rect 310716 229066 310928 229094
rect 309876 228540 309928 228546
rect 309876 228482 309928 228488
rect 310428 227044 310480 227050
rect 310428 226986 310480 226992
rect 309232 220380 309284 220386
rect 309232 220322 309284 220328
rect 308220 219428 308272 219434
rect 308876 219406 308996 219434
rect 309060 219428 309192 219434
rect 309060 219406 309140 219428
rect 308220 219370 308272 219376
rect 307668 218068 307720 218074
rect 307668 218010 307720 218016
rect 308232 217138 308260 219370
rect 308968 217274 308996 219406
rect 309140 219370 309192 219376
rect 310440 218074 310468 226986
rect 310704 222148 310756 222154
rect 310704 222090 310756 222096
rect 309876 218068 309928 218074
rect 309876 218010 309928 218016
rect 310428 218068 310480 218074
rect 310428 218010 310480 218016
rect 308968 217246 309042 217274
rect 305702 217110 305776 217138
rect 306530 217110 306604 217138
rect 307358 217110 307432 217138
rect 308186 217110 308260 217138
rect 305702 216988 305730 217110
rect 306530 216988 306558 217110
rect 307358 216988 307386 217110
rect 308186 216988 308214 217110
rect 309014 216988 309042 217246
rect 309888 217138 309916 218010
rect 310716 217274 310744 222090
rect 310900 221882 310928 229066
rect 311176 224126 311204 231676
rect 311820 227730 311848 231676
rect 311992 230444 312044 230450
rect 311992 230386 312044 230392
rect 312004 229906 312032 230386
rect 311992 229900 312044 229906
rect 311992 229842 312044 229848
rect 311808 227724 311860 227730
rect 311808 227666 311860 227672
rect 311532 224800 311584 224806
rect 311532 224742 311584 224748
rect 311164 224120 311216 224126
rect 311164 224062 311216 224068
rect 310888 221876 310940 221882
rect 310888 221818 310940 221824
rect 311544 217274 311572 224742
rect 312464 224670 312492 231676
rect 313108 230450 313136 231676
rect 313292 231662 313766 231690
rect 313936 231662 314410 231690
rect 313096 230444 313148 230450
rect 313096 230386 313148 230392
rect 312636 229900 312688 229906
rect 312636 229842 312688 229848
rect 312452 224664 312504 224670
rect 312452 224606 312504 224612
rect 312648 222154 312676 229842
rect 313292 226030 313320 231662
rect 313936 229094 313964 231662
rect 313936 229066 314056 229094
rect 313832 228540 313884 228546
rect 313832 228482 313884 228488
rect 313280 226024 313332 226030
rect 313280 225966 313332 225972
rect 312912 223440 312964 223446
rect 312912 223382 312964 223388
rect 312636 222148 312688 222154
rect 312636 222090 312688 222096
rect 312924 218074 312952 223382
rect 313188 221876 313240 221882
rect 313188 221818 313240 221824
rect 312360 218068 312412 218074
rect 312360 218010 312412 218016
rect 312912 218068 312964 218074
rect 312912 218010 312964 218016
rect 309842 217110 309916 217138
rect 310670 217246 310744 217274
rect 311498 217246 311572 217274
rect 309842 216988 309870 217110
rect 310670 216988 310698 217246
rect 311498 216988 311526 217246
rect 312372 217138 312400 218010
rect 313200 217274 313228 221818
rect 313844 219298 313872 228482
rect 314028 222018 314056 229066
rect 315040 223038 315068 231676
rect 315684 229090 315712 231676
rect 315672 229084 315724 229090
rect 315672 229026 315724 229032
rect 315672 225752 315724 225758
rect 315672 225694 315724 225700
rect 315028 223032 315080 223038
rect 315028 222974 315080 222980
rect 314016 222012 314068 222018
rect 314016 221954 314068 221960
rect 314844 220380 314896 220386
rect 314844 220322 314896 220328
rect 314016 219428 314068 219434
rect 314016 219370 314068 219376
rect 313832 219292 313884 219298
rect 313832 219234 313884 219240
rect 312326 217110 312400 217138
rect 313154 217246 313228 217274
rect 312326 216988 312354 217110
rect 313154 216988 313182 217246
rect 314028 217138 314056 219370
rect 314856 217274 314884 220322
rect 315684 217274 315712 225694
rect 316328 222902 316356 231676
rect 316512 231662 316986 231690
rect 316316 222896 316368 222902
rect 316316 222838 316368 222844
rect 316512 220250 316540 231662
rect 317616 227186 317644 231676
rect 318260 229770 318288 231676
rect 318248 229764 318300 229770
rect 318248 229706 318300 229712
rect 318064 229628 318116 229634
rect 318064 229570 318116 229576
rect 317604 227180 317656 227186
rect 317604 227122 317656 227128
rect 316684 223032 316736 223038
rect 316684 222974 316736 222980
rect 316500 220244 316552 220250
rect 316500 220186 316552 220192
rect 316500 220108 316552 220114
rect 316500 220050 316552 220056
rect 316512 217274 316540 220050
rect 316696 218482 316724 222974
rect 318076 219434 318104 229570
rect 318904 228410 318932 231676
rect 318892 228404 318944 228410
rect 318892 228346 318944 228352
rect 319548 223990 319576 231676
rect 320192 225622 320220 231676
rect 320836 228546 320864 231676
rect 321112 231662 321494 231690
rect 320824 228540 320876 228546
rect 320824 228482 320876 228488
rect 320180 225616 320232 225622
rect 320180 225558 320232 225564
rect 319812 224664 319864 224670
rect 319812 224606 319864 224612
rect 319536 223984 319588 223990
rect 319536 223926 319588 223932
rect 319628 223712 319680 223718
rect 319628 223654 319680 223660
rect 318248 222012 318300 222018
rect 318248 221954 318300 221960
rect 318260 219434 318288 221954
rect 317984 219406 318104 219434
rect 318168 219406 318288 219434
rect 316684 218476 316736 218482
rect 316684 218418 316736 218424
rect 317984 218074 318012 219406
rect 317328 218068 317380 218074
rect 317328 218010 317380 218016
rect 317972 218068 318024 218074
rect 317972 218010 318024 218016
rect 313982 217110 314056 217138
rect 314810 217246 314884 217274
rect 315638 217246 315712 217274
rect 316466 217246 316540 217274
rect 313982 216988 314010 217110
rect 314810 216988 314838 217246
rect 315638 216988 315666 217246
rect 316466 216988 316494 217246
rect 317340 217138 317368 218010
rect 318168 217274 318196 219406
rect 319640 218074 319668 223654
rect 318984 218068 319036 218074
rect 318984 218010 319036 218016
rect 319628 218068 319680 218074
rect 319628 218010 319680 218016
rect 317294 217110 317368 217138
rect 318122 217246 318196 217274
rect 317294 216988 317322 217110
rect 318122 216988 318150 217246
rect 318996 217138 319024 218010
rect 319824 217274 319852 224606
rect 319996 224528 320048 224534
rect 319996 224470 320048 224476
rect 320008 223718 320036 224470
rect 319996 223712 320048 223718
rect 319996 223654 320048 223660
rect 321112 223174 321140 231662
rect 322124 226302 322152 231676
rect 322400 231662 322782 231690
rect 322112 226296 322164 226302
rect 322112 226238 322164 226244
rect 321376 226024 321428 226030
rect 321376 225966 321428 225972
rect 321100 223168 321152 223174
rect 321100 223110 321152 223116
rect 320640 219156 320692 219162
rect 320640 219098 320692 219104
rect 318950 217110 319024 217138
rect 319778 217246 319852 217274
rect 318950 216988 318978 217110
rect 319778 216988 319806 217246
rect 320652 217138 320680 219098
rect 321388 217274 321416 225966
rect 321652 220244 321704 220250
rect 321652 220186 321704 220192
rect 321664 218754 321692 220186
rect 322400 219978 322428 231662
rect 323412 230314 323440 231676
rect 323688 231662 324070 231690
rect 324516 231662 324714 231690
rect 324976 231662 325358 231690
rect 325896 231662 326002 231690
rect 326264 231662 326646 231690
rect 323400 230308 323452 230314
rect 323400 230250 323452 230256
rect 322848 227180 322900 227186
rect 322848 227122 322900 227128
rect 322388 219972 322440 219978
rect 322388 219914 322440 219920
rect 321652 218748 321704 218754
rect 321652 218690 321704 218696
rect 322860 218074 322888 227122
rect 323688 224262 323716 231662
rect 323676 224256 323728 224262
rect 323676 224198 323728 224204
rect 323952 224256 324004 224262
rect 323952 224198 324004 224204
rect 322296 218068 322348 218074
rect 322296 218010 322348 218016
rect 322848 218068 322900 218074
rect 322848 218010 322900 218016
rect 323124 218068 323176 218074
rect 323124 218010 323176 218016
rect 321388 217246 321462 217274
rect 320606 217110 320680 217138
rect 320606 216988 320634 217110
rect 321434 216988 321462 217246
rect 322308 217138 322336 218010
rect 323136 217138 323164 218010
rect 323964 217274 323992 224198
rect 324136 222896 324188 222902
rect 324136 222838 324188 222844
rect 324148 218074 324176 222838
rect 324516 220250 324544 231662
rect 324976 226914 325004 231662
rect 325424 228540 325476 228546
rect 325424 228482 325476 228488
rect 324964 226908 325016 226914
rect 324964 226850 325016 226856
rect 324504 220244 324556 220250
rect 324504 220186 324556 220192
rect 325436 218074 325464 228482
rect 325896 220658 325924 231662
rect 326264 221474 326292 231662
rect 326896 229084 326948 229090
rect 326896 229026 326948 229032
rect 326252 221468 326304 221474
rect 326252 221410 326304 221416
rect 325884 220652 325936 220658
rect 325884 220594 325936 220600
rect 325608 220108 325660 220114
rect 325608 220050 325660 220056
rect 324136 218068 324188 218074
rect 324136 218010 324188 218016
rect 324780 218068 324832 218074
rect 324780 218010 324832 218016
rect 325424 218068 325476 218074
rect 325424 218010 325476 218016
rect 322262 217110 322336 217138
rect 323090 217110 323164 217138
rect 323918 217246 323992 217274
rect 322262 216988 322290 217110
rect 323090 216988 323118 217110
rect 323918 216988 323946 217246
rect 324792 217138 324820 218010
rect 325620 217274 325648 220050
rect 326908 218074 326936 229026
rect 327276 223038 327304 231676
rect 327920 225894 327948 231676
rect 327908 225888 327960 225894
rect 327908 225830 327960 225836
rect 327724 225004 327776 225010
rect 327724 224946 327776 224952
rect 327264 223032 327316 223038
rect 327264 222974 327316 222980
rect 327736 218890 327764 224946
rect 328564 223310 328592 231676
rect 329208 228682 329236 231676
rect 329852 230042 329880 231676
rect 329840 230036 329892 230042
rect 329840 229978 329892 229984
rect 330496 228818 330524 231676
rect 330944 230036 330996 230042
rect 330944 229978 330996 229984
rect 330956 229094 330984 229978
rect 330956 229066 331076 229094
rect 330484 228812 330536 228818
rect 330484 228754 330536 228760
rect 329196 228676 329248 228682
rect 329196 228618 329248 228624
rect 330484 228404 330536 228410
rect 330484 228346 330536 228352
rect 329748 225888 329800 225894
rect 329748 225830 329800 225836
rect 328552 223304 328604 223310
rect 328552 223246 328604 223252
rect 328092 223032 328144 223038
rect 328092 222974 328144 222980
rect 327724 218884 327776 218890
rect 327724 218826 327776 218832
rect 327264 218748 327316 218754
rect 327264 218690 327316 218696
rect 326436 218068 326488 218074
rect 326436 218010 326488 218016
rect 326896 218068 326948 218074
rect 326896 218010 326948 218016
rect 324746 217110 324820 217138
rect 325574 217246 325648 217274
rect 324746 216988 324774 217110
rect 325574 216988 325602 217246
rect 326448 217138 326476 218010
rect 327276 217138 327304 218690
rect 328104 217274 328132 222974
rect 328920 218204 328972 218210
rect 328920 218146 328972 218152
rect 326402 217110 326476 217138
rect 327230 217110 327304 217138
rect 328058 217246 328132 217274
rect 326402 216988 326430 217110
rect 327230 216988 327258 217110
rect 328058 216988 328086 217246
rect 328932 217138 328960 218146
rect 329760 217274 329788 225830
rect 330300 219428 330352 219434
rect 330300 219370 330352 219376
rect 330312 219026 330340 219370
rect 330300 219020 330352 219026
rect 330300 218962 330352 218968
rect 330496 218210 330524 228346
rect 330484 218204 330536 218210
rect 330484 218146 330536 218152
rect 331048 218074 331076 229066
rect 331140 228970 331168 231676
rect 331140 228954 331260 228970
rect 331140 228948 331272 228954
rect 331140 228942 331220 228948
rect 331220 228890 331272 228896
rect 331784 224398 331812 231676
rect 332060 231662 332442 231690
rect 332796 231662 333086 231690
rect 332060 225010 332088 231662
rect 332232 225616 332284 225622
rect 332232 225558 332284 225564
rect 332048 225004 332100 225010
rect 332048 224946 332100 224952
rect 331772 224392 331824 224398
rect 331772 224334 331824 224340
rect 331404 222148 331456 222154
rect 331404 222090 331456 222096
rect 330576 218068 330628 218074
rect 330576 218010 330628 218016
rect 331036 218068 331088 218074
rect 331036 218010 331088 218016
rect 328886 217110 328960 217138
rect 329714 217246 329788 217274
rect 328886 216988 328914 217110
rect 329714 216988 329742 217246
rect 330588 217138 330616 218010
rect 331416 217274 331444 222090
rect 332244 217274 332272 225558
rect 332796 221746 332824 231662
rect 333716 227458 333744 231676
rect 334084 231662 334374 231690
rect 333704 227452 333756 227458
rect 333704 227394 333756 227400
rect 333888 227452 333940 227458
rect 333888 227394 333940 227400
rect 332784 221740 332836 221746
rect 332784 221682 332836 221688
rect 332692 220584 332744 220590
rect 332692 220526 332744 220532
rect 332704 218890 332732 220526
rect 333704 219428 333756 219434
rect 333704 219370 333756 219376
rect 332692 218884 332744 218890
rect 332692 218826 332744 218832
rect 333060 218068 333112 218074
rect 333060 218010 333112 218016
rect 330542 217110 330616 217138
rect 331370 217246 331444 217274
rect 332198 217246 332272 217274
rect 330542 216988 330570 217110
rect 331370 216988 331398 217246
rect 332198 216988 332226 217246
rect 333072 217138 333100 218010
rect 333716 217274 333744 219370
rect 333900 218074 333928 227394
rect 334084 220794 334112 231662
rect 335004 230178 335032 231676
rect 334992 230172 335044 230178
rect 334992 230114 335044 230120
rect 335176 230172 335228 230178
rect 335176 230114 335228 230120
rect 335188 229094 335216 230114
rect 335004 229066 335216 229094
rect 335004 224262 335032 229066
rect 335176 224392 335228 224398
rect 335176 224334 335228 224340
rect 334992 224256 335044 224262
rect 334992 224198 335044 224204
rect 334072 220788 334124 220794
rect 334072 220730 334124 220736
rect 335188 218074 335216 224334
rect 335648 223582 335676 231676
rect 336292 226166 336320 231676
rect 336464 228676 336516 228682
rect 336464 228618 336516 228624
rect 336280 226160 336332 226166
rect 336280 226102 336332 226108
rect 335636 223576 335688 223582
rect 335636 223518 335688 223524
rect 336004 223372 336056 223378
rect 336004 223314 336056 223320
rect 336016 219026 336044 223314
rect 336476 219434 336504 228618
rect 336936 227322 336964 231676
rect 337212 231662 337594 231690
rect 336924 227316 336976 227322
rect 336924 227258 336976 227264
rect 337212 220590 337240 231662
rect 338224 227050 338252 231676
rect 338212 227044 338264 227050
rect 338212 226986 338264 226992
rect 338672 227044 338724 227050
rect 338672 226986 338724 226992
rect 337200 220584 337252 220590
rect 337200 220526 337252 220532
rect 338028 220516 338080 220522
rect 338028 220458 338080 220464
rect 336384 219406 336504 219434
rect 336004 219020 336056 219026
rect 336004 218962 336056 218968
rect 333888 218068 333940 218074
rect 333888 218010 333940 218016
rect 334716 218068 334768 218074
rect 334716 218010 334768 218016
rect 335176 218068 335228 218074
rect 335176 218010 335228 218016
rect 335544 218068 335596 218074
rect 335544 218010 335596 218016
rect 333716 217246 333882 217274
rect 333026 217110 333100 217138
rect 333026 216988 333054 217110
rect 333854 216988 333882 217246
rect 334728 217138 334756 218010
rect 335556 217138 335584 218010
rect 336384 217274 336412 219406
rect 337200 219020 337252 219026
rect 337200 218962 337252 218968
rect 334682 217110 334756 217138
rect 335510 217110 335584 217138
rect 336338 217246 336412 217274
rect 334682 216988 334710 217110
rect 335510 216988 335538 217110
rect 336338 216988 336366 217246
rect 337212 217138 337240 218962
rect 338040 217274 338068 220458
rect 338684 218074 338712 226986
rect 338868 224806 338896 231676
rect 339526 231662 339724 231690
rect 338856 224800 338908 224806
rect 338856 224742 338908 224748
rect 339408 224256 339460 224262
rect 339408 224198 339460 224204
rect 339420 218074 339448 224198
rect 339696 221610 339724 231662
rect 340156 229906 340184 231676
rect 340432 231662 340814 231690
rect 341076 231662 341458 231690
rect 340144 229900 340196 229906
rect 340144 229842 340196 229848
rect 340432 221882 340460 231662
rect 340696 227316 340748 227322
rect 340696 227258 340748 227264
rect 340420 221876 340472 221882
rect 340420 221818 340472 221824
rect 339684 221604 339736 221610
rect 339684 221546 339736 221552
rect 340512 218884 340564 218890
rect 340512 218826 340564 218832
rect 338672 218068 338724 218074
rect 338672 218010 338724 218016
rect 338856 218068 338908 218074
rect 338856 218010 338908 218016
rect 339408 218068 339460 218074
rect 339408 218010 339460 218016
rect 339684 218068 339736 218074
rect 339684 218010 339736 218016
rect 337166 217110 337240 217138
rect 337994 217246 338068 217274
rect 337166 216988 337194 217110
rect 337994 216988 338022 217246
rect 338868 217138 338896 218010
rect 339696 217138 339724 218010
rect 340524 217138 340552 218826
rect 340708 218074 340736 227258
rect 341076 220386 341104 231662
rect 342088 223514 342116 231676
rect 342272 231662 342746 231690
rect 342916 231662 343390 231690
rect 343836 231662 344034 231690
rect 342076 223508 342128 223514
rect 342076 223450 342128 223456
rect 342272 223378 342300 231662
rect 342916 229094 342944 231662
rect 342640 229066 342944 229094
rect 342260 223372 342312 223378
rect 342260 223314 342312 223320
rect 341340 221604 341392 221610
rect 341340 221546 341392 221552
rect 341064 220380 341116 220386
rect 341064 220322 341116 220328
rect 340696 218068 340748 218074
rect 340696 218010 340748 218016
rect 341352 217274 341380 221546
rect 342168 221468 342220 221474
rect 342168 221410 342220 221416
rect 342180 217274 342208 221410
rect 342640 220250 342668 229066
rect 342812 223440 342864 223446
rect 342812 223382 342864 223388
rect 342628 220244 342680 220250
rect 342628 220186 342680 220192
rect 342824 219162 342852 223382
rect 343836 222018 343864 231662
rect 344664 225758 344692 231676
rect 345308 229770 345336 231676
rect 345664 229900 345716 229906
rect 345664 229842 345716 229848
rect 345296 229764 345348 229770
rect 345296 229706 345348 229712
rect 344652 225752 344704 225758
rect 344652 225694 344704 225700
rect 344652 223168 344704 223174
rect 344652 223110 344704 223116
rect 343824 222012 343876 222018
rect 343824 221954 343876 221960
rect 342996 220380 343048 220386
rect 342996 220322 343048 220328
rect 342812 219156 342864 219162
rect 342812 219098 342864 219104
rect 343008 217274 343036 220322
rect 343824 219156 343876 219162
rect 343824 219098 343876 219104
rect 338822 217110 338896 217138
rect 339650 217110 339724 217138
rect 340478 217110 340552 217138
rect 341306 217246 341380 217274
rect 342134 217246 342208 217274
rect 342962 217246 343036 217274
rect 338822 216988 338850 217110
rect 339650 216988 339678 217110
rect 340478 216988 340506 217110
rect 341306 216988 341334 217246
rect 342134 216988 342162 217246
rect 342962 216988 342990 217246
rect 343836 217138 343864 219098
rect 344664 217274 344692 223110
rect 345676 219026 345704 229842
rect 345952 224670 345980 231676
rect 346596 226030 346624 231676
rect 346584 226024 346636 226030
rect 346584 225966 346636 225972
rect 347044 225752 347096 225758
rect 347044 225694 347096 225700
rect 345940 224664 345992 224670
rect 345940 224606 345992 224612
rect 346216 224664 346268 224670
rect 346216 224606 346268 224612
rect 345664 219020 345716 219026
rect 345664 218962 345716 218968
rect 345480 218068 345532 218074
rect 345480 218010 345532 218016
rect 343790 217110 343864 217138
rect 344618 217246 344692 217274
rect 343790 216988 343818 217110
rect 344618 216988 344646 217246
rect 345492 217138 345520 218010
rect 346228 217274 346256 224606
rect 347056 218074 347084 225694
rect 347240 224534 347268 231676
rect 347228 224528 347280 224534
rect 347228 224470 347280 224476
rect 347884 223446 347912 231676
rect 347872 223440 347924 223446
rect 347872 223382 347924 223388
rect 347228 223304 347280 223310
rect 347228 223246 347280 223252
rect 347240 219434 347268 223246
rect 348528 222902 348556 231676
rect 349172 228546 349200 231676
rect 349160 228540 349212 228546
rect 349160 228482 349212 228488
rect 349816 227186 349844 231676
rect 350460 230178 350488 231676
rect 350448 230172 350500 230178
rect 350448 230114 350500 230120
rect 351104 229090 351132 231676
rect 351472 231662 351762 231690
rect 352116 231662 352406 231690
rect 351092 229084 351144 229090
rect 351092 229026 351144 229032
rect 350448 228540 350500 228546
rect 350448 228482 350500 228488
rect 349804 227180 349856 227186
rect 349804 227122 349856 227128
rect 350264 226364 350316 226370
rect 350264 226306 350316 226312
rect 348516 222896 348568 222902
rect 348516 222838 348568 222844
rect 349068 222896 349120 222902
rect 349068 222838 349120 222844
rect 348792 220244 348844 220250
rect 348792 220186 348844 220192
rect 347228 219428 347280 219434
rect 347228 219370 347280 219376
rect 347228 219020 347280 219026
rect 347228 218962 347280 218968
rect 347044 218068 347096 218074
rect 347044 218010 347096 218016
rect 347240 217274 347268 218962
rect 347964 218068 348016 218074
rect 347964 218010 348016 218016
rect 346228 217246 346302 217274
rect 345446 217110 345520 217138
rect 345446 216988 345474 217110
rect 346274 216988 346302 217246
rect 347102 217246 347268 217274
rect 347102 216988 347130 217246
rect 347976 217138 348004 218010
rect 348804 217274 348832 220186
rect 349080 218074 349108 222838
rect 350276 219434 350304 226306
rect 350460 219434 350488 228482
rect 351092 226500 351144 226506
rect 351092 226442 351144 226448
rect 349620 219428 349672 219434
rect 350276 219406 350396 219434
rect 350460 219428 350592 219434
rect 350460 219406 350540 219428
rect 349620 219370 349672 219376
rect 349068 218068 349120 218074
rect 349068 218010 349120 218016
rect 347930 217110 348004 217138
rect 348758 217246 348832 217274
rect 347930 216988 347958 217110
rect 348758 216988 348786 217246
rect 349632 217138 349660 219370
rect 350368 217274 350396 219406
rect 350540 219370 350592 219376
rect 351104 218754 351132 226442
rect 351472 223038 351500 231662
rect 351736 229764 351788 229770
rect 351736 229706 351788 229712
rect 351748 226370 351776 229706
rect 351736 226364 351788 226370
rect 351736 226306 351788 226312
rect 351460 223032 351512 223038
rect 351460 222974 351512 222980
rect 351276 221876 351328 221882
rect 351276 221818 351328 221824
rect 351092 218748 351144 218754
rect 351092 218690 351144 218696
rect 351288 217274 351316 221818
rect 352116 220114 352144 231662
rect 353036 226506 353064 231676
rect 353024 226500 353076 226506
rect 353024 226442 353076 226448
rect 352932 226024 352984 226030
rect 352932 225966 352984 225972
rect 352104 220108 352156 220114
rect 352104 220050 352156 220056
rect 352104 219428 352156 219434
rect 352104 219370 352156 219376
rect 350368 217246 350442 217274
rect 349586 217110 349660 217138
rect 349586 216988 349614 217110
rect 350414 216988 350442 217246
rect 351242 217246 351316 217274
rect 351242 216988 351270 217246
rect 352116 217138 352144 219370
rect 352944 217274 352972 225966
rect 353680 225894 353708 231676
rect 353864 231662 354338 231690
rect 353668 225888 353720 225894
rect 353668 225830 353720 225836
rect 353864 223122 353892 231662
rect 354968 228410 354996 231676
rect 355612 230042 355640 231676
rect 355600 230036 355652 230042
rect 355600 229978 355652 229984
rect 354956 228404 355008 228410
rect 354956 228346 355008 228352
rect 355324 228404 355376 228410
rect 355324 228346 355376 228352
rect 354588 225888 354640 225894
rect 354588 225830 354640 225836
rect 353772 223094 353892 223122
rect 353772 222154 353800 223094
rect 353944 223032 353996 223038
rect 353944 222974 353996 222980
rect 353760 222148 353812 222154
rect 353760 222090 353812 222096
rect 353956 219162 353984 222974
rect 353944 219156 353996 219162
rect 353944 219098 353996 219104
rect 353760 218748 353812 218754
rect 353760 218690 353812 218696
rect 352070 217110 352144 217138
rect 352898 217246 352972 217274
rect 352070 216988 352098 217110
rect 352898 216988 352926 217246
rect 353772 217138 353800 218690
rect 354600 217274 354628 225830
rect 355336 219434 355364 228346
rect 356256 227458 356284 231676
rect 356244 227452 356296 227458
rect 356244 227394 356296 227400
rect 355876 227180 355928 227186
rect 355876 227122 355928 227128
rect 355324 219428 355376 219434
rect 355324 219370 355376 219376
rect 355888 218074 355916 227122
rect 356900 224398 356928 231676
rect 357072 227452 357124 227458
rect 357072 227394 357124 227400
rect 356888 224392 356940 224398
rect 356888 224334 356940 224340
rect 357084 222034 357112 227394
rect 357544 225622 357572 231676
rect 357912 231662 358202 231690
rect 357532 225616 357584 225622
rect 357532 225558 357584 225564
rect 357912 223310 357940 231662
rect 358832 228682 358860 231676
rect 359016 231662 359490 231690
rect 358820 228676 358872 228682
rect 358820 228618 358872 228624
rect 358084 224256 358136 224262
rect 358084 224198 358136 224204
rect 357900 223304 357952 223310
rect 357900 223246 357952 223252
rect 356992 222006 357112 222034
rect 356992 218074 357020 222006
rect 357164 221740 357216 221746
rect 357164 221682 357216 221688
rect 355416 218068 355468 218074
rect 355416 218010 355468 218016
rect 355876 218068 355928 218074
rect 355876 218010 355928 218016
rect 356244 218068 356296 218074
rect 356244 218010 356296 218016
rect 356980 218068 357032 218074
rect 356980 218010 357032 218016
rect 353726 217110 353800 217138
rect 354554 217246 354628 217274
rect 353726 216988 353754 217110
rect 354554 216988 354582 217246
rect 355428 217138 355456 218010
rect 356256 217138 356284 218010
rect 357176 217274 357204 221682
rect 357900 220652 357952 220658
rect 357900 220594 357952 220600
rect 357912 217274 357940 220594
rect 358096 218890 358124 224198
rect 359016 220522 359044 231662
rect 359924 228676 359976 228682
rect 359924 228618 359976 228624
rect 359004 220516 359056 220522
rect 359004 220458 359056 220464
rect 358820 220108 358872 220114
rect 358820 220050 358872 220056
rect 358832 219434 358860 220050
rect 358740 219406 358860 219434
rect 359936 219434 359964 228618
rect 360120 227050 360148 231676
rect 360764 229906 360792 231676
rect 360752 229900 360804 229906
rect 360752 229842 360804 229848
rect 361212 229900 361264 229906
rect 361212 229842 361264 229848
rect 361224 229094 361252 229842
rect 361040 229066 361252 229094
rect 360108 227044 360160 227050
rect 360108 226986 360160 226992
rect 359936 219406 360148 219434
rect 358084 218884 358136 218890
rect 358084 218826 358136 218832
rect 358740 217274 358768 219406
rect 360120 218074 360148 219406
rect 361040 218074 361068 229066
rect 361408 227322 361436 231676
rect 361776 231662 362066 231690
rect 362328 231662 362710 231690
rect 362972 231662 363354 231690
rect 363524 231662 363998 231690
rect 361396 227316 361448 227322
rect 361396 227258 361448 227264
rect 361212 224392 361264 224398
rect 361212 224334 361264 224340
rect 359556 218068 359608 218074
rect 359556 218010 359608 218016
rect 360108 218068 360160 218074
rect 360108 218010 360160 218016
rect 360384 218068 360436 218074
rect 360384 218010 360436 218016
rect 361028 218068 361080 218074
rect 361028 218010 361080 218016
rect 355382 217110 355456 217138
rect 356210 217110 356284 217138
rect 357038 217246 357204 217274
rect 357866 217246 357940 217274
rect 358694 217246 358768 217274
rect 355382 216988 355410 217110
rect 356210 216988 356238 217110
rect 357038 216988 357066 217246
rect 357866 216988 357894 217246
rect 358694 216988 358722 217246
rect 359568 217138 359596 218010
rect 360396 217138 360424 218010
rect 361224 217274 361252 224334
rect 361776 221610 361804 231662
rect 362328 224126 362356 231662
rect 362776 227044 362828 227050
rect 362776 226986 362828 226992
rect 362316 224120 362368 224126
rect 362316 224062 362368 224068
rect 361764 221604 361816 221610
rect 361764 221546 361816 221552
rect 362040 219428 362092 219434
rect 362040 219370 362092 219376
rect 359522 217110 359596 217138
rect 360350 217110 360424 217138
rect 361178 217246 361252 217274
rect 359522 216988 359550 217110
rect 360350 216988 360378 217110
rect 361178 216988 361206 217246
rect 362052 217138 362080 219370
rect 362788 217274 362816 226986
rect 362972 224262 363000 231662
rect 363524 229094 363552 231662
rect 363340 229066 363552 229094
rect 362960 224256 363012 224262
rect 362960 224198 363012 224204
rect 363340 220386 363368 229066
rect 363512 224528 363564 224534
rect 363512 224470 363564 224476
rect 363328 220380 363380 220386
rect 363328 220322 363380 220328
rect 363524 219026 363552 224470
rect 364628 223174 364656 231676
rect 364812 231662 365286 231690
rect 364616 223168 364668 223174
rect 364616 223110 364668 223116
rect 364812 221474 364840 231662
rect 365536 223168 365588 223174
rect 365536 223110 365588 223116
rect 364800 221468 364852 221474
rect 364800 221410 364852 221416
rect 363696 219156 363748 219162
rect 363696 219098 363748 219104
rect 363512 219020 363564 219026
rect 363512 218962 363564 218968
rect 362788 217246 362862 217274
rect 362006 217110 362080 217138
rect 362006 216988 362034 217110
rect 362834 216988 362862 217246
rect 363708 217138 363736 219098
rect 365352 218204 365404 218210
rect 365352 218146 365404 218152
rect 364524 218068 364576 218074
rect 364524 218010 364576 218016
rect 364536 217138 364564 218010
rect 365364 217138 365392 218146
rect 365548 218074 365576 223110
rect 365916 223038 365944 231676
rect 366560 224738 366588 231676
rect 366548 224732 366600 224738
rect 366548 224674 366600 224680
rect 366732 224256 366784 224262
rect 366732 224198 366784 224204
rect 365904 223032 365956 223038
rect 365904 222974 365956 222980
rect 366744 218074 366772 224198
rect 366916 223032 366968 223038
rect 366916 222974 366968 222980
rect 365536 218068 365588 218074
rect 365536 218010 365588 218016
rect 366180 218068 366232 218074
rect 366180 218010 366232 218016
rect 366732 218068 366784 218074
rect 366732 218010 366784 218016
rect 366192 217138 366220 218010
rect 366928 217274 366956 222974
rect 367204 222902 367232 231676
rect 367848 225758 367876 231676
rect 367836 225752 367888 225758
rect 367836 225694 367888 225700
rect 368492 224534 368520 231676
rect 369136 228546 369164 231676
rect 369320 231662 369794 231690
rect 369964 231662 370438 231690
rect 369124 228540 369176 228546
rect 369124 228482 369176 228488
rect 369124 225004 369176 225010
rect 369124 224946 369176 224952
rect 368480 224528 368532 224534
rect 368480 224470 368532 224476
rect 367192 222896 367244 222902
rect 367192 222838 367244 222844
rect 368388 222896 368440 222902
rect 368388 222838 368440 222844
rect 367652 222012 367704 222018
rect 367652 221954 367704 221960
rect 367664 219434 367692 221954
rect 367652 219428 367704 219434
rect 367652 219370 367704 219376
rect 368400 218074 368428 222838
rect 368664 219020 368716 219026
rect 368664 218962 368716 218968
rect 367836 218068 367888 218074
rect 367836 218010 367888 218016
rect 368388 218068 368440 218074
rect 368388 218010 368440 218016
rect 366928 217246 367002 217274
rect 363662 217110 363736 217138
rect 364490 217110 364564 217138
rect 365318 217110 365392 217138
rect 366146 217110 366220 217138
rect 363662 216988 363690 217110
rect 364490 216988 364518 217110
rect 365318 216988 365346 217110
rect 366146 216988 366174 217110
rect 366974 216988 367002 217246
rect 367848 217138 367876 218010
rect 368676 217138 368704 218962
rect 369136 218754 369164 224946
rect 369320 221882 369348 231662
rect 369308 221876 369360 221882
rect 369308 221818 369360 221824
rect 369492 221604 369544 221610
rect 369492 221546 369544 221552
rect 369124 218748 369176 218754
rect 369124 218690 369176 218696
rect 369504 217274 369532 221546
rect 369964 220250 369992 231662
rect 371068 229770 371096 231676
rect 371056 229764 371108 229770
rect 371056 229706 371108 229712
rect 371056 228540 371108 228546
rect 371056 228482 371108 228488
rect 369952 220244 370004 220250
rect 369952 220186 370004 220192
rect 370504 220244 370556 220250
rect 370504 220186 370556 220192
rect 370516 219162 370544 220186
rect 370504 219156 370556 219162
rect 370504 219098 370556 219104
rect 370320 218748 370372 218754
rect 370320 218690 370372 218696
rect 370332 217274 370360 218690
rect 367802 217110 367876 217138
rect 368630 217110 368704 217138
rect 369458 217246 369532 217274
rect 370286 217246 370360 217274
rect 371068 217274 371096 228482
rect 371712 226030 371740 231676
rect 371700 226024 371752 226030
rect 371700 225966 371752 225972
rect 372356 225894 372384 231676
rect 373000 228410 373028 231676
rect 372988 228404 373040 228410
rect 372988 228346 373040 228352
rect 373448 228404 373500 228410
rect 373448 228346 373500 228352
rect 372344 225888 372396 225894
rect 372344 225830 372396 225836
rect 371792 225752 371844 225758
rect 371792 225694 371844 225700
rect 371804 218210 371832 225694
rect 372528 225616 372580 225622
rect 372528 225558 372580 225564
rect 371792 218204 371844 218210
rect 371792 218146 371844 218152
rect 372540 218074 372568 225558
rect 373460 218074 373488 228346
rect 373644 225010 373672 231676
rect 374288 227458 374316 231676
rect 374472 231662 374946 231690
rect 374276 227452 374328 227458
rect 374276 227394 374328 227400
rect 373816 225888 373868 225894
rect 373816 225830 373868 225836
rect 373632 225004 373684 225010
rect 373632 224946 373684 224952
rect 373828 219434 373856 225830
rect 374472 220658 374500 231662
rect 374644 230444 374696 230450
rect 374644 230386 374696 230392
rect 374656 221746 374684 230386
rect 375576 227186 375604 231676
rect 376220 230450 376248 231676
rect 376208 230444 376260 230450
rect 376208 230386 376260 230392
rect 376024 228812 376076 228818
rect 376024 228754 376076 228760
rect 375564 227180 375616 227186
rect 375564 227122 375616 227128
rect 374644 221740 374696 221746
rect 374644 221682 374696 221688
rect 375288 221468 375340 221474
rect 375288 221410 375340 221416
rect 374460 220652 374512 220658
rect 374460 220594 374512 220600
rect 373644 219406 373856 219434
rect 371976 218068 372028 218074
rect 371976 218010 372028 218016
rect 372528 218068 372580 218074
rect 372528 218010 372580 218016
rect 372804 218068 372856 218074
rect 372804 218010 372856 218016
rect 373448 218068 373500 218074
rect 373448 218010 373500 218016
rect 371068 217246 371142 217274
rect 367802 216988 367830 217110
rect 368630 216988 368658 217110
rect 369458 216988 369486 217246
rect 370286 216988 370314 217246
rect 371114 216988 371142 217246
rect 371988 217138 372016 218010
rect 372816 217138 372844 218010
rect 373644 217274 373672 219406
rect 374460 218204 374512 218210
rect 374460 218146 374512 218152
rect 371942 217110 372016 217138
rect 372770 217110 372844 217138
rect 373598 217246 373672 217274
rect 371942 216988 371970 217110
rect 372770 216988 372798 217110
rect 373598 216988 373626 217246
rect 374472 217138 374500 218146
rect 375300 217274 375328 221410
rect 376036 218210 376064 228754
rect 376864 228682 376892 231676
rect 376852 228676 376904 228682
rect 376852 228618 376904 228624
rect 376668 227180 376720 227186
rect 376668 227122 376720 227128
rect 376024 218204 376076 218210
rect 376024 218146 376076 218152
rect 376680 218074 376708 227122
rect 377508 224398 377536 231676
rect 378166 231662 378364 231690
rect 377680 229764 377732 229770
rect 377680 229706 377732 229712
rect 377692 225894 377720 229706
rect 377680 225888 377732 225894
rect 377680 225830 377732 225836
rect 377864 225888 377916 225894
rect 377864 225830 377916 225836
rect 377496 224392 377548 224398
rect 377496 224334 377548 224340
rect 377404 224120 377456 224126
rect 377404 224062 377456 224068
rect 377416 219026 377444 224062
rect 377876 219434 377904 225830
rect 378336 220114 378364 231662
rect 378796 229906 378824 231676
rect 378784 229900 378836 229906
rect 378784 229842 378836 229848
rect 379440 227050 379468 231676
rect 379624 231662 380098 231690
rect 380268 231662 380742 231690
rect 381096 231662 381386 231690
rect 381648 231662 382030 231690
rect 382384 231662 382674 231690
rect 382844 231662 383318 231690
rect 379428 227044 379480 227050
rect 379428 226986 379480 226992
rect 379244 224392 379296 224398
rect 379244 224334 379296 224340
rect 378324 220108 378376 220114
rect 378324 220050 378376 220056
rect 377784 219406 377904 219434
rect 377404 219020 377456 219026
rect 377404 218962 377456 218968
rect 376944 218884 376996 218890
rect 376944 218826 376996 218832
rect 376116 218068 376168 218074
rect 376116 218010 376168 218016
rect 376668 218068 376720 218074
rect 376668 218010 376720 218016
rect 374426 217110 374500 217138
rect 375254 217246 375328 217274
rect 374426 216988 374454 217110
rect 375254 216988 375282 217246
rect 376128 217138 376156 218010
rect 376956 217138 376984 218826
rect 377784 217274 377812 219406
rect 379256 218074 379284 224334
rect 379624 223174 379652 231662
rect 379612 223168 379664 223174
rect 379612 223110 379664 223116
rect 380072 223168 380124 223174
rect 380072 223110 380124 223116
rect 379428 220108 379480 220114
rect 379428 220050 379480 220056
rect 378600 218068 378652 218074
rect 378600 218010 378652 218016
rect 379244 218068 379296 218074
rect 379244 218010 379296 218016
rect 376082 217110 376156 217138
rect 376910 217110 376984 217138
rect 377738 217246 377812 217274
rect 376082 216988 376110 217110
rect 376910 216988 376938 217110
rect 377738 216988 377766 217246
rect 378612 217138 378640 218010
rect 379440 217274 379468 220050
rect 380084 218754 380112 223110
rect 380268 222018 380296 231662
rect 380256 222012 380308 222018
rect 380256 221954 380308 221960
rect 381096 220250 381124 231662
rect 381648 224262 381676 231662
rect 382096 227316 382148 227322
rect 382096 227258 382148 227264
rect 381636 224256 381688 224262
rect 381636 224198 381688 224204
rect 381084 220244 381136 220250
rect 381084 220186 381136 220192
rect 380256 219428 380308 219434
rect 380256 219370 380308 219376
rect 380072 218748 380124 218754
rect 380072 218690 380124 218696
rect 378566 217110 378640 217138
rect 379394 217246 379468 217274
rect 378566 216988 378594 217110
rect 379394 216988 379422 217246
rect 380268 217138 380296 219370
rect 381912 218204 381964 218210
rect 381912 218146 381964 218152
rect 381084 218068 381136 218074
rect 381084 218010 381136 218016
rect 381096 217138 381124 218010
rect 381924 217138 381952 218146
rect 382108 218074 382136 227258
rect 382384 222902 382412 231662
rect 382844 229094 382872 231662
rect 383948 229094 383976 231676
rect 384132 231662 384606 231690
rect 384132 229094 384160 231662
rect 382752 229066 382872 229094
rect 383856 229066 383976 229094
rect 384040 229066 384160 229094
rect 382752 225758 382780 229066
rect 382740 225752 382792 225758
rect 382740 225694 382792 225700
rect 382924 225752 382976 225758
rect 382924 225694 382976 225700
rect 382372 222896 382424 222902
rect 382372 222838 382424 222844
rect 382740 218884 382792 218890
rect 382740 218826 382792 218832
rect 382096 218068 382148 218074
rect 382096 218010 382148 218016
rect 382752 217138 382780 218826
rect 382936 218210 382964 225694
rect 383856 223038 383884 229066
rect 383844 223032 383896 223038
rect 383844 222974 383896 222980
rect 383476 222896 383528 222902
rect 383476 222838 383528 222844
rect 383488 218890 383516 222838
rect 384040 221610 384068 229066
rect 385236 228546 385264 231676
rect 385224 228540 385276 228546
rect 385224 228482 385276 228488
rect 385880 224126 385908 231676
rect 386052 228540 386104 228546
rect 386052 228482 386104 228488
rect 385868 224120 385920 224126
rect 385868 224062 385920 224068
rect 384212 223032 384264 223038
rect 384212 222974 384264 222980
rect 384028 221604 384080 221610
rect 384028 221546 384080 221552
rect 384224 219434 384252 222974
rect 384396 221604 384448 221610
rect 384396 221546 384448 221552
rect 384212 219428 384264 219434
rect 384212 219370 384264 219376
rect 383476 218884 383528 218890
rect 383476 218826 383528 218832
rect 383568 218748 383620 218754
rect 383568 218690 383620 218696
rect 382924 218204 382976 218210
rect 382924 218146 382976 218152
rect 383580 217138 383608 218690
rect 384408 217274 384436 221546
rect 385224 220788 385276 220794
rect 385224 220730 385276 220736
rect 385236 217274 385264 220730
rect 386064 217274 386092 228482
rect 386524 223174 386552 231676
rect 387168 228410 387196 231676
rect 387432 230376 387484 230382
rect 387432 230318 387484 230324
rect 387156 228404 387208 228410
rect 387156 228346 387208 228352
rect 387444 225622 387472 230318
rect 387812 228818 387840 231676
rect 388456 230382 388484 231676
rect 388444 230376 388496 230382
rect 388444 230318 388496 230324
rect 389100 229770 389128 231676
rect 389088 229764 389140 229770
rect 389088 229706 389140 229712
rect 388628 229628 388680 229634
rect 388628 229570 388680 229576
rect 388640 229094 388668 229570
rect 388640 229066 388760 229094
rect 387800 228812 387852 228818
rect 387800 228754 387852 228760
rect 388536 226364 388588 226370
rect 388536 226306 388588 226312
rect 387432 225616 387484 225622
rect 387432 225558 387484 225564
rect 387708 224528 387760 224534
rect 387708 224470 387760 224476
rect 386512 223168 386564 223174
rect 386512 223110 386564 223116
rect 386880 219020 386932 219026
rect 386880 218962 386932 218968
rect 380222 217110 380296 217138
rect 381050 217110 381124 217138
rect 381878 217110 381952 217138
rect 382706 217110 382780 217138
rect 383534 217110 383608 217138
rect 384362 217246 384436 217274
rect 385190 217246 385264 217274
rect 386018 217246 386092 217274
rect 380222 216988 380250 217110
rect 381050 216988 381078 217110
rect 381878 216988 381906 217110
rect 382706 216988 382734 217110
rect 383534 216988 383562 217110
rect 384362 216988 384390 217246
rect 385190 216988 385218 217246
rect 386018 216988 386046 217246
rect 386892 217138 386920 218962
rect 387720 217274 387748 224470
rect 388548 218890 388576 226306
rect 388732 220794 388760 229066
rect 389744 227186 389772 231676
rect 390008 228404 390060 228410
rect 390008 228346 390060 228352
rect 389732 227180 389784 227186
rect 389732 227122 389784 227128
rect 388720 220788 388772 220794
rect 388720 220730 388772 220736
rect 388720 220244 388772 220250
rect 388720 220186 388772 220192
rect 388536 218884 388588 218890
rect 388536 218826 388588 218832
rect 388732 217274 388760 220186
rect 390020 218074 390048 228346
rect 390388 225894 390416 231676
rect 390756 231662 391046 231690
rect 390376 225888 390428 225894
rect 390376 225830 390428 225836
rect 390192 225616 390244 225622
rect 390192 225558 390244 225564
rect 389364 218068 389416 218074
rect 389364 218010 389416 218016
rect 390008 218068 390060 218074
rect 390008 218010 390060 218016
rect 386846 217110 386920 217138
rect 387674 217246 387748 217274
rect 388502 217246 388760 217274
rect 386846 216988 386874 217110
rect 387674 216988 387702 217246
rect 388502 216988 388530 217246
rect 389376 217138 389404 218010
rect 390204 217274 390232 225558
rect 390756 221474 390784 231662
rect 391676 226370 391704 231676
rect 392136 231662 392334 231690
rect 391848 227044 391900 227050
rect 391848 226986 391900 226992
rect 391664 226364 391716 226370
rect 391664 226306 391716 226312
rect 391020 221740 391072 221746
rect 391020 221682 391072 221688
rect 390744 221468 390796 221474
rect 390744 221410 390796 221416
rect 391032 217274 391060 221682
rect 391860 219434 391888 226986
rect 392136 220114 392164 231662
rect 392964 227322 392992 231676
rect 392952 227316 393004 227322
rect 392952 227258 393004 227264
rect 393136 227180 393188 227186
rect 393136 227122 393188 227128
rect 392124 220108 392176 220114
rect 392124 220050 392176 220056
rect 389330 217110 389404 217138
rect 390158 217246 390232 217274
rect 390986 217246 391060 217274
rect 391768 219406 391888 219434
rect 391768 217274 391796 219406
rect 393148 218074 393176 227122
rect 393608 224398 393636 231676
rect 393976 231662 394266 231690
rect 393596 224392 393648 224398
rect 393596 224334 393648 224340
rect 393976 223038 394004 231662
rect 394332 225888 394384 225894
rect 394332 225830 394384 225836
rect 393964 223032 394016 223038
rect 393964 222974 394016 222980
rect 392676 218068 392728 218074
rect 392676 218010 392728 218016
rect 393136 218068 393188 218074
rect 393136 218010 393188 218016
rect 393504 218068 393556 218074
rect 393504 218010 393556 218016
rect 391768 217246 391842 217274
rect 389330 216988 389358 217110
rect 390158 216988 390186 217246
rect 390986 216988 391014 217246
rect 391814 216988 391842 217246
rect 392688 217138 392716 218010
rect 393516 217138 393544 218010
rect 394344 217274 394372 225830
rect 394516 224256 394568 224262
rect 394516 224198 394568 224204
rect 394528 218074 394556 224198
rect 394896 222902 394924 231676
rect 395172 231662 395554 231690
rect 394884 222896 394936 222902
rect 394884 222838 394936 222844
rect 395172 221610 395200 231662
rect 396184 225758 396212 231676
rect 396368 231662 396842 231690
rect 396172 225752 396224 225758
rect 396172 225694 396224 225700
rect 395804 222896 395856 222902
rect 395804 222838 395856 222844
rect 395160 221604 395212 221610
rect 395160 221546 395212 221552
rect 395816 218074 395844 222838
rect 395988 220108 396040 220114
rect 395988 220050 396040 220056
rect 394516 218068 394568 218074
rect 394516 218010 394568 218016
rect 395160 218068 395212 218074
rect 395160 218010 395212 218016
rect 395804 218068 395856 218074
rect 395804 218010 395856 218016
rect 392642 217110 392716 217138
rect 393470 217110 393544 217138
rect 394298 217246 394372 217274
rect 392642 216988 392670 217110
rect 393470 216988 393498 217110
rect 394298 216988 394326 217246
rect 395172 217138 395200 218010
rect 396000 217274 396028 220050
rect 396368 219434 396396 231662
rect 397472 228546 397500 231676
rect 397840 231662 398130 231690
rect 397460 228540 397512 228546
rect 397460 228482 397512 228488
rect 397840 224534 397868 231662
rect 398104 230376 398156 230382
rect 398104 230318 398156 230324
rect 397828 224528 397880 224534
rect 397828 224470 397880 224476
rect 396816 221468 396868 221474
rect 396816 221410 396868 221416
rect 396276 219406 396396 219434
rect 396276 218754 396304 219406
rect 396264 218748 396316 218754
rect 396264 218690 396316 218696
rect 396828 217274 396856 221410
rect 398116 219026 398144 230318
rect 398760 229634 398788 231676
rect 399404 230382 399432 231676
rect 399392 230376 399444 230382
rect 399392 230318 399444 230324
rect 399852 229764 399904 229770
rect 399852 229706 399904 229712
rect 398748 229628 398800 229634
rect 398748 229570 398800 229576
rect 399864 219434 399892 229706
rect 400048 228410 400076 231676
rect 400232 231662 400706 231690
rect 400968 231662 401350 231690
rect 400232 229094 400260 231662
rect 400232 229066 400352 229094
rect 400036 228404 400088 228410
rect 400036 228346 400088 228352
rect 400128 228132 400180 228138
rect 400128 228074 400180 228080
rect 400140 219434 400168 228074
rect 400324 221746 400352 229066
rect 400312 221740 400364 221746
rect 400312 221682 400364 221688
rect 400772 221604 400824 221610
rect 400772 221546 400824 221552
rect 399300 219428 399352 219434
rect 399864 219406 400076 219434
rect 400140 219428 400272 219434
rect 400140 219406 400220 219428
rect 399300 219370 399352 219376
rect 398104 219020 398156 219026
rect 398104 218962 398156 218968
rect 398472 218612 398524 218618
rect 398472 218554 398524 218560
rect 397644 218068 397696 218074
rect 397644 218010 397696 218016
rect 395126 217110 395200 217138
rect 395954 217246 396028 217274
rect 396782 217246 396856 217274
rect 395126 216988 395154 217110
rect 395954 216988 395982 217246
rect 396782 216988 396810 217246
rect 397656 217138 397684 218010
rect 398484 217138 398512 218554
rect 399312 217138 399340 219370
rect 400048 217274 400076 219406
rect 400220 219370 400272 219376
rect 400784 218074 400812 221546
rect 400968 220250 400996 231662
rect 401980 225622 402008 231676
rect 402624 227322 402652 231676
rect 402796 228404 402848 228410
rect 402796 228346 402848 228352
rect 402612 227316 402664 227322
rect 402612 227258 402664 227264
rect 402244 227180 402296 227186
rect 402244 227122 402296 227128
rect 401968 225616 402020 225622
rect 401968 225558 402020 225564
rect 400956 220244 401008 220250
rect 400956 220186 401008 220192
rect 401784 218204 401836 218210
rect 401784 218146 401836 218152
rect 400772 218068 400824 218074
rect 400772 218010 400824 218016
rect 400956 218068 401008 218074
rect 400956 218010 401008 218016
rect 400048 217246 400122 217274
rect 397610 217110 397684 217138
rect 398438 217110 398512 217138
rect 399266 217110 399340 217138
rect 397610 216988 397638 217110
rect 398438 216988 398466 217110
rect 399266 216988 399294 217110
rect 400094 216988 400122 217246
rect 400968 217138 400996 218010
rect 401796 217138 401824 218146
rect 402256 218074 402284 227122
rect 402612 218884 402664 218890
rect 402612 218826 402664 218832
rect 402244 218068 402296 218074
rect 402244 218010 402296 218016
rect 402624 217138 402652 218826
rect 402808 218210 402836 228346
rect 403268 225894 403296 231676
rect 403544 231662 403926 231690
rect 403544 227050 403572 231662
rect 403532 227044 403584 227050
rect 403532 226986 403584 226992
rect 403992 226500 404044 226506
rect 403992 226442 404044 226448
rect 403256 225888 403308 225894
rect 403256 225830 403308 225836
rect 402796 218204 402848 218210
rect 402796 218146 402848 218152
rect 404004 218074 404032 226442
rect 404176 225004 404228 225010
rect 404176 224946 404228 224952
rect 403440 218068 403492 218074
rect 403440 218010 403492 218016
rect 403992 218068 404044 218074
rect 403992 218010 404044 218016
rect 403452 217138 403480 218010
rect 404188 217274 404216 224946
rect 404556 224262 404584 231676
rect 404740 231662 405214 231690
rect 405752 231662 405858 231690
rect 404544 224256 404596 224262
rect 404544 224198 404596 224204
rect 404740 220114 404768 231662
rect 405556 224256 405608 224262
rect 405556 224198 405608 224204
rect 404728 220108 404780 220114
rect 404728 220050 404780 220056
rect 405568 218074 405596 224198
rect 405752 221610 405780 231662
rect 406488 222902 406516 231676
rect 407146 231662 407344 231690
rect 406752 223576 406804 223582
rect 406752 223518 406804 223524
rect 406476 222896 406528 222902
rect 406476 222838 406528 222844
rect 405740 221604 405792 221610
rect 405740 221546 405792 221552
rect 405924 219496 405976 219502
rect 405924 219438 405976 219444
rect 405096 218068 405148 218074
rect 405096 218010 405148 218016
rect 405556 218068 405608 218074
rect 405556 218010 405608 218016
rect 404188 217246 404262 217274
rect 400922 217110 400996 217138
rect 401750 217110 401824 217138
rect 402578 217110 402652 217138
rect 403406 217110 403480 217138
rect 400922 216988 400950 217110
rect 401750 216988 401778 217110
rect 402578 216988 402606 217110
rect 403406 216988 403434 217110
rect 404234 216988 404262 217246
rect 405108 217138 405136 218010
rect 405936 217274 405964 219438
rect 406764 217274 406792 223518
rect 407316 221474 407344 231662
rect 407776 228546 407804 231676
rect 407764 228540 407816 228546
rect 407764 228482 407816 228488
rect 408420 227186 408448 231676
rect 408696 231662 409078 231690
rect 408408 227180 408460 227186
rect 408408 227122 408460 227128
rect 408696 226370 408724 231662
rect 409708 229770 409736 231676
rect 409696 229764 409748 229770
rect 409696 229706 409748 229712
rect 409788 228540 409840 228546
rect 409788 228482 409840 228488
rect 409052 227792 409104 227798
rect 409052 227734 409104 227740
rect 407764 226364 407816 226370
rect 407764 226306 407816 226312
rect 408684 226364 408736 226370
rect 408684 226306 408736 226312
rect 407304 221468 407356 221474
rect 407304 221410 407356 221416
rect 407776 218618 407804 226306
rect 408408 221468 408460 221474
rect 408408 221410 408460 221416
rect 407764 218612 407816 218618
rect 407764 218554 407816 218560
rect 407580 218204 407632 218210
rect 407580 218146 407632 218152
rect 405062 217110 405136 217138
rect 405890 217246 405964 217274
rect 406718 217246 406792 217274
rect 405062 216988 405090 217110
rect 405890 216988 405918 217246
rect 406718 216988 406746 217246
rect 407592 217138 407620 218146
rect 408420 217274 408448 221410
rect 409064 218890 409092 227734
rect 409052 218884 409104 218890
rect 409052 218826 409104 218832
rect 409800 218074 409828 228482
rect 410352 227798 410380 231676
rect 410720 231662 411010 231690
rect 410720 229094 410748 231662
rect 410892 229764 410944 229770
rect 410892 229706 410944 229712
rect 410904 229094 410932 229706
rect 410628 229066 410748 229094
rect 410812 229066 410932 229094
rect 410340 227792 410392 227798
rect 410340 227734 410392 227740
rect 410628 225010 410656 229066
rect 410616 225004 410668 225010
rect 410616 224946 410668 224952
rect 410812 219434 410840 229066
rect 411640 228410 411668 231676
rect 411628 228404 411680 228410
rect 411628 228346 411680 228352
rect 411904 227792 411956 227798
rect 411904 227734 411956 227740
rect 410984 225616 411036 225622
rect 410984 225558 411036 225564
rect 410996 219434 411024 225558
rect 410720 219406 410840 219434
rect 410904 219406 411024 219434
rect 410720 218074 410748 219406
rect 409236 218068 409288 218074
rect 409236 218010 409288 218016
rect 409788 218068 409840 218074
rect 409788 218010 409840 218016
rect 410064 218068 410116 218074
rect 410064 218010 410116 218016
rect 410708 218068 410760 218074
rect 410708 218010 410760 218016
rect 407546 217110 407620 217138
rect 408374 217246 408448 217274
rect 407546 216988 407574 217110
rect 408374 216988 408402 217246
rect 409248 217138 409276 218010
rect 410076 217138 410104 218010
rect 410904 217274 410932 219406
rect 411720 218884 411772 218890
rect 411720 218826 411772 218832
rect 409202 217110 409276 217138
rect 410030 217110 410104 217138
rect 410858 217246 410932 217274
rect 409202 216988 409230 217110
rect 410030 216988 410058 217110
rect 410858 216988 410886 217246
rect 411732 217138 411760 218826
rect 411916 218210 411944 227734
rect 412284 226506 412312 231676
rect 412744 231662 412942 231690
rect 412548 227044 412600 227050
rect 412548 226986 412600 226992
rect 412272 226500 412324 226506
rect 412272 226442 412324 226448
rect 412560 218890 412588 226986
rect 412744 219502 412772 231662
rect 413572 227798 413600 231676
rect 413836 229356 413888 229362
rect 413836 229298 413888 229304
rect 413560 227792 413612 227798
rect 413560 227734 413612 227740
rect 412732 219496 412784 219502
rect 412732 219438 412784 219444
rect 412548 218884 412600 218890
rect 412548 218826 412600 218832
rect 412548 218748 412600 218754
rect 412548 218690 412600 218696
rect 411904 218204 411956 218210
rect 411904 218146 411956 218152
rect 412560 217138 412588 218690
rect 413848 218074 413876 229298
rect 414216 224262 414244 231676
rect 414204 224256 414256 224262
rect 414204 224198 414256 224204
rect 414860 223582 414888 231676
rect 415504 228546 415532 231676
rect 415492 228540 415544 228546
rect 415492 228482 415544 228488
rect 415032 228064 415084 228070
rect 415032 228006 415084 228012
rect 414848 223576 414900 223582
rect 414848 223518 414900 223524
rect 414204 220788 414256 220794
rect 414204 220730 414256 220736
rect 413376 218068 413428 218074
rect 413376 218010 413428 218016
rect 413836 218068 413888 218074
rect 413836 218010 413888 218016
rect 413388 217138 413416 218010
rect 414216 217274 414244 220730
rect 415044 217274 415072 228006
rect 416148 225622 416176 231676
rect 416792 229094 416820 231676
rect 417436 229770 417464 231676
rect 417712 231662 418094 231690
rect 418356 231662 418738 231690
rect 417424 229764 417476 229770
rect 417424 229706 417476 229712
rect 417712 229094 417740 231662
rect 416792 229066 416912 229094
rect 416688 227928 416740 227934
rect 416688 227870 416740 227876
rect 416136 225616 416188 225622
rect 416136 225558 416188 225564
rect 416504 225004 416556 225010
rect 416504 224946 416556 224952
rect 416516 219434 416544 224946
rect 416700 219434 416728 227870
rect 416884 221474 416912 229066
rect 417160 229066 417740 229094
rect 416872 221468 416924 221474
rect 416872 221410 416924 221416
rect 415860 219428 415912 219434
rect 416516 219406 416636 219434
rect 416700 219428 416832 219434
rect 416700 219406 416780 219428
rect 415860 219370 415912 219376
rect 411686 217110 411760 217138
rect 412514 217110 412588 217138
rect 413342 217110 413416 217138
rect 414170 217246 414244 217274
rect 414998 217246 415072 217274
rect 411686 216988 411714 217110
rect 412514 216988 412542 217110
rect 413342 216988 413370 217110
rect 414170 216988 414198 217246
rect 414998 216988 415026 217246
rect 415872 217138 415900 219370
rect 416608 217274 416636 219406
rect 416780 219370 416832 219376
rect 417160 218754 417188 229066
rect 418356 224954 418384 231662
rect 419368 227050 419396 231676
rect 420012 229362 420040 231676
rect 420000 229356 420052 229362
rect 420000 229298 420052 229304
rect 420656 227934 420684 231676
rect 421024 231662 421314 231690
rect 420644 227928 420696 227934
rect 420644 227870 420696 227876
rect 420644 227792 420696 227798
rect 420644 227734 420696 227740
rect 419356 227044 419408 227050
rect 419356 226986 419408 226992
rect 418172 224926 418384 224954
rect 418172 220794 418200 224926
rect 418344 220856 418396 220862
rect 418344 220798 418396 220804
rect 418160 220788 418212 220794
rect 418160 220730 418212 220736
rect 417516 219428 417568 219434
rect 417516 219370 417568 219376
rect 417148 218748 417200 218754
rect 417148 218690 417200 218696
rect 416608 217246 416682 217274
rect 415826 217110 415900 217138
rect 415826 216988 415854 217110
rect 416654 216988 416682 217246
rect 417528 217138 417556 219370
rect 418356 217274 418384 220798
rect 420656 219434 420684 227734
rect 420828 222896 420880 222902
rect 420828 222838 420880 222844
rect 420656 219406 420776 219434
rect 419172 219292 419224 219298
rect 419172 219234 419224 219240
rect 419184 217274 419212 219234
rect 420000 218068 420052 218074
rect 420000 218010 420052 218016
rect 417482 217110 417556 217138
rect 418310 217246 418384 217274
rect 419138 217246 419212 217274
rect 417482 216988 417510 217110
rect 418310 216988 418338 217246
rect 419138 216988 419166 217246
rect 420012 217138 420040 218010
rect 420748 217274 420776 219406
rect 420840 218090 420868 222838
rect 421024 219502 421052 231662
rect 421944 228070 421972 231676
rect 422312 231662 422602 231690
rect 422864 231662 423246 231690
rect 422312 229094 422340 231662
rect 422220 229066 422340 229094
rect 421932 228064 421984 228070
rect 421932 228006 421984 228012
rect 422220 225010 422248 229066
rect 422208 225004 422260 225010
rect 422208 224946 422260 224952
rect 421656 220108 421708 220114
rect 421656 220050 421708 220056
rect 421012 219496 421064 219502
rect 421012 219438 421064 219444
rect 420840 218074 420960 218090
rect 420840 218068 420972 218074
rect 420840 218062 420920 218068
rect 420920 218010 420972 218016
rect 421668 217274 421696 220050
rect 422864 219434 422892 231662
rect 423496 229152 423548 229158
rect 423496 229094 423548 229100
rect 423508 219434 423536 229094
rect 423876 227798 423904 231676
rect 424060 231662 424534 231690
rect 423864 227792 423916 227798
rect 423864 227734 423916 227740
rect 424060 220862 424088 231662
rect 425164 222902 425192 231676
rect 425440 231662 425822 231690
rect 425152 222896 425204 222902
rect 425152 222838 425204 222844
rect 424968 222148 425020 222154
rect 424968 222090 425020 222096
rect 424048 220856 424100 220862
rect 424048 220798 424100 220804
rect 422680 219406 422892 219434
rect 423324 219406 423536 219434
rect 422680 219298 422708 219406
rect 422668 219292 422720 219298
rect 422668 219234 422720 219240
rect 422484 218204 422536 218210
rect 422484 218146 422536 218152
rect 420748 217246 420822 217274
rect 419966 217110 420040 217138
rect 419966 216988 419994 217110
rect 420794 216988 420822 217246
rect 421622 217246 421696 217274
rect 421622 216988 421650 217246
rect 422496 217138 422524 218146
rect 423324 217274 423352 219406
rect 424140 218068 424192 218074
rect 424140 218010 424192 218016
rect 422450 217110 422524 217138
rect 423278 217246 423352 217274
rect 422450 216988 422478 217110
rect 423278 216988 423306 217246
rect 424152 217138 424180 218010
rect 424980 217274 425008 222090
rect 425440 218210 425468 231662
rect 426452 224330 426480 231676
rect 426820 231662 427110 231690
rect 426440 224324 426492 224330
rect 426440 224266 426492 224272
rect 426820 220114 426848 231662
rect 427740 229158 427768 231676
rect 427728 229152 427780 229158
rect 427728 229094 427780 229100
rect 428384 229094 428412 231676
rect 428752 231662 429042 231690
rect 429304 231662 429686 231690
rect 429948 231662 430330 231690
rect 430684 231662 430974 231690
rect 431236 231662 431618 231690
rect 432064 231662 432262 231690
rect 432708 231662 432906 231690
rect 428384 229066 428504 229094
rect 426992 224324 427044 224330
rect 426992 224266 427044 224272
rect 426808 220108 426860 220114
rect 426808 220050 426860 220056
rect 426624 218340 426676 218346
rect 426624 218282 426676 218288
rect 425428 218204 425480 218210
rect 425428 218146 425480 218152
rect 425796 218204 425848 218210
rect 425796 218146 425848 218152
rect 424106 217110 424180 217138
rect 424934 217246 425008 217274
rect 424106 216988 424134 217110
rect 424934 216988 424962 217246
rect 425808 217138 425836 218146
rect 426636 217138 426664 218282
rect 427004 218074 427032 224266
rect 427912 224256 427964 224262
rect 427912 224198 427964 224204
rect 427924 218074 427952 224198
rect 428280 219428 428332 219434
rect 428280 219370 428332 219376
rect 426992 218068 427044 218074
rect 426992 218010 427044 218016
rect 427452 218068 427504 218074
rect 427452 218010 427504 218016
rect 427912 218068 427964 218074
rect 427912 218010 427964 218016
rect 427464 217138 427492 218010
rect 428292 217138 428320 219370
rect 428476 218210 428504 229066
rect 428752 224262 428780 231662
rect 428740 224256 428792 224262
rect 428740 224198 428792 224204
rect 429304 222154 429332 231662
rect 429292 222148 429344 222154
rect 429292 222090 429344 222096
rect 429948 219434 429976 231662
rect 430684 219434 430712 231662
rect 431236 219434 431264 231662
rect 432064 219570 432092 231662
rect 432236 220244 432288 220250
rect 432236 220186 432288 220192
rect 432052 219564 432104 219570
rect 432052 219506 432104 219512
rect 432248 219434 432276 220186
rect 429580 219406 429976 219434
rect 430592 219406 430712 219434
rect 430776 219406 431264 219434
rect 431972 219406 432276 219434
rect 429580 218346 429608 219406
rect 429936 218612 429988 218618
rect 429936 218554 429988 218560
rect 429568 218340 429620 218346
rect 429568 218282 429620 218288
rect 428464 218204 428516 218210
rect 428464 218146 428516 218152
rect 429108 218068 429160 218074
rect 429108 218010 429160 218016
rect 429120 217138 429148 218010
rect 429948 217138 429976 218554
rect 430592 218074 430620 219406
rect 430580 218068 430632 218074
rect 430580 218010 430632 218016
rect 430776 217274 430804 219406
rect 431972 218090 432000 219406
rect 432708 218618 432736 231662
rect 433536 230602 433564 231676
rect 433536 230574 433656 230602
rect 433432 230444 433484 230450
rect 433432 230386 433484 230392
rect 433444 229094 433472 230386
rect 433628 229094 433656 230574
rect 434180 230450 434208 231676
rect 434168 230444 434220 230450
rect 434168 230386 434220 230392
rect 433444 229066 433564 229094
rect 433628 229066 433748 229094
rect 432696 218612 432748 218618
rect 432696 218554 432748 218560
rect 433248 218204 433300 218210
rect 433248 218146 433300 218152
rect 425762 217110 425836 217138
rect 426590 217110 426664 217138
rect 427418 217110 427492 217138
rect 428246 217110 428320 217138
rect 429074 217110 429148 217138
rect 429902 217110 429976 217138
rect 430730 217246 430804 217274
rect 431604 218062 432000 218090
rect 432420 218068 432472 218074
rect 425762 216988 425790 217110
rect 426590 216988 426618 217110
rect 427418 216988 427446 217110
rect 428246 216988 428274 217110
rect 429074 216988 429102 217110
rect 429902 216988 429930 217110
rect 430730 216988 430758 217246
rect 431604 217138 431632 218062
rect 432420 218010 432472 218016
rect 432432 217138 432460 218010
rect 433260 217138 433288 218146
rect 433536 217274 433564 229066
rect 433720 218074 433748 229066
rect 434824 220250 434852 231676
rect 435284 231662 435482 231690
rect 436126 231662 436324 231690
rect 434812 220244 434864 220250
rect 434812 220186 434864 220192
rect 434904 218340 434956 218346
rect 434904 218282 434956 218288
rect 433708 218068 433760 218074
rect 433708 218010 433760 218016
rect 433536 217246 434070 217274
rect 431558 217110 431632 217138
rect 432386 217110 432460 217138
rect 433214 217110 433288 217138
rect 431558 216988 431586 217110
rect 432386 216988 432414 217110
rect 433214 216988 433242 217110
rect 434042 216988 434070 217246
rect 434916 217138 434944 218282
rect 435284 218210 435312 231662
rect 436100 230376 436152 230382
rect 436100 230318 436152 230324
rect 435272 218204 435324 218210
rect 435272 218146 435324 218152
rect 435732 218068 435784 218074
rect 435732 218010 435784 218016
rect 435744 217138 435772 218010
rect 436112 217258 436140 230318
rect 436296 218074 436324 231662
rect 436756 230382 436784 231676
rect 436940 231662 437414 231690
rect 437584 231662 438058 231690
rect 436744 230376 436796 230382
rect 436744 230318 436796 230324
rect 436940 219434 436968 231662
rect 437584 219434 437612 231662
rect 438688 230382 438716 231676
rect 439332 230586 439360 231676
rect 439516 231662 439990 231690
rect 440344 231662 440634 231690
rect 439320 230580 439372 230586
rect 439320 230522 439372 230528
rect 439516 230466 439544 231662
rect 438964 230438 439544 230466
rect 438676 230376 438728 230382
rect 438676 230318 438728 230324
rect 438964 219434 438992 230438
rect 439320 230376 439372 230382
rect 439320 230318 439372 230324
rect 439332 219434 439360 230318
rect 436664 219406 436968 219434
rect 437492 219406 437612 219434
rect 438872 219406 438992 219434
rect 439056 219406 439360 219434
rect 436664 218346 436692 219406
rect 436652 218340 436704 218346
rect 436652 218282 436704 218288
rect 437492 218074 437520 219406
rect 438872 218074 438900 219406
rect 436284 218068 436336 218074
rect 436284 218010 436336 218016
rect 436560 218068 436612 218074
rect 436560 218010 436612 218016
rect 437480 218068 437532 218074
rect 437480 218010 437532 218016
rect 438216 218068 438268 218074
rect 438216 218010 438268 218016
rect 438860 218068 438912 218074
rect 438860 218010 438912 218016
rect 436100 217252 436152 217258
rect 436100 217194 436152 217200
rect 436572 217138 436600 218010
rect 437342 217252 437394 217258
rect 437342 217194 437394 217200
rect 434870 217110 434944 217138
rect 435698 217110 435772 217138
rect 436526 217110 436600 217138
rect 434870 216988 434898 217110
rect 435698 216988 435726 217110
rect 436526 216988 436554 217110
rect 437354 216988 437382 217194
rect 438228 217138 438256 218010
rect 439056 217274 439084 219406
rect 440344 218074 440372 231662
rect 440700 230444 440752 230450
rect 440700 230386 440752 230392
rect 439872 218068 439924 218074
rect 439872 218010 439924 218016
rect 440332 218068 440384 218074
rect 440332 218010 440384 218016
rect 438182 217110 438256 217138
rect 439010 217246 439084 217274
rect 438182 216988 438210 217110
rect 439010 216988 439038 217246
rect 439884 217138 439912 218010
rect 440712 217274 440740 230386
rect 441264 229158 441292 231676
rect 441908 230450 441936 231676
rect 442092 231662 442566 231690
rect 443104 231662 443210 231690
rect 441896 230444 441948 230450
rect 441896 230386 441948 230392
rect 442092 230330 442120 231662
rect 441724 230302 442120 230330
rect 441252 229152 441304 229158
rect 441252 229094 441304 229100
rect 441724 219434 441752 230302
rect 442080 229152 442132 229158
rect 442080 229094 442132 229100
rect 442092 229066 442304 229094
rect 441632 219406 441752 219434
rect 441632 218090 441660 219406
rect 439838 217110 439912 217138
rect 440666 217246 440740 217274
rect 441540 218062 441660 218090
rect 439838 216988 439866 217110
rect 440666 216988 440694 217246
rect 441540 217138 441568 218062
rect 442276 217274 442304 229066
rect 443104 217274 443132 231662
rect 443460 230444 443512 230450
rect 443460 230386 443512 230392
rect 443472 229094 443500 230386
rect 443840 230382 443868 231676
rect 443828 230376 443880 230382
rect 443828 230318 443880 230324
rect 444484 230246 444512 231676
rect 444668 231662 445142 231690
rect 444472 230240 444524 230246
rect 444472 230182 444524 230188
rect 444668 229094 444696 231662
rect 444932 230376 444984 230382
rect 444932 230318 444984 230324
rect 444944 229094 444972 230318
rect 445772 229094 445800 231676
rect 446416 229294 446444 231676
rect 446404 229288 446456 229294
rect 446404 229230 446456 229236
rect 443472 229066 443960 229094
rect 444668 229066 444788 229094
rect 444944 229066 445616 229094
rect 445772 229066 446444 229094
rect 443932 217274 443960 229066
rect 444760 217274 444788 229066
rect 445588 217274 445616 229066
rect 446416 217274 446444 229066
rect 447060 227934 447088 231676
rect 447244 231662 447718 231690
rect 447048 227928 447100 227934
rect 447048 227870 447100 227876
rect 447244 219434 447272 231662
rect 447600 230240 447652 230246
rect 447600 230182 447652 230188
rect 447612 219434 447640 230182
rect 448348 230042 448376 231676
rect 449006 231662 449296 231690
rect 448336 230036 448388 230042
rect 448336 229978 448388 229984
rect 448980 230036 449032 230042
rect 448980 229978 449032 229984
rect 448612 229288 448664 229294
rect 448612 229230 448664 229236
rect 448624 229094 448652 229230
rect 448992 229094 449020 229978
rect 449268 229566 449296 231662
rect 449636 229906 449664 231676
rect 449624 229900 449676 229906
rect 449624 229842 449676 229848
rect 449256 229560 449308 229566
rect 449256 229502 449308 229508
rect 450280 229294 450308 231676
rect 450544 229900 450596 229906
rect 450544 229842 450596 229848
rect 450268 229288 450320 229294
rect 450268 229230 450320 229236
rect 450556 229094 450584 229842
rect 450924 229158 450952 231676
rect 451568 230450 451596 231676
rect 452226 231662 452608 231690
rect 451556 230444 451608 230450
rect 451556 230386 451608 230392
rect 451924 229560 451976 229566
rect 451924 229502 451976 229508
rect 451740 229288 451792 229294
rect 451740 229230 451792 229236
rect 450912 229152 450964 229158
rect 450912 229094 450964 229100
rect 448624 229066 448928 229094
rect 448992 229066 449756 229094
rect 450556 229066 450768 229094
rect 447152 219406 447272 219434
rect 447336 219406 447640 219434
rect 442276 217246 442350 217274
rect 443104 217246 443178 217274
rect 443932 217246 444006 217274
rect 444760 217246 444834 217274
rect 445588 217246 445662 217274
rect 446416 217246 446490 217274
rect 447152 217258 447180 219406
rect 447336 217274 447364 219406
rect 441494 217110 441568 217138
rect 441494 216988 441522 217110
rect 442322 216988 442350 217246
rect 443150 216988 443178 217246
rect 443978 216988 444006 217246
rect 444806 216988 444834 217246
rect 445634 216988 445662 217246
rect 446462 216988 446490 217246
rect 447140 217252 447192 217258
rect 447140 217194 447192 217200
rect 447290 217246 447364 217274
rect 448900 217274 448928 229066
rect 449728 217274 449756 229066
rect 450544 227928 450596 227934
rect 450544 227870 450596 227876
rect 450556 217274 450584 227870
rect 450740 218346 450768 229066
rect 451752 219434 451780 229230
rect 451936 229094 451964 229502
rect 451936 229066 452240 229094
rect 451476 219406 451780 219434
rect 450728 218340 450780 218346
rect 450728 218282 450780 218288
rect 451476 217274 451504 219406
rect 448106 217252 448158 217258
rect 447290 216988 447318 217246
rect 448900 217246 448974 217274
rect 449728 217246 449802 217274
rect 450556 217246 450630 217274
rect 448106 217194 448158 217200
rect 448118 216988 448146 217194
rect 448946 216988 448974 217246
rect 449774 216988 449802 217246
rect 450602 216988 450630 217246
rect 451430 217246 451504 217274
rect 452212 217274 452240 229066
rect 452580 222154 452608 231662
rect 452856 230246 452884 231676
rect 453304 230444 453356 230450
rect 453304 230386 453356 230392
rect 452844 230240 452896 230246
rect 452844 230182 452896 230188
rect 452752 229152 452804 229158
rect 452752 229094 452804 229100
rect 452764 229066 453068 229094
rect 452568 222148 452620 222154
rect 452568 222090 452620 222096
rect 453040 217274 453068 229066
rect 453316 218074 453344 230386
rect 453500 229974 453528 231676
rect 454144 230110 454172 231676
rect 454316 230240 454368 230246
rect 454316 230182 454368 230188
rect 454132 230104 454184 230110
rect 454132 230046 454184 230052
rect 453488 229968 453540 229974
rect 453488 229910 453540 229916
rect 454328 229094 454356 230182
rect 454788 229094 454816 231676
rect 455432 230382 455460 231676
rect 455420 230376 455472 230382
rect 455420 230318 455472 230324
rect 455328 230104 455380 230110
rect 455328 230046 455380 230052
rect 454328 229066 454724 229094
rect 454788 229066 454908 229094
rect 453856 218340 453908 218346
rect 453856 218282 453908 218288
rect 453304 218068 453356 218074
rect 453304 218010 453356 218016
rect 452212 217246 452286 217274
rect 453040 217246 453114 217274
rect 451430 216988 451458 217246
rect 452258 216988 452286 217246
rect 453086 216988 453114 217246
rect 453868 217138 453896 218282
rect 454696 217274 454724 229066
rect 454880 223582 454908 229066
rect 454868 223576 454920 223582
rect 454868 223518 454920 223524
rect 455340 220794 455368 230046
rect 455788 229968 455840 229974
rect 455788 229910 455840 229916
rect 455604 222148 455656 222154
rect 455604 222090 455656 222096
rect 455328 220788 455380 220794
rect 455328 220730 455380 220736
rect 455616 218074 455644 222090
rect 455800 219434 455828 229910
rect 456076 224534 456104 231676
rect 456064 224528 456116 224534
rect 456064 224470 456116 224476
rect 456720 220930 456748 231676
rect 457168 230376 457220 230382
rect 457168 230318 457220 230324
rect 456708 220924 456760 220930
rect 456708 220866 456760 220872
rect 457180 219434 457208 230318
rect 457364 229770 457392 231676
rect 457352 229764 457404 229770
rect 457352 229706 457404 229712
rect 458008 229094 458036 231676
rect 458008 229066 458128 229094
rect 455800 219406 456380 219434
rect 457180 219406 458036 219434
rect 455420 218068 455472 218074
rect 455420 218010 455472 218016
rect 455604 218068 455656 218074
rect 455604 218010 455656 218016
rect 455432 217274 455460 218010
rect 456352 217274 456380 219406
rect 457168 218068 457220 218074
rect 457168 218010 457220 218016
rect 454696 217246 454770 217274
rect 455432 217246 455598 217274
rect 456352 217246 456426 217274
rect 453868 217110 453942 217138
rect 453914 216988 453942 217110
rect 454742 216988 454770 217246
rect 455570 216988 455598 217246
rect 456398 216988 456426 217246
rect 457180 217138 457208 218010
rect 458008 217274 458036 219406
rect 458100 218498 458128 229066
rect 458652 226302 458680 231676
rect 459310 231662 459508 231690
rect 458640 226296 458692 226302
rect 458640 226238 458692 226244
rect 458824 220788 458876 220794
rect 458824 220730 458876 220736
rect 458100 218470 458220 218498
rect 458192 218414 458220 218470
rect 458180 218408 458232 218414
rect 458180 218350 458232 218356
rect 458836 217274 458864 220730
rect 459480 220250 459508 231662
rect 459744 224528 459796 224534
rect 459744 224470 459796 224476
rect 459468 220244 459520 220250
rect 459468 220186 459520 220192
rect 459756 217274 459784 224470
rect 459940 222902 459968 231676
rect 460584 224942 460612 231676
rect 461242 231662 461716 231690
rect 461886 231662 462176 231690
rect 461688 229094 461716 231662
rect 461688 229066 461992 229094
rect 460572 224936 460624 224942
rect 460572 224878 460624 224884
rect 460480 223576 460532 223582
rect 460480 223518 460532 223524
rect 459928 222896 459980 222902
rect 459928 222838 459980 222844
rect 458008 217246 458082 217274
rect 458836 217246 458910 217274
rect 457180 217110 457254 217138
rect 457226 216988 457254 217110
rect 458054 216988 458082 217246
rect 458882 216988 458910 217246
rect 459710 217246 459784 217274
rect 460492 217274 460520 223518
rect 461308 218340 461360 218346
rect 461308 218282 461360 218288
rect 460492 217246 460566 217274
rect 459710 216988 459738 217246
rect 460538 216988 460566 217246
rect 461320 217138 461348 218282
rect 461964 218210 461992 229066
rect 462148 222154 462176 231662
rect 462516 224806 462544 231676
rect 462964 226296 463016 226302
rect 462964 226238 463016 226244
rect 462504 224800 462556 224806
rect 462504 224742 462556 224748
rect 462136 222148 462188 222154
rect 462136 222090 462188 222096
rect 462136 220856 462188 220862
rect 462136 220798 462188 220804
rect 461952 218204 462004 218210
rect 461952 218146 462004 218152
rect 462148 217274 462176 220798
rect 462976 217274 463004 226238
rect 463160 225418 463188 231676
rect 463804 230382 463832 231676
rect 464462 231662 465028 231690
rect 465106 231662 465488 231690
rect 465750 231662 465948 231690
rect 463792 230376 463844 230382
rect 463792 230318 463844 230324
rect 463884 229764 463936 229770
rect 463884 229706 463936 229712
rect 463148 225412 463200 225418
rect 463148 225354 463200 225360
rect 463148 224936 463200 224942
rect 463148 224878 463200 224884
rect 463160 218074 463188 224878
rect 463148 218068 463200 218074
rect 463148 218010 463200 218016
rect 463896 217274 463924 229706
rect 465000 219638 465028 231662
rect 465460 229770 465488 231662
rect 465724 230376 465776 230382
rect 465724 230318 465776 230324
rect 465448 229764 465500 229770
rect 465448 229706 465500 229712
rect 465736 220794 465764 230318
rect 465920 227662 465948 231662
rect 466104 231662 466394 231690
rect 465908 227656 465960 227662
rect 465908 227598 465960 227604
rect 466104 220930 466132 231662
rect 467024 229906 467052 231676
rect 467012 229900 467064 229906
rect 467012 229842 467064 229848
rect 467472 229764 467524 229770
rect 467472 229706 467524 229712
rect 467288 225412 467340 225418
rect 467288 225354 467340 225360
rect 467104 222896 467156 222902
rect 467104 222838 467156 222844
rect 466092 220924 466144 220930
rect 466092 220866 466144 220872
rect 465724 220788 465776 220794
rect 465724 220730 465776 220736
rect 465448 220244 465500 220250
rect 465448 220186 465500 220192
rect 464988 219632 465040 219638
rect 464988 219574 465040 219580
rect 464620 218068 464672 218074
rect 464620 218010 464672 218016
rect 462148 217246 462222 217274
rect 462976 217246 463050 217274
rect 461320 217110 461394 217138
rect 461366 216988 461394 217110
rect 462194 216988 462222 217246
rect 463022 216988 463050 217246
rect 463850 217246 463924 217274
rect 463850 216988 463878 217246
rect 464632 217138 464660 218010
rect 465460 217274 465488 220186
rect 466276 218204 466328 218210
rect 466276 218146 466328 218152
rect 465460 217246 465534 217274
rect 464632 217110 464706 217138
rect 464678 216988 464706 217110
rect 465506 216988 465534 217246
rect 466288 217138 466316 218146
rect 467116 217274 467144 222838
rect 467300 218074 467328 225354
rect 467484 222902 467512 229706
rect 467668 225622 467696 231676
rect 468312 230246 468340 231676
rect 468300 230240 468352 230246
rect 468300 230182 468352 230188
rect 467656 225616 467708 225622
rect 467656 225558 467708 225564
rect 467472 222896 467524 222902
rect 467472 222838 467524 222844
rect 468760 222148 468812 222154
rect 468760 222090 468812 222096
rect 467288 218068 467340 218074
rect 467288 218010 467340 218016
rect 467932 218068 467984 218074
rect 467932 218010 467984 218016
rect 467116 217246 467190 217274
rect 466288 217110 466362 217138
rect 466334 216988 466362 217110
rect 467162 216988 467190 217246
rect 467944 217138 467972 218010
rect 468772 217274 468800 222090
rect 468956 221474 468984 231676
rect 469128 230240 469180 230246
rect 469128 230182 469180 230188
rect 468944 221468 468996 221474
rect 468944 221410 468996 221416
rect 469140 220522 469168 230182
rect 469600 229770 469628 231676
rect 469588 229764 469640 229770
rect 469588 229706 469640 229712
rect 469864 227656 469916 227662
rect 469864 227598 469916 227604
rect 469312 224800 469364 224806
rect 469312 224742 469364 224748
rect 469128 220516 469180 220522
rect 469128 220458 469180 220464
rect 468772 217246 468846 217274
rect 469324 217258 469352 224742
rect 469588 220788 469640 220794
rect 469588 220730 469640 220736
rect 469600 217274 469628 220730
rect 469876 218618 469904 227598
rect 470244 224262 470272 231676
rect 470888 230382 470916 231676
rect 470876 230376 470928 230382
rect 470876 230318 470928 230324
rect 471532 227798 471560 231676
rect 471888 230376 471940 230382
rect 471888 230318 471940 230324
rect 471520 227792 471572 227798
rect 471520 227734 471572 227740
rect 470232 224256 470284 224262
rect 470232 224198 470284 224204
rect 471900 222154 471928 230318
rect 472176 229362 472204 231676
rect 472834 231662 473216 231690
rect 472164 229356 472216 229362
rect 472164 229298 472216 229304
rect 472992 229356 473044 229362
rect 472992 229298 473044 229304
rect 471888 222148 471940 222154
rect 471888 222090 471940 222096
rect 471428 220924 471480 220930
rect 471428 220866 471480 220872
rect 469864 218612 469916 218618
rect 469864 218554 469916 218560
rect 471244 218612 471296 218618
rect 471244 218554 471296 218560
rect 467944 217110 468018 217138
rect 467990 216988 468018 217110
rect 468818 216988 468846 217246
rect 469312 217252 469364 217258
rect 469600 217246 469674 217274
rect 469312 217194 469364 217200
rect 469646 216988 469674 217246
rect 470462 217252 470514 217258
rect 470462 217194 470514 217200
rect 470474 216988 470502 217194
rect 471256 217138 471284 218554
rect 471440 218074 471468 220866
rect 473004 220386 473032 229298
rect 472992 220380 473044 220386
rect 472992 220322 473044 220328
rect 473188 220250 473216 231662
rect 473464 223582 473492 231676
rect 474122 231662 474504 231690
rect 474004 229900 474056 229906
rect 474004 229842 474056 229848
rect 473452 223576 473504 223582
rect 473452 223518 473504 223524
rect 473728 222896 473780 222902
rect 473728 222838 473780 222844
rect 473176 220244 473228 220250
rect 473176 220186 473228 220192
rect 472072 219632 472124 219638
rect 472072 219574 472124 219580
rect 471428 218068 471480 218074
rect 471428 218010 471480 218016
rect 472084 217274 472112 219574
rect 472900 218068 472952 218074
rect 472900 218010 472952 218016
rect 472084 217246 472158 217274
rect 471256 217110 471330 217138
rect 471302 216988 471330 217110
rect 472130 216988 472158 217246
rect 472912 217138 472940 218010
rect 473740 217274 473768 222838
rect 474016 220794 474044 229842
rect 474476 228410 474504 231662
rect 474464 228404 474516 228410
rect 474464 228346 474516 228352
rect 474752 226506 474780 231676
rect 475410 231662 475884 231690
rect 474740 226500 474792 226506
rect 474740 226442 474792 226448
rect 475568 223576 475620 223582
rect 475568 223518 475620 223524
rect 474004 220788 474056 220794
rect 474004 220730 474056 220736
rect 475384 220788 475436 220794
rect 475384 220730 475436 220736
rect 474556 220516 474608 220522
rect 474556 220458 474608 220464
rect 474568 217274 474596 220458
rect 475396 217274 475424 220730
rect 475580 218618 475608 223518
rect 475856 221746 475884 231662
rect 476040 230382 476068 231676
rect 476028 230376 476080 230382
rect 476028 230318 476080 230324
rect 476684 229906 476712 231676
rect 476672 229900 476724 229906
rect 476672 229842 476724 229848
rect 476764 229764 476816 229770
rect 476764 229706 476816 229712
rect 476580 225616 476632 225622
rect 476580 225558 476632 225564
rect 475844 221740 475896 221746
rect 475844 221682 475896 221688
rect 476212 221468 476264 221474
rect 476212 221410 476264 221416
rect 475568 218612 475620 218618
rect 475568 218554 475620 218560
rect 476224 217274 476252 221410
rect 476592 217274 476620 225558
rect 476776 220794 476804 229706
rect 477328 225622 477356 231676
rect 477986 231662 478368 231690
rect 478630 231662 478828 231690
rect 477316 225616 477368 225622
rect 477316 225558 477368 225564
rect 477868 222148 477920 222154
rect 477868 222090 477920 222096
rect 476764 220788 476816 220794
rect 476764 220730 476816 220736
rect 477880 217274 477908 222090
rect 478340 220114 478368 231662
rect 478604 230376 478656 230382
rect 478604 230318 478656 230324
rect 478616 227186 478644 230318
rect 478800 229094 478828 231662
rect 479260 229770 479288 231676
rect 479248 229764 479300 229770
rect 479248 229706 479300 229712
rect 478800 229066 478920 229094
rect 478892 228818 478920 229066
rect 478880 228812 478932 228818
rect 478880 228754 478932 228760
rect 479524 227792 479576 227798
rect 479524 227734 479576 227740
rect 478604 227180 478656 227186
rect 478604 227122 478656 227128
rect 478696 220788 478748 220794
rect 478696 220730 478748 220736
rect 478328 220108 478380 220114
rect 478328 220050 478380 220056
rect 478708 217274 478736 220730
rect 479536 217274 479564 227734
rect 479904 222902 479932 231676
rect 480548 224398 480576 231676
rect 480824 231662 481206 231690
rect 480536 224392 480588 224398
rect 480536 224334 480588 224340
rect 480444 224256 480496 224262
rect 480444 224198 480496 224204
rect 479892 222896 479944 222902
rect 479892 222838 479944 222844
rect 480456 217274 480484 224198
rect 480824 221610 480852 231662
rect 481836 229906 481864 231676
rect 482494 231662 482968 231690
rect 481640 229900 481692 229906
rect 481640 229842 481692 229848
rect 481824 229900 481876 229906
rect 481824 229842 481876 229848
rect 481652 226370 481680 229842
rect 482744 226500 482796 226506
rect 482744 226442 482796 226448
rect 481640 226364 481692 226370
rect 481640 226306 481692 226312
rect 482756 222766 482784 226442
rect 482744 222760 482796 222766
rect 482744 222702 482796 222708
rect 480812 221604 480864 221610
rect 480812 221546 480864 221552
rect 481180 220380 481232 220386
rect 481180 220322 481232 220328
rect 473740 217246 473814 217274
rect 474568 217246 474642 217274
rect 475396 217246 475470 217274
rect 476224 217246 476298 217274
rect 476592 217246 477126 217274
rect 477880 217246 477954 217274
rect 478708 217246 478782 217274
rect 479536 217246 479610 217274
rect 472912 217110 472986 217138
rect 472958 216988 472986 217110
rect 473786 216988 473814 217246
rect 474614 216988 474642 217246
rect 475442 216988 475470 217246
rect 476270 216988 476298 217246
rect 477098 216988 477126 217246
rect 477926 216988 477954 217246
rect 478754 216988 478782 217246
rect 479582 216988 479610 217246
rect 480410 217246 480484 217274
rect 481192 217274 481220 220322
rect 482008 220244 482060 220250
rect 482008 220186 482060 220192
rect 482020 217274 482048 220186
rect 482756 218754 482784 222702
rect 482940 220250 482968 231662
rect 483124 223310 483152 231676
rect 483768 225894 483796 231676
rect 484412 230042 484440 231676
rect 484400 230036 484452 230042
rect 484400 229978 484452 229984
rect 485056 228546 485084 231676
rect 485700 228682 485728 231676
rect 486358 231662 486648 231690
rect 485688 228676 485740 228682
rect 485688 228618 485740 228624
rect 485044 228540 485096 228546
rect 485044 228482 485096 228488
rect 484492 228404 484544 228410
rect 484492 228346 484544 228352
rect 483756 225888 483808 225894
rect 483756 225830 483808 225836
rect 483112 223304 483164 223310
rect 483112 223246 483164 223252
rect 484504 222358 484532 228346
rect 486620 224262 486648 231662
rect 486792 227180 486844 227186
rect 486792 227122 486844 227128
rect 486804 224954 486832 227122
rect 486988 227050 487016 231676
rect 487632 230246 487660 231676
rect 488290 231662 488488 231690
rect 488460 230330 488488 231662
rect 488460 230302 488672 230330
rect 487620 230240 487672 230246
rect 487620 230182 487672 230188
rect 488448 230240 488500 230246
rect 488448 230182 488500 230188
rect 486976 227044 487028 227050
rect 486976 226986 487028 226992
rect 487804 226364 487856 226370
rect 487804 226306 487856 226312
rect 486804 224926 487016 224954
rect 486608 224256 486660 224262
rect 486608 224198 486660 224204
rect 484492 222352 484544 222358
rect 484492 222294 484544 222300
rect 483756 221468 483808 221474
rect 483756 221410 483808 221416
rect 482928 220244 482980 220250
rect 482928 220186 482980 220192
rect 482744 218748 482796 218754
rect 482744 218690 482796 218696
rect 482836 218612 482888 218618
rect 482836 218554 482888 218560
rect 481192 217246 481266 217274
rect 482020 217246 482094 217274
rect 480410 216988 480438 217246
rect 481238 216988 481266 217246
rect 482066 216988 482094 217246
rect 482848 217138 482876 218554
rect 483768 217274 483796 221410
rect 483722 217246 483796 217274
rect 484504 217274 484532 222294
rect 486148 221740 486200 221746
rect 486148 221682 486200 221688
rect 485320 218748 485372 218754
rect 485320 218690 485372 218696
rect 484504 217246 484578 217274
rect 482848 217110 482922 217138
rect 482894 216988 482922 217110
rect 483722 216988 483750 217246
rect 484550 216988 484578 217246
rect 485332 217138 485360 218690
rect 486160 217138 486188 221682
rect 486988 220289 487016 224926
rect 486974 220280 487030 220289
rect 486974 220215 487030 220224
rect 486988 217274 487016 220215
rect 487816 218113 487844 226306
rect 488460 220522 488488 230182
rect 488644 223174 488672 230302
rect 488920 225758 488948 231676
rect 489564 227186 489592 231676
rect 489920 229764 489972 229770
rect 489920 229706 489972 229712
rect 489552 227180 489604 227186
rect 489552 227122 489604 227128
rect 488908 225752 488960 225758
rect 488908 225694 488960 225700
rect 488816 225616 488868 225622
rect 488816 225558 488868 225564
rect 488632 223168 488684 223174
rect 488632 223110 488684 223116
rect 488448 220516 488500 220522
rect 488448 220458 488500 220464
rect 487802 218104 487858 218113
rect 487802 218039 487858 218048
rect 487816 217274 487844 218039
rect 488828 217274 488856 225558
rect 489932 222494 489960 229706
rect 490208 228410 490236 231676
rect 490866 231662 491248 231690
rect 491220 229094 491248 231662
rect 491496 230110 491524 231676
rect 491484 230104 491536 230110
rect 491484 230046 491536 230052
rect 492140 229770 492168 231676
rect 492798 231662 493088 231690
rect 492496 230104 492548 230110
rect 492496 230046 492548 230052
rect 492128 229764 492180 229770
rect 492128 229706 492180 229712
rect 491220 229066 491340 229094
rect 490380 228812 490432 228818
rect 490380 228754 490432 228760
rect 490196 228404 490248 228410
rect 490196 228346 490248 228352
rect 489920 222488 489972 222494
rect 489920 222430 489972 222436
rect 489460 220108 489512 220114
rect 489460 220050 489512 220056
rect 486988 217246 487062 217274
rect 487816 217246 487890 217274
rect 485332 217110 485406 217138
rect 486160 217110 486234 217138
rect 485378 216988 485406 217110
rect 486206 216988 486234 217110
rect 487034 216988 487062 217246
rect 487862 216988 487890 217246
rect 488690 217246 488856 217274
rect 488690 216988 488718 217246
rect 488828 217161 488856 217246
rect 488814 217152 488870 217161
rect 489472 217138 489500 220050
rect 490392 218074 490420 228754
rect 491312 224534 491340 229066
rect 491300 224528 491352 224534
rect 491300 224470 491352 224476
rect 491944 222896 491996 222902
rect 491944 222838 491996 222844
rect 491116 222488 491168 222494
rect 491116 222430 491168 222436
rect 490380 218068 490432 218074
rect 490380 218010 490432 218016
rect 490392 217274 490420 218010
rect 490346 217246 490420 217274
rect 489472 217110 489546 217138
rect 488814 217087 488870 217096
rect 489518 216988 489546 217110
rect 490346 216988 490374 217246
rect 491128 217138 491156 222430
rect 491956 218210 491984 222838
rect 492508 220114 492536 230046
rect 492772 224392 492824 224398
rect 492772 224334 492824 224340
rect 492496 220108 492548 220114
rect 492496 220050 492548 220056
rect 491944 218204 491996 218210
rect 491944 218146 491996 218152
rect 491956 217138 491984 218146
rect 492784 217138 492812 224334
rect 493060 223038 493088 231662
rect 493428 230382 493456 231676
rect 493416 230376 493468 230382
rect 493416 230318 493468 230324
rect 493600 229900 493652 229906
rect 493600 229842 493652 229848
rect 493612 225010 493640 229842
rect 494072 225622 494100 231676
rect 494716 227322 494744 231676
rect 495164 230240 495216 230246
rect 495164 230182 495216 230188
rect 494704 227316 494756 227322
rect 494704 227258 494756 227264
rect 494060 225616 494112 225622
rect 494060 225558 494112 225564
rect 495176 225010 495204 230182
rect 495360 229294 495388 231676
rect 496004 229906 496032 231676
rect 496188 231662 496662 231690
rect 495992 229900 496044 229906
rect 495992 229842 496044 229848
rect 495348 229288 495400 229294
rect 495348 229230 495400 229236
rect 496188 229094 496216 231662
rect 497292 230382 497320 231676
rect 497476 231662 497950 231690
rect 496360 230376 496412 230382
rect 496360 230318 496412 230324
rect 497280 230376 497332 230382
rect 497280 230318 497332 230324
rect 496372 229094 496400 230318
rect 496188 229066 496308 229094
rect 496372 229066 496492 229094
rect 493600 225004 493652 225010
rect 493600 224946 493652 224952
rect 494704 225004 494756 225010
rect 494704 224946 494756 224952
rect 495164 225004 495216 225010
rect 495164 224946 495216 224952
rect 493048 223032 493100 223038
rect 493048 222974 493100 222980
rect 492956 221604 493008 221610
rect 492956 221546 493008 221552
rect 492968 219745 492996 221546
rect 492954 219736 493010 219745
rect 492954 219671 493010 219680
rect 493690 219736 493746 219745
rect 493690 219671 493746 219680
rect 493704 217138 493732 219671
rect 494716 218385 494744 224946
rect 495176 222086 495204 224946
rect 496084 223304 496136 223310
rect 496084 223246 496136 223252
rect 495164 222080 495216 222086
rect 495164 222022 495216 222028
rect 495256 220244 495308 220250
rect 495256 220186 495308 220192
rect 494702 218376 494758 218385
rect 494532 218334 494702 218362
rect 494532 217274 494560 218334
rect 494702 218311 494758 218320
rect 495268 217274 495296 220186
rect 496096 217274 496124 223246
rect 496280 221746 496308 229066
rect 496268 221740 496320 221746
rect 496268 221682 496320 221688
rect 496464 220386 496492 229066
rect 497280 225888 497332 225894
rect 497280 225830 497332 225836
rect 496452 220380 496504 220386
rect 496452 220322 496504 220328
rect 497292 219434 497320 225830
rect 497476 221610 497504 231662
rect 498108 230376 498160 230382
rect 498108 230318 498160 230324
rect 498120 226030 498148 230318
rect 498580 228682 498608 231676
rect 498292 228676 498344 228682
rect 498292 228618 498344 228624
rect 498568 228676 498620 228682
rect 498568 228618 498620 228624
rect 498108 226024 498160 226030
rect 498108 225966 498160 225972
rect 497740 222080 497792 222086
rect 497740 222022 497792 222028
rect 497464 221604 497516 221610
rect 497464 221546 497516 221552
rect 497292 219406 497504 219434
rect 497476 218346 497504 219406
rect 497464 218340 497516 218346
rect 497464 218282 497516 218288
rect 497476 218074 497504 218282
rect 497004 218068 497056 218074
rect 497004 218010 497056 218016
rect 497464 218068 497516 218074
rect 497464 218010 497516 218016
rect 497016 217274 497044 218010
rect 491128 217110 491202 217138
rect 491956 217110 492030 217138
rect 492784 217110 492858 217138
rect 491174 216988 491202 217110
rect 492002 216988 492030 217110
rect 492830 216988 492858 217110
rect 493658 217110 493732 217138
rect 494486 217246 494560 217274
rect 495176 217246 495342 217274
rect 496096 217246 496170 217274
rect 493658 216988 493686 217110
rect 494486 216988 494514 217246
rect 495176 217161 495204 217246
rect 495162 217152 495218 217161
rect 495162 217087 495218 217096
rect 495314 216988 495342 217246
rect 496142 216988 496170 217246
rect 496970 217246 497044 217274
rect 497752 217274 497780 222022
rect 498304 219434 498332 228618
rect 498660 228540 498712 228546
rect 498660 228482 498712 228488
rect 498212 219406 498332 219434
rect 497752 217246 497826 217274
rect 498212 217258 498240 219406
rect 498672 217274 498700 228482
rect 499224 224398 499252 231676
rect 499868 228818 499896 231676
rect 500526 231662 500816 231690
rect 500224 229288 500276 229294
rect 500224 229230 500276 229236
rect 499856 228812 499908 228818
rect 499856 228754 499908 228760
rect 499212 224392 499264 224398
rect 499212 224334 499264 224340
rect 500236 220658 500264 229230
rect 500408 224256 500460 224262
rect 500408 224198 500460 224204
rect 500224 220652 500276 220658
rect 500224 220594 500276 220600
rect 500420 218754 500448 224198
rect 500788 222902 500816 231662
rect 500960 227044 501012 227050
rect 500960 226986 501012 226992
rect 500776 222896 500828 222902
rect 500776 222838 500828 222844
rect 500972 220368 501000 226986
rect 501156 225894 501184 231676
rect 501340 231662 501814 231690
rect 501144 225888 501196 225894
rect 501144 225830 501196 225836
rect 500972 220340 501184 220368
rect 501156 219570 501184 220340
rect 501340 220250 501368 231662
rect 502444 228546 502472 231676
rect 503102 231662 503392 231690
rect 502432 228540 502484 228546
rect 502432 228482 502484 228488
rect 503364 223310 503392 231662
rect 503732 229158 503760 231676
rect 503720 229152 503772 229158
rect 503720 229094 503772 229100
rect 504180 227180 504232 227186
rect 504180 227122 504232 227128
rect 503628 225752 503680 225758
rect 503628 225694 503680 225700
rect 503352 223304 503404 223310
rect 503352 223246 503404 223252
rect 503168 223168 503220 223174
rect 503168 223110 503220 223116
rect 501880 220516 501932 220522
rect 501880 220458 501932 220464
rect 501328 220244 501380 220250
rect 501328 220186 501380 220192
rect 501144 219564 501196 219570
rect 501144 219506 501196 219512
rect 500408 218748 500460 218754
rect 500408 218690 500460 218696
rect 500420 217274 500448 218690
rect 501156 217274 501184 219506
rect 496970 216988 496998 217246
rect 497798 216988 497826 217246
rect 498200 217252 498252 217258
rect 498200 217194 498252 217200
rect 498626 217246 498700 217274
rect 499442 217252 499494 217258
rect 498626 217122 498654 217246
rect 499442 217194 499494 217200
rect 500282 217246 500448 217274
rect 501110 217246 501184 217274
rect 501892 217274 501920 220458
rect 503180 218482 503208 223110
rect 503640 219910 503668 225694
rect 503628 219904 503680 219910
rect 503628 219846 503680 219852
rect 502800 218476 502852 218482
rect 502800 218418 502852 218424
rect 503168 218476 503220 218482
rect 503168 218418 503220 218424
rect 502248 218204 502300 218210
rect 502248 218146 502300 218152
rect 502260 217297 502288 218146
rect 502246 217288 502302 217297
rect 501892 217246 501966 217274
rect 498614 217116 498666 217122
rect 498614 217058 498666 217064
rect 498626 216988 498654 217058
rect 499454 216988 499482 217194
rect 500282 216988 500310 217246
rect 501110 216988 501138 217246
rect 501938 216988 501966 217246
rect 502246 217223 502302 217232
rect 502812 217138 502840 218418
rect 503640 217274 503668 219846
rect 504192 219434 504220 227122
rect 504376 224262 504404 231676
rect 505020 227050 505048 231676
rect 505664 229294 505692 231676
rect 506216 231662 506322 231690
rect 505652 229288 505704 229294
rect 505652 229230 505704 229236
rect 505192 228404 505244 228410
rect 505192 228346 505244 228352
rect 505008 227044 505060 227050
rect 505008 226986 505060 226992
rect 505204 224670 505232 228346
rect 506216 227186 506244 231662
rect 506388 229900 506440 229906
rect 506388 229842 506440 229848
rect 506400 228954 506428 229842
rect 506388 228948 506440 228954
rect 506388 228890 506440 228896
rect 506204 227180 506256 227186
rect 506204 227122 506256 227128
rect 506952 224806 506980 231676
rect 507596 229906 507624 231676
rect 507584 229900 507636 229906
rect 507584 229842 507636 229848
rect 507124 229764 507176 229770
rect 507124 229706 507176 229712
rect 506940 224800 506992 224806
rect 506940 224742 506992 224748
rect 505192 224664 505244 224670
rect 505192 224606 505244 224612
rect 504364 224256 504416 224262
rect 504364 224198 504416 224204
rect 504364 222488 504416 222494
rect 504364 222430 504416 222436
rect 504376 222222 504404 222430
rect 504364 222216 504416 222222
rect 504364 222158 504416 222164
rect 504192 219406 504404 219434
rect 502766 217110 502840 217138
rect 503594 217246 503668 217274
rect 504376 217274 504404 219406
rect 505204 217274 505232 224606
rect 506112 224528 506164 224534
rect 506112 224470 506164 224476
rect 506124 217326 506152 224470
rect 506848 220108 506900 220114
rect 506848 220050 506900 220056
rect 506112 217320 506164 217326
rect 504376 217246 504450 217274
rect 505204 217246 505278 217274
rect 506112 217262 506164 217268
rect 506860 217274 506888 220050
rect 507136 218210 507164 229706
rect 508240 223174 508268 231676
rect 508884 225758 508912 231676
rect 509528 229702 509556 231676
rect 509516 229696 509568 229702
rect 509516 229638 509568 229644
rect 509884 229152 509936 229158
rect 509884 229094 509936 229100
rect 508872 225752 508924 225758
rect 508872 225694 508924 225700
rect 509700 225616 509752 225622
rect 509700 225558 509752 225564
rect 509712 223922 509740 225558
rect 509700 223916 509752 223922
rect 509700 223858 509752 223864
rect 508228 223168 508280 223174
rect 508228 223110 508280 223116
rect 508504 223032 508556 223038
rect 508504 222974 508556 222980
rect 508044 218748 508096 218754
rect 508044 218690 508096 218696
rect 507676 218612 507728 218618
rect 507676 218554 507728 218560
rect 507688 218210 507716 218554
rect 508056 218482 508084 218690
rect 507860 218476 507912 218482
rect 507860 218418 507912 218424
rect 508044 218476 508096 218482
rect 508044 218418 508096 218424
rect 507872 218210 507900 218418
rect 507124 218204 507176 218210
rect 507124 218146 507176 218152
rect 507676 218204 507728 218210
rect 507676 218146 507728 218152
rect 507860 218204 507912 218210
rect 507860 218146 507912 218152
rect 502766 216988 502794 217110
rect 503594 216988 503622 217246
rect 504422 216988 504450 217246
rect 505250 216988 505278 217246
rect 506124 217138 506152 217262
rect 506860 217246 506934 217274
rect 506078 217110 506152 217138
rect 506078 216988 506106 217110
rect 506906 216988 506934 217246
rect 507688 217138 507716 218146
rect 508516 217274 508544 222974
rect 509896 221882 509924 229094
rect 510172 225622 510200 231676
rect 510816 230382 510844 231676
rect 510804 230376 510856 230382
rect 510804 230318 510856 230324
rect 511460 230246 511488 231676
rect 511908 230376 511960 230382
rect 511908 230318 511960 230324
rect 511448 230240 511500 230246
rect 511448 230182 511500 230188
rect 510620 229288 510672 229294
rect 510620 229230 510672 229236
rect 510632 227322 510660 229230
rect 511920 229094 511948 230318
rect 511828 229066 511948 229094
rect 510620 227316 510672 227322
rect 510620 227258 510672 227264
rect 510988 226908 511040 226914
rect 510988 226850 511040 226856
rect 510160 225616 510212 225622
rect 510160 225558 510212 225564
rect 510160 223916 510212 223922
rect 510160 223858 510212 223864
rect 509884 221876 509936 221882
rect 509884 221818 509936 221824
rect 509332 220380 509384 220386
rect 509332 220322 509384 220328
rect 509344 217274 509372 220322
rect 510172 217274 510200 223858
rect 511000 217569 511028 226850
rect 511828 220794 511856 229066
rect 512104 228410 512132 231676
rect 512762 231662 513144 231690
rect 512736 228948 512788 228954
rect 512736 228890 512788 228896
rect 512092 228404 512144 228410
rect 512092 228346 512144 228352
rect 511816 220788 511868 220794
rect 511816 220730 511868 220736
rect 511816 220652 511868 220658
rect 511816 220594 511868 220600
rect 510986 217560 511042 217569
rect 510986 217495 511042 217504
rect 508516 217246 508590 217274
rect 509344 217246 509418 217274
rect 510172 217246 510246 217274
rect 508562 217190 508590 217246
rect 508550 217184 508602 217190
rect 507688 217110 507762 217138
rect 508550 217126 508602 217132
rect 507734 216988 507762 217110
rect 508562 216988 508590 217126
rect 509390 216988 509418 217246
rect 510218 216988 510246 217246
rect 511000 217138 511028 217495
rect 511828 217274 511856 220594
rect 512748 218890 512776 228890
rect 513116 220114 513144 231662
rect 513392 229294 513420 231676
rect 513380 229288 513432 229294
rect 513380 229230 513432 229236
rect 514036 227458 514064 231676
rect 514024 227452 514076 227458
rect 514024 227394 514076 227400
rect 514300 226024 514352 226030
rect 514300 225966 514352 225972
rect 513564 221740 513616 221746
rect 513564 221682 513616 221688
rect 513576 221513 513604 221682
rect 513562 221504 513618 221513
rect 513562 221439 513618 221448
rect 513104 220108 513156 220114
rect 513104 220050 513156 220056
rect 512736 218884 512788 218890
rect 512736 218826 512788 218832
rect 512748 217274 512776 218826
rect 513576 217274 513604 221439
rect 511828 217246 511902 217274
rect 511000 217110 511074 217138
rect 511046 216988 511074 217110
rect 511874 216988 511902 217246
rect 512702 217246 512776 217274
rect 513530 217246 513604 217274
rect 514312 217274 514340 225966
rect 514680 223310 514708 231676
rect 515324 229158 515352 231676
rect 515496 229696 515548 229702
rect 515496 229638 515548 229644
rect 515312 229152 515364 229158
rect 515312 229094 515364 229100
rect 514668 223304 514720 223310
rect 514668 223246 514720 223252
rect 515508 222086 515536 229638
rect 515772 228676 515824 228682
rect 515772 228618 515824 228624
rect 515496 222080 515548 222086
rect 515496 222022 515548 222028
rect 515128 221604 515180 221610
rect 515128 221546 515180 221552
rect 515140 220017 515168 221546
rect 515784 221241 515812 228618
rect 515968 224534 515996 231676
rect 516612 226030 516640 231676
rect 517256 230042 517284 231676
rect 517520 230240 517572 230246
rect 517520 230182 517572 230188
rect 517244 230036 517296 230042
rect 517244 229978 517296 229984
rect 516784 229900 516836 229906
rect 516784 229842 516836 229848
rect 516796 229094 516824 229842
rect 516796 229066 517008 229094
rect 516600 226024 516652 226030
rect 516600 225966 516652 225972
rect 515956 224528 516008 224534
rect 515956 224470 516008 224476
rect 516784 224392 516836 224398
rect 516784 224334 516836 224340
rect 515770 221232 515826 221241
rect 515770 221167 515826 221176
rect 515126 220008 515182 220017
rect 515126 219943 515182 219952
rect 515140 217274 515168 219943
rect 515784 219434 515812 221167
rect 515784 219406 516088 219434
rect 516060 217274 516088 219406
rect 514312 217246 514386 217274
rect 515140 217246 515214 217274
rect 512702 216988 512730 217246
rect 513530 216988 513558 217246
rect 514358 216988 514386 217246
rect 515186 216988 515214 217246
rect 516014 217246 516088 217274
rect 516796 217274 516824 224334
rect 516980 220386 517008 229066
rect 517532 223446 517560 230182
rect 517900 228682 517928 231676
rect 518544 228818 518572 231676
rect 519188 229906 519216 231676
rect 519176 229900 519228 229906
rect 519176 229842 519228 229848
rect 519176 229288 519228 229294
rect 519176 229230 519228 229236
rect 519188 229094 519216 229230
rect 519096 229066 519216 229094
rect 518164 228812 518216 228818
rect 518164 228754 518216 228760
rect 518532 228812 518584 228818
rect 518532 228754 518584 228760
rect 517888 228676 517940 228682
rect 517888 228618 517940 228624
rect 517520 223440 517572 223446
rect 517520 223382 517572 223388
rect 517520 222896 517572 222902
rect 517520 222838 517572 222844
rect 517532 220862 517560 222838
rect 517520 220856 517572 220862
rect 517520 220798 517572 220804
rect 516968 220380 517020 220386
rect 516968 220322 517020 220328
rect 518176 218754 518204 228754
rect 519096 224126 519124 229066
rect 519268 225888 519320 225894
rect 519268 225830 519320 225836
rect 519084 224120 519136 224126
rect 519084 224062 519136 224068
rect 518532 220856 518584 220862
rect 518532 220798 518584 220804
rect 517704 218748 517756 218754
rect 517704 218690 517756 218696
rect 518164 218748 518216 218754
rect 518164 218690 518216 218696
rect 517716 217274 517744 218690
rect 518544 217274 518572 220798
rect 516796 217246 516870 217274
rect 516014 216988 516042 217246
rect 516842 216988 516870 217246
rect 517670 217246 517744 217274
rect 518498 217246 518572 217274
rect 519280 217274 519308 225830
rect 519832 222902 519860 231676
rect 520476 224398 520504 231676
rect 521120 230382 521148 231676
rect 521108 230376 521160 230382
rect 521108 230318 521160 230324
rect 520924 229152 520976 229158
rect 520924 229094 520976 229100
rect 520464 224392 520516 224398
rect 520464 224334 520516 224340
rect 519820 222896 519872 222902
rect 519820 222838 519872 222844
rect 520936 220658 520964 229094
rect 521108 228540 521160 228546
rect 521108 228482 521160 228488
rect 521120 221134 521148 228482
rect 521764 225894 521792 231676
rect 522422 231662 522896 231690
rect 521752 225888 521804 225894
rect 521752 225830 521804 225836
rect 521752 223168 521804 223174
rect 521752 223110 521804 223116
rect 521108 221128 521160 221134
rect 521108 221070 521160 221076
rect 520924 220652 520976 220658
rect 520924 220594 520976 220600
rect 520188 220244 520240 220250
rect 520188 220186 520240 220192
rect 520200 219473 520228 220186
rect 520186 219464 520242 219473
rect 521120 219434 521148 221070
rect 520186 219399 520242 219408
rect 521028 219406 521148 219434
rect 520004 218748 520056 218754
rect 520004 218690 520056 218696
rect 520016 217569 520044 218690
rect 520002 217560 520058 217569
rect 520002 217495 520058 217504
rect 520200 217274 520228 219399
rect 521028 217274 521056 219406
rect 519280 217246 519354 217274
rect 517670 216988 517698 217246
rect 518498 216988 518526 217246
rect 519326 216988 519354 217246
rect 520154 217246 520228 217274
rect 520982 217246 521056 217274
rect 521764 217274 521792 223110
rect 522672 221876 522724 221882
rect 522672 221818 522724 221824
rect 522684 220969 522712 221818
rect 522868 221746 522896 231662
rect 523052 229770 523080 231676
rect 523040 229764 523092 229770
rect 523040 229706 523092 229712
rect 523696 227050 523724 231676
rect 524248 231662 524354 231690
rect 523040 227044 523092 227050
rect 523040 226986 523092 226992
rect 523684 227044 523736 227050
rect 523684 226986 523736 226992
rect 522856 221740 522908 221746
rect 522856 221682 522908 221688
rect 522670 220960 522726 220969
rect 522670 220895 522726 220904
rect 522684 217274 522712 220895
rect 523052 217870 523080 226986
rect 523500 224256 523552 224262
rect 523500 224198 523552 224204
rect 523512 221338 523540 224198
rect 523684 222488 523736 222494
rect 523684 222430 523736 222436
rect 523696 222222 523724 222430
rect 523684 222216 523736 222222
rect 523684 222158 523736 222164
rect 524248 221610 524276 231662
rect 524604 230036 524656 230042
rect 524604 229978 524656 229984
rect 524616 227594 524644 229978
rect 524984 229158 525012 231676
rect 524972 229152 525024 229158
rect 524972 229094 525024 229100
rect 524604 227588 524656 227594
rect 524604 227530 524656 227536
rect 524420 227316 524472 227322
rect 524420 227258 524472 227264
rect 524432 223786 524460 227258
rect 525628 224262 525656 231676
rect 526272 227322 526300 231676
rect 526444 230376 526496 230382
rect 526444 230318 526496 230324
rect 526456 228954 526484 230318
rect 526916 229634 526944 231676
rect 526904 229628 526956 229634
rect 526904 229570 526956 229576
rect 526444 228948 526496 228954
rect 526444 228890 526496 228896
rect 527560 228546 527588 231676
rect 528218 231662 528416 231690
rect 527548 228540 527600 228546
rect 527548 228482 527600 228488
rect 526260 227316 526312 227322
rect 526260 227258 526312 227264
rect 525984 227180 526036 227186
rect 525984 227122 526036 227128
rect 525616 224256 525668 224262
rect 525616 224198 525668 224204
rect 524420 223780 524472 223786
rect 524420 223722 524472 223728
rect 525064 223780 525116 223786
rect 525064 223722 525116 223728
rect 524236 221604 524288 221610
rect 524236 221546 524288 221552
rect 523500 221332 523552 221338
rect 523500 221274 523552 221280
rect 523040 217864 523092 217870
rect 523040 217806 523092 217812
rect 523512 217274 523540 221274
rect 524236 217864 524288 217870
rect 524236 217806 524288 217812
rect 521764 217246 521838 217274
rect 520154 216988 520182 217246
rect 520982 216988 521010 217246
rect 521810 216988 521838 217246
rect 522638 217246 522712 217274
rect 523466 217246 523540 217274
rect 522638 216988 522666 217246
rect 523466 216988 523494 217246
rect 524248 217138 524276 217806
rect 525076 217274 525104 223722
rect 525996 220998 526024 227122
rect 526720 224800 526772 224806
rect 526720 224742 526772 224748
rect 525984 220992 526036 220998
rect 525984 220934 526036 220940
rect 525996 217274 526024 220934
rect 525076 217246 525150 217274
rect 524248 217110 524322 217138
rect 524294 216988 524322 217110
rect 525122 216988 525150 217246
rect 525950 217246 526024 217274
rect 526732 217274 526760 224742
rect 527824 223032 527876 223038
rect 527824 222974 527876 222980
rect 527548 220380 527600 220386
rect 527548 220322 527600 220328
rect 527560 219638 527588 220322
rect 527548 219632 527600 219638
rect 527548 219574 527600 219580
rect 527560 217274 527588 219574
rect 527836 217462 527864 222974
rect 528388 220250 528416 231662
rect 528848 230110 528876 231676
rect 528836 230104 528888 230110
rect 528836 230046 528888 230052
rect 528560 229900 528612 229906
rect 528560 229842 528612 229848
rect 528572 226166 528600 229842
rect 528560 226160 528612 226166
rect 528560 226102 528612 226108
rect 529204 225752 529256 225758
rect 529204 225694 529256 225700
rect 528376 220244 528428 220250
rect 528376 220186 528428 220192
rect 527824 217456 527876 217462
rect 527824 217398 527876 217404
rect 528468 217456 528520 217462
rect 528468 217398 528520 217404
rect 526732 217246 526806 217274
rect 527560 217246 527634 217274
rect 525950 216988 525978 217246
rect 526778 216988 526806 217246
rect 527606 216988 527634 217246
rect 528480 217138 528508 217398
rect 529216 217274 529244 225694
rect 529492 223038 529520 231676
rect 530136 230382 530164 231676
rect 530124 230376 530176 230382
rect 530124 230318 530176 230324
rect 530780 230246 530808 231676
rect 531136 230376 531188 230382
rect 531136 230318 531188 230324
rect 530768 230240 530820 230246
rect 530768 230182 530820 230188
rect 529940 229152 529992 229158
rect 529940 229094 529992 229100
rect 531148 229094 531176 230318
rect 529952 224806 529980 229094
rect 531148 229066 531268 229094
rect 531044 225616 531096 225622
rect 531044 225558 531096 225564
rect 529940 224800 529992 224806
rect 529940 224742 529992 224748
rect 530860 224528 530912 224534
rect 530860 224470 530912 224476
rect 530872 224126 530900 224470
rect 530676 224120 530728 224126
rect 530676 224062 530728 224068
rect 530860 224120 530912 224126
rect 530860 224062 530912 224068
rect 530688 223650 530716 224062
rect 530676 223644 530728 223650
rect 530676 223586 530728 223592
rect 529480 223032 529532 223038
rect 529480 222974 529532 222980
rect 529848 222488 529900 222494
rect 529848 222430 529900 222436
rect 529860 222086 529888 222430
rect 529848 222080 529900 222086
rect 529848 222022 529900 222028
rect 529860 221320 529888 222022
rect 529860 221292 530072 221320
rect 530044 217274 530072 221292
rect 531056 219434 531084 225558
rect 531240 220386 531268 229066
rect 531424 225622 531452 231676
rect 531412 225616 531464 225622
rect 531412 225558 531464 225564
rect 531504 223440 531556 223446
rect 531504 223382 531556 223388
rect 531228 220380 531280 220386
rect 531228 220322 531280 220328
rect 530964 219406 531084 219434
rect 530964 217598 530992 219406
rect 530952 217592 531004 217598
rect 531516 217569 531544 223382
rect 532068 223174 532096 231676
rect 532516 230444 532568 230450
rect 532516 230386 532568 230392
rect 532528 230110 532556 230386
rect 532712 230178 532740 231676
rect 532700 230172 532752 230178
rect 532700 230114 532752 230120
rect 532516 230104 532568 230110
rect 532516 230046 532568 230052
rect 532976 228404 533028 228410
rect 532976 228346 533028 228352
rect 532700 224256 532752 224262
rect 532700 224198 532752 224204
rect 532712 223786 532740 224198
rect 532700 223780 532752 223786
rect 532700 223722 532752 223728
rect 532056 223168 532108 223174
rect 532056 223110 532108 223116
rect 531688 220516 531740 220522
rect 531688 220458 531740 220464
rect 530952 217534 531004 217540
rect 531502 217560 531558 217569
rect 529216 217246 529290 217274
rect 530044 217246 530118 217274
rect 528434 217110 528508 217138
rect 528434 216988 528462 217110
rect 529262 216988 529290 217246
rect 530090 216988 530118 217246
rect 530964 217138 530992 217534
rect 531502 217495 531558 217504
rect 531700 217274 531728 220458
rect 532988 219434 533016 228346
rect 533356 227186 533384 231676
rect 533344 227180 533396 227186
rect 533344 227122 533396 227128
rect 534000 222086 534028 231676
rect 534644 230042 534672 231676
rect 534632 230036 534684 230042
rect 534632 229978 534684 229984
rect 534724 229764 534776 229770
rect 534724 229706 534776 229712
rect 534540 224800 534592 224806
rect 534540 224742 534592 224748
rect 534552 224126 534580 224742
rect 534356 224120 534408 224126
rect 534356 224062 534408 224068
rect 534540 224120 534592 224126
rect 534540 224062 534592 224068
rect 534368 223650 534396 224062
rect 534356 223644 534408 223650
rect 534356 223586 534408 223592
rect 534736 223446 534764 229706
rect 535288 224670 535316 231676
rect 535736 227452 535788 227458
rect 535736 227394 535788 227400
rect 535276 224664 535328 224670
rect 535276 224606 535328 224612
rect 535000 223780 535052 223786
rect 535000 223722 535052 223728
rect 534724 223440 534776 223446
rect 534724 223382 534776 223388
rect 533988 222080 534040 222086
rect 533250 222048 533306 222057
rect 533988 222022 534040 222028
rect 533250 221983 533306 221992
rect 533264 221474 533292 221983
rect 533620 221604 533672 221610
rect 533620 221546 533672 221552
rect 533252 221468 533304 221474
rect 533252 221410 533304 221416
rect 533160 221332 533212 221338
rect 533632 221320 533660 221546
rect 533212 221292 533660 221320
rect 533160 221274 533212 221280
rect 534172 220108 534224 220114
rect 534172 220050 534224 220056
rect 532988 219406 533476 219434
rect 533448 217734 533476 219406
rect 533436 217728 533488 217734
rect 533436 217670 533488 217676
rect 532514 217560 532570 217569
rect 532514 217495 532570 217504
rect 531700 217246 531774 217274
rect 530918 217110 530992 217138
rect 530918 216988 530946 217110
rect 531746 216988 531774 217246
rect 532528 217138 532556 217495
rect 533448 217138 533476 217670
rect 532528 217110 532602 217138
rect 532574 216988 532602 217110
rect 533402 217110 533476 217138
rect 534184 217138 534212 220050
rect 535012 217138 535040 223722
rect 535748 221785 535776 227394
rect 535932 225758 535960 231676
rect 536576 229906 536604 231676
rect 536564 229900 536616 229906
rect 536564 229842 536616 229848
rect 536104 229628 536156 229634
rect 536104 229570 536156 229576
rect 535920 225752 535972 225758
rect 535920 225694 535972 225700
rect 536116 221950 536144 229570
rect 537220 228410 537248 231676
rect 537878 231662 538168 231690
rect 537208 228404 537260 228410
rect 537208 228346 537260 228352
rect 536288 223304 536340 223310
rect 536288 223246 536340 223252
rect 536104 221944 536156 221950
rect 536104 221886 536156 221892
rect 535734 221776 535790 221785
rect 535734 221711 535790 221720
rect 535748 217274 535776 221711
rect 536300 221388 536328 223246
rect 536208 221360 536328 221388
rect 536208 219298 536236 221360
rect 537484 220652 537536 220658
rect 537484 220594 537536 220600
rect 536196 219292 536248 219298
rect 536196 219234 536248 219240
rect 536656 219292 536708 219298
rect 536656 219234 536708 219240
rect 535748 217246 535914 217274
rect 534184 217110 534258 217138
rect 535012 217110 535086 217138
rect 533402 216988 533430 217110
rect 534230 216988 534258 217110
rect 535058 216988 535086 217110
rect 535886 216988 535914 217246
rect 536668 217138 536696 219234
rect 537496 218754 537524 220594
rect 538140 220114 538168 231662
rect 538312 230444 538364 230450
rect 538312 230386 538364 230392
rect 538324 227458 538352 230386
rect 538508 229770 538536 231676
rect 538784 231662 539166 231690
rect 538496 229764 538548 229770
rect 538496 229706 538548 229712
rect 538784 229094 538812 231662
rect 539600 230308 539652 230314
rect 539600 230250 539652 230256
rect 538508 229066 538812 229094
rect 538312 227452 538364 227458
rect 538312 227394 538364 227400
rect 538312 223644 538364 223650
rect 538312 223586 538364 223592
rect 538324 220590 538352 223586
rect 538508 222057 538536 229066
rect 539612 228682 539640 230250
rect 547144 230172 547196 230178
rect 547144 230114 547196 230120
rect 544016 228948 544068 228954
rect 544016 228890 544068 228896
rect 541532 228812 541584 228818
rect 541532 228754 541584 228760
rect 539416 228676 539468 228682
rect 539416 228618 539468 228624
rect 539600 228676 539652 228682
rect 539600 228618 539652 228624
rect 539428 228274 539456 228618
rect 539416 228268 539468 228274
rect 539416 228210 539468 228216
rect 540796 228268 540848 228274
rect 540796 228210 540848 228216
rect 539968 227588 540020 227594
rect 539968 227530 540020 227536
rect 538680 226024 538732 226030
rect 538680 225966 538732 225972
rect 538692 224954 538720 225966
rect 538692 224926 539180 224954
rect 538494 222048 538550 222057
rect 538494 221983 538550 221992
rect 538678 221776 538734 221785
rect 538678 221711 538734 221720
rect 538692 221406 538720 221711
rect 538680 221400 538732 221406
rect 538680 221342 538732 221348
rect 538312 220584 538364 220590
rect 538312 220526 538364 220532
rect 538128 220108 538180 220114
rect 538128 220050 538180 220056
rect 537484 218748 537536 218754
rect 537484 218690 537536 218696
rect 537496 217138 537524 218690
rect 538324 217138 538352 220526
rect 539152 217274 539180 224926
rect 539980 223650 540008 227530
rect 539968 223644 540020 223650
rect 539968 223586 540020 223592
rect 539980 217274 540008 223586
rect 540808 219638 540836 228210
rect 541544 224954 541572 228754
rect 543004 226160 543056 226166
rect 543004 226102 543056 226108
rect 541544 224926 541664 224954
rect 540796 219632 540848 219638
rect 540796 219574 540848 219580
rect 540808 217274 540836 219574
rect 541636 217274 541664 224926
rect 542360 222896 542412 222902
rect 542360 222838 542412 222844
rect 542372 217598 542400 222838
rect 543016 219162 543044 226102
rect 544028 224954 544056 228890
rect 545764 225888 545816 225894
rect 545764 225830 545816 225836
rect 543936 224926 544056 224954
rect 543738 224496 543794 224505
rect 543738 224431 543794 224440
rect 543752 224126 543780 224431
rect 543740 224120 543792 224126
rect 543740 224062 543792 224068
rect 543936 224058 543964 224926
rect 544108 224528 544160 224534
rect 544292 224528 544344 224534
rect 544108 224470 544160 224476
rect 544290 224496 544292 224505
rect 544344 224496 544346 224505
rect 543924 224052 543976 224058
rect 543924 223994 543976 224000
rect 543832 222896 543884 222902
rect 543832 222838 543884 222844
rect 543844 222034 543872 222838
rect 543706 222006 543872 222034
rect 543706 221950 543734 222006
rect 543694 221944 543746 221950
rect 543694 221886 543746 221892
rect 543648 221264 543700 221270
rect 543648 221206 543700 221212
rect 543832 221264 543884 221270
rect 543832 221206 543884 221212
rect 543660 220726 543688 221206
rect 543648 220720 543700 220726
rect 543648 220662 543700 220668
rect 543844 220590 543872 221206
rect 543832 220584 543884 220590
rect 543832 220526 543884 220532
rect 542544 219156 542596 219162
rect 542544 219098 542596 219104
rect 543004 219156 543056 219162
rect 543004 219098 543056 219104
rect 542360 217592 542412 217598
rect 542360 217534 542412 217540
rect 539152 217246 539226 217274
rect 539980 217246 540054 217274
rect 540808 217246 540882 217274
rect 541636 217246 541710 217274
rect 536668 217110 536742 217138
rect 537496 217110 537570 217138
rect 538324 217110 538398 217138
rect 536714 216988 536742 217110
rect 537542 216988 537570 217110
rect 538370 216988 538398 217110
rect 539198 216988 539226 217246
rect 540026 216988 540054 217246
rect 540854 216988 540882 217246
rect 541682 216988 541710 217246
rect 542556 217138 542584 219098
rect 543280 217592 543332 217598
rect 543280 217534 543332 217540
rect 542510 217110 542584 217138
rect 543292 217138 543320 217534
rect 544120 217274 544148 224470
rect 544290 224431 544346 224440
rect 545028 224052 545080 224058
rect 545028 223994 545080 224000
rect 544120 217246 544194 217274
rect 543292 217110 543366 217138
rect 542510 216988 542538 217110
rect 543338 216988 543366 217110
rect 544166 216988 544194 217246
rect 545040 217138 545068 223994
rect 545776 221785 545804 225830
rect 547156 221882 547184 230114
rect 550548 230036 550600 230042
rect 550548 229978 550600 229984
rect 548340 227044 548392 227050
rect 548340 226986 548392 226992
rect 547420 223440 547472 223446
rect 547420 223382 547472 223388
rect 546592 221876 546644 221882
rect 546592 221818 546644 221824
rect 547144 221876 547196 221882
rect 547144 221818 547196 221824
rect 545762 221776 545818 221785
rect 545762 221711 545818 221720
rect 545776 217274 545804 221711
rect 545776 217246 545850 217274
rect 544994 217110 545068 217138
rect 544994 216988 545022 217110
rect 545822 216988 545850 217246
rect 546604 217138 546632 221818
rect 547432 218890 547460 223382
rect 548352 219586 548380 226986
rect 550560 224618 550588 229978
rect 553308 228540 553360 228546
rect 553308 228482 553360 228488
rect 550916 227316 550968 227322
rect 550916 227258 550968 227264
rect 550928 224954 550956 227258
rect 550928 224926 551600 224954
rect 550560 224590 551232 224618
rect 551204 224534 551232 224590
rect 549996 224528 550048 224534
rect 549996 224470 550048 224476
rect 550364 224528 550416 224534
rect 551192 224528 551244 224534
rect 550364 224470 550416 224476
rect 549258 221776 549314 221785
rect 549258 221711 549260 221720
rect 549312 221711 549314 221720
rect 549260 221682 549312 221688
rect 548892 221400 548944 221406
rect 548536 221348 548892 221354
rect 548536 221342 548944 221348
rect 548536 221326 548932 221342
rect 548536 221270 548564 221326
rect 548524 221264 548576 221270
rect 548524 221206 548576 221212
rect 549076 220720 549128 220726
rect 549076 220662 549128 220668
rect 548708 220244 548760 220250
rect 548708 220186 548760 220192
rect 548720 219774 548748 220186
rect 548708 219768 548760 219774
rect 548708 219710 548760 219716
rect 548892 219768 548944 219774
rect 548892 219710 548944 219716
rect 548904 219586 548932 219710
rect 548352 219558 548932 219586
rect 547420 218884 547472 218890
rect 547420 218826 547472 218832
rect 547432 217138 547460 218826
rect 548352 217274 548380 219558
rect 548892 219292 548944 219298
rect 548892 219234 548944 219240
rect 548708 219020 548760 219026
rect 548708 218962 548760 218968
rect 548720 218618 548748 218962
rect 548904 218618 548932 219234
rect 548708 218612 548760 218618
rect 548708 218554 548760 218560
rect 548892 218612 548944 218618
rect 548892 218554 548944 218560
rect 548306 217246 548380 217274
rect 546604 217110 546678 217138
rect 547432 217110 547506 217138
rect 546650 216988 546678 217110
rect 547478 216988 547506 217110
rect 548306 216988 548334 217246
rect 549088 217138 549116 220662
rect 550008 217138 550036 224470
rect 550376 224210 550404 224470
rect 550652 224454 551048 224482
rect 551192 224470 551244 224476
rect 550652 224398 550680 224454
rect 550640 224392 550692 224398
rect 550640 224334 550692 224340
rect 550824 224392 550876 224398
rect 550824 224334 550876 224340
rect 550836 224210 550864 224334
rect 550376 224182 550864 224210
rect 551020 220658 551048 224454
rect 551008 220652 551060 220658
rect 551008 220594 551060 220600
rect 551020 219178 551048 220594
rect 550836 219150 551048 219178
rect 550836 217274 550864 219150
rect 549088 217110 549162 217138
rect 549134 216988 549162 217110
rect 549962 217110 550036 217138
rect 550790 217246 550864 217274
rect 551572 217274 551600 224926
rect 552480 222896 552532 222902
rect 552480 222838 552532 222844
rect 551572 217246 551646 217274
rect 549962 216988 549990 217110
rect 550790 216988 550818 217246
rect 551618 216988 551646 217246
rect 552492 217138 552520 222838
rect 553320 221785 553348 228482
rect 554056 223310 554084 249047
rect 555424 244316 555476 244322
rect 555424 244258 555476 244264
rect 554502 240408 554558 240417
rect 554502 240343 554558 240352
rect 554516 240174 554544 240343
rect 554504 240168 554556 240174
rect 554504 240110 554556 240116
rect 554320 238740 554372 238746
rect 554320 238682 554372 238688
rect 554332 238241 554360 238682
rect 554318 238232 554374 238241
rect 554318 238167 554374 238176
rect 554412 234592 554464 234598
rect 554412 234534 554464 234540
rect 554424 233889 554452 234534
rect 554410 233880 554466 233889
rect 554410 233815 554466 233824
rect 555436 227050 555464 244258
rect 556816 228546 556844 251194
rect 556988 228676 557040 228682
rect 556988 228618 557040 228624
rect 556804 228540 556856 228546
rect 556804 228482 556856 228488
rect 556068 227452 556120 227458
rect 556068 227394 556120 227400
rect 555424 227044 555476 227050
rect 555424 226986 555476 226992
rect 556080 224505 556108 227394
rect 554870 224496 554926 224505
rect 554870 224431 554926 224440
rect 556066 224496 556122 224505
rect 556066 224431 556122 224440
rect 554044 223304 554096 223310
rect 554044 223246 554096 223252
rect 553306 221776 553362 221785
rect 553306 221711 553362 221720
rect 553320 217274 553348 221711
rect 554228 220652 554280 220658
rect 554228 220594 554280 220600
rect 554240 220386 554268 220594
rect 554044 220380 554096 220386
rect 554044 220322 554096 220328
rect 554228 220380 554280 220386
rect 554228 220322 554280 220328
rect 552446 217110 552520 217138
rect 553274 217246 553348 217274
rect 554056 217274 554084 220322
rect 554884 217274 554912 224431
rect 555700 223032 555752 223038
rect 555700 222974 555752 222980
rect 555712 220658 555740 222974
rect 556802 222048 556858 222057
rect 556802 221983 556858 221992
rect 556816 221882 556844 221983
rect 556804 221876 556856 221882
rect 556804 221818 556856 221824
rect 555700 220652 555752 220658
rect 555700 220594 555752 220600
rect 555712 217274 555740 220594
rect 556528 220516 556580 220522
rect 556528 220458 556580 220464
rect 556540 217274 556568 220458
rect 557000 219434 557028 228618
rect 558196 225894 558224 255546
rect 559564 246356 559616 246362
rect 559564 246298 559616 246304
rect 559576 236842 559604 246298
rect 559564 236836 559616 236842
rect 559564 236778 559616 236784
rect 560956 230110 560984 256702
rect 562324 252612 562376 252618
rect 562324 252554 562376 252560
rect 560944 230104 560996 230110
rect 560944 230046 560996 230052
rect 559564 229900 559616 229906
rect 559564 229842 559616 229848
rect 558184 225888 558236 225894
rect 558184 225830 558236 225836
rect 558276 225616 558328 225622
rect 558276 225558 558328 225564
rect 557184 224862 557534 224890
rect 557184 224534 557212 224862
rect 557356 224800 557408 224806
rect 557356 224742 557408 224748
rect 557506 224754 557534 224862
rect 557630 224768 557686 224777
rect 557368 224618 557396 224742
rect 557506 224726 557630 224754
rect 557630 224703 557686 224712
rect 557816 224664 557868 224670
rect 557368 224612 557816 224618
rect 557368 224606 557868 224612
rect 557368 224590 557856 224606
rect 557172 224528 557224 224534
rect 557172 224470 557224 224476
rect 557630 224496 557686 224505
rect 557686 224454 557856 224482
rect 557630 224431 557686 224440
rect 557828 224398 557856 224454
rect 557816 224392 557868 224398
rect 557816 224334 557868 224340
rect 557540 222624 557592 222630
rect 557540 222566 557592 222572
rect 557552 222057 557580 222566
rect 557538 222048 557594 222057
rect 557538 221983 557594 221992
rect 557172 221944 557224 221950
rect 557172 221886 557224 221892
rect 557184 221785 557212 221886
rect 557170 221776 557226 221785
rect 557170 221711 557226 221720
rect 558288 220386 558316 225558
rect 559012 223168 559064 223174
rect 559012 223110 559064 223116
rect 558276 220380 558328 220386
rect 558276 220322 558328 220328
rect 557000 219406 557396 219434
rect 557368 219298 557396 219406
rect 557356 219292 557408 219298
rect 557356 219234 557408 219240
rect 557368 217274 557396 219234
rect 558288 217274 558316 220322
rect 554056 217246 554130 217274
rect 554884 217246 554958 217274
rect 555712 217246 555786 217274
rect 556540 217246 556614 217274
rect 557368 217246 557442 217274
rect 552446 216988 552474 217110
rect 553274 216988 553302 217246
rect 554102 216988 554130 217246
rect 554930 216988 554958 217246
rect 555758 216988 555786 217246
rect 556586 216988 556614 217246
rect 557414 216988 557442 217246
rect 558242 217246 558316 217274
rect 559024 217274 559052 223110
rect 559380 223032 559432 223038
rect 559380 222974 559432 222980
rect 559392 222222 559420 222974
rect 559380 222216 559432 222222
rect 559380 222158 559432 222164
rect 559576 222154 559604 229842
rect 560944 227180 560996 227186
rect 560944 227122 560996 227128
rect 559840 223168 559892 223174
rect 559840 223110 559892 223116
rect 559852 222630 559880 223110
rect 559840 222624 559892 222630
rect 559840 222566 559892 222572
rect 559564 222148 559616 222154
rect 559564 222090 559616 222096
rect 559380 222080 559432 222086
rect 559378 222048 559380 222057
rect 559432 222048 559434 222057
rect 559378 221983 559434 221992
rect 559852 217274 559880 222566
rect 560956 217569 560984 227122
rect 562336 224806 562364 252554
rect 563716 225010 563744 259422
rect 568120 230104 568172 230110
rect 568120 230046 568172 230052
rect 566832 229764 566884 229770
rect 566832 229706 566884 229712
rect 565636 228404 565688 228410
rect 565636 228346 565688 228352
rect 563980 225752 564032 225758
rect 563980 225694 564032 225700
rect 563704 225004 563756 225010
rect 563704 224946 563756 224952
rect 562140 224800 562192 224806
rect 561954 224768 562010 224777
rect 561954 224703 562010 224712
rect 562138 224768 562140 224777
rect 562324 224800 562376 224806
rect 562192 224768 562194 224777
rect 562324 224742 562376 224748
rect 563702 224768 563758 224777
rect 562138 224703 562194 224712
rect 563702 224703 563758 224712
rect 561968 223446 561996 224703
rect 561956 223440 562008 223446
rect 561956 223382 562008 223388
rect 561968 222442 561996 223382
rect 562508 223304 562560 223310
rect 562508 223246 562560 223252
rect 562520 222902 562548 223246
rect 562324 222896 562376 222902
rect 562324 222838 562376 222844
rect 562508 222896 562560 222902
rect 562508 222838 562560 222844
rect 562336 222630 562364 222838
rect 562324 222624 562376 222630
rect 562324 222566 562376 222572
rect 561968 222414 562364 222442
rect 561494 222048 561550 222057
rect 561494 221983 561550 221992
rect 561312 219156 561364 219162
rect 561312 219098 561364 219104
rect 561324 217841 561352 219098
rect 561310 217832 561366 217841
rect 561310 217767 561366 217776
rect 560758 217560 560814 217569
rect 560758 217495 560814 217504
rect 560942 217560 560998 217569
rect 560942 217495 560998 217504
rect 559024 217246 559098 217274
rect 559852 217246 559926 217274
rect 558242 216988 558270 217246
rect 559070 216988 559098 217246
rect 559898 216988 559926 217246
rect 560772 217138 560800 217495
rect 561508 217274 561536 221983
rect 561770 220552 561826 220561
rect 561770 220487 561826 220496
rect 562140 220516 562192 220522
rect 561784 220386 561812 220487
rect 562140 220458 562192 220464
rect 561772 220380 561824 220386
rect 561772 220322 561824 220328
rect 561772 220108 561824 220114
rect 561772 220050 561824 220056
rect 561784 218793 561812 220050
rect 562152 220046 562180 220458
rect 562140 220040 562192 220046
rect 562140 219982 562192 219988
rect 562048 219360 562100 219366
rect 562048 219302 562100 219308
rect 562060 219201 562088 219302
rect 562046 219192 562102 219201
rect 562046 219127 562102 219136
rect 561770 218784 561826 218793
rect 561770 218719 561826 218728
rect 562336 217274 562364 222414
rect 563716 221785 563744 224703
rect 563702 221776 563758 221785
rect 563702 221711 563758 221720
rect 563058 220688 563114 220697
rect 562876 220652 562928 220658
rect 563058 220623 563060 220632
rect 562876 220594 562928 220600
rect 563112 220623 563114 220632
rect 563060 220594 563112 220600
rect 562888 220250 562916 220594
rect 562876 220244 562928 220250
rect 562876 220186 562928 220192
rect 562598 219192 562654 219201
rect 562598 219127 562654 219136
rect 562612 218890 562640 219127
rect 563164 219026 563376 219042
rect 563152 219020 563388 219026
rect 563204 219014 563336 219020
rect 563152 218962 563204 218968
rect 563336 218962 563388 218968
rect 563520 219020 563572 219026
rect 563520 218962 563572 218968
rect 562600 218884 562652 218890
rect 562600 218826 562652 218832
rect 562968 218884 563020 218890
rect 563336 218884 563388 218890
rect 563020 218844 563336 218872
rect 562968 218826 563020 218832
rect 563336 218826 563388 218832
rect 563532 218770 563560 218962
rect 562888 218742 563560 218770
rect 562600 218612 562652 218618
rect 562888 218600 562916 218742
rect 562652 218572 562916 218600
rect 563058 218648 563114 218657
rect 563058 218583 563114 218592
rect 562600 218554 562652 218560
rect 563072 218210 563100 218583
rect 563060 218204 563112 218210
rect 563060 218146 563112 218152
rect 563336 218000 563388 218006
rect 563072 217948 563336 217954
rect 563072 217942 563388 217948
rect 563072 217926 563376 217942
rect 561508 217246 561582 217274
rect 562336 217246 562410 217274
rect 560726 217110 560800 217138
rect 560726 216988 560754 217110
rect 561554 216988 561582 217246
rect 562382 216988 562410 217246
rect 563072 217190 563100 217926
rect 563716 217682 563744 221711
rect 563164 217654 563744 217682
rect 563164 217274 563192 217654
rect 563334 217560 563390 217569
rect 563334 217495 563390 217504
rect 563348 217326 563376 217495
rect 563336 217320 563388 217326
rect 563164 217246 563238 217274
rect 563336 217262 563388 217268
rect 563992 217274 564020 225694
rect 564808 222148 564860 222154
rect 564808 222090 564860 222096
rect 564820 219065 564848 222090
rect 565648 220561 565676 228346
rect 566844 223310 566872 229706
rect 567016 225140 567068 225146
rect 567016 225082 567068 225088
rect 567028 224806 567056 225082
rect 567016 224800 567068 224806
rect 567016 224742 567068 224748
rect 567844 224800 567896 224806
rect 567844 224742 567896 224748
rect 567856 223650 567884 224742
rect 567844 223644 567896 223650
rect 567844 223586 567896 223592
rect 566832 223304 566884 223310
rect 566832 223246 566884 223252
rect 565634 220552 565690 220561
rect 565634 220487 565690 220496
rect 564806 219056 564862 219065
rect 564806 218991 564862 219000
rect 564162 218648 564218 218657
rect 564162 218583 564164 218592
rect 564216 218583 564218 218592
rect 564164 218554 564216 218560
rect 563992 217246 564066 217274
rect 563060 217184 563112 217190
rect 563060 217126 563112 217132
rect 563210 216988 563238 217246
rect 564038 216988 564066 217246
rect 564820 217138 564848 218991
rect 565648 217274 565676 220487
rect 566844 220386 566872 223246
rect 567660 223168 567712 223174
rect 567660 223110 567712 223116
rect 567672 222222 567700 223110
rect 567660 222216 567712 222222
rect 567660 222158 567712 222164
rect 566832 220380 566884 220386
rect 566832 220322 566884 220328
rect 567292 220380 567344 220386
rect 567292 220322 567344 220328
rect 566462 218784 566518 218793
rect 566462 218719 566518 218728
rect 565648 217246 565722 217274
rect 564820 217110 564894 217138
rect 564866 216988 564894 217110
rect 565694 216988 565722 217246
rect 566476 217172 566504 218719
rect 567304 217274 567332 220322
rect 568132 217274 568160 230046
rect 568304 223644 568356 223650
rect 568304 223586 568356 223592
rect 568316 223310 568344 223586
rect 568304 223304 568356 223310
rect 568304 223246 568356 223252
rect 568304 223032 568356 223038
rect 568304 222974 568356 222980
rect 568316 222358 568344 222974
rect 568304 222352 568356 222358
rect 568304 222294 568356 222300
rect 568592 220522 568620 260850
rect 570616 234598 570644 261462
rect 596824 245676 596876 245682
rect 596824 245618 596876 245624
rect 576124 242208 576176 242214
rect 576124 242150 576176 242156
rect 576136 238746 576164 242150
rect 577504 240168 577556 240174
rect 577504 240110 577556 240116
rect 576124 238740 576176 238746
rect 576124 238682 576176 238688
rect 570604 234592 570656 234598
rect 570604 234534 570656 234540
rect 570604 228540 570656 228546
rect 570604 228482 570656 228488
rect 568948 224936 569000 224942
rect 568948 224878 569000 224884
rect 568764 223440 568816 223446
rect 568764 223382 568816 223388
rect 568776 222358 568804 223382
rect 568764 222352 568816 222358
rect 568764 222294 568816 222300
rect 568580 220516 568632 220522
rect 568580 220458 568632 220464
rect 567304 217246 567378 217274
rect 568132 217246 568206 217274
rect 566476 217144 566550 217172
rect 566522 216988 566550 217144
rect 567350 216988 567378 217246
rect 568178 216988 568206 217246
rect 568960 217138 568988 224878
rect 569776 220516 569828 220522
rect 569776 220458 569828 220464
rect 569788 217138 569816 220458
rect 570616 217274 570644 228482
rect 571984 225888 572036 225894
rect 571984 225830 572036 225836
rect 571432 225140 571484 225146
rect 571432 225082 571484 225088
rect 571444 217274 571472 225082
rect 571996 224954 572024 225830
rect 571996 224926 572208 224954
rect 571982 217560 572038 217569
rect 571982 217495 572038 217504
rect 571996 217326 572024 217495
rect 571984 217320 572036 217326
rect 570616 217246 570690 217274
rect 571444 217246 571518 217274
rect 571984 217262 572036 217268
rect 572180 217274 572208 224926
rect 572626 221776 572682 221785
rect 572626 221711 572682 221720
rect 572640 220538 572668 221711
rect 574742 220552 574798 220561
rect 572640 220522 572714 220538
rect 572640 220516 572726 220522
rect 572640 220510 572674 220516
rect 574742 220487 574798 220496
rect 572674 220458 572726 220464
rect 574756 220386 574784 220487
rect 572352 220380 572404 220386
rect 572352 220322 572404 220328
rect 574744 220380 574796 220386
rect 574744 220322 574796 220328
rect 572364 219450 572392 220322
rect 572364 219422 572714 219450
rect 572536 219360 572588 219366
rect 572536 219302 572588 219308
rect 572352 219020 572404 219026
rect 572352 218962 572404 218968
rect 572364 218657 572392 218962
rect 572548 218770 572576 219302
rect 572686 219298 572714 219422
rect 572674 219292 572726 219298
rect 572674 219234 572726 219240
rect 574560 219156 574612 219162
rect 574560 219098 574612 219104
rect 572672 219056 572728 219065
rect 572672 218991 572674 219000
rect 572726 218991 572728 219000
rect 572674 218962 572726 218968
rect 572548 218742 572714 218770
rect 572350 218648 572406 218657
rect 572686 218618 572714 218742
rect 574374 218648 574430 218657
rect 572350 218583 572406 218592
rect 572536 218612 572588 218618
rect 572536 218554 572588 218560
rect 572674 218612 572726 218618
rect 574374 218583 574430 218592
rect 572674 218554 572726 218560
rect 572548 218226 572576 218554
rect 572548 218210 572714 218226
rect 572548 218204 572726 218210
rect 572548 218198 572674 218204
rect 572674 218146 572726 218152
rect 572352 218000 572404 218006
rect 572404 217948 572576 217954
rect 572352 217942 572576 217948
rect 572364 217926 572576 217942
rect 572180 217246 572300 217274
rect 568960 217110 569034 217138
rect 569788 217110 569862 217138
rect 569006 216988 569034 217110
rect 569834 216988 569862 217110
rect 570662 216988 570690 217246
rect 571490 216988 571518 217246
rect 572272 217138 572300 217246
rect 572548 217138 572576 217926
rect 574190 217560 574246 217569
rect 574190 217495 574246 217504
rect 572674 217184 572726 217190
rect 572272 217110 572346 217138
rect 572548 217132 572674 217138
rect 572548 217126 572726 217132
rect 572548 217110 572714 217126
rect 572318 216988 572346 217110
rect 574204 217054 574232 217495
rect 574192 217048 574244 217054
rect 574192 216990 574244 216996
rect 52458 215112 52514 215121
rect 52458 215047 52514 215056
rect 53286 215112 53342 215121
rect 53286 215047 53342 215056
rect 52472 214305 52500 215047
rect 574388 214742 574416 218583
rect 574376 214736 574428 214742
rect 574376 214678 574428 214684
rect 574572 214606 574600 219098
rect 574742 217832 574798 217841
rect 574742 217767 574798 217776
rect 574756 214878 574784 217767
rect 575478 216744 575534 216753
rect 575478 216679 575534 216688
rect 574744 214872 574796 214878
rect 574744 214814 574796 214820
rect 574560 214600 574612 214606
rect 574560 214542 574612 214548
rect 52458 214296 52514 214305
rect 52458 214231 52514 214240
rect 575492 213246 575520 216679
rect 575480 213240 575532 213246
rect 575480 213182 575532 213188
rect 577516 99142 577544 240110
rect 596836 224954 596864 245618
rect 629944 241528 629996 241534
rect 629944 241470 629996 241476
rect 629956 229094 629984 241470
rect 629956 229066 630076 229094
rect 596836 224926 597048 224954
rect 591486 224224 591542 224233
rect 591486 224159 591542 224168
rect 586980 223304 587032 223310
rect 586980 223246 587032 223252
rect 586992 222766 587020 223246
rect 587164 223032 587216 223038
rect 587164 222974 587216 222980
rect 587176 222766 587204 222974
rect 586980 222760 587032 222766
rect 586980 222702 587032 222708
rect 587164 222760 587216 222766
rect 587164 222702 587216 222708
rect 582378 220688 582434 220697
rect 587530 220688 587586 220697
rect 582378 220623 582434 220632
rect 587348 220652 587400 220658
rect 582392 219502 582420 220623
rect 587530 220623 587532 220632
rect 587348 220594 587400 220600
rect 587584 220623 587586 220632
rect 587532 220594 587584 220600
rect 587360 220114 587388 220594
rect 587348 220108 587400 220114
rect 587348 220050 587400 220056
rect 586980 219904 587032 219910
rect 586980 219846 587032 219852
rect 582380 219496 582432 219502
rect 582380 219438 582432 219444
rect 586992 219230 587020 219846
rect 586980 219224 587032 219230
rect 586980 219166 587032 219172
rect 578882 214024 578938 214033
rect 578882 213959 578938 213968
rect 578514 211712 578570 211721
rect 578514 211647 578570 211656
rect 578528 211206 578556 211647
rect 578516 211200 578568 211206
rect 578516 211142 578568 211148
rect 578896 208350 578924 213959
rect 591304 212696 591356 212702
rect 591304 212638 591356 212644
rect 580908 211200 580960 211206
rect 580908 211142 580960 211148
rect 579528 209840 579580 209846
rect 579526 209808 579528 209817
rect 579580 209808 579582 209817
rect 579526 209743 579582 209752
rect 578884 208344 578936 208350
rect 578884 208286 578936 208292
rect 579526 207496 579582 207505
rect 579582 207454 579752 207482
rect 579526 207431 579582 207440
rect 579526 205864 579582 205873
rect 579526 205799 579528 205808
rect 579580 205799 579582 205808
rect 579528 205770 579580 205776
rect 579724 204270 579752 207454
rect 580920 206922 580948 211142
rect 582288 209840 582340 209846
rect 582288 209782 582340 209788
rect 581644 208616 581696 208622
rect 581644 208558 581696 208564
rect 580908 206916 580960 206922
rect 580908 206858 580960 206864
rect 581000 205828 581052 205834
rect 581000 205770 581052 205776
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578330 203280 578386 203289
rect 578330 203215 578386 203224
rect 578344 202910 578372 203215
rect 578332 202904 578384 202910
rect 578332 202846 578384 202852
rect 580264 202904 580316 202910
rect 580264 202846 580316 202852
rect 578790 200832 578846 200841
rect 578790 200767 578846 200776
rect 578804 200190 578832 200767
rect 578792 200184 578844 200190
rect 578792 200126 578844 200132
rect 580276 200054 580304 202846
rect 581012 202842 581040 205770
rect 581000 202836 581052 202842
rect 581000 202778 581052 202784
rect 580264 200048 580316 200054
rect 580264 199990 580316 199996
rect 579526 198928 579582 198937
rect 579526 198863 579582 198872
rect 579540 198762 579568 198863
rect 579528 198756 579580 198762
rect 579528 198698 579580 198704
rect 578514 196480 578570 196489
rect 578514 196415 578570 196424
rect 578528 196042 578556 196415
rect 578516 196036 578568 196042
rect 578516 195978 578568 195984
rect 579526 194984 579582 194993
rect 579526 194919 579582 194928
rect 579540 194614 579568 194919
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 579526 192264 579582 192273
rect 579526 192199 579582 192208
rect 579540 191894 579568 192199
rect 579528 191888 579580 191894
rect 579528 191830 579580 191836
rect 579526 190768 579582 190777
rect 579526 190703 579582 190712
rect 579540 190534 579568 190703
rect 579528 190528 579580 190534
rect 579528 190470 579580 190476
rect 579526 188048 579582 188057
rect 579526 187983 579582 187992
rect 579540 187746 579568 187983
rect 579528 187740 579580 187746
rect 579528 187682 579580 187688
rect 579528 186312 579580 186318
rect 579526 186280 579528 186289
rect 579580 186280 579582 186289
rect 579526 186215 579582 186224
rect 579528 184884 579580 184890
rect 579528 184826 579580 184832
rect 579540 184385 579568 184826
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 579528 182164 579580 182170
rect 579528 182106 579580 182112
rect 579540 181937 579568 182106
rect 579526 181928 579582 181937
rect 579526 181863 579582 181872
rect 578792 180804 578844 180810
rect 578792 180746 578844 180752
rect 578804 180169 578832 180746
rect 578790 180160 578846 180169
rect 578790 180095 578846 180104
rect 578792 178084 578844 178090
rect 578792 178026 578844 178032
rect 578804 175137 578832 178026
rect 579528 177948 579580 177954
rect 579528 177890 579580 177896
rect 579540 177721 579568 177890
rect 579526 177712 579582 177721
rect 579526 177647 579582 177656
rect 579988 175296 580040 175302
rect 579988 175238 580040 175244
rect 578790 175128 578846 175137
rect 578790 175063 578846 175072
rect 578424 174548 578476 174554
rect 578424 174490 578476 174496
rect 578436 173505 578464 174490
rect 578422 173496 578478 173505
rect 578422 173431 578478 173440
rect 580000 172922 580028 175238
rect 578240 172916 578292 172922
rect 578240 172858 578292 172864
rect 579988 172916 580040 172922
rect 579988 172858 580040 172864
rect 578252 171057 578280 172858
rect 580908 172576 580960 172582
rect 580908 172518 580960 172524
rect 580264 171148 580316 171154
rect 580264 171090 580316 171096
rect 578238 171048 578294 171057
rect 578238 170983 578294 170992
rect 578700 169788 578752 169794
rect 578700 169730 578752 169736
rect 578712 169289 578740 169730
rect 578698 169280 578754 169289
rect 578698 169215 578754 169224
rect 580276 167346 580304 171090
rect 580920 169794 580948 172518
rect 580908 169788 580960 169794
rect 580908 169730 580960 169736
rect 578240 167340 578292 167346
rect 578240 167282 578292 167288
rect 580264 167340 580316 167346
rect 580264 167282 580316 167288
rect 578252 166977 578280 167282
rect 579988 167068 580040 167074
rect 579988 167010 580040 167016
rect 578238 166968 578294 166977
rect 578238 166903 578294 166912
rect 579528 166320 579580 166326
rect 579528 166262 579580 166268
rect 579344 165232 579396 165238
rect 579344 165174 579396 165180
rect 578240 163668 578292 163674
rect 578240 163610 578292 163616
rect 578252 159905 578280 163610
rect 579356 162761 579384 165174
rect 579540 164529 579568 166262
rect 579526 164520 579582 164529
rect 579526 164455 579582 164464
rect 580000 163674 580028 167010
rect 579988 163668 580040 163674
rect 579988 163610 580040 163616
rect 580908 162920 580960 162926
rect 580908 162862 580960 162868
rect 579342 162752 579398 162761
rect 578424 162716 578476 162722
rect 579342 162687 579398 162696
rect 578424 162658 578476 162664
rect 578238 159896 578294 159905
rect 578238 159831 578294 159840
rect 578436 158409 578464 162658
rect 580540 161492 580592 161498
rect 580540 161434 580592 161440
rect 578884 158772 578936 158778
rect 578884 158714 578936 158720
rect 578422 158400 578478 158409
rect 578422 158335 578478 158344
rect 578896 155961 578924 158714
rect 578882 155952 578938 155961
rect 578882 155887 578938 155896
rect 580552 154834 580580 161434
rect 580724 160132 580776 160138
rect 580724 160074 580776 160080
rect 578332 154828 578384 154834
rect 578332 154770 578384 154776
rect 580540 154828 580592 154834
rect 580540 154770 580592 154776
rect 578344 153649 578372 154770
rect 578330 153640 578386 153649
rect 578330 153575 578386 153584
rect 580736 152794 580764 160074
rect 580920 158778 580948 162862
rect 580908 158772 580960 158778
rect 580908 158714 580960 158720
rect 578240 152788 578292 152794
rect 578240 152730 578292 152736
rect 580724 152788 580776 152794
rect 580724 152730 580776 152736
rect 578252 151745 578280 152730
rect 580264 151836 580316 151842
rect 580264 151778 580316 151784
rect 578238 151736 578294 151745
rect 578238 151671 578294 151680
rect 578884 150612 578936 150618
rect 578884 150554 578936 150560
rect 578896 149705 578924 150554
rect 578882 149696 578938 149705
rect 578882 149631 578938 149640
rect 579528 148368 579580 148374
rect 579528 148310 579580 148316
rect 579540 147529 579568 148310
rect 579526 147520 579582 147529
rect 579526 147455 579582 147464
rect 578884 146328 578936 146334
rect 578884 146270 578936 146276
rect 578608 140752 578660 140758
rect 578608 140694 578660 140700
rect 578620 140593 578648 140694
rect 578606 140584 578662 140593
rect 578606 140519 578662 140528
rect 578608 139324 578660 139330
rect 578608 139266 578660 139272
rect 578620 138825 578648 139266
rect 578606 138816 578662 138825
rect 578606 138751 578662 138760
rect 578896 136649 578924 146270
rect 579252 144696 579304 144702
rect 579250 144664 579252 144673
rect 579304 144664 579306 144673
rect 579250 144599 579306 144608
rect 579528 143472 579580 143478
rect 579528 143414 579580 143420
rect 579540 143041 579568 143414
rect 579526 143032 579582 143041
rect 579526 142967 579582 142976
rect 580276 140758 580304 151778
rect 580448 140820 580500 140826
rect 580448 140762 580500 140768
rect 580264 140752 580316 140758
rect 580264 140694 580316 140700
rect 579528 138712 579580 138718
rect 579528 138654 579580 138660
rect 579068 137352 579120 137358
rect 579068 137294 579120 137300
rect 578882 136640 578938 136649
rect 578882 136575 578938 136584
rect 579080 132297 579108 137294
rect 579540 134473 579568 138654
rect 580264 134564 580316 134570
rect 580264 134506 580316 134512
rect 579526 134464 579582 134473
rect 579526 134399 579582 134408
rect 579066 132288 579122 132297
rect 579066 132223 579122 132232
rect 578884 131164 578936 131170
rect 578884 131106 578936 131112
rect 578896 129713 578924 131106
rect 578882 129704 578938 129713
rect 578882 129639 578938 129648
rect 579528 129056 579580 129062
rect 579528 128998 579580 129004
rect 579540 127945 579568 128998
rect 579526 127936 579582 127945
rect 579526 127871 579582 127880
rect 579068 127016 579120 127022
rect 579068 126958 579120 126964
rect 578332 125656 578384 125662
rect 578332 125598 578384 125604
rect 578344 125361 578372 125598
rect 578330 125352 578386 125361
rect 578330 125287 578386 125296
rect 578424 123616 578476 123622
rect 578422 123584 578424 123593
rect 578476 123584 578478 123593
rect 578422 123519 578478 123528
rect 578884 122188 578936 122194
rect 578884 122130 578936 122136
rect 578896 121417 578924 122130
rect 578882 121408 578938 121417
rect 578882 121343 578938 121352
rect 578516 118448 578568 118454
rect 578514 118416 578516 118425
rect 578568 118416 578570 118425
rect 578514 118351 578570 118360
rect 578332 108724 578384 108730
rect 578332 108666 578384 108672
rect 578344 108361 578372 108666
rect 578330 108352 578386 108361
rect 578330 108287 578386 108296
rect 578884 107636 578936 107642
rect 578884 107578 578936 107584
rect 578608 99272 578660 99278
rect 578606 99240 578608 99249
rect 578660 99240 578662 99249
rect 578606 99175 578662 99184
rect 577504 99136 577556 99142
rect 577504 99078 577556 99084
rect 578332 97980 578384 97986
rect 578332 97922 578384 97928
rect 578344 97481 578372 97922
rect 578330 97472 578386 97481
rect 578330 97407 578386 97416
rect 578516 93492 578568 93498
rect 578516 93434 578568 93440
rect 578528 93129 578556 93434
rect 578514 93120 578570 93129
rect 578514 93055 578570 93064
rect 578896 80073 578924 107578
rect 579080 105913 579108 126958
rect 580276 118454 580304 134506
rect 580460 125662 580488 140762
rect 580448 125656 580500 125662
rect 580448 125598 580500 125604
rect 580448 124228 580500 124234
rect 580448 124170 580500 124176
rect 580264 118448 580316 118454
rect 580264 118390 580316 118396
rect 579528 116952 579580 116958
rect 579526 116920 579528 116929
rect 579580 116920 579582 116929
rect 579526 116855 579582 116864
rect 579252 114504 579304 114510
rect 579250 114472 579252 114481
rect 579304 114472 579306 114481
rect 579250 114407 579306 114416
rect 579528 112872 579580 112878
rect 579528 112814 579580 112820
rect 579540 112577 579568 112814
rect 579526 112568 579582 112577
rect 579526 112503 579582 112512
rect 579344 110152 579396 110158
rect 579342 110120 579344 110129
rect 579396 110120 579398 110129
rect 579342 110055 579398 110064
rect 579066 105904 579122 105913
rect 579066 105839 579122 105848
rect 580264 104916 580316 104922
rect 580264 104858 580316 104864
rect 579528 103488 579580 103494
rect 579528 103430 579580 103436
rect 579540 103329 579568 103430
rect 579526 103320 579582 103329
rect 579526 103255 579582 103264
rect 579528 101856 579580 101862
rect 579528 101798 579580 101804
rect 579540 101697 579568 101798
rect 579526 101688 579582 101697
rect 579526 101623 579582 101632
rect 579068 99408 579120 99414
rect 579068 99350 579120 99356
rect 579080 90953 579108 99350
rect 579528 95056 579580 95062
rect 579526 95024 579528 95033
rect 579580 95024 579582 95033
rect 579526 94959 579582 94968
rect 579344 91112 579396 91118
rect 579344 91054 579396 91060
rect 579066 90944 579122 90953
rect 579066 90879 579122 90888
rect 579356 86465 579384 91054
rect 579528 88120 579580 88126
rect 579526 88088 579528 88097
rect 579580 88088 579582 88097
rect 579526 88023 579582 88032
rect 579342 86456 579398 86465
rect 579342 86391 579398 86400
rect 579160 84176 579212 84182
rect 579160 84118 579212 84124
rect 579172 84017 579200 84118
rect 579158 84008 579214 84017
rect 579158 83943 579214 83952
rect 579068 82408 579120 82414
rect 579068 82350 579120 82356
rect 579080 82249 579108 82350
rect 579066 82240 579122 82249
rect 579066 82175 579122 82184
rect 579528 82136 579580 82142
rect 579528 82078 579580 82084
rect 578882 80064 578938 80073
rect 578882 79999 578938 80008
rect 579068 79348 579120 79354
rect 579068 79290 579120 79296
rect 578240 75880 578292 75886
rect 578240 75822 578292 75828
rect 578252 75585 578280 75822
rect 578238 75576 578294 75585
rect 578238 75511 578294 75520
rect 579080 73137 579108 79290
rect 579540 77897 579568 82078
rect 579526 77888 579582 77897
rect 579526 77823 579582 77832
rect 580276 75886 580304 104858
rect 580460 99278 580488 124170
rect 580632 122052 580684 122058
rect 580632 121994 580684 122000
rect 580644 108730 580672 121994
rect 581656 114510 581684 208558
rect 582300 205562 582328 209782
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208049 589504 208286
rect 589462 208040 589518 208049
rect 589462 207975 589518 207984
rect 589464 206916 589516 206922
rect 589464 206858 589516 206864
rect 589476 206417 589504 206858
rect 589462 206408 589518 206417
rect 589462 206343 589518 206352
rect 582288 205556 582340 205562
rect 582288 205498 582340 205504
rect 589464 205556 589516 205562
rect 589464 205498 589516 205504
rect 589476 204785 589504 205498
rect 589462 204776 589518 204785
rect 589462 204711 589518 204720
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203153 589504 204206
rect 589462 203144 589518 203153
rect 589462 203079 589518 203088
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 201521 589504 202778
rect 589462 201512 589518 201521
rect 589462 201447 589518 201456
rect 590384 200184 590436 200190
rect 590384 200126 590436 200132
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 589464 198756 589516 198762
rect 589464 198698 589516 198704
rect 589476 196625 589504 198698
rect 590396 198257 590424 200126
rect 590382 198248 590438 198257
rect 590382 198183 590438 198192
rect 589462 196616 589518 196625
rect 589462 196551 589518 196560
rect 589280 196036 589332 196042
rect 589280 195978 589332 195984
rect 589292 194993 589320 195978
rect 589278 194984 589334 194993
rect 589278 194919 589334 194928
rect 589464 194608 589516 194614
rect 589464 194550 589516 194556
rect 589476 193361 589504 194550
rect 589462 193352 589518 193361
rect 589462 193287 589518 193296
rect 589464 191888 589516 191894
rect 589464 191830 589516 191836
rect 589476 191729 589504 191830
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 590568 190528 590620 190534
rect 590568 190470 590620 190476
rect 590580 190097 590608 190470
rect 590566 190088 590622 190097
rect 590566 190023 590622 190032
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 589464 187740 589516 187746
rect 589464 187682 589516 187688
rect 589476 186833 589504 187682
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 589660 186318 589688 188391
rect 589648 186312 589700 186318
rect 589648 186254 589700 186260
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184890 589504 185127
rect 589464 184884 589516 184890
rect 589464 184826 589516 184832
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182170 589504 183495
rect 589464 182164 589516 182170
rect 589464 182106 589516 182112
rect 590566 181928 590622 181937
rect 590566 181863 590622 181872
rect 590580 180810 590608 181863
rect 590568 180804 590620 180810
rect 590568 180746 590620 180752
rect 589646 180296 589702 180305
rect 589646 180231 589702 180240
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 589660 177954 589688 180231
rect 589648 177948 589700 177954
rect 589648 177890 589700 177896
rect 589646 177032 589702 177041
rect 589646 176967 589702 176976
rect 589462 175400 589518 175409
rect 589462 175335 589464 175344
rect 589516 175335 589518 175344
rect 589464 175306 589516 175312
rect 589660 174554 589688 176967
rect 589648 174548 589700 174554
rect 589648 174490 589700 174496
rect 589462 173768 589518 173777
rect 589462 173703 589518 173712
rect 589476 172582 589504 173703
rect 589464 172576 589516 172582
rect 589464 172518 589516 172524
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 589646 170504 589702 170513
rect 589646 170439 589702 170448
rect 589462 168872 589518 168881
rect 589462 168807 589518 168816
rect 589476 168434 589504 168807
rect 582380 168428 582432 168434
rect 582380 168370 582432 168376
rect 589464 168428 589516 168434
rect 589464 168370 589516 168376
rect 582392 165238 582420 168370
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 589660 166326 589688 170439
rect 589648 166320 589700 166326
rect 589648 166262 589700 166268
rect 589462 165608 589518 165617
rect 589462 165543 589518 165552
rect 582380 165232 582432 165238
rect 582380 165174 582432 165180
rect 589476 164286 589504 165543
rect 582472 164280 582524 164286
rect 582472 164222 582524 164228
rect 589464 164280 589516 164286
rect 589464 164222 589516 164228
rect 582484 162722 582512 164222
rect 589462 163976 589518 163985
rect 589462 163911 589518 163920
rect 589476 162926 589504 163911
rect 589464 162920 589516 162926
rect 589464 162862 589516 162868
rect 582472 162716 582524 162722
rect 582472 162658 582524 162664
rect 589462 162344 589518 162353
rect 589462 162279 589518 162288
rect 589476 161498 589504 162279
rect 589464 161492 589516 161498
rect 589464 161434 589516 161440
rect 589462 160712 589518 160721
rect 589462 160647 589518 160656
rect 589476 160138 589504 160647
rect 589464 160132 589516 160138
rect 589464 160074 589516 160080
rect 589462 159080 589518 159089
rect 589462 159015 589518 159024
rect 589476 158778 589504 159015
rect 585784 158772 585836 158778
rect 585784 158714 585836 158720
rect 589464 158772 589516 158778
rect 589464 158714 589516 158720
rect 584404 154624 584456 154630
rect 584404 154566 584456 154572
rect 583024 153264 583076 153270
rect 583024 153206 583076 153212
rect 583036 143478 583064 153206
rect 584416 144702 584444 154566
rect 585796 150618 585824 158714
rect 589278 157448 589334 157457
rect 587164 157412 587216 157418
rect 589278 157383 589280 157392
rect 587164 157354 587216 157360
rect 589332 157383 589334 157392
rect 589280 157354 589332 157360
rect 585784 150612 585836 150618
rect 585784 150554 585836 150560
rect 585140 149116 585192 149122
rect 585140 149058 585192 149064
rect 585152 146334 585180 149058
rect 587176 148374 587204 157354
rect 589462 155816 589518 155825
rect 589462 155751 589518 155760
rect 589476 154630 589504 155751
rect 589464 154624 589516 154630
rect 589464 154566 589516 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589462 152552 589518 152561
rect 589462 152487 589518 152496
rect 589476 151842 589504 152487
rect 589464 151836 589516 151842
rect 589464 151778 589516 151784
rect 590014 150920 590070 150929
rect 590014 150855 590070 150864
rect 589462 149288 589518 149297
rect 589462 149223 589518 149232
rect 589476 149122 589504 149223
rect 589464 149116 589516 149122
rect 589464 149058 589516 149064
rect 587164 148368 587216 148374
rect 587164 148310 587216 148316
rect 588542 147656 588598 147665
rect 588542 147591 588598 147600
rect 585140 146328 585192 146334
rect 585140 146270 585192 146276
rect 584772 144968 584824 144974
rect 584772 144910 584824 144916
rect 584404 144696 584456 144702
rect 584404 144638 584456 144644
rect 583024 143472 583076 143478
rect 583024 143414 583076 143420
rect 583024 139460 583076 139466
rect 583024 139402 583076 139408
rect 581828 131300 581880 131306
rect 581828 131242 581880 131248
rect 581644 114504 581696 114510
rect 581644 114446 581696 114452
rect 581644 110492 581696 110498
rect 581644 110434 581696 110440
rect 580632 108724 580684 108730
rect 580632 108666 580684 108672
rect 580448 99272 580500 99278
rect 580448 99214 580500 99220
rect 581656 84182 581684 110434
rect 581840 110158 581868 131242
rect 583036 123622 583064 139402
rect 584784 137358 584812 144910
rect 585968 143608 586020 143614
rect 585968 143550 586020 143556
rect 584772 137352 584824 137358
rect 584772 137294 584824 137300
rect 584588 136672 584640 136678
rect 584588 136614 584640 136620
rect 583208 129192 583260 129198
rect 583208 129134 583260 129140
rect 583024 123616 583076 123622
rect 583024 123558 583076 123564
rect 583220 116958 583248 129134
rect 584404 122868 584456 122874
rect 584404 122810 584456 122816
rect 583208 116952 583260 116958
rect 583208 116894 583260 116900
rect 583208 115252 583260 115258
rect 583208 115194 583260 115200
rect 583024 113212 583076 113218
rect 583024 113154 583076 113160
rect 581828 110152 581880 110158
rect 581828 110094 581880 110100
rect 581644 84176 581696 84182
rect 581644 84118 581696 84124
rect 583036 82414 583064 113154
rect 583220 95062 583248 115194
rect 584416 101862 584444 122810
rect 584600 122194 584628 136614
rect 585784 132524 585836 132530
rect 585784 132466 585836 132472
rect 584588 122188 584640 122194
rect 584588 122130 584640 122136
rect 585796 112878 585824 132466
rect 585980 131170 586008 143550
rect 587164 142452 587216 142458
rect 587164 142394 587216 142400
rect 585968 131164 586020 131170
rect 585968 131106 586020 131112
rect 587176 129062 587204 142394
rect 588556 138718 588584 147591
rect 589462 146024 589518 146033
rect 589462 145959 589518 145968
rect 589476 144974 589504 145959
rect 589464 144968 589516 144974
rect 589464 144910 589516 144916
rect 589462 144392 589518 144401
rect 589462 144327 589518 144336
rect 589476 143614 589504 144327
rect 589464 143608 589516 143614
rect 589464 143550 589516 143556
rect 589830 142760 589886 142769
rect 589830 142695 589886 142704
rect 589844 142458 589872 142695
rect 589832 142452 589884 142458
rect 589832 142394 589884 142400
rect 590028 142154 590056 150855
rect 589936 142126 590056 142154
rect 589462 141128 589518 141137
rect 589462 141063 589518 141072
rect 589476 140826 589504 141063
rect 589464 140820 589516 140826
rect 589464 140762 589516 140768
rect 589462 139496 589518 139505
rect 589462 139431 589464 139440
rect 589516 139431 589518 139440
rect 589464 139402 589516 139408
rect 589936 139330 589964 142126
rect 589924 139324 589976 139330
rect 589924 139266 589976 139272
rect 588544 138712 588596 138718
rect 588544 138654 588596 138660
rect 589462 137864 589518 137873
rect 589462 137799 589518 137808
rect 589476 136678 589504 137799
rect 589464 136672 589516 136678
rect 589464 136614 589516 136620
rect 589462 136232 589518 136241
rect 589462 136167 589518 136176
rect 589476 134570 589504 136167
rect 590382 134600 590438 134609
rect 589464 134564 589516 134570
rect 590382 134535 590438 134544
rect 589464 134506 589516 134512
rect 589462 132968 589518 132977
rect 589462 132903 589518 132912
rect 589476 132530 589504 132903
rect 589464 132524 589516 132530
rect 589464 132466 589516 132472
rect 589462 131336 589518 131345
rect 589462 131271 589464 131280
rect 589516 131271 589518 131280
rect 589464 131242 589516 131248
rect 588542 129704 588598 129713
rect 588542 129639 588598 129648
rect 587164 129056 587216 129062
rect 587164 128998 587216 129004
rect 587348 118720 587400 118726
rect 587348 118662 587400 118668
rect 586152 116000 586204 116006
rect 586152 115942 586204 115948
rect 585784 112872 585836 112878
rect 585784 112814 585836 112820
rect 585968 112464 586020 112470
rect 585968 112406 586020 112412
rect 584588 109064 584640 109070
rect 584588 109006 584640 109012
rect 584404 101856 584456 101862
rect 584404 101798 584456 101804
rect 584404 100156 584456 100162
rect 584404 100098 584456 100104
rect 583208 95056 583260 95062
rect 583208 94998 583260 95004
rect 583024 82408 583076 82414
rect 583024 82350 583076 82356
rect 581642 77888 581698 77897
rect 581642 77823 581698 77832
rect 580264 75880 580316 75886
rect 580264 75822 580316 75828
rect 579066 73128 579122 73137
rect 579066 73063 579122 73072
rect 578884 72480 578936 72486
rect 578884 72422 578936 72428
rect 577504 60036 577556 60042
rect 577504 59978 577556 59984
rect 576124 58676 576176 58682
rect 576124 58618 576176 58624
rect 574928 57248 574980 57254
rect 574928 57190 574980 57196
rect 574560 56024 574612 56030
rect 574560 55966 574612 55972
rect 574572 53990 574600 55966
rect 574744 55888 574796 55894
rect 574744 55830 574796 55836
rect 574756 54126 574784 55830
rect 574744 54120 574796 54126
rect 574744 54062 574796 54068
rect 574560 53984 574612 53990
rect 574560 53926 574612 53932
rect 574940 53854 574968 57190
rect 576136 55049 576164 58618
rect 576122 55040 576178 55049
rect 576122 54975 576178 54984
rect 577516 54233 577544 59978
rect 578896 54505 578924 72422
rect 579068 71392 579120 71398
rect 579068 71334 579120 71340
rect 579080 71233 579108 71334
rect 579066 71224 579122 71233
rect 579066 71159 579122 71168
rect 580264 68332 580316 68338
rect 580264 68274 580316 68280
rect 580276 54777 580304 68274
rect 580262 54768 580318 54777
rect 580262 54703 580318 54712
rect 578882 54496 578938 54505
rect 578882 54431 578938 54440
rect 581656 54262 581684 77823
rect 584416 71398 584444 100098
rect 584600 91118 584628 109006
rect 585980 93498 586008 112406
rect 586164 99414 586192 115942
rect 587164 106344 587216 106350
rect 587164 106286 587216 106292
rect 586152 99408 586204 99414
rect 586152 99350 586204 99356
rect 585968 93492 586020 93498
rect 585968 93434 586020 93440
rect 584588 91112 584640 91118
rect 584588 91054 584640 91060
rect 585140 89004 585192 89010
rect 585140 88946 585192 88952
rect 585152 88126 585180 88946
rect 585140 88120 585192 88126
rect 585140 88062 585192 88068
rect 587176 82142 587204 106286
rect 587360 97986 587388 118662
rect 588556 103494 588584 129639
rect 590396 129198 590424 134535
rect 590384 129192 590436 129198
rect 590384 129134 590436 129140
rect 589462 128072 589518 128081
rect 589462 128007 589518 128016
rect 589476 127022 589504 128007
rect 589464 127016 589516 127022
rect 589464 126958 589516 126964
rect 589922 126440 589978 126449
rect 589922 126375 589978 126384
rect 589462 124808 589518 124817
rect 589462 124743 589518 124752
rect 589476 124234 589504 124743
rect 589464 124228 589516 124234
rect 589464 124170 589516 124176
rect 589462 123176 589518 123185
rect 589462 123111 589518 123120
rect 589476 122874 589504 123111
rect 589464 122868 589516 122874
rect 589464 122810 589516 122816
rect 589936 122058 589964 126375
rect 589924 122052 589976 122058
rect 589924 121994 589976 122000
rect 590014 121544 590070 121553
rect 590014 121479 590070 121488
rect 589646 119912 589702 119921
rect 589646 119847 589702 119856
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 589660 115258 589688 119847
rect 590028 118726 590056 121479
rect 590016 118720 590068 118726
rect 590016 118662 590068 118668
rect 590106 118280 590162 118289
rect 590106 118215 590162 118224
rect 589648 115252 589700 115258
rect 589648 115194 589700 115200
rect 589462 113384 589518 113393
rect 589462 113319 589518 113328
rect 589476 113218 589504 113319
rect 589464 113212 589516 113218
rect 589464 113154 589516 113160
rect 590120 112470 590148 118215
rect 590290 115016 590346 115025
rect 590290 114951 590346 114960
rect 590108 112464 590160 112470
rect 590108 112406 590160 112412
rect 589462 111752 589518 111761
rect 589462 111687 589518 111696
rect 589476 110498 589504 111687
rect 589464 110492 589516 110498
rect 589464 110434 589516 110440
rect 589278 110120 589334 110129
rect 589278 110055 589334 110064
rect 589292 109070 589320 110055
rect 589280 109064 589332 109070
rect 589280 109006 589332 109012
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589830 106856 589886 106865
rect 589830 106791 589886 106800
rect 589844 106350 589872 106791
rect 589832 106344 589884 106350
rect 589832 106286 589884 106292
rect 589462 105224 589518 105233
rect 589462 105159 589518 105168
rect 589476 104922 589504 105159
rect 589464 104916 589516 104922
rect 589464 104858 589516 104864
rect 588726 103592 588782 103601
rect 588726 103527 588782 103536
rect 588544 103488 588596 103494
rect 588544 103430 588596 103436
rect 587348 97980 587400 97986
rect 587348 97922 587400 97928
rect 587164 82136 587216 82142
rect 587164 82078 587216 82084
rect 588740 79354 588768 103527
rect 590304 103514 590332 114951
rect 589936 103486 590332 103514
rect 589462 101960 589518 101969
rect 589462 101895 589518 101904
rect 589476 100162 589504 101895
rect 589464 100156 589516 100162
rect 589464 100098 589516 100104
rect 589936 89010 589964 103486
rect 589924 89004 589976 89010
rect 589924 88946 589976 88952
rect 588728 79348 588780 79354
rect 588728 79290 588780 79296
rect 584404 71392 584456 71398
rect 584404 71334 584456 71340
rect 581644 54256 581696 54262
rect 577502 54224 577558 54233
rect 581644 54198 581696 54204
rect 577502 54159 577558 54168
rect 574928 53848 574980 53854
rect 574928 53790 574980 53796
rect 459834 53680 459890 53689
rect 459834 53615 459890 53624
rect 460754 53680 460810 53689
rect 460754 53615 460810 53624
rect 461674 53680 461730 53689
rect 461674 53615 461730 53624
rect 462594 53680 462650 53689
rect 462594 53615 462650 53624
rect 463240 53644 463292 53650
rect 459468 53508 459520 53514
rect 459468 53450 459520 53456
rect 50528 53236 50580 53242
rect 50528 53178 50580 53184
rect 130384 53236 130436 53242
rect 130384 53178 130436 53184
rect 50344 51876 50396 51882
rect 50344 51818 50396 51824
rect 129004 51876 129056 51882
rect 129004 51818 129056 51824
rect 129648 51876 129700 51882
rect 129648 51818 129700 51824
rect 128820 51740 128872 51746
rect 128820 51682 128872 51688
rect 49148 49156 49200 49162
rect 49148 49098 49200 49104
rect 45468 49020 45520 49026
rect 45468 48962 45520 48968
rect 128832 44810 128860 51682
rect 128820 44804 128872 44810
rect 128820 44746 128872 44752
rect 129016 44470 129044 51818
rect 129280 49156 129332 49162
rect 129280 49098 129332 49104
rect 129292 44946 129320 49098
rect 129464 49020 129516 49026
rect 129464 48962 129516 48968
rect 129476 45422 129504 48962
rect 129464 45416 129516 45422
rect 129464 45358 129516 45364
rect 129660 45082 129688 51818
rect 129648 45076 129700 45082
rect 129648 45018 129700 45024
rect 129280 44940 129332 44946
rect 129280 44882 129332 44888
rect 129004 44464 129056 44470
rect 129004 44406 129056 44412
rect 43628 44328 43680 44334
rect 130396 44305 130424 53178
rect 312360 53168 312412 53174
rect 312018 53116 312360 53122
rect 312018 53110 312412 53116
rect 313740 53168 313792 53174
rect 316316 53168 316368 53174
rect 313792 53116 314042 53122
rect 313740 53110 314042 53116
rect 130568 53100 130620 53106
rect 312018 53094 312400 53110
rect 313752 53108 314042 53110
rect 316020 53116 316316 53122
rect 316020 53110 316368 53116
rect 317696 53168 317748 53174
rect 317748 53116 318380 53122
rect 317696 53110 318380 53116
rect 313752 53094 314056 53108
rect 316020 53094 316356 53110
rect 317708 53094 318380 53110
rect 130568 53042 130620 53048
rect 130580 46102 130608 53042
rect 130752 52012 130804 52018
rect 130752 51954 130804 51960
rect 130568 46096 130620 46102
rect 130568 46038 130620 46044
rect 130764 45558 130792 51954
rect 314028 50386 314056 53094
rect 318352 50522 318380 53094
rect 459480 52578 459508 53450
rect 459848 52578 459876 53615
rect 460386 53408 460442 53417
rect 460386 53343 460442 53352
rect 460400 52578 460428 53343
rect 460768 52578 460796 53615
rect 461308 52964 461360 52970
rect 461308 52906 461360 52912
rect 461320 52578 461348 52906
rect 461688 52578 461716 53615
rect 461906 52828 461958 52834
rect 461906 52770 461958 52776
rect 459172 52550 459508 52578
rect 459632 52550 459876 52578
rect 460092 52550 460428 52578
rect 460552 52550 460796 52578
rect 461012 52550 461348 52578
rect 461472 52550 461716 52578
rect 461918 52564 461946 52770
rect 462608 52578 462636 53615
rect 463240 53586 463292 53592
rect 464068 53644 464120 53650
rect 464068 53586 464120 53592
rect 464252 53644 464304 53650
rect 464252 53586 464304 53592
rect 465264 53644 465316 53650
rect 465264 53586 465316 53592
rect 465448 53644 465500 53650
rect 465448 53586 465500 53592
rect 466368 53644 466420 53650
rect 466368 53586 466420 53592
rect 467104 53644 467156 53650
rect 467104 53586 467156 53592
rect 471060 53644 471112 53650
rect 471060 53586 471112 53592
rect 463056 53372 463108 53378
rect 463056 53314 463108 53320
rect 463068 52578 463096 53314
rect 463252 53242 463280 53586
rect 463240 53236 463292 53242
rect 463240 53178 463292 53184
rect 463792 53236 463844 53242
rect 463792 53178 463844 53184
rect 463608 53100 463660 53106
rect 463608 53042 463660 53048
rect 463620 52578 463648 53042
rect 463804 52578 463832 53178
rect 462392 52550 462636 52578
rect 462852 52550 463096 52578
rect 463312 52550 463648 52578
rect 463772 52550 463832 52578
rect 464080 52578 464108 53586
rect 464264 53106 464292 53586
rect 464988 53508 465040 53514
rect 464988 53450 465040 53456
rect 464252 53100 464304 53106
rect 464252 53042 464304 53048
rect 465000 52578 465028 53450
rect 465276 53224 465304 53586
rect 465460 53417 465488 53586
rect 465446 53408 465502 53417
rect 465446 53343 465502 53352
rect 465276 53196 465672 53224
rect 465448 53100 465500 53106
rect 465448 53042 465500 53048
rect 465460 52578 465488 53042
rect 465644 52578 465672 53196
rect 466380 53106 466408 53586
rect 466368 53100 466420 53106
rect 466368 53042 466420 53048
rect 467116 52834 467144 53586
rect 471072 52970 471100 53586
rect 471060 52964 471112 52970
rect 471060 52906 471112 52912
rect 467104 52828 467156 52834
rect 467104 52770 467156 52776
rect 464080 52550 464232 52578
rect 464692 52550 465028 52578
rect 465152 52550 465488 52578
rect 465612 52550 465672 52578
rect 318340 50516 318392 50522
rect 318340 50458 318392 50464
rect 458180 50516 458232 50522
rect 458180 50458 458232 50464
rect 131028 50380 131080 50386
rect 131028 50322 131080 50328
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 130752 45552 130804 45558
rect 130752 45494 130804 45500
rect 43628 44270 43680 44276
rect 130382 44296 130438 44305
rect 130382 44231 130438 44240
rect 43444 44192 43496 44198
rect 43444 44134 43496 44140
rect 131040 44062 131068 50322
rect 458192 47025 458220 50458
rect 544028 50386 544056 53108
rect 545684 53094 546020 53122
rect 547892 53094 548044 53122
rect 458364 50380 458416 50386
rect 458364 50322 458416 50328
rect 522948 50380 523000 50386
rect 522948 50322 523000 50328
rect 544016 50380 544068 50386
rect 544016 50322 544068 50328
rect 458178 47016 458234 47025
rect 458178 46951 458234 46960
rect 458376 46753 458404 50322
rect 522960 47841 522988 50322
rect 522946 47832 523002 47841
rect 522946 47767 523002 47776
rect 459172 47654 459232 47682
rect 459632 47654 459968 47682
rect 460092 47654 460152 47682
rect 460552 47654 460796 47682
rect 458362 46744 458418 46753
rect 142370 46702 142660 46730
rect 132316 46096 132368 46102
rect 132316 46038 132368 46044
rect 131672 44668 131724 44674
rect 131672 44610 131724 44616
rect 131684 44198 131712 44610
rect 132328 44292 132356 46038
rect 132592 45552 132644 45558
rect 132592 45494 132644 45500
rect 132604 44422 132632 45494
rect 132592 44416 132644 44422
rect 132592 44358 132644 44364
rect 132500 44304 132552 44310
rect 132776 44305 132828 44310
rect 142632 44305 142660 46702
rect 458362 46679 458418 46688
rect 132328 44264 132500 44292
rect 132500 44246 132552 44252
rect 132774 44304 132830 44305
rect 132774 44296 132776 44304
rect 132828 44296 132830 44304
rect 132774 44231 132830 44240
rect 142618 44296 142674 44305
rect 142618 44231 142674 44240
rect 131672 44192 131724 44198
rect 131672 44134 131724 44140
rect 255870 44160 255926 44169
rect 255870 44095 255926 44104
rect 131028 44056 131080 44062
rect 131028 43998 131080 44004
rect 255884 42838 255912 44095
rect 419722 43888 419778 43897
rect 419722 43823 419778 43832
rect 440238 43888 440294 43897
rect 440238 43823 440240 43832
rect 187332 42832 187384 42838
rect 187332 42774 187384 42780
rect 255872 42832 255924 42838
rect 255872 42774 255924 42780
rect 187344 42092 187372 42774
rect 307300 42764 307352 42770
rect 307300 42706 307352 42712
rect 307312 42106 307340 42706
rect 310428 42628 310480 42634
rect 310428 42570 310480 42576
rect 310440 42106 310468 42570
rect 419736 42364 419764 43823
rect 440292 43823 440294 43832
rect 441066 43888 441122 43897
rect 441066 43823 441068 43832
rect 440240 43794 440292 43800
rect 441120 43823 441122 43832
rect 441068 43794 441120 43800
rect 431224 42764 431276 42770
rect 431224 42706 431276 42712
rect 441068 42764 441120 42770
rect 441068 42706 441120 42712
rect 449164 42764 449216 42770
rect 449164 42706 449216 42712
rect 453580 42764 453632 42770
rect 453580 42706 453632 42712
rect 427084 42628 427136 42634
rect 427084 42570 427136 42576
rect 404452 42356 404504 42362
rect 404452 42298 404504 42304
rect 405188 42356 405240 42362
rect 405188 42298 405240 42304
rect 420736 42356 420788 42362
rect 420736 42298 420788 42304
rect 426900 42356 426952 42362
rect 426900 42298 426952 42304
rect 307004 42078 307340 42106
rect 310132 42078 310468 42106
rect 361946 41848 362002 41857
rect 361790 41806 361946 41834
rect 365166 41848 365222 41857
rect 364918 41806 365166 41834
rect 361946 41783 362002 41792
rect 365166 41783 365222 41792
rect 404464 41478 404492 42298
rect 405200 42106 405228 42298
rect 416686 42256 416742 42265
rect 416686 42191 416742 42200
rect 415582 42120 415638 42129
rect 405200 42078 405582 42106
rect 415426 42078 415582 42106
rect 416700 42106 416728 42191
rect 416622 42078 416728 42106
rect 415582 42055 415638 42064
rect 420748 41478 420776 42298
rect 426912 41478 426940 42298
rect 427096 42022 427124 42570
rect 431236 42022 431264 42706
rect 441080 42022 441108 42706
rect 441252 42628 441304 42634
rect 441252 42570 441304 42576
rect 446404 42628 446456 42634
rect 446404 42570 446456 42576
rect 427084 42016 427136 42022
rect 427084 41958 427136 41964
rect 431224 42016 431276 42022
rect 431224 41958 431276 41964
rect 441068 42016 441120 42022
rect 441068 41958 441120 41964
rect 441264 41886 441292 42570
rect 446218 42256 446274 42265
rect 446218 42191 446274 42200
rect 441252 41880 441304 41886
rect 441252 41822 441304 41828
rect 446232 41585 446260 42191
rect 446416 42022 446444 42570
rect 446404 42016 446456 42022
rect 446404 41958 446456 41964
rect 449176 41886 449204 42706
rect 453592 41886 453620 42706
rect 454500 42492 454552 42498
rect 454500 42434 454552 42440
rect 454512 42022 454540 42434
rect 454500 42016 454552 42022
rect 454500 41958 454552 41964
rect 449164 41880 449216 41886
rect 449164 41822 449216 41828
rect 453580 41880 453632 41886
rect 453580 41822 453632 41828
rect 446218 41576 446274 41585
rect 446218 41511 446274 41520
rect 459204 41478 459232 47654
rect 459940 42106 459968 47654
rect 460124 44169 460152 47654
rect 460110 44160 460166 44169
rect 460110 44095 460166 44104
rect 460768 43489 460796 47654
rect 460998 47410 461026 47668
rect 461472 47654 461808 47682
rect 461932 47654 461992 47682
rect 462392 47654 462728 47682
rect 462852 47654 462912 47682
rect 460952 47382 461026 47410
rect 460754 43480 460810 43489
rect 460754 43415 460810 43424
rect 460952 42401 460980 47382
rect 461780 42945 461808 47654
rect 461964 44305 461992 47654
rect 461950 44296 462006 44305
rect 461950 44231 462006 44240
rect 462700 43217 462728 47654
rect 462884 44033 462912 47654
rect 463068 47654 463312 47682
rect 462870 44024 462926 44033
rect 462870 43959 462926 43968
rect 462686 43208 462742 43217
rect 462686 43143 462742 43152
rect 461766 42936 461822 42945
rect 461766 42871 461822 42880
rect 463068 42498 463096 47654
rect 463758 47410 463786 47668
rect 464218 47410 464246 47668
rect 464692 47654 464752 47682
rect 463712 47382 463786 47410
rect 464172 47382 464246 47410
rect 463712 44305 463740 47382
rect 463698 44296 463754 44305
rect 463698 44231 463754 44240
rect 463974 42936 464030 42945
rect 463974 42871 464030 42880
rect 463988 42514 464016 42871
rect 464172 42770 464200 47382
rect 464724 44305 464752 47654
rect 465138 47410 465166 47668
rect 465092 47382 465166 47410
rect 465276 47654 465612 47682
rect 465092 47025 465120 47382
rect 465078 47016 465134 47025
rect 465078 46951 465134 46960
rect 465276 46753 465304 47654
rect 545684 47297 545712 53094
rect 547892 47569 547920 53094
rect 550008 48929 550036 53108
rect 549994 48920 550050 48929
rect 549994 48855 550050 48864
rect 552032 47841 552060 53108
rect 553688 53094 554024 53122
rect 553688 48113 553716 53094
rect 591316 51882 591344 212638
rect 591500 101697 591528 224159
rect 593972 223304 594024 223310
rect 593972 223246 594024 223252
rect 592040 222080 592092 222086
rect 592040 222022 592092 222028
rect 592052 221218 592080 222022
rect 591960 221190 592080 221218
rect 591960 221134 591988 221190
rect 591948 221128 592000 221134
rect 591948 221070 592000 221076
rect 592132 221128 592184 221134
rect 592132 221070 592184 221076
rect 592144 220946 592172 221070
rect 592052 220918 592172 220946
rect 592052 220862 592080 220918
rect 592040 220856 592092 220862
rect 592040 220798 592092 220804
rect 592684 212560 592736 212566
rect 592684 212502 592736 212508
rect 591486 101688 591542 101697
rect 591486 101623 591542 101632
rect 591304 51876 591356 51882
rect 591304 51818 591356 51824
rect 592696 51746 592724 212502
rect 593984 210202 594012 223246
rect 596640 222080 596692 222086
rect 596640 222022 596692 222028
rect 596824 222080 596876 222086
rect 596824 222022 596876 222028
rect 596652 220946 596680 222022
rect 596836 221406 596864 222022
rect 597020 221474 597048 224926
rect 610452 224874 611032 224890
rect 610452 224868 611044 224874
rect 610452 224862 610992 224868
rect 610452 224670 610480 224862
rect 610992 224810 611044 224816
rect 614948 224868 615000 224874
rect 614948 224810 615000 224816
rect 610808 224800 610860 224806
rect 610808 224742 610860 224748
rect 610440 224664 610492 224670
rect 610440 224606 610492 224612
rect 610624 224664 610676 224670
rect 610624 224606 610676 224612
rect 610636 223922 610664 224606
rect 610820 223922 610848 224742
rect 610624 223916 610676 223922
rect 610624 223858 610676 223864
rect 610808 223916 610860 223922
rect 610808 223858 610860 223864
rect 605012 222080 605064 222086
rect 605012 222022 605064 222028
rect 601976 221604 602028 221610
rect 601976 221546 602028 221552
rect 599490 221504 599546 221513
rect 597008 221468 597060 221474
rect 599490 221439 599546 221448
rect 597008 221410 597060 221416
rect 596824 221400 596876 221406
rect 596824 221342 596876 221348
rect 596652 220918 596956 220946
rect 596928 220862 596956 220918
rect 596916 220856 596968 220862
rect 596916 220798 596968 220804
rect 596732 220788 596784 220794
rect 596732 220730 596784 220736
rect 595628 219768 595680 219774
rect 595628 219710 595680 219716
rect 595640 219366 595668 219710
rect 595628 219360 595680 219366
rect 595628 219302 595680 219308
rect 595996 218340 596048 218346
rect 595996 218282 596048 218288
rect 595166 217288 595222 217297
rect 595166 217223 595222 217232
rect 594800 213240 594852 213246
rect 594800 213182 594852 213188
rect 594812 210202 594840 213182
rect 595180 210202 595208 217223
rect 595718 217016 595774 217025
rect 595718 216951 595774 216960
rect 595732 210202 595760 216951
rect 596008 216782 596036 218282
rect 596548 217184 596600 217190
rect 596548 217126 596600 217132
rect 596560 216918 596588 217126
rect 596364 216912 596416 216918
rect 596364 216854 596416 216860
rect 596548 216912 596600 216918
rect 596548 216854 596600 216860
rect 595996 216776 596048 216782
rect 595996 216718 596048 216724
rect 596376 210202 596404 216854
rect 596744 210202 596772 220730
rect 597560 219224 597612 219230
rect 597560 219166 597612 219172
rect 596916 217456 596968 217462
rect 596916 217398 596968 217404
rect 596928 217190 596956 217398
rect 596916 217184 596968 217190
rect 596916 217126 596968 217132
rect 597572 210202 597600 219166
rect 598112 218748 598164 218754
rect 598112 218690 598164 218696
rect 598124 217326 598152 218690
rect 597928 217320 597980 217326
rect 597928 217262 597980 217268
rect 598112 217320 598164 217326
rect 598112 217262 598164 217268
rect 597940 210202 597968 217262
rect 598480 216912 598532 216918
rect 598480 216854 598532 216860
rect 598492 210202 598520 216854
rect 599030 215656 599086 215665
rect 599030 215591 599086 215600
rect 599044 210202 599072 215591
rect 599504 210202 599532 221439
rect 600870 221232 600926 221241
rect 600870 221167 600926 221176
rect 600412 221128 600464 221134
rect 600412 221070 600464 221076
rect 600424 210458 600452 221070
rect 600688 220856 600740 220862
rect 600688 220798 600740 220804
rect 600700 213178 600728 220798
rect 600688 213172 600740 213178
rect 600688 213114 600740 213120
rect 600412 210452 600464 210458
rect 600412 210394 600464 210400
rect 600884 210202 600912 221167
rect 601792 220992 601844 220998
rect 601792 220934 601844 220940
rect 601804 214470 601832 220934
rect 601792 214464 601844 214470
rect 601792 214406 601844 214412
rect 601240 213172 601292 213178
rect 601240 213114 601292 213120
rect 601010 210452 601062 210458
rect 601010 210394 601062 210400
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596376 210174 596620 210202
rect 596744 210174 597172 210202
rect 597572 210174 597724 210202
rect 597940 210174 598276 210202
rect 598492 210174 598828 210202
rect 599044 210174 599380 210202
rect 599504 210174 599932 210202
rect 600484 210174 600912 210202
rect 601022 210188 601050 210394
rect 601252 210202 601280 213114
rect 601988 210202 602016 221546
rect 604644 221264 604696 221270
rect 604644 221206 604696 221212
rect 603080 219020 603132 219026
rect 603080 218962 603132 218968
rect 603092 217462 603120 218962
rect 604460 218476 604512 218482
rect 604460 218418 604512 218424
rect 604000 217864 604052 217870
rect 604000 217806 604052 217812
rect 603448 217728 603500 217734
rect 603448 217670 603500 217676
rect 603080 217456 603132 217462
rect 603080 217398 603132 217404
rect 603080 217184 603132 217190
rect 603080 217126 603132 217132
rect 602344 214464 602396 214470
rect 602344 214406 602396 214412
rect 602356 210202 602384 214406
rect 603092 210202 603120 217126
rect 603460 210202 603488 217670
rect 604012 210202 604040 217806
rect 604472 217734 604500 218418
rect 604460 217728 604512 217734
rect 604460 217670 604512 217676
rect 604656 210202 604684 221206
rect 605024 210202 605052 222022
rect 608600 221944 608652 221950
rect 608600 221886 608652 221892
rect 606668 221740 606720 221746
rect 606668 221682 606720 221688
rect 606024 219768 606076 219774
rect 606024 219710 606076 219716
rect 606036 210202 606064 219710
rect 606208 217592 606260 217598
rect 606208 217534 606260 217540
rect 601252 210174 601588 210202
rect 601988 210174 602140 210202
rect 602356 210174 602692 210202
rect 603092 210174 603244 210202
rect 603460 210174 603796 210202
rect 604012 210174 604348 210202
rect 604656 210174 604900 210202
rect 605024 210174 605452 210202
rect 606004 210174 606064 210202
rect 606220 210202 606248 217534
rect 606680 210202 606708 221682
rect 607312 219904 607364 219910
rect 607312 219846 607364 219852
rect 607324 214606 607352 219846
rect 607496 219496 607548 219502
rect 607496 219438 607548 219444
rect 607312 214600 607364 214606
rect 607312 214542 607364 214548
rect 607508 210202 607536 219438
rect 607864 214600 607916 214606
rect 607864 214542 607916 214548
rect 607876 210202 607904 214542
rect 608612 210202 608640 221886
rect 610532 220516 610584 220522
rect 610532 220458 610584 220464
rect 608968 220244 609020 220250
rect 608968 220186 609020 220192
rect 608784 220108 608836 220114
rect 608784 220050 608836 220056
rect 608796 214606 608824 220050
rect 608784 214600 608836 214606
rect 608784 214542 608836 214548
rect 608980 210202 609008 220186
rect 610072 217048 610124 217054
rect 610072 216990 610124 216996
rect 609520 214600 609572 214606
rect 609520 214542 609572 214548
rect 609532 210202 609560 214542
rect 610084 210202 610112 216990
rect 610544 210202 610572 220458
rect 611452 220380 611504 220386
rect 611452 220322 611504 220328
rect 610716 218612 610768 218618
rect 610716 218554 610768 218560
rect 610728 216782 610756 218554
rect 610716 216776 610768 216782
rect 610716 216718 610768 216724
rect 611464 210202 611492 220322
rect 611634 220280 611690 220289
rect 611634 220215 611690 220224
rect 611648 210202 611676 220215
rect 612738 219736 612794 219745
rect 612738 219671 612794 219680
rect 612280 218000 612332 218006
rect 612280 217942 612332 217948
rect 612292 210202 612320 217942
rect 612752 210202 612780 219671
rect 614120 218884 614172 218890
rect 614120 218826 614172 218832
rect 614132 217598 614160 218826
rect 614488 218000 614540 218006
rect 614488 217942 614540 217948
rect 614304 217728 614356 217734
rect 614304 217670 614356 217676
rect 614120 217592 614172 217598
rect 614120 217534 614172 217540
rect 613384 216912 613436 216918
rect 613384 216854 613436 216860
rect 613396 210202 613424 216854
rect 614316 210202 614344 217670
rect 606220 210174 606556 210202
rect 606680 210174 607108 210202
rect 607508 210174 607660 210202
rect 607876 210174 608212 210202
rect 608612 210174 608764 210202
rect 608980 210174 609316 210202
rect 609532 210174 609868 210202
rect 610084 210174 610420 210202
rect 610544 210174 610972 210202
rect 611464 210174 611524 210202
rect 611648 210174 612076 210202
rect 612292 210174 612628 210202
rect 612752 210174 613180 210202
rect 613396 210174 613732 210202
rect 614284 210174 614344 210202
rect 614500 210202 614528 217942
rect 614960 210202 614988 224810
rect 616052 224664 616104 224670
rect 616052 224606 616104 224612
rect 615684 216776 615736 216782
rect 615684 216718 615736 216724
rect 615696 210202 615724 216718
rect 616064 210202 616092 224606
rect 625252 224528 625304 224534
rect 625252 224470 625304 224476
rect 619640 224256 619692 224262
rect 619640 224198 619692 224204
rect 617340 223032 617392 223038
rect 617340 222974 617392 222980
rect 617352 222630 617380 222974
rect 617340 222624 617392 222630
rect 617340 222566 617392 222572
rect 618258 220960 618314 220969
rect 618258 220895 618314 220904
rect 617154 220008 617210 220017
rect 617154 219943 617210 219952
rect 616880 214872 616932 214878
rect 616880 214814 616932 214820
rect 616892 210202 616920 214814
rect 617168 210202 617196 219943
rect 617798 215928 617854 215937
rect 617798 215863 617854 215872
rect 617812 210202 617840 215863
rect 618272 214606 618300 220895
rect 618442 219464 618498 219473
rect 618442 219399 618498 219408
rect 618260 214600 618312 214606
rect 618260 214542 618312 214548
rect 618456 210202 618484 219399
rect 618904 214600 618956 214606
rect 618904 214542 618956 214548
rect 618916 210202 618944 214542
rect 619652 210202 619680 224198
rect 623780 224052 623832 224058
rect 623780 223994 623832 224000
rect 622676 223916 622728 223922
rect 622676 223858 622728 223864
rect 621572 223780 621624 223786
rect 621572 223722 621624 223728
rect 620652 223168 620704 223174
rect 620652 223110 620704 223116
rect 620468 222760 620520 222766
rect 620468 222702 620520 222708
rect 619916 222488 619968 222494
rect 619916 222430 619968 222436
rect 619928 214606 619956 222430
rect 620480 222222 620508 222702
rect 620664 222222 620692 223110
rect 620468 222216 620520 222222
rect 620468 222158 620520 222164
rect 620652 222216 620704 222222
rect 620652 222158 620704 222164
rect 620100 219632 620152 219638
rect 620100 219574 620152 219580
rect 619916 214600 619968 214606
rect 619916 214542 619968 214548
rect 620112 210202 620140 219574
rect 621110 215384 621166 215393
rect 621110 215319 621166 215328
rect 620560 214600 620612 214606
rect 620560 214542 620612 214548
rect 620572 210202 620600 214542
rect 621124 210202 621152 215319
rect 621584 210202 621612 223722
rect 622400 217320 622452 217326
rect 622400 217262 622452 217268
rect 622412 210202 622440 217262
rect 622688 210202 622716 223858
rect 623320 214736 623372 214742
rect 623320 214678 623372 214684
rect 623332 210202 623360 214678
rect 623792 210202 623820 223994
rect 623962 218104 624018 218113
rect 623962 218039 624018 218048
rect 623976 214606 624004 218039
rect 623964 214600 624016 214606
rect 623964 214542 624016 214548
rect 624424 214464 624476 214470
rect 624424 214406 624476 214412
rect 624436 210202 624464 214406
rect 625264 210202 625292 224470
rect 625436 224392 625488 224398
rect 625436 224334 625488 224340
rect 625448 214606 625476 224334
rect 628748 223644 628800 223650
rect 628748 223586 628800 223592
rect 625620 223032 625672 223038
rect 625620 222974 625672 222980
rect 625436 214600 625488 214606
rect 625436 214542 625488 214548
rect 625632 210202 625660 222974
rect 627092 222760 627144 222766
rect 627092 222702 627144 222708
rect 626632 217592 626684 217598
rect 626632 217534 626684 217540
rect 626080 214600 626132 214606
rect 626080 214542 626132 214548
rect 626092 210202 626120 214542
rect 626644 210202 626672 217534
rect 627104 210202 627132 222702
rect 627920 222352 627972 222358
rect 627920 222294 627972 222300
rect 627932 210202 627960 222294
rect 628288 217456 628340 217462
rect 628288 217398 628340 217404
rect 628300 210202 628328 217398
rect 628760 210202 628788 223586
rect 629852 222624 629904 222630
rect 629852 222566 629904 222572
rect 629392 214464 629444 214470
rect 629392 214406 629444 214412
rect 629404 210202 629432 214406
rect 629864 210202 629892 222566
rect 630048 214606 630076 229066
rect 633716 227044 633768 227050
rect 633716 226986 633768 226992
rect 630864 225004 630916 225010
rect 630864 224946 630916 224952
rect 630678 218376 630734 218385
rect 630678 218311 630734 218320
rect 630036 214600 630088 214606
rect 630036 214542 630088 214548
rect 630692 210202 630720 218311
rect 630876 210338 630904 224946
rect 632704 222896 632756 222902
rect 632704 222838 632756 222844
rect 631508 222216 631560 222222
rect 631508 222158 631560 222164
rect 630876 210310 630996 210338
rect 630968 210202 630996 210310
rect 631520 210202 631548 222158
rect 632716 213042 632744 222838
rect 633440 221468 633492 221474
rect 633440 221410 633492 221416
rect 632888 214600 632940 214606
rect 632888 214542 632940 214548
rect 632704 213036 632756 213042
rect 632704 212978 632756 212984
rect 632900 210202 632928 214542
rect 633452 210202 633480 221410
rect 633728 210202 633756 226986
rect 634360 213036 634412 213042
rect 634360 212978 634412 212984
rect 634372 210202 634400 212978
rect 635016 210202 635044 278258
rect 635568 272814 635596 278052
rect 636200 277636 636252 277642
rect 636200 277578 636252 277584
rect 635556 272808 635608 272814
rect 635556 272750 635608 272756
rect 636212 229094 636240 277578
rect 636764 275466 636792 278052
rect 636752 275460 636804 275466
rect 636752 275402 636804 275408
rect 637592 269822 637620 278310
rect 637764 278180 637816 278186
rect 637764 278122 637816 278128
rect 637580 269816 637632 269822
rect 637580 269758 637632 269764
rect 637776 229094 637804 278122
rect 639156 273970 639184 278052
rect 639144 273964 639196 273970
rect 639144 273906 639196 273912
rect 640352 272678 640380 278052
rect 640536 278038 641470 278066
rect 641732 278038 642666 278066
rect 640340 272672 640392 272678
rect 640340 272614 640392 272620
rect 640536 269958 640564 278038
rect 640524 269952 640576 269958
rect 640524 269894 640576 269900
rect 641732 268394 641760 278038
rect 643848 275330 643876 278052
rect 643836 275324 643888 275330
rect 643836 275266 643888 275272
rect 645044 271318 645072 278052
rect 645872 278038 646254 278066
rect 647252 278038 647450 278066
rect 645032 271312 645084 271318
rect 645032 271254 645084 271260
rect 641720 268388 641772 268394
rect 641720 268330 641772 268336
rect 645872 261526 645900 278038
rect 645860 261520 645912 261526
rect 645860 261462 645912 261468
rect 647252 246362 647280 278038
rect 647240 246356 647292 246362
rect 647240 246298 647292 246304
rect 648632 242214 648660 278052
rect 650656 277778 650684 509866
rect 660316 491366 660344 550598
rect 661696 534138 661724 594798
rect 663064 549908 663116 549914
rect 663064 549850 663116 549856
rect 661684 534132 661736 534138
rect 661684 534074 661736 534080
rect 663076 491502 663104 549850
rect 664456 535498 664484 596158
rect 665088 564460 665140 564466
rect 665088 564402 665140 564408
rect 664444 535492 664496 535498
rect 664444 535434 664496 535440
rect 663064 491496 663116 491502
rect 663064 491438 663116 491444
rect 660304 491360 660356 491366
rect 660304 491302 660356 491308
rect 665100 485858 665128 564402
rect 665824 552696 665876 552702
rect 665824 552638 665876 552644
rect 665836 491638 665864 552638
rect 665824 491632 665876 491638
rect 665824 491574 665876 491580
rect 665088 485852 665140 485858
rect 665088 485794 665140 485800
rect 665180 480412 665232 480418
rect 665180 480354 665232 480360
rect 665192 476202 665220 480354
rect 659660 476196 659712 476202
rect 659660 476138 659712 476144
rect 665180 476196 665232 476202
rect 665180 476138 665232 476144
rect 659672 473482 659700 476138
rect 656164 473476 656216 473482
rect 656164 473418 656216 473424
rect 659660 473476 659712 473482
rect 659660 473418 659712 473424
rect 656176 470626 656204 473418
rect 650828 470620 650880 470626
rect 650828 470562 650880 470568
rect 656164 470620 656216 470626
rect 656164 470562 656216 470568
rect 650840 277914 650868 470562
rect 667032 456618 667060 703802
rect 667662 698320 667718 698329
rect 667662 698255 667718 698264
rect 667204 686520 667256 686526
rect 667204 686462 667256 686468
rect 667216 625734 667244 686462
rect 667478 645824 667534 645833
rect 667478 645759 667534 645768
rect 667204 625728 667256 625734
rect 667204 625670 667256 625676
rect 667294 600944 667350 600953
rect 667294 600879 667350 600888
rect 667308 529990 667336 600879
rect 667492 574122 667520 645759
rect 667676 621654 667704 698255
rect 667664 621648 667716 621654
rect 667664 621590 667716 621596
rect 667664 608660 667716 608666
rect 667664 608602 667716 608608
rect 667480 574116 667532 574122
rect 667480 574058 667532 574064
rect 667676 531894 667704 608602
rect 667664 531888 667716 531894
rect 667664 531830 667716 531836
rect 667296 529984 667348 529990
rect 667296 529926 667348 529932
rect 667020 456612 667072 456618
rect 667020 456554 667072 456560
rect 667860 456006 667888 705162
rect 668398 689480 668454 689489
rect 668398 689415 668454 689424
rect 668214 687848 668270 687857
rect 668214 687783 668270 687792
rect 668228 617982 668256 687783
rect 668216 617976 668268 617982
rect 668216 617918 668268 617924
rect 668412 616894 668440 689415
rect 668596 671158 668624 733382
rect 668858 730144 668914 730153
rect 668858 730079 668914 730088
rect 668584 671152 668636 671158
rect 668584 671094 668636 671100
rect 668872 660142 668900 730079
rect 669056 709374 669084 782478
rect 669044 709368 669096 709374
rect 669044 709310 669096 709316
rect 669240 708286 669268 784110
rect 670424 777028 670476 777034
rect 670424 776970 670476 776976
rect 669964 775600 670016 775606
rect 669964 775542 670016 775548
rect 669596 735616 669648 735622
rect 669596 735558 669648 735564
rect 669410 728784 669466 728793
rect 669410 728719 669466 728728
rect 669228 708280 669280 708286
rect 669228 708222 669280 708228
rect 669042 690568 669098 690577
rect 669042 690503 669098 690512
rect 668860 660136 668912 660142
rect 668860 660078 668912 660084
rect 668584 640348 668636 640354
rect 668584 640290 668636 640296
rect 668400 616888 668452 616894
rect 668400 616830 668452 616836
rect 668398 593464 668454 593473
rect 668398 593399 668454 593408
rect 668412 529174 668440 593399
rect 668596 580310 668624 640290
rect 669056 620430 669084 690503
rect 669424 663950 669452 728719
rect 669608 665310 669636 735558
rect 669976 715766 670004 775542
rect 669964 715760 670016 715766
rect 669964 715702 670016 715708
rect 670436 705362 670464 776970
rect 670620 709238 670648 784246
rect 670896 728142 670924 886858
rect 670884 728136 670936 728142
rect 670884 728078 670936 728084
rect 671080 715358 671108 894406
rect 671896 894328 671948 894334
rect 671896 894270 671948 894276
rect 671436 773424 671488 773430
rect 671436 773366 671488 773372
rect 671250 733816 671306 733825
rect 671250 733751 671306 733760
rect 671068 715352 671120 715358
rect 671068 715294 671120 715300
rect 671068 713244 671120 713250
rect 671068 713186 671120 713192
rect 670608 709232 670660 709238
rect 670608 709174 670660 709180
rect 670424 705356 670476 705362
rect 670424 705298 670476 705304
rect 670882 694920 670938 694929
rect 670882 694855 670938 694864
rect 669964 687268 670016 687274
rect 669964 687210 670016 687216
rect 669778 683904 669834 683913
rect 669778 683839 669834 683848
rect 669596 665304 669648 665310
rect 669596 665246 669648 665252
rect 669412 663944 669464 663950
rect 669412 663886 669464 663892
rect 669228 661156 669280 661162
rect 669228 661098 669280 661104
rect 669044 620424 669096 620430
rect 669044 620366 669096 620372
rect 669042 594824 669098 594833
rect 669042 594759 669098 594768
rect 668584 580304 668636 580310
rect 668584 580246 668636 580252
rect 668766 562320 668822 562329
rect 668766 562255 668822 562264
rect 668400 529168 668452 529174
rect 668400 529110 668452 529116
rect 668584 524476 668636 524482
rect 668584 524418 668636 524424
rect 668596 518226 668624 524418
rect 668584 518220 668636 518226
rect 668584 518162 668636 518168
rect 668780 484430 668808 562255
rect 669056 524618 669084 594759
rect 669044 524612 669096 524618
rect 669044 524554 669096 524560
rect 669056 524482 669084 524554
rect 669044 524476 669096 524482
rect 669044 524418 669096 524424
rect 668768 484424 668820 484430
rect 668768 484366 668820 484372
rect 667848 456000 667900 456006
rect 667848 455942 667900 455948
rect 669240 455666 669268 661098
rect 669594 644328 669650 644337
rect 669594 644263 669650 644272
rect 669412 623892 669464 623898
rect 669412 623834 669464 623840
rect 669424 578950 669452 623834
rect 669412 578944 669464 578950
rect 669412 578886 669464 578892
rect 669412 576904 669464 576910
rect 669412 576846 669464 576852
rect 669424 532574 669452 576846
rect 669608 571402 669636 644263
rect 669792 619886 669820 683839
rect 669976 626006 670004 687210
rect 670606 684992 670662 685001
rect 670606 684927 670662 684936
rect 670240 669656 670292 669662
rect 670240 669598 670292 669604
rect 669964 626000 670016 626006
rect 669964 625942 670016 625948
rect 670252 625054 670280 669598
rect 670240 625048 670292 625054
rect 670240 624990 670292 624996
rect 670240 624708 670292 624714
rect 670240 624650 670292 624656
rect 669780 619880 669832 619886
rect 669780 619822 669832 619828
rect 669964 597576 670016 597582
rect 669964 597518 670016 597524
rect 669596 571396 669648 571402
rect 669596 571338 669648 571344
rect 669780 568608 669832 568614
rect 669780 568550 669832 568556
rect 669596 553444 669648 553450
rect 669596 553386 669648 553392
rect 669608 552265 669636 553386
rect 669594 552256 669650 552265
rect 669594 552191 669650 552200
rect 669412 532568 669464 532574
rect 669412 532510 669464 532516
rect 669228 455660 669280 455666
rect 669228 455602 669280 455608
rect 669792 455433 669820 568550
rect 669976 535974 670004 597518
rect 670252 580038 670280 624650
rect 670424 623076 670476 623082
rect 670424 623018 670476 623024
rect 670240 580032 670292 580038
rect 670240 579974 670292 579980
rect 670240 577652 670292 577658
rect 670240 577594 670292 577600
rect 669964 535968 670016 535974
rect 669964 535910 670016 535916
rect 670252 533322 670280 577594
rect 670436 577454 670464 623018
rect 670620 615534 670648 684927
rect 670896 620702 670924 694855
rect 671080 668574 671108 713186
rect 671068 668568 671120 668574
rect 671068 668510 671120 668516
rect 671068 668160 671120 668166
rect 671068 668102 671120 668108
rect 671080 623558 671108 668102
rect 671264 661638 671292 733751
rect 671448 710054 671476 773366
rect 671908 743834 671936 894270
rect 672540 892900 672592 892906
rect 672540 892842 672592 892848
rect 672552 746594 672580 892842
rect 672736 866658 672764 895630
rect 675850 895520 675906 895529
rect 675850 895455 675906 895464
rect 675864 894470 675892 895455
rect 676034 894704 676090 894713
rect 676034 894639 676090 894648
rect 675852 894464 675904 894470
rect 675852 894406 675904 894412
rect 676048 894334 676076 894639
rect 676036 894328 676088 894334
rect 676036 894270 676088 894276
rect 675850 893888 675906 893897
rect 675850 893823 675906 893832
rect 672908 893036 672960 893042
rect 672908 892978 672960 892984
rect 672724 866652 672776 866658
rect 672724 866594 672776 866600
rect 672724 775668 672776 775674
rect 672724 775610 672776 775616
rect 672736 746594 672764 775610
rect 672552 746566 672672 746594
rect 672736 746566 672856 746594
rect 671908 743806 672028 743834
rect 671804 742212 671856 742218
rect 671804 742154 671856 742160
rect 671620 741192 671672 741198
rect 671620 741134 671672 741140
rect 671436 710048 671488 710054
rect 671436 709990 671488 709996
rect 671632 673454 671660 741134
rect 671816 734174 671844 742154
rect 672000 734174 672028 743806
rect 672264 738472 672316 738478
rect 672264 738414 672316 738420
rect 671540 673426 671660 673454
rect 671724 734146 671844 734174
rect 671908 734146 672028 734174
rect 671540 668137 671568 673426
rect 671526 668128 671582 668137
rect 671526 668063 671582 668072
rect 671436 667956 671488 667962
rect 671436 667898 671488 667904
rect 671252 661632 671304 661638
rect 671252 661574 671304 661580
rect 671448 654134 671476 667898
rect 671724 664426 671752 734146
rect 671908 714542 671936 734146
rect 672080 732760 672132 732766
rect 672080 732702 672132 732708
rect 671896 714536 671948 714542
rect 671896 714478 671948 714484
rect 671896 712428 671948 712434
rect 671896 712370 671948 712376
rect 671908 666942 671936 712370
rect 671896 666936 671948 666942
rect 671896 666878 671948 666884
rect 671896 666596 671948 666602
rect 671896 666538 671948 666544
rect 671712 664420 671764 664426
rect 671712 664362 671764 664368
rect 671448 654106 671568 654134
rect 671342 638752 671398 638761
rect 671342 638687 671398 638696
rect 671356 628538 671384 638687
rect 671540 637574 671568 654106
rect 671710 647864 671766 647873
rect 671710 647799 671766 647808
rect 671540 637546 671660 637574
rect 671632 636194 671660 637546
rect 671540 636166 671660 636194
rect 671540 628794 671568 636166
rect 671528 628788 671580 628794
rect 671528 628730 671580 628736
rect 671356 628510 671660 628538
rect 671344 628448 671396 628454
rect 671344 628390 671396 628396
rect 671356 626534 671384 628390
rect 671356 626506 671476 626534
rect 671448 624374 671476 626506
rect 671436 624368 671488 624374
rect 671436 624310 671488 624316
rect 671068 623552 671120 623558
rect 671068 623494 671120 623500
rect 671436 622260 671488 622266
rect 671436 622202 671488 622208
rect 670884 620696 670936 620702
rect 670884 620638 670936 620644
rect 670608 615528 670660 615534
rect 670608 615470 670660 615476
rect 670608 614916 670660 614922
rect 670608 614858 670660 614864
rect 670424 577448 670476 577454
rect 670424 577390 670476 577396
rect 670422 549672 670478 549681
rect 670422 549607 670478 549616
rect 670240 533316 670292 533322
rect 670240 533258 670292 533264
rect 670436 480418 670464 549607
rect 670424 480412 670476 480418
rect 670424 480354 670476 480360
rect 669778 455424 669834 455433
rect 669778 455359 669834 455368
rect 670620 455161 670648 614858
rect 671158 608560 671214 608569
rect 671158 608495 671214 608504
rect 670792 578264 670844 578270
rect 670792 578206 670844 578212
rect 670974 578232 671030 578241
rect 670804 534750 670832 578206
rect 670974 578167 671030 578176
rect 670988 535022 671016 578167
rect 670976 535016 671028 535022
rect 670976 534958 671028 534964
rect 670792 534744 670844 534750
rect 670792 534686 670844 534692
rect 670974 534032 671030 534041
rect 670974 533967 671030 533976
rect 670792 532772 670844 532778
rect 670792 532714 670844 532720
rect 670804 489326 670832 532714
rect 670988 490958 671016 533967
rect 671172 529446 671200 608495
rect 671448 577182 671476 622202
rect 671436 577176 671488 577182
rect 671436 577118 671488 577124
rect 671632 574598 671660 628510
rect 671724 601694 671752 647799
rect 671908 622742 671936 666538
rect 672092 662454 672120 732702
rect 672276 665174 672304 738414
rect 672448 714876 672500 714882
rect 672448 714818 672500 714824
rect 672460 670614 672488 714818
rect 672644 713726 672672 746566
rect 672632 713720 672684 713726
rect 672632 713662 672684 713668
rect 672828 713538 672856 746566
rect 672736 713510 672856 713538
rect 672736 711657 672764 713510
rect 672920 712881 672948 892978
rect 675864 892906 675892 893823
rect 676034 893072 676090 893081
rect 676034 893007 676036 893016
rect 676088 893007 676090 893016
rect 676036 892978 676088 892984
rect 675852 892900 675904 892906
rect 675852 892842 675904 892848
rect 676034 892664 676090 892673
rect 676090 892622 676444 892650
rect 676034 892599 676090 892608
rect 676034 891440 676090 891449
rect 676034 891375 676090 891384
rect 675206 891032 675262 891041
rect 675206 890967 675262 890976
rect 675024 890384 675076 890390
rect 675024 890326 675076 890332
rect 674656 888956 674708 888962
rect 674656 888898 674708 888904
rect 674668 888734 674696 888898
rect 674576 888706 674696 888734
rect 674380 888548 674432 888554
rect 674380 888490 674432 888496
rect 674196 887324 674248 887330
rect 674196 887266 674248 887272
rect 673092 885692 673144 885698
rect 673092 885634 673144 885640
rect 673104 728346 673132 885634
rect 674208 868766 674236 887266
rect 674392 872166 674420 888490
rect 674576 879074 674604 888706
rect 675036 879646 675064 890326
rect 675024 879640 675076 879646
rect 675024 879582 675076 879588
rect 674748 879232 674800 879238
rect 674748 879174 674800 879180
rect 674760 879084 674788 879174
rect 674576 879046 674696 879074
rect 674760 879056 674880 879084
rect 674380 872160 674432 872166
rect 674380 872102 674432 872108
rect 674668 869802 674696 879046
rect 674852 878370 674880 879056
rect 675220 878830 675248 890967
rect 676048 890390 676076 891375
rect 676036 890384 676088 890390
rect 676036 890326 676088 890332
rect 676034 890216 676090 890225
rect 676090 890186 676260 890202
rect 676090 890180 676272 890186
rect 676090 890174 676220 890180
rect 676034 890151 676090 890160
rect 676220 890122 676272 890128
rect 676034 889400 676090 889409
rect 676090 889358 676260 889386
rect 676034 889335 676090 889344
rect 676034 888992 676090 889001
rect 676034 888927 676036 888936
rect 676088 888927 676090 888936
rect 676036 888898 676088 888904
rect 676232 888758 676260 889358
rect 676220 888752 676272 888758
rect 676220 888694 676272 888700
rect 676034 888584 676090 888593
rect 676034 888519 676036 888528
rect 676088 888519 676090 888528
rect 676036 888490 676088 888496
rect 676034 887360 676090 887369
rect 676034 887295 676036 887304
rect 676088 887295 676090 887304
rect 676036 887266 676088 887272
rect 676034 886952 676090 886961
rect 676034 886887 676036 886896
rect 676088 886887 676090 886896
rect 676036 886858 676088 886864
rect 676034 885728 676090 885737
rect 676034 885663 676036 885672
rect 676088 885663 676090 885672
rect 676036 885634 676088 885640
rect 675392 880388 675444 880394
rect 675392 880330 675444 880336
rect 675404 878914 675432 880330
rect 675944 879368 675996 879374
rect 675944 879310 675996 879316
rect 675760 879096 675812 879102
rect 675760 879038 675812 879044
rect 675404 878886 675616 878914
rect 675208 878824 675260 878830
rect 675208 878766 675260 878772
rect 675392 878824 675444 878830
rect 675392 878766 675444 878772
rect 675404 878642 675432 878766
rect 674806 878342 674880 878370
rect 675312 878614 675432 878642
rect 674806 878098 674834 878342
rect 674932 878212 674984 878218
rect 674932 878154 674984 878160
rect 674806 878070 674880 878098
rect 674852 874206 674880 878070
rect 674944 874698 674972 878154
rect 675312 878098 675340 878614
rect 675128 878070 675340 878098
rect 675588 878084 675616 878886
rect 675772 878529 675800 879038
rect 675758 878520 675814 878529
rect 675956 878490 675984 879310
rect 676416 878626 676444 892622
rect 679622 891848 679678 891857
rect 679622 891783 679678 891792
rect 676864 890180 676916 890186
rect 676864 890122 676916 890128
rect 676876 879374 676904 890122
rect 678242 889808 678298 889817
rect 678242 889743 678298 889752
rect 677048 888752 677100 888758
rect 677048 888694 677100 888700
rect 677060 879510 677088 888694
rect 677048 879504 677100 879510
rect 677048 879446 677100 879452
rect 676864 879368 676916 879374
rect 676864 879310 676916 879316
rect 678256 879102 678284 889743
rect 678244 879096 678296 879102
rect 678244 879038 678296 879044
rect 676404 878620 676456 878626
rect 676404 878562 676456 878568
rect 679636 878529 679664 891783
rect 681002 890624 681058 890633
rect 681002 890559 681058 890568
rect 681016 880705 681044 890559
rect 683118 888176 683174 888185
rect 683118 888111 683174 888120
rect 681002 880696 681058 880705
rect 681002 880631 681058 880640
rect 683132 880433 683160 888111
rect 683118 880424 683174 880433
rect 683118 880359 683174 880368
rect 679622 878520 679678 878529
rect 675758 878455 675814 878464
rect 675944 878484 675996 878490
rect 679622 878455 679678 878464
rect 675944 878426 675996 878432
rect 675128 877962 675156 878070
rect 675036 877934 675156 877962
rect 675390 877976 675446 877985
rect 675036 876194 675064 877934
rect 675390 877911 675446 877920
rect 675208 877804 675260 877810
rect 675208 877746 675260 877752
rect 675220 876262 675248 877746
rect 675404 877694 675432 877911
rect 675312 877666 675432 877694
rect 675312 877418 675340 877666
rect 675404 877418 675432 877540
rect 675312 877390 675432 877418
rect 675484 877260 675536 877266
rect 675484 877202 675536 877208
rect 675496 876860 675524 877202
rect 675220 876234 675418 876262
rect 675036 876166 675156 876194
rect 675128 874698 675156 876166
rect 674944 874670 675064 874698
rect 675128 874670 675340 874698
rect 674840 874200 674892 874206
rect 674840 874142 674892 874148
rect 675036 873474 675064 874670
rect 675312 874290 675340 874670
rect 675404 874290 675432 874412
rect 675312 874262 675432 874290
rect 675300 874200 675352 874206
rect 675300 874142 675352 874148
rect 675574 874168 675630 874177
rect 675036 873446 675156 873474
rect 675128 872174 675156 873446
rect 675312 873202 675340 874142
rect 675574 874103 675630 874112
rect 675588 873868 675616 874103
rect 675312 873174 675418 873202
rect 675758 872808 675814 872817
rect 675758 872743 675814 872752
rect 675772 872576 675800 872743
rect 674840 872160 674892 872166
rect 675036 872146 675156 872174
rect 674892 872108 674972 872114
rect 674840 872102 674972 872108
rect 674852 872086 674972 872102
rect 674944 869802 674972 872086
rect 675036 870482 675064 872146
rect 675036 870454 675432 870482
rect 675404 870060 675432 870454
rect 675758 869816 675814 869825
rect 674668 869774 674880 869802
rect 674944 869774 675248 869802
rect 674852 869258 674880 869774
rect 675024 869440 675076 869446
rect 675076 869388 675156 869394
rect 675024 869382 675156 869388
rect 675036 869366 675156 869382
rect 674852 869230 675064 869258
rect 674196 868760 674248 868766
rect 674196 868702 674248 868708
rect 674840 868080 674892 868086
rect 674840 868022 674892 868028
rect 674852 865858 674880 868022
rect 675036 867049 675064 869230
rect 675128 867694 675156 869366
rect 675220 868889 675248 869774
rect 675758 869751 675814 869760
rect 675772 869516 675800 869751
rect 675220 868861 675418 868889
rect 675300 868760 675352 868766
rect 675300 868702 675352 868708
rect 675312 868238 675340 868702
rect 675312 868210 675418 868238
rect 675128 867666 675418 867694
rect 675036 867021 675418 867049
rect 674852 865830 675418 865858
rect 675298 865736 675354 865745
rect 675298 865671 675354 865680
rect 675312 863818 675340 865671
rect 675758 865464 675814 865473
rect 675758 865399 675814 865408
rect 675772 865195 675800 865399
rect 675666 864920 675722 864929
rect 675666 864855 675722 864864
rect 675680 864552 675708 864855
rect 675312 863790 675432 863818
rect 675404 863328 675432 863790
rect 675392 790832 675444 790838
rect 675392 790774 675444 790780
rect 675404 788868 675432 790774
rect 675772 788089 675800 788324
rect 675758 788080 675814 788089
rect 675758 788015 675814 788024
rect 675128 787665 675418 787693
rect 675128 786729 675156 787665
rect 675404 786729 675432 787032
rect 675114 786720 675170 786729
rect 675114 786655 675170 786664
rect 675390 786720 675446 786729
rect 675390 786655 675446 786664
rect 674852 785182 675418 785210
rect 673736 782672 673788 782678
rect 673736 782614 673788 782620
rect 673274 777472 673330 777481
rect 673274 777407 673330 777416
rect 673092 728340 673144 728346
rect 673092 728282 673144 728288
rect 673090 714096 673146 714105
rect 673090 714031 673146 714040
rect 672906 712872 672962 712881
rect 672906 712807 672962 712816
rect 672722 711648 672778 711657
rect 672722 711583 672778 711592
rect 673104 702434 673132 714031
rect 673288 708393 673316 777407
rect 673552 738676 673604 738682
rect 673552 738618 673604 738624
rect 673564 736934 673592 738618
rect 673564 736906 673684 736934
rect 673458 734224 673514 734233
rect 673458 734159 673514 734168
rect 673274 708384 673330 708393
rect 673274 708319 673330 708328
rect 672644 702406 673132 702434
rect 672448 670608 672500 670614
rect 672448 670550 672500 670556
rect 672644 669905 672672 702406
rect 673182 696960 673238 696969
rect 673182 696895 673238 696904
rect 673000 688832 673052 688838
rect 672998 688800 673000 688809
rect 673052 688800 673054 688809
rect 672998 688735 673054 688744
rect 672814 685672 672870 685681
rect 672814 685607 672870 685616
rect 672630 669896 672686 669905
rect 672630 669831 672686 669840
rect 672264 665168 672316 665174
rect 672264 665110 672316 665116
rect 672080 662448 672132 662454
rect 672080 662390 672132 662396
rect 672170 652488 672226 652497
rect 672170 652423 672226 652432
rect 672184 652338 672212 652423
rect 672000 652310 672212 652338
rect 672000 622962 672028 652310
rect 672630 649224 672686 649233
rect 672630 649159 672686 649168
rect 672644 640334 672672 649159
rect 672644 640306 672764 640334
rect 672736 630674 672764 640306
rect 672644 630646 672764 630674
rect 672000 622934 672120 622962
rect 671896 622736 671948 622742
rect 671896 622678 671948 622684
rect 672092 622554 672120 622934
rect 672000 622526 672120 622554
rect 671724 601666 671844 601694
rect 671620 574592 671672 574598
rect 671620 574534 671672 574540
rect 671816 571606 671844 601666
rect 672000 574326 672028 622526
rect 672644 621014 672672 630646
rect 672828 621489 672856 685607
rect 672998 648816 673054 648825
rect 672998 648751 673054 648760
rect 672814 621480 672870 621489
rect 672814 621415 672870 621424
rect 672644 620986 672764 621014
rect 672540 620696 672592 620702
rect 672538 620664 672540 620673
rect 672592 620664 672594 620673
rect 672538 620599 672594 620608
rect 672170 609104 672226 609113
rect 672170 609039 672226 609048
rect 671988 574320 672040 574326
rect 671988 574262 672040 574268
rect 671804 571600 671856 571606
rect 671804 571542 671856 571548
rect 671344 571124 671396 571130
rect 671344 571066 671396 571072
rect 671160 529440 671212 529446
rect 671160 529382 671212 529388
rect 670976 490952 671028 490958
rect 670976 490894 671028 490900
rect 670792 489320 670844 489326
rect 670792 489262 670844 489268
rect 670606 455152 670662 455161
rect 670606 455087 670662 455096
rect 657542 403336 657598 403345
rect 657542 403271 657598 403280
rect 652022 400888 652078 400897
rect 652022 400823 652078 400832
rect 651472 373992 651524 373998
rect 651472 373934 651524 373940
rect 651484 373289 651512 373934
rect 651470 373280 651526 373289
rect 651470 373215 651526 373224
rect 652036 372201 652064 400823
rect 652206 396672 652262 396681
rect 652206 396607 652262 396616
rect 652220 373969 652248 396607
rect 654782 382936 654838 382945
rect 654782 382871 654838 382880
rect 652206 373960 652262 373969
rect 652206 373895 652262 373904
rect 652022 372192 652078 372201
rect 652022 372127 652078 372136
rect 654796 371006 654824 382871
rect 657556 373998 657584 403271
rect 670514 392592 670570 392601
rect 670514 392527 670570 392536
rect 657544 373992 657596 373998
rect 657544 373934 657596 373940
rect 668582 371240 668638 371249
rect 668582 371175 668638 371184
rect 651472 371000 651524 371006
rect 651472 370942 651524 370948
rect 654784 371000 654836 371006
rect 654784 370942 654836 370948
rect 651484 370705 651512 370942
rect 651470 370696 651526 370705
rect 651470 370631 651526 370640
rect 668596 365022 668624 371175
rect 655520 365016 655572 365022
rect 655520 364958 655572 364964
rect 668584 365016 668636 365022
rect 668584 364958 668636 364964
rect 655532 361622 655560 364958
rect 651012 361616 651064 361622
rect 651012 361558 651064 361564
rect 655520 361616 655572 361622
rect 655520 361558 655572 361564
rect 651024 278458 651052 361558
rect 654782 358592 654838 358601
rect 654782 358527 654838 358536
rect 652022 356688 652078 356697
rect 652022 356623 652078 356632
rect 651380 328296 651432 328302
rect 651380 328238 651432 328244
rect 651392 328137 651420 328238
rect 651378 328128 651434 328137
rect 651378 328063 651434 328072
rect 652036 326913 652064 356623
rect 652390 351112 652446 351121
rect 652390 351047 652446 351056
rect 652404 329769 652432 351047
rect 653402 338736 653458 338745
rect 653402 338671 653458 338680
rect 652390 329760 652446 329769
rect 652390 329695 652446 329704
rect 652022 326904 652078 326913
rect 652022 326839 652078 326848
rect 651378 325680 651434 325689
rect 653416 325650 653444 338671
rect 654796 328302 654824 358527
rect 669410 347304 669466 347313
rect 669410 347239 669466 347248
rect 654784 328296 654836 328302
rect 654784 328238 654836 328244
rect 651378 325615 651380 325624
rect 651432 325615 651434 325624
rect 653404 325644 653456 325650
rect 651380 325586 651432 325592
rect 653404 325586 653456 325592
rect 653402 313304 653458 313313
rect 653402 313239 653458 313248
rect 652298 309904 652354 309913
rect 652298 309839 652354 309848
rect 651380 303544 651432 303550
rect 651380 303486 651432 303492
rect 651392 303385 651420 303486
rect 651378 303376 651434 303385
rect 651378 303311 651434 303320
rect 652312 302161 652340 309839
rect 653416 303550 653444 313239
rect 660302 311944 660358 311953
rect 660302 311879 660358 311888
rect 653404 303544 653456 303550
rect 653404 303486 653456 303492
rect 652298 302152 652354 302161
rect 652298 302087 652354 302096
rect 660316 300830 660344 311879
rect 651472 300824 651524 300830
rect 651472 300766 651524 300772
rect 660304 300824 660356 300830
rect 660304 300766 660356 300772
rect 651484 300665 651512 300766
rect 651470 300656 651526 300665
rect 651470 300591 651526 300600
rect 652574 298616 652630 298625
rect 652630 298574 652800 298602
rect 652574 298551 652630 298560
rect 652114 297528 652170 297537
rect 652114 297463 652170 297472
rect 651930 296848 651986 296857
rect 651930 296783 651932 296792
rect 651984 296783 651986 296792
rect 651932 296754 651984 296760
rect 652128 296714 652156 297463
rect 652036 296686 652156 296714
rect 652772 296714 652800 298574
rect 665824 296744 665876 296750
rect 652772 296686 652892 296714
rect 665824 296686 665876 296692
rect 651654 295352 651710 295361
rect 651654 295287 651710 295296
rect 651470 294264 651526 294273
rect 651470 294199 651526 294208
rect 651484 294030 651512 294199
rect 651472 294024 651524 294030
rect 651472 293966 651524 293972
rect 651470 291680 651526 291689
rect 651470 291615 651526 291624
rect 651484 291242 651512 291615
rect 651472 291236 651524 291242
rect 651472 291178 651524 291184
rect 651668 290465 651696 295287
rect 651378 290456 651434 290465
rect 651378 290391 651380 290400
rect 651432 290391 651434 290400
rect 651654 290456 651710 290465
rect 651654 290391 651710 290400
rect 651380 290362 651432 290368
rect 651470 288688 651526 288697
rect 651470 288623 651526 288632
rect 651484 288454 651512 288623
rect 651472 288448 651524 288454
rect 651472 288390 651524 288396
rect 651470 287464 651526 287473
rect 651470 287399 651526 287408
rect 651484 287094 651512 287399
rect 651472 287088 651524 287094
rect 651472 287030 651524 287036
rect 651470 285968 651526 285977
rect 651470 285903 651526 285912
rect 651484 285734 651512 285903
rect 651472 285728 651524 285734
rect 651472 285670 651524 285676
rect 651470 284744 651526 284753
rect 651470 284679 651526 284688
rect 651484 284374 651512 284679
rect 651472 284368 651524 284374
rect 651472 284310 651524 284316
rect 652036 283529 652064 296686
rect 652864 293865 652892 296686
rect 664444 294024 664496 294030
rect 664444 293966 664496 293972
rect 652850 293856 652906 293865
rect 652850 293791 652906 293800
rect 652390 292768 652446 292777
rect 652390 292703 652446 292712
rect 652206 289232 652262 289241
rect 652206 289167 652262 289176
rect 652022 283520 652078 283529
rect 652022 283455 652078 283464
rect 651470 283248 651526 283257
rect 651470 283183 651526 283192
rect 651484 282198 651512 283183
rect 651472 282192 651524 282198
rect 651472 282134 651524 282140
rect 652022 282160 652078 282169
rect 652022 282095 652078 282104
rect 651470 280936 651526 280945
rect 651470 280871 651526 280880
rect 651484 280226 651512 280871
rect 651472 280220 651524 280226
rect 651472 280162 651524 280168
rect 651012 278452 651064 278458
rect 651012 278394 651064 278400
rect 650828 277908 650880 277914
rect 650828 277850 650880 277856
rect 650644 277772 650696 277778
rect 650644 277714 650696 277720
rect 648620 242208 648672 242214
rect 648620 242150 648672 242156
rect 636212 229066 636516 229094
rect 637776 229066 638172 229094
rect 636488 210202 636516 229066
rect 638144 210202 638172 229066
rect 651288 224256 651340 224262
rect 651288 224198 651340 224204
rect 649814 221504 649870 221513
rect 649814 221439 649870 221448
rect 646042 219872 646098 219881
rect 646042 219807 646098 219816
rect 644940 218068 644992 218074
rect 644940 218010 644992 218016
rect 643836 213240 643888 213246
rect 643836 213182 643888 213188
rect 639880 212696 639932 212702
rect 639880 212638 639932 212644
rect 639892 210202 639920 212638
rect 641720 212560 641772 212566
rect 641720 212502 641772 212508
rect 641732 210202 641760 212502
rect 643848 210202 643876 213182
rect 644952 210202 644980 218010
rect 646056 213926 646084 219807
rect 648526 218648 648582 218657
rect 648526 218583 648582 218592
rect 646320 216096 646372 216102
rect 646320 216038 646372 216044
rect 646044 213920 646096 213926
rect 646044 213862 646096 213868
rect 645492 213784 645544 213790
rect 645492 213726 645544 213732
rect 645504 210202 645532 213726
rect 646332 210202 646360 216038
rect 648252 214600 648304 214606
rect 648252 214542 648304 214548
rect 646504 213920 646556 213926
rect 646504 213862 646556 213868
rect 614500 210174 614836 210202
rect 614960 210174 615388 210202
rect 615696 210174 615940 210202
rect 616064 210174 616492 210202
rect 616892 210174 617044 210202
rect 617168 210174 617596 210202
rect 617812 210174 618148 210202
rect 618456 210174 618700 210202
rect 618916 210174 619252 210202
rect 619652 210174 619804 210202
rect 620112 210174 620356 210202
rect 620572 210174 620908 210202
rect 621124 210174 621460 210202
rect 621584 210174 622012 210202
rect 622412 210174 622564 210202
rect 622688 210174 623116 210202
rect 623332 210174 623668 210202
rect 623792 210174 624220 210202
rect 624436 210174 624772 210202
rect 625264 210174 625324 210202
rect 625632 210174 625876 210202
rect 626092 210174 626428 210202
rect 626644 210174 626980 210202
rect 627104 210174 627532 210202
rect 627932 210174 628084 210202
rect 628300 210174 628636 210202
rect 628760 210174 629188 210202
rect 629404 210174 629740 210202
rect 629864 210174 630292 210202
rect 630692 210174 630844 210202
rect 630968 210174 631396 210202
rect 631520 210174 631948 210202
rect 632900 210174 633052 210202
rect 633452 210174 633604 210202
rect 633728 210174 634156 210202
rect 634372 210174 634708 210202
rect 635016 210174 635260 210202
rect 636488 210174 636916 210202
rect 638144 210174 638572 210202
rect 639892 210174 640228 210202
rect 641732 210174 641884 210202
rect 643540 210174 643876 210202
rect 644644 210174 644980 210202
rect 645196 210174 645532 210202
rect 646300 210174 646360 210202
rect 646516 210202 646544 213862
rect 648264 210202 648292 214542
rect 648540 210202 648568 218583
rect 649632 215960 649684 215966
rect 649632 215902 649684 215908
rect 649644 210202 649672 215902
rect 649828 213790 649856 221439
rect 651102 217288 651158 217297
rect 651102 217223 651158 217232
rect 649816 213784 649868 213790
rect 649816 213726 649868 213732
rect 650460 212764 650512 212770
rect 650460 212706 650512 212712
rect 650472 210202 650500 212706
rect 646516 210174 646852 210202
rect 647956 210174 648292 210202
rect 648508 210174 648568 210202
rect 649612 210174 649672 210202
rect 650164 210174 650500 210202
rect 651116 210202 651144 217223
rect 651300 212770 651328 224198
rect 651470 221776 651526 221785
rect 651470 221711 651526 221720
rect 651288 212764 651340 212770
rect 651288 212706 651340 212712
rect 651484 210202 651512 221711
rect 651116 210174 651268 210202
rect 651484 210174 651820 210202
rect 652036 209574 652064 282095
rect 652220 228585 652248 289167
rect 652404 233918 652432 292703
rect 663064 291236 663116 291242
rect 663064 291178 663116 291184
rect 653404 290420 653456 290426
rect 653404 290362 653456 290368
rect 652574 280392 652630 280401
rect 652574 280327 652630 280336
rect 652392 233912 652444 233918
rect 652392 233854 652444 233860
rect 652206 228576 652262 228585
rect 652206 228511 652262 228520
rect 652588 226953 652616 280327
rect 653416 232558 653444 290362
rect 663076 232694 663104 291178
rect 664456 248033 664484 293966
rect 665836 268569 665864 296686
rect 667572 287088 667624 287094
rect 667572 287030 667624 287036
rect 667388 285728 667440 285734
rect 667388 285670 667440 285676
rect 666560 282192 666612 282198
rect 666560 282134 666612 282140
rect 665822 268560 665878 268569
rect 665822 268495 665878 268504
rect 664442 248024 664498 248033
rect 664442 247959 664498 247968
rect 666572 245721 666600 282134
rect 667204 280220 667256 280226
rect 667204 280162 667256 280168
rect 666558 245712 666614 245721
rect 666558 245647 666614 245656
rect 663064 232688 663116 232694
rect 663064 232630 663116 232636
rect 653404 232552 653456 232558
rect 653404 232494 653456 232500
rect 666284 231600 666336 231606
rect 666284 231542 666336 231548
rect 665088 231192 665140 231198
rect 665088 231134 665140 231140
rect 663890 229800 663946 229809
rect 663708 229764 663760 229770
rect 663890 229735 663946 229744
rect 663708 229706 663760 229712
rect 660948 229288 661000 229294
rect 660948 229230 661000 229236
rect 652574 226944 652630 226953
rect 652574 226879 652630 226888
rect 653586 226400 653642 226409
rect 653586 226335 653642 226344
rect 653402 222864 653458 222873
rect 653402 222799 653458 222808
rect 653220 213920 653272 213926
rect 653220 213862 653272 213868
rect 653232 210202 653260 213862
rect 653416 213246 653444 222799
rect 653600 218074 653628 226335
rect 659106 225584 659162 225593
rect 659106 225519 659162 225528
rect 654782 225040 654838 225049
rect 654782 224975 654838 224984
rect 658188 225004 658240 225010
rect 654138 220824 654194 220833
rect 654138 220759 654194 220768
rect 653588 218068 653640 218074
rect 653588 218010 653640 218016
rect 653770 217560 653826 217569
rect 653770 217495 653826 217504
rect 653404 213240 653456 213246
rect 653404 213182 653456 213188
rect 653784 210202 653812 217495
rect 654152 213790 654180 220759
rect 654796 216102 654824 224975
rect 658188 224946 658240 224952
rect 658200 224262 658228 224946
rect 658188 224256 658240 224262
rect 658188 224198 658240 224204
rect 656162 223952 656218 223961
rect 656162 223887 656218 223896
rect 654784 216096 654836 216102
rect 654784 216038 654836 216044
rect 656176 213926 656204 223887
rect 657542 223680 657598 223689
rect 657542 223615 657598 223624
rect 656714 218920 656770 218929
rect 656714 218855 656770 218864
rect 656164 213920 656216 213926
rect 656164 213862 656216 213868
rect 654140 213784 654192 213790
rect 654140 213726 654192 213732
rect 654784 213784 654836 213790
rect 654784 213726 654836 213732
rect 654600 213308 654652 213314
rect 654600 213250 654652 213256
rect 654612 210202 654640 213250
rect 652924 210174 653260 210202
rect 653476 210174 653812 210202
rect 654580 210174 654640 210202
rect 654796 210202 654824 213726
rect 656532 212560 656584 212566
rect 656532 212502 656584 212508
rect 656544 210202 656572 212502
rect 654796 210174 655132 210202
rect 656236 210174 656572 210202
rect 656728 210202 656756 218855
rect 657556 213314 657584 223615
rect 658922 222320 658978 222329
rect 658922 222255 658978 222264
rect 657910 215384 657966 215393
rect 657910 215319 657966 215328
rect 657544 213308 657596 213314
rect 657544 213250 657596 213256
rect 657924 212566 657952 215319
rect 658738 213480 658794 213489
rect 658738 213415 658794 213424
rect 658188 212900 658240 212906
rect 658188 212842 658240 212848
rect 657912 212560 657964 212566
rect 657912 212502 657964 212508
rect 658200 210202 658228 212842
rect 658752 210202 658780 213415
rect 658936 212906 658964 222255
rect 659120 215966 659148 225519
rect 659108 215960 659160 215966
rect 659108 215902 659160 215908
rect 660394 214568 660450 214577
rect 660394 214503 660450 214512
rect 658924 212900 658976 212906
rect 658924 212842 658976 212848
rect 659568 212696 659620 212702
rect 659568 212638 659620 212644
rect 659580 210202 659608 212638
rect 660408 210202 660436 214503
rect 660960 210202 660988 229230
rect 662328 229152 662380 229158
rect 662328 229094 662380 229100
rect 662052 227792 662104 227798
rect 662052 227734 662104 227740
rect 661498 213208 661554 213217
rect 661498 213143 661554 213152
rect 661512 210202 661540 213143
rect 662064 210202 662092 227734
rect 662340 219434 662368 229094
rect 656728 210174 656788 210202
rect 657892 210174 658228 210202
rect 658444 210174 658780 210202
rect 659548 210174 659608 210202
rect 660100 210174 660436 210202
rect 660652 210174 660988 210202
rect 661204 210174 661540 210202
rect 661756 210174 662092 210202
rect 662248 219406 662368 219434
rect 662248 210202 662276 219406
rect 662418 215656 662474 215665
rect 662418 215591 662474 215600
rect 662432 212702 662460 215591
rect 663156 213784 663208 213790
rect 663156 213726 663208 213732
rect 662420 212696 662472 212702
rect 662420 212638 662472 212644
rect 663168 210202 663196 213726
rect 663720 210202 663748 229706
rect 663904 227798 663932 229735
rect 663892 227792 663944 227798
rect 663892 227734 663944 227740
rect 664442 225856 664498 225865
rect 664442 225791 664498 225800
rect 664456 214606 664484 225791
rect 664444 214600 664496 214606
rect 664444 214542 664496 214548
rect 664812 214600 664864 214606
rect 664812 214542 664864 214548
rect 664260 213036 664312 213042
rect 664260 212978 664312 212984
rect 664272 210202 664300 212978
rect 664824 210202 664852 214542
rect 665100 213042 665128 231134
rect 665822 230480 665878 230489
rect 665822 230415 665878 230424
rect 665836 213790 665864 230415
rect 666006 230208 666062 230217
rect 666006 230143 666062 230152
rect 666020 214606 666048 230143
rect 666296 229294 666324 231542
rect 666468 230988 666520 230994
rect 666468 230930 666520 230936
rect 666284 229288 666336 229294
rect 666284 229230 666336 229236
rect 666480 229158 666508 230930
rect 666468 229152 666520 229158
rect 666468 229094 666520 229100
rect 667020 224120 667072 224126
rect 667020 224062 667072 224068
rect 667032 223689 667060 224062
rect 667018 223680 667074 223689
rect 667018 223615 667074 223624
rect 666652 223508 666704 223514
rect 666652 223450 666704 223456
rect 666664 218929 666692 223450
rect 667020 223168 667072 223174
rect 667020 223110 667072 223116
rect 667032 222329 667060 223110
rect 667018 222320 667074 222329
rect 667018 222255 667074 222264
rect 666650 218920 666706 218929
rect 666650 218855 666706 218864
rect 666650 217832 666706 217841
rect 666650 217767 666706 217776
rect 666008 214600 666060 214606
rect 666008 214542 666060 214548
rect 665824 213784 665876 213790
rect 665824 213726 665876 213732
rect 665088 213036 665140 213042
rect 665088 212978 665140 212984
rect 662248 210174 662308 210202
rect 662860 210174 663196 210202
rect 663412 210174 663748 210202
rect 663964 210174 664300 210202
rect 664516 210174 664852 210202
rect 632152 209568 632204 209574
rect 652024 209568 652076 209574
rect 632204 209516 632500 209522
rect 632152 209510 632500 209516
rect 652024 209510 652076 209516
rect 632164 209494 632500 209510
rect 666664 188873 666692 217767
rect 666834 215656 666890 215665
rect 666834 215591 666890 215600
rect 666848 198529 666876 215591
rect 667020 209092 667072 209098
rect 667020 209034 667072 209040
rect 666834 198520 666890 198529
rect 666834 198455 666890 198464
rect 666650 188864 666706 188873
rect 666650 188799 666706 188808
rect 667032 132705 667060 209034
rect 667216 134609 667244 280162
rect 667400 178809 667428 285670
rect 667584 181393 667612 287030
rect 667940 278044 667992 278050
rect 667940 277986 667992 277992
rect 667756 224460 667808 224466
rect 667756 224402 667808 224408
rect 667768 224233 667796 224402
rect 667754 224224 667810 224233
rect 667754 224159 667810 224168
rect 667756 223984 667808 223990
rect 667756 223926 667808 223932
rect 667768 220833 667796 223926
rect 667754 220824 667810 220833
rect 667754 220759 667810 220768
rect 667754 219464 667810 219473
rect 667754 219399 667810 219408
rect 667570 181384 667626 181393
rect 667570 181319 667626 181328
rect 667386 178800 667442 178809
rect 667386 178735 667442 178744
rect 667768 175001 667796 219399
rect 667952 184521 667980 277986
rect 668124 264376 668176 264382
rect 668124 264318 668176 264324
rect 668136 194313 668164 264318
rect 669228 264240 669280 264246
rect 669228 264182 669280 264188
rect 668674 232520 668730 232529
rect 668674 232455 668730 232464
rect 668306 231160 668362 231169
rect 668306 231095 668362 231104
rect 668320 204105 668348 231095
rect 668688 229094 668716 232455
rect 668860 231328 668912 231334
rect 668860 231270 668912 231276
rect 668872 229094 668900 231270
rect 669240 230474 669268 264182
rect 669056 230446 669268 230474
rect 669424 230466 669452 347239
rect 669962 302016 670018 302025
rect 669962 301951 670018 301960
rect 669780 234592 669832 234598
rect 669780 234534 669832 234540
rect 669596 234184 669648 234190
rect 669596 234126 669648 234132
rect 669608 230474 669636 234126
rect 669792 230474 669820 234534
rect 669976 230474 670004 301951
rect 670330 263800 670386 263809
rect 670330 263735 670386 263744
rect 670146 258496 670202 258505
rect 670146 258431 670202 258440
rect 670160 230474 670188 258431
rect 670344 238649 670372 263735
rect 670330 238640 670386 238649
rect 670330 238575 670386 238584
rect 670332 233096 670384 233102
rect 670332 233038 670384 233044
rect 668688 229066 668808 229094
rect 668872 229066 668992 229094
rect 668584 226976 668636 226982
rect 668584 226918 668636 226924
rect 668596 224890 668624 226918
rect 668596 224862 668716 224890
rect 668492 224732 668544 224738
rect 668492 224674 668544 224680
rect 668504 223938 668532 224674
rect 668412 223910 668532 223938
rect 668412 222170 668440 223910
rect 668412 222142 668532 222170
rect 668504 221785 668532 222142
rect 668490 221776 668546 221785
rect 668490 221711 668546 221720
rect 668688 219434 668716 224862
rect 668596 219406 668716 219434
rect 668306 204096 668362 204105
rect 668306 204031 668362 204040
rect 668398 198792 668454 198801
rect 668398 198727 668454 198736
rect 668122 194304 668178 194313
rect 668122 194239 668178 194248
rect 667938 184512 667994 184521
rect 667938 184447 667994 184456
rect 668216 178016 668268 178022
rect 668214 177984 668216 177993
rect 668268 177984 668270 177993
rect 668214 177919 668270 177928
rect 667754 174992 667810 175001
rect 667754 174927 667810 174936
rect 667940 174752 667992 174758
rect 667938 174720 667940 174729
rect 667992 174720 667994 174729
rect 667938 174655 667994 174664
rect 667940 169720 667992 169726
rect 667938 169688 667940 169697
rect 667992 169688 667994 169697
rect 667938 169623 667994 169632
rect 668032 164960 668084 164966
rect 668030 164928 668032 164937
rect 668084 164928 668086 164937
rect 668030 164863 668086 164872
rect 668216 160064 668268 160070
rect 668214 160032 668216 160041
rect 668268 160032 668270 160041
rect 668214 159967 668270 159976
rect 668216 155168 668268 155174
rect 668214 155136 668216 155145
rect 668268 155136 668270 155145
rect 668214 155071 668270 155080
rect 668412 143721 668440 198727
rect 668398 143712 668454 143721
rect 668398 143647 668454 143656
rect 668596 138825 668624 219406
rect 668780 163305 668808 229066
rect 668964 199209 668992 229066
rect 669056 220538 669084 230446
rect 669332 230438 669452 230466
rect 669516 230446 669636 230474
rect 669700 230446 669820 230474
rect 669884 230446 670004 230474
rect 670068 230446 670188 230474
rect 669332 229094 669360 230438
rect 669516 229094 669544 230446
rect 669240 229066 669360 229094
rect 669424 229066 669544 229094
rect 669700 229094 669728 230446
rect 669700 229066 669820 229094
rect 669240 220674 669268 229066
rect 669424 220930 669452 229066
rect 669792 221406 669820 229066
rect 669884 222194 669912 230446
rect 670068 222850 670096 230446
rect 670344 224641 670372 233038
rect 670330 224632 670386 224641
rect 670330 224567 670386 224576
rect 670528 223961 670556 392527
rect 670974 296304 671030 296313
rect 670974 296239 671030 296248
rect 670988 293865 671016 296239
rect 670974 293856 671030 293865
rect 670974 293791 671030 293800
rect 671356 278730 671384 571066
rect 671988 569968 672040 569974
rect 671988 569910 672040 569916
rect 671802 557560 671858 557569
rect 671802 557495 671858 557504
rect 671620 532024 671672 532030
rect 671620 531966 671672 531972
rect 671632 488510 671660 531966
rect 671620 488504 671672 488510
rect 671620 488446 671672 488452
rect 671816 483206 671844 557495
rect 671804 483200 671856 483206
rect 671804 483142 671856 483148
rect 672000 454866 672028 569910
rect 672184 530942 672212 609039
rect 672354 604344 672410 604353
rect 672354 604279 672410 604288
rect 672172 530936 672224 530942
rect 672172 530878 672224 530884
rect 672368 528902 672396 604279
rect 672538 597408 672594 597417
rect 672538 597343 672594 597352
rect 672356 528896 672408 528902
rect 672356 528838 672408 528844
rect 672552 528086 672580 597343
rect 672736 573617 672764 620986
rect 672722 573608 672778 573617
rect 672722 573543 672778 573552
rect 673012 572801 673040 648751
rect 673196 619449 673224 696895
rect 673472 682417 673500 734159
rect 673656 721754 673684 736906
rect 673564 721726 673684 721754
rect 673564 698294 673592 721726
rect 673748 707577 673776 782614
rect 673920 780020 673972 780026
rect 673920 779962 673972 779968
rect 673932 760394 673960 779962
rect 674852 779714 674880 785182
rect 675128 784638 675418 784666
rect 675128 784310 675156 784638
rect 675116 784304 675168 784310
rect 675116 784246 675168 784252
rect 675392 784168 675444 784174
rect 675392 784110 675444 784116
rect 675404 783972 675432 784110
rect 675128 783346 675418 783374
rect 675128 782678 675156 783346
rect 675116 782672 675168 782678
rect 675116 782614 675168 782620
rect 675300 782536 675352 782542
rect 675300 782478 675352 782484
rect 675312 781402 675340 782478
rect 675312 781374 675432 781402
rect 675024 781108 675076 781114
rect 675024 781050 675076 781056
rect 675036 780994 675064 781050
rect 674944 780966 675064 780994
rect 674944 779906 674972 780966
rect 675404 780844 675432 781374
rect 675312 780422 675432 780450
rect 675312 780314 675340 780422
rect 675128 780286 675340 780314
rect 675404 780300 675432 780422
rect 675128 780026 675156 780286
rect 675116 780020 675168 780026
rect 675116 779962 675168 779968
rect 674944 779878 675248 779906
rect 675220 779714 675248 779878
rect 674852 779686 675156 779714
rect 675220 779686 675340 779714
rect 674378 779376 674434 779385
rect 674378 779311 674434 779320
rect 673840 760366 673960 760394
rect 673840 721562 673868 760366
rect 674010 735040 674066 735049
rect 674010 734975 674066 734984
rect 674024 721721 674052 734975
rect 674392 726442 674420 779311
rect 674562 778832 674618 778841
rect 674562 778767 674618 778776
rect 674576 726782 674604 778767
rect 674932 778388 674984 778394
rect 674932 778330 674984 778336
rect 674944 777073 674972 778330
rect 674930 777064 674986 777073
rect 674930 776999 674986 777008
rect 674930 775704 674986 775713
rect 674930 775639 674932 775648
rect 674984 775639 674986 775648
rect 674932 775610 674984 775616
rect 675128 750734 675156 779686
rect 675312 778478 675340 779686
rect 675496 779385 675524 779688
rect 675482 779376 675538 779385
rect 675482 779311 675538 779320
rect 675496 778841 675524 779008
rect 675482 778832 675538 778841
rect 675482 778767 675538 778776
rect 675312 778450 675418 778478
rect 675404 777481 675432 777852
rect 675390 777472 675446 777481
rect 675390 777407 675446 777416
rect 675482 777064 675538 777073
rect 675300 777028 675352 777034
rect 675482 776999 675538 777008
rect 675300 776970 675352 776976
rect 675312 776914 675340 776970
rect 675220 776886 675340 776914
rect 675220 775350 675248 776886
rect 675496 776628 675524 776999
rect 675404 775713 675432 776016
rect 675390 775704 675446 775713
rect 675390 775639 675446 775648
rect 675220 775322 675418 775350
rect 675404 773650 675432 774180
rect 675312 773622 675432 773650
rect 675312 773430 675340 773622
rect 675300 773424 675352 773430
rect 675300 773366 675352 773372
rect 674852 750706 675156 750734
rect 674852 734174 674880 750706
rect 675392 746632 675444 746638
rect 675392 746574 675444 746580
rect 675404 743852 675432 746574
rect 675114 743336 675170 743345
rect 675170 743294 675418 743322
rect 675114 743271 675170 743280
rect 675404 742218 675432 742696
rect 675392 742212 675444 742218
rect 675392 742154 675444 742160
rect 675312 742070 675432 742098
rect 675312 742030 675340 742070
rect 675128 742002 675340 742030
rect 675404 742016 675432 742070
rect 675128 741198 675156 742002
rect 675116 741192 675168 741198
rect 675116 741134 675168 741140
rect 674668 734146 674880 734174
rect 674944 740166 675418 740194
rect 674668 729722 674696 734146
rect 674944 731134 674972 740166
rect 675128 739622 675418 739650
rect 675128 738478 675156 739622
rect 675404 738682 675432 739024
rect 675392 738676 675444 738682
rect 675392 738618 675444 738624
rect 675116 738472 675168 738478
rect 675116 738414 675168 738420
rect 675128 738330 675418 738358
rect 675128 738177 675156 738330
rect 675114 738168 675170 738177
rect 675114 738103 675170 738112
rect 675128 735882 675340 735910
rect 675128 735622 675156 735882
rect 675312 735842 675340 735882
rect 675404 735842 675432 735896
rect 675312 735814 675432 735842
rect 675300 735752 675352 735758
rect 675300 735694 675352 735700
rect 675116 735616 675168 735622
rect 675116 735558 675168 735564
rect 675116 734256 675168 734262
rect 675116 734198 675168 734204
rect 675128 731898 675156 734198
rect 675312 733493 675340 735694
rect 675496 735049 675524 735319
rect 675482 735040 675538 735049
rect 675482 734975 675538 734984
rect 675496 734233 675524 734672
rect 675482 734224 675538 734233
rect 675482 734159 675538 734168
rect 675496 733825 675524 734031
rect 675482 733816 675538 733825
rect 675482 733751 675538 733760
rect 675312 733465 675418 733493
rect 675312 732822 675418 732850
rect 675312 732766 675340 732822
rect 675300 732760 675352 732766
rect 675300 732702 675352 732708
rect 675128 731870 675432 731898
rect 675404 731612 675432 731870
rect 674932 731128 674984 731134
rect 674932 731070 674984 731076
rect 674944 730986 675418 731014
rect 674668 729694 674788 729722
rect 674564 726776 674616 726782
rect 674564 726718 674616 726724
rect 674760 726578 674788 729694
rect 674748 726572 674800 726578
rect 674748 726514 674800 726520
rect 674380 726436 674432 726442
rect 674380 726378 674432 726384
rect 674944 721721 674972 730986
rect 675116 730924 675168 730930
rect 675116 730866 675168 730872
rect 675128 729881 675156 730866
rect 675298 730824 675354 730833
rect 675298 730759 675354 730768
rect 675114 729872 675170 729881
rect 675114 729807 675170 729816
rect 675312 727274 675340 730759
rect 675496 730153 675524 730351
rect 675482 730144 675538 730153
rect 675482 730079 675538 730088
rect 675496 728793 675524 729164
rect 675482 728784 675538 728793
rect 675482 728719 675538 728728
rect 675220 727246 675340 727274
rect 675220 726730 675248 727246
rect 683396 726776 683448 726782
rect 675220 726702 675340 726730
rect 683396 726718 683448 726724
rect 675312 721750 675340 726702
rect 682382 726608 682438 726617
rect 681004 726572 681056 726578
rect 682382 726543 682438 726552
rect 681004 726514 681056 726520
rect 675300 721744 675352 721750
rect 674010 721712 674066 721721
rect 674010 721647 674066 721656
rect 674930 721712 674986 721721
rect 675300 721686 675352 721692
rect 674930 721647 674986 721656
rect 673840 721534 673960 721562
rect 673932 721070 673960 721534
rect 675300 721268 675352 721274
rect 675300 721210 675352 721216
rect 673920 721064 673972 721070
rect 673920 721006 673972 721012
rect 675312 720866 675340 721210
rect 675300 720860 675352 720866
rect 675300 720802 675352 720808
rect 674472 720520 674524 720526
rect 674472 720462 674524 720468
rect 675300 720520 675352 720526
rect 675300 720462 675352 720468
rect 674010 719808 674066 719817
rect 673840 719766 674010 719794
rect 673840 707690 673868 719766
rect 674010 719743 674066 719752
rect 674288 716508 674340 716514
rect 674288 716450 674340 716456
rect 674300 716394 674328 716450
rect 674024 716366 674328 716394
rect 674024 716310 674052 716366
rect 674012 716304 674064 716310
rect 674012 716246 674064 716252
rect 674012 715760 674064 715766
rect 674010 715728 674012 715737
rect 674064 715728 674066 715737
rect 674010 715663 674066 715672
rect 674012 715352 674064 715358
rect 674010 715320 674012 715329
rect 674064 715320 674066 715329
rect 674010 715255 674066 715264
rect 674288 715080 674340 715086
rect 674024 715028 674288 715034
rect 674024 715022 674340 715028
rect 674024 715018 674328 715022
rect 674012 715012 674328 715018
rect 674064 715006 674328 715012
rect 674012 714954 674064 714960
rect 674288 714944 674340 714950
rect 674024 714892 674288 714898
rect 674024 714886 674340 714892
rect 674024 714882 674328 714886
rect 674012 714876 674328 714882
rect 674064 714870 674328 714876
rect 674012 714818 674064 714824
rect 674012 714536 674064 714542
rect 674010 714504 674012 714513
rect 674064 714504 674066 714513
rect 674010 714439 674066 714448
rect 674012 713720 674064 713726
rect 674010 713688 674012 713697
rect 674064 713688 674066 713697
rect 674010 713623 674066 713632
rect 674010 713280 674066 713289
rect 674010 713215 674012 713224
rect 674064 713215 674066 713224
rect 674012 713186 674064 713192
rect 674010 712464 674066 712473
rect 674010 712399 674012 712408
rect 674064 712399 674066 712408
rect 674012 712370 674064 712376
rect 674012 710048 674064 710054
rect 674010 710016 674012 710025
rect 674064 710016 674066 710025
rect 674010 709951 674066 709960
rect 674288 709776 674340 709782
rect 674024 709724 674288 709730
rect 674024 709718 674340 709724
rect 674024 709702 674328 709718
rect 674024 709374 674052 709702
rect 674012 709368 674064 709374
rect 674012 709310 674064 709316
rect 674012 709232 674064 709238
rect 674010 709200 674012 709209
rect 674064 709200 674066 709209
rect 674010 709135 674066 709144
rect 674288 708756 674340 708762
rect 674288 708698 674340 708704
rect 674300 708642 674328 708698
rect 674024 708614 674328 708642
rect 674024 708286 674052 708614
rect 674012 708280 674064 708286
rect 674012 708222 674064 708228
rect 673840 707662 674052 707690
rect 673734 707568 673790 707577
rect 673734 707503 673790 707512
rect 674024 707418 674052 707662
rect 673840 707390 674052 707418
rect 673840 702434 673868 707390
rect 674484 707198 674512 720462
rect 675312 712065 675340 720462
rect 676034 716544 676090 716553
rect 676034 716479 676036 716488
rect 676088 716479 676090 716488
rect 676036 716450 676088 716456
rect 676034 716136 676090 716145
rect 676034 716071 676090 716080
rect 676048 715086 676076 716071
rect 676036 715080 676088 715086
rect 676036 715022 676088 715028
rect 676036 714944 676088 714950
rect 676034 714912 676036 714921
rect 676088 714912 676090 714921
rect 676034 714847 676090 714856
rect 675298 712056 675354 712065
rect 675298 711991 675354 712000
rect 681016 710841 681044 726514
rect 682396 711249 682424 726543
rect 682382 711240 682438 711249
rect 682382 711175 682438 711184
rect 681002 710832 681058 710841
rect 681002 710767 681058 710776
rect 676034 710424 676090 710433
rect 676034 710359 676090 710368
rect 676048 709782 676076 710359
rect 676036 709776 676088 709782
rect 676036 709718 676088 709724
rect 676034 708792 676090 708801
rect 676034 708727 676036 708736
rect 676088 708727 676090 708736
rect 676036 708698 676088 708704
rect 674472 707192 674524 707198
rect 676036 707192 676088 707198
rect 674472 707134 674524 707140
rect 676034 707160 676036 707169
rect 676088 707160 676090 707169
rect 676034 707095 676090 707104
rect 683408 706761 683436 726718
rect 684040 726436 684092 726442
rect 684040 726378 684092 726384
rect 684052 707985 684080 726378
rect 684222 726336 684278 726345
rect 684222 726271 684278 726280
rect 684236 709617 684264 726271
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 684222 709608 684278 709617
rect 684222 709543 684278 709552
rect 684038 707976 684094 707985
rect 684038 707911 684094 707920
rect 683394 706752 683450 706761
rect 683394 706687 683450 706696
rect 675850 706344 675906 706353
rect 675850 706279 675906 706288
rect 674012 705356 674064 705362
rect 674288 705356 674340 705362
rect 674064 705316 674288 705344
rect 674012 705298 674064 705304
rect 674288 705298 674340 705304
rect 675864 705226 675892 706279
rect 683118 705528 683174 705537
rect 683118 705463 683174 705472
rect 683132 705362 683160 705463
rect 683120 705356 683172 705362
rect 683120 705298 683172 705304
rect 674012 705220 674064 705226
rect 674288 705220 674340 705226
rect 674064 705168 674288 705194
rect 674012 705166 674340 705168
rect 674012 705162 674064 705166
rect 674288 705162 674340 705166
rect 675852 705220 675904 705226
rect 675852 705162 675904 705168
rect 676034 705120 676090 705129
rect 676034 705055 676090 705064
rect 676048 703934 676076 705055
rect 674288 703928 674340 703934
rect 674024 703876 674288 703882
rect 674024 703870 674340 703876
rect 676036 703928 676088 703934
rect 676036 703870 676088 703876
rect 674024 703866 674328 703870
rect 674012 703860 674328 703866
rect 674064 703854 674328 703860
rect 674012 703802 674064 703808
rect 673840 702406 673960 702434
rect 673736 701208 673788 701214
rect 673734 701176 673736 701185
rect 673788 701176 673790 701185
rect 673734 701111 673790 701120
rect 673564 698266 673684 698294
rect 673458 682408 673514 682417
rect 673458 682343 673514 682352
rect 673656 682258 673684 698266
rect 673932 695534 673960 702406
rect 675114 701176 675170 701185
rect 675114 701111 675170 701120
rect 675128 698889 675156 701111
rect 675128 698861 675418 698889
rect 675128 698329 675418 698337
rect 675114 698320 675418 698329
rect 675170 698309 675418 698320
rect 675114 698255 675170 698264
rect 675128 697666 675418 697694
rect 675128 696969 675156 697666
rect 675114 696960 675170 696969
rect 675114 696895 675170 696904
rect 675496 696833 675524 697035
rect 675482 696824 675538 696833
rect 675482 696759 675538 696768
rect 673932 695506 674236 695534
rect 674010 693016 674066 693025
rect 674010 692951 674066 692960
rect 674024 690418 674052 692951
rect 673472 682230 673684 682258
rect 673748 690390 674052 690418
rect 673472 682145 673500 682230
rect 673458 682136 673514 682145
rect 673458 682071 673514 682080
rect 673550 671392 673606 671401
rect 673550 671327 673552 671336
rect 673604 671327 673606 671336
rect 673552 671298 673604 671304
rect 673552 671152 673604 671158
rect 673552 671094 673604 671100
rect 673564 670993 673592 671094
rect 673550 670984 673606 670993
rect 673550 670919 673606 670928
rect 673368 670608 673420 670614
rect 673368 670550 673420 670556
rect 673550 670576 673606 670585
rect 673380 670177 673408 670550
rect 673550 670511 673606 670520
rect 673366 670168 673422 670177
rect 673366 670103 673422 670112
rect 673368 669656 673420 669662
rect 673368 669598 673420 669604
rect 673380 669497 673408 669598
rect 673564 669526 673592 670511
rect 673552 669520 673604 669526
rect 673366 669488 673422 669497
rect 673552 669462 673604 669468
rect 673366 669423 673422 669432
rect 673550 668944 673606 668953
rect 673550 668879 673606 668888
rect 673564 668710 673592 668879
rect 673552 668704 673604 668710
rect 673552 668646 673604 668652
rect 673552 668568 673604 668574
rect 673550 668536 673552 668545
rect 673604 668536 673606 668545
rect 673550 668471 673606 668480
rect 673552 668160 673604 668166
rect 673550 668128 673552 668137
rect 673604 668128 673606 668137
rect 673550 668063 673606 668072
rect 673550 667720 673606 667729
rect 673550 667655 673606 667664
rect 673564 666942 673592 667655
rect 673552 666936 673604 666942
rect 673552 666878 673604 666884
rect 673550 666768 673606 666777
rect 673550 666703 673606 666712
rect 673564 666602 673592 666703
rect 673552 666596 673604 666602
rect 673552 666538 673604 666544
rect 673552 665304 673604 665310
rect 673550 665272 673552 665281
rect 673604 665272 673606 665281
rect 673550 665207 673606 665216
rect 673368 665168 673420 665174
rect 673368 665110 673420 665116
rect 673380 664057 673408 665110
rect 673550 664456 673606 664465
rect 673550 664391 673552 664400
rect 673604 664391 673606 664400
rect 673552 664362 673604 664368
rect 673366 664048 673422 664057
rect 673366 663983 673422 663992
rect 673552 663944 673604 663950
rect 673552 663886 673604 663892
rect 673564 663785 673592 663886
rect 673550 663776 673606 663785
rect 673550 663711 673606 663720
rect 673552 663400 673604 663406
rect 673552 663342 673604 663348
rect 673564 662017 673592 663342
rect 673550 662008 673606 662017
rect 673550 661943 673606 661952
rect 673366 659696 673422 659705
rect 673366 659631 673422 659640
rect 673182 619440 673238 619449
rect 673182 619375 673238 619384
rect 673184 608660 673236 608666
rect 673184 608602 673236 608608
rect 673196 608297 673224 608602
rect 673182 608288 673238 608297
rect 673182 608223 673238 608232
rect 673184 599004 673236 599010
rect 673184 598946 673236 598952
rect 673196 598097 673224 598946
rect 673182 598088 673238 598097
rect 673182 598023 673238 598032
rect 673182 581088 673238 581097
rect 673182 581023 673184 581032
rect 673236 581023 673238 581032
rect 673184 580994 673236 581000
rect 673184 580304 673236 580310
rect 673182 580272 673184 580281
rect 673236 580272 673238 580281
rect 673182 580207 673238 580216
rect 673184 580032 673236 580038
rect 673182 580000 673184 580009
rect 673236 580000 673238 580009
rect 673182 579935 673238 579944
rect 673182 579728 673238 579737
rect 673182 579663 673184 579672
rect 673236 579663 673238 579672
rect 673184 579634 673236 579640
rect 673184 578944 673236 578950
rect 673182 578912 673184 578921
rect 673236 578912 673238 578921
rect 673182 578847 673238 578856
rect 673184 578264 673236 578270
rect 673184 578206 673236 578212
rect 673196 577969 673224 578206
rect 673182 577960 673238 577969
rect 673182 577895 673238 577904
rect 673182 577688 673238 577697
rect 673182 577623 673184 577632
rect 673236 577623 673238 577632
rect 673184 577594 673236 577600
rect 673184 577448 673236 577454
rect 673182 577416 673184 577425
rect 673236 577416 673238 577425
rect 673182 577351 673238 577360
rect 673184 577176 673236 577182
rect 673182 577144 673184 577153
rect 673236 577144 673238 577153
rect 673182 577079 673238 577088
rect 673184 576904 673236 576910
rect 673182 576872 673184 576881
rect 673236 576872 673238 576881
rect 673182 576807 673238 576816
rect 672998 572792 673054 572801
rect 672998 572727 673054 572736
rect 673090 559056 673146 559065
rect 673090 558991 673146 559000
rect 672906 555248 672962 555257
rect 672906 555183 672962 555192
rect 672722 554840 672778 554849
rect 672722 554775 672724 554784
rect 672776 554775 672778 554784
rect 672724 554746 672776 554752
rect 672722 533624 672778 533633
rect 672722 533559 672778 533568
rect 672540 528080 672592 528086
rect 672540 528022 672592 528028
rect 672540 490748 672592 490754
rect 672540 490690 672592 490696
rect 672552 489954 672580 490690
rect 672736 490113 672764 533559
rect 672920 490754 672948 555183
rect 672908 490748 672960 490754
rect 672908 490690 672960 490696
rect 672906 490512 672962 490521
rect 672906 490447 672962 490456
rect 672722 490104 672778 490113
rect 672722 490039 672778 490048
rect 672552 489926 672672 489954
rect 672448 489660 672500 489666
rect 672448 489602 672500 489608
rect 672000 454850 672120 454866
rect 672000 454844 672132 454850
rect 672000 454838 672080 454844
rect 672080 454786 672132 454792
rect 672264 453960 672316 453966
rect 672262 453928 672264 453937
rect 672316 453928 672318 453937
rect 672262 453863 672318 453872
rect 672460 401985 672488 489602
rect 672644 486062 672672 489926
rect 672632 486056 672684 486062
rect 672632 485998 672684 486004
rect 672920 485774 672948 490447
rect 672644 485746 672948 485774
rect 672644 402529 672672 485746
rect 673104 484809 673132 558991
rect 673090 484800 673146 484809
rect 673090 484735 673146 484744
rect 673380 455870 673408 659631
rect 673552 626000 673604 626006
rect 673550 625968 673552 625977
rect 673604 625968 673606 625977
rect 673550 625903 673606 625912
rect 673748 621014 673776 690390
rect 674010 690296 674066 690305
rect 674010 690231 674012 690240
rect 674064 690231 674066 690240
rect 674012 690202 674064 690208
rect 674208 689466 674236 695506
rect 675128 695181 675418 695209
rect 675128 694929 675156 695181
rect 675114 694920 675170 694929
rect 675114 694855 675170 694864
rect 675312 694742 675432 694770
rect 675114 694648 675170 694657
rect 675312 694634 675340 694742
rect 675170 694606 675340 694634
rect 675404 694620 675432 694742
rect 675114 694583 675170 694592
rect 674668 693994 675418 694022
rect 674472 690056 674524 690062
rect 674472 689998 674524 690004
rect 673932 689438 674236 689466
rect 673932 663406 673960 689438
rect 674484 688634 674512 689998
rect 674668 689330 674696 693994
rect 675496 693025 675524 693328
rect 675482 693016 675538 693025
rect 675482 692951 675538 692960
rect 675128 690866 675418 690894
rect 675128 690577 675156 690866
rect 675114 690568 675170 690577
rect 675114 690503 675170 690512
rect 675128 690322 675340 690350
rect 674930 690296 674986 690305
rect 674930 690231 674986 690240
rect 674116 688606 674512 688634
rect 674576 689302 674696 689330
rect 673920 663400 673972 663406
rect 673920 663342 673972 663348
rect 673918 663232 673974 663241
rect 673918 663167 673974 663176
rect 673932 662454 673960 663167
rect 673920 662448 673972 662454
rect 673920 662390 673972 662396
rect 673920 661632 673972 661638
rect 673918 661600 673920 661609
rect 673972 661600 673974 661609
rect 673918 661535 673974 661544
rect 673918 661192 673974 661201
rect 673918 661127 673920 661136
rect 673972 661127 673974 661136
rect 673920 661098 673972 661104
rect 673920 660136 673972 660142
rect 673918 660104 673920 660113
rect 673972 660104 673974 660113
rect 673918 660039 673974 660048
rect 673918 655616 673974 655625
rect 673918 655551 673920 655560
rect 673972 655551 673974 655560
rect 673920 655522 673972 655528
rect 674116 654134 674144 688606
rect 674576 685874 674604 689302
rect 674944 689042 674972 690231
rect 675128 690062 675156 690322
rect 675312 690282 675340 690322
rect 675404 690282 675432 690336
rect 675312 690254 675432 690282
rect 675116 690056 675168 690062
rect 675116 689998 675168 690004
rect 675312 689710 675432 689738
rect 675312 689670 675340 689710
rect 675128 689642 675340 689670
rect 675404 689656 675432 689710
rect 675128 689489 675156 689642
rect 675114 689480 675170 689489
rect 675114 689415 675170 689424
rect 674932 689036 674984 689042
rect 674932 688978 674984 688984
rect 675220 689030 675418 689058
rect 675220 688922 675248 689030
rect 674484 685846 674604 685874
rect 674668 688894 675248 688922
rect 674288 684004 674340 684010
rect 674288 683946 674340 683952
rect 674300 676214 674328 683946
rect 674484 676214 674512 685846
rect 674668 684010 674696 688894
rect 675116 688832 675168 688838
rect 674930 688800 674986 688809
rect 675116 688774 675168 688780
rect 674930 688735 674986 688744
rect 674944 686678 674972 688735
rect 675128 688514 675156 688774
rect 675128 688486 675340 688514
rect 675312 688378 675340 688486
rect 675404 688378 675432 688500
rect 675312 688350 675432 688378
rect 675114 687848 675170 687857
rect 675170 687806 675418 687834
rect 675114 687783 675170 687792
rect 674944 686650 675340 686678
rect 675312 686610 675340 686650
rect 675404 686610 675432 686664
rect 675312 686582 675432 686610
rect 675298 686216 675354 686225
rect 675298 686151 675354 686160
rect 675022 685944 675078 685953
rect 675022 685879 675078 685888
rect 674656 684004 674708 684010
rect 674656 683946 674708 683952
rect 674748 682440 674800 682446
rect 674746 682408 674748 682417
rect 674800 682408 674802 682417
rect 674746 682343 674802 682352
rect 675036 676433 675064 685879
rect 675022 676424 675078 676433
rect 675022 676359 675078 676368
rect 674300 676186 674420 676214
rect 674484 676186 674696 676214
rect 674116 654106 674328 654134
rect 674012 645924 674064 645930
rect 674012 645866 674064 645872
rect 674024 645561 674052 645866
rect 674010 645552 674066 645561
rect 674010 645487 674066 645496
rect 674010 643512 674066 643521
rect 674010 643447 674066 643456
rect 674024 643226 674052 643447
rect 674024 643198 674236 643226
rect 674012 643136 674064 643142
rect 674010 643104 674012 643113
rect 674064 643104 674066 643113
rect 674010 643039 674066 643048
rect 673918 641744 673974 641753
rect 673918 641679 673974 641688
rect 673932 640334 673960 641679
rect 673472 620986 673776 621014
rect 673840 640306 673960 640334
rect 673472 619290 673500 620986
rect 673644 620424 673696 620430
rect 673644 620366 673696 620372
rect 673656 620265 673684 620366
rect 673642 620256 673698 620265
rect 673642 620191 673698 620200
rect 673644 619880 673696 619886
rect 673642 619848 673644 619857
rect 673696 619848 673698 619857
rect 673642 619783 673698 619792
rect 673472 619262 673684 619290
rect 673656 619177 673684 619262
rect 673642 619168 673698 619177
rect 673642 619103 673698 619112
rect 673642 618216 673698 618225
rect 673642 618151 673698 618160
rect 673656 617982 673684 618151
rect 673644 617976 673696 617982
rect 673644 617918 673696 617924
rect 673642 617808 673698 617817
rect 673642 617743 673698 617752
rect 673656 616894 673684 617743
rect 673644 616888 673696 616894
rect 673644 616830 673696 616836
rect 673644 615528 673696 615534
rect 673642 615496 673644 615505
rect 673696 615496 673698 615505
rect 673642 615431 673698 615440
rect 673642 614952 673698 614961
rect 673642 614887 673644 614896
rect 673696 614887 673698 614896
rect 673644 614858 673696 614864
rect 673642 611416 673698 611425
rect 673642 611351 673644 611360
rect 673696 611351 673698 611360
rect 673644 611322 673696 611328
rect 673840 600681 673868 640306
rect 674208 639826 674236 643198
rect 674024 639798 674236 639826
rect 674024 627914 674052 639798
rect 674300 637498 674328 654106
rect 674392 637650 674420 676186
rect 674668 649994 674696 676186
rect 674838 669896 674894 669905
rect 674838 669831 674894 669840
rect 674852 669526 674880 669831
rect 674840 669520 674892 669526
rect 674840 669462 674892 669468
rect 674838 667448 674894 667457
rect 674838 667383 674894 667392
rect 674852 667078 674880 667383
rect 674840 667072 674892 667078
rect 674840 667014 674892 667020
rect 675312 666505 675340 686151
rect 675496 685681 675524 685984
rect 675482 685672 675538 685681
rect 675482 685607 675538 685616
rect 675496 685001 675524 685372
rect 675482 684992 675538 685001
rect 675482 684927 675538 684936
rect 675496 683913 675524 684148
rect 675482 683904 675538 683913
rect 675482 683839 675538 683848
rect 684130 682680 684186 682689
rect 684130 682615 684186 682624
rect 675484 682576 675536 682582
rect 675484 682518 675536 682524
rect 683212 682576 683264 682582
rect 683212 682518 683264 682524
rect 675496 682145 675524 682518
rect 675482 682136 675538 682145
rect 675482 682071 675538 682080
rect 676496 669520 676548 669526
rect 676494 669488 676496 669497
rect 676548 669488 676550 669497
rect 676494 669423 676550 669432
rect 676496 667072 676548 667078
rect 676494 667040 676496 667049
rect 676548 667040 676550 667049
rect 676494 666975 676550 666984
rect 675298 666496 675354 666505
rect 675298 666431 675354 666440
rect 676034 664864 676090 664873
rect 676034 664799 676090 664808
rect 676048 663814 676076 664799
rect 674840 663808 674892 663814
rect 674838 663776 674840 663785
rect 676036 663808 676088 663814
rect 674892 663776 674894 663785
rect 683224 663785 683252 682518
rect 683488 682440 683540 682446
rect 683488 682382 683540 682388
rect 676036 663750 676088 663756
rect 683210 663776 683266 663785
rect 674838 663711 674894 663720
rect 683210 663711 683266 663720
rect 683500 662969 683528 682382
rect 684144 666233 684172 682615
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 684130 666224 684186 666233
rect 684130 666159 684186 666168
rect 683486 662960 683542 662969
rect 683486 662895 683542 662904
rect 674838 660104 674894 660113
rect 674838 660039 674894 660048
rect 683118 660104 683174 660113
rect 683118 660039 683174 660048
rect 674852 659870 674880 660039
rect 683132 659870 683160 660039
rect 674840 659864 674892 659870
rect 674840 659806 674892 659812
rect 683120 659864 683172 659870
rect 683120 659806 683172 659812
rect 675114 655616 675170 655625
rect 675114 655551 675170 655560
rect 675128 653698 675156 655551
rect 675128 653670 675418 653698
rect 675404 652905 675432 653140
rect 675390 652896 675446 652905
rect 675390 652831 675446 652840
rect 675312 652582 675432 652610
rect 675114 652488 675170 652497
rect 675312 652474 675340 652582
rect 675170 652446 675340 652474
rect 675404 652460 675432 652582
rect 675114 652423 675170 652432
rect 674852 651834 675418 651862
rect 674668 649966 674788 649994
rect 674564 644632 674616 644638
rect 674564 644574 674616 644580
rect 674392 637622 674512 637650
rect 674288 637492 674340 637498
rect 674288 637434 674340 637440
rect 674484 636194 674512 637622
rect 674576 636970 674604 644574
rect 674760 642649 674788 649966
rect 674852 642818 674880 651834
rect 675128 649998 675340 650026
rect 675128 649994 675156 649998
rect 674944 649966 675156 649994
rect 675312 649994 675340 649998
rect 675404 649994 675432 650012
rect 675312 649966 675432 649994
rect 674944 647234 674972 649966
rect 675404 649233 675432 649468
rect 675390 649224 675446 649233
rect 675390 649159 675446 649168
rect 675114 648816 675170 648825
rect 675170 648774 675418 648802
rect 675114 648751 675170 648760
rect 675404 647873 675432 648176
rect 675390 647864 675446 647873
rect 675390 647799 675446 647808
rect 674944 647206 675064 647234
rect 675036 646105 675064 647206
rect 675022 646096 675078 646105
rect 675022 646031 675078 646040
rect 675114 645824 675170 645833
rect 675114 645759 675170 645768
rect 675128 645674 675156 645759
rect 675128 645646 675418 645674
rect 675114 645552 675170 645561
rect 675114 645487 675170 645496
rect 675128 643294 675156 645487
rect 675312 645102 675418 645130
rect 675312 644638 675340 645102
rect 675300 644632 675352 644638
rect 675300 644574 675352 644580
rect 675312 644461 675418 644489
rect 675312 644337 675340 644461
rect 675298 644328 675354 644337
rect 675298 644263 675354 644272
rect 675312 643810 675418 643838
rect 675312 643521 675340 643810
rect 675298 643512 675354 643521
rect 675298 643447 675354 643456
rect 675128 643266 675418 643294
rect 675114 643104 675170 643113
rect 675114 643039 675170 643048
rect 674852 642790 675064 642818
rect 674668 642621 674788 642649
rect 674668 642410 674696 642621
rect 674668 642382 674788 642410
rect 674760 641102 674788 642382
rect 674748 641096 674800 641102
rect 674748 641038 674800 641044
rect 674748 640892 674800 640898
rect 674748 640834 674800 640840
rect 674760 640336 674788 640834
rect 674668 640308 674788 640336
rect 674668 639690 674696 640308
rect 674838 640248 674894 640257
rect 674838 640183 674840 640192
rect 674892 640183 674894 640192
rect 674840 640154 674892 640160
rect 675036 640166 675064 642790
rect 675128 641458 675156 643039
rect 675312 642621 675418 642649
rect 675312 641753 675340 642621
rect 675298 641744 675354 641753
rect 675298 641679 675354 641688
rect 675128 641430 675418 641458
rect 675220 640781 675418 640809
rect 675220 640286 675248 640781
rect 675208 640280 675260 640286
rect 675208 640222 675260 640228
rect 675036 640138 675248 640166
rect 675024 639940 675076 639946
rect 675024 639882 675076 639888
rect 674840 639804 674892 639810
rect 674840 639746 674892 639752
rect 674668 639662 674788 639690
rect 674760 637770 674788 639662
rect 674852 637922 674880 639746
rect 674852 637894 674972 637922
rect 674748 637764 674800 637770
rect 674748 637706 674800 637712
rect 674748 637628 674800 637634
rect 674748 637570 674800 637576
rect 674760 637090 674788 637570
rect 674748 637084 674800 637090
rect 674748 637026 674800 637032
rect 674576 636942 674788 636970
rect 674392 636166 674512 636194
rect 674024 627886 674236 627914
rect 674010 626376 674066 626385
rect 674010 626311 674066 626320
rect 674024 625734 674052 626311
rect 674012 625728 674064 625734
rect 674012 625670 674064 625676
rect 674010 625560 674066 625569
rect 674010 625495 674066 625504
rect 674024 625190 674052 625495
rect 674012 625184 674064 625190
rect 674012 625126 674064 625132
rect 674012 625048 674064 625054
rect 674010 625016 674012 625025
rect 674064 625016 674066 625025
rect 674010 624951 674066 624960
rect 674010 624744 674066 624753
rect 674010 624679 674012 624688
rect 674064 624679 674066 624688
rect 674012 624650 674064 624656
rect 674012 624368 674064 624374
rect 674010 624336 674012 624345
rect 674064 624336 674066 624345
rect 674010 624271 674066 624280
rect 674010 623928 674066 623937
rect 674010 623863 674012 623872
rect 674064 623863 674066 623872
rect 674012 623834 674064 623840
rect 674012 623552 674064 623558
rect 674010 623520 674012 623529
rect 674064 623520 674066 623529
rect 674010 623455 674066 623464
rect 674010 623112 674066 623121
rect 674010 623047 674012 623056
rect 674064 623047 674066 623056
rect 674012 623018 674064 623024
rect 674012 622736 674064 622742
rect 674010 622704 674012 622713
rect 674064 622704 674066 622713
rect 674010 622639 674066 622648
rect 674010 622296 674066 622305
rect 674010 622231 674012 622240
rect 674064 622231 674066 622240
rect 674012 622202 674064 622208
rect 674012 621648 674064 621654
rect 674012 621590 674064 621596
rect 674024 621217 674052 621590
rect 674010 621208 674066 621217
rect 674010 621143 674066 621152
rect 674208 621014 674236 627886
rect 674392 623082 674420 636166
rect 674760 627914 674788 636942
rect 674944 635526 674972 637894
rect 675036 637650 675064 639882
rect 675036 637622 675156 637650
rect 674932 635520 674984 635526
rect 674932 635462 674984 635468
rect 674576 627886 674788 627914
rect 674380 623076 674432 623082
rect 674380 623018 674432 623024
rect 674576 621014 674604 627886
rect 674746 625968 674802 625977
rect 674746 625903 674802 625912
rect 674760 625734 674788 625903
rect 674748 625728 674800 625734
rect 674748 625670 674800 625676
rect 673932 620986 674236 621014
rect 674484 620986 674604 621014
rect 673932 601694 673960 620986
rect 674286 619168 674342 619177
rect 674286 619103 674342 619112
rect 674300 617574 674328 619103
rect 674288 617568 674340 617574
rect 674288 617510 674340 617516
rect 674288 615528 674340 615534
rect 674286 615496 674288 615505
rect 674340 615496 674342 615505
rect 674286 615431 674342 615440
rect 674286 609104 674342 609113
rect 674286 609039 674342 609048
rect 674300 608394 674328 609039
rect 674288 608388 674340 608394
rect 674288 608330 674340 608336
rect 674288 603288 674340 603294
rect 674288 603230 674340 603236
rect 674300 601694 674328 603230
rect 673932 601666 674052 601694
rect 673826 600672 673882 600681
rect 673826 600607 673882 600616
rect 673828 600432 673880 600438
rect 673826 600400 673828 600409
rect 673880 600400 673882 600409
rect 673826 600335 673882 600344
rect 673734 599856 673790 599865
rect 673734 599791 673790 599800
rect 673550 598632 673606 598641
rect 673550 598567 673606 598576
rect 673564 550634 673592 598567
rect 673748 598210 673776 599791
rect 673656 598182 673776 598210
rect 673656 592034 673684 598182
rect 673656 592006 673776 592034
rect 673472 550606 673592 550634
rect 673472 539050 673500 550606
rect 673748 550497 673776 592006
rect 674024 586514 674052 601666
rect 674116 601666 674328 601694
rect 674484 601694 674512 620986
rect 675128 611354 675156 637622
rect 675220 630674 675248 640138
rect 675404 639826 675432 640152
rect 675312 639798 675432 639826
rect 675312 631394 675340 639798
rect 675496 638761 675524 638928
rect 675482 638752 675538 638761
rect 675482 638687 675538 638696
rect 679622 637528 679678 637537
rect 675484 637492 675536 637498
rect 679622 637463 679678 637472
rect 675484 637434 675536 637440
rect 675496 636886 675524 637434
rect 675484 636880 675536 636886
rect 675484 636822 675536 636828
rect 675668 635520 675720 635526
rect 675668 635462 675720 635468
rect 675680 631417 675708 635462
rect 675482 631408 675538 631417
rect 675312 631366 675482 631394
rect 675482 631343 675538 631352
rect 675666 631408 675722 631417
rect 675666 631343 675722 631352
rect 675220 630646 675340 630674
rect 675312 617137 675340 630646
rect 676496 625728 676548 625734
rect 676494 625696 676496 625705
rect 676548 625696 676550 625705
rect 676494 625631 676550 625640
rect 679636 622033 679664 637463
rect 683212 637084 683264 637090
rect 683212 637026 683264 637032
rect 679622 622024 679678 622033
rect 679622 621959 679678 621968
rect 683224 618769 683252 637026
rect 683396 636880 683448 636886
rect 683396 636822 683448 636828
rect 683408 634814 683436 636822
rect 683408 634786 683620 634814
rect 683396 623076 683448 623082
rect 683396 623018 683448 623024
rect 683210 618760 683266 618769
rect 683210 618695 683266 618704
rect 676220 617568 676272 617574
rect 676218 617536 676220 617545
rect 676272 617536 676274 617545
rect 676218 617471 676274 617480
rect 675298 617128 675354 617137
rect 675298 617063 675354 617072
rect 683408 616729 683436 623018
rect 683592 617137 683620 634786
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683578 617128 683634 617137
rect 683578 617063 683634 617072
rect 683394 616720 683450 616729
rect 683394 616655 683450 616664
rect 683120 615528 683172 615534
rect 683118 615496 683120 615505
rect 683172 615496 683174 615505
rect 683118 615431 683174 615440
rect 674852 611326 675156 611354
rect 675298 611416 675354 611425
rect 675298 611351 675354 611360
rect 674852 608410 674880 611326
rect 675312 608682 675340 611351
rect 675312 608654 675418 608682
rect 675022 608560 675078 608569
rect 675022 608495 675078 608504
rect 674760 608382 674880 608410
rect 675036 608410 675064 608495
rect 675036 608382 675156 608410
rect 674760 608138 674788 608382
rect 674930 608288 674986 608297
rect 674930 608223 674986 608232
rect 674760 608110 674880 608138
rect 674484 601666 674696 601694
rect 674116 592034 674144 601666
rect 674286 600672 674342 600681
rect 674286 600607 674342 600616
rect 674300 592686 674328 600607
rect 674472 599004 674524 599010
rect 674472 598946 674524 598952
rect 674288 592680 674340 592686
rect 674288 592622 674340 592628
rect 674484 592034 674512 598946
rect 674116 592006 674236 592034
rect 674208 591410 674236 592006
rect 673932 586486 674052 586514
rect 674116 591382 674236 591410
rect 674392 592006 674512 592034
rect 673932 574841 673960 586486
rect 673918 574832 673974 574841
rect 673918 574767 673974 574776
rect 673920 574592 673972 574598
rect 673918 574560 673920 574569
rect 673972 574560 673974 574569
rect 673918 574495 673974 574504
rect 673920 574320 673972 574326
rect 673920 574262 673972 574268
rect 673932 574161 673960 574262
rect 673918 574152 673974 574161
rect 673918 574087 673974 574096
rect 673920 573912 673972 573918
rect 673918 573880 673920 573889
rect 673972 573880 673974 573889
rect 673918 573815 673974 573824
rect 673918 572112 673974 572121
rect 673918 572047 673974 572056
rect 673932 571606 673960 572047
rect 673920 571600 673972 571606
rect 673920 571542 673972 571548
rect 673918 571432 673974 571441
rect 673918 571367 673920 571376
rect 673972 571367 673974 571376
rect 673920 571338 673972 571344
rect 673918 571160 673974 571169
rect 673918 571095 673920 571104
rect 673972 571095 673974 571104
rect 673920 571066 673972 571072
rect 673918 570888 673974 570897
rect 673918 570823 673974 570832
rect 673932 569974 673960 570823
rect 673920 569968 673972 569974
rect 673920 569910 673972 569916
rect 673918 569664 673974 569673
rect 673918 569599 673974 569608
rect 673932 568614 673960 569599
rect 673920 568608 673972 568614
rect 673920 568550 673972 568556
rect 673920 565888 673972 565894
rect 673918 565856 673920 565865
rect 673972 565856 673974 565865
rect 673918 565791 673974 565800
rect 673918 564496 673974 564505
rect 673918 564431 673920 564440
rect 673972 564431 673974 564440
rect 673920 564402 673972 564408
rect 673918 558376 673974 558385
rect 673918 558311 673974 558320
rect 673932 554933 673960 558311
rect 673840 554905 673960 554933
rect 673840 550634 673868 554905
rect 674116 554169 674144 591382
rect 674392 586514 674420 592006
rect 674668 588606 674696 601666
rect 674852 591530 674880 608110
rect 674944 606846 674972 608223
rect 675128 607493 675156 608382
rect 675484 608388 675536 608394
rect 675484 608330 675536 608336
rect 675496 608124 675524 608330
rect 675128 607465 675418 607493
rect 674944 606818 675418 606846
rect 674944 604982 675418 605010
rect 674944 593178 674972 604982
rect 675128 604438 675418 604466
rect 675128 604353 675156 604438
rect 675114 604344 675170 604353
rect 675114 604279 675170 604288
rect 675312 603894 675432 603922
rect 675312 603786 675340 603894
rect 675128 603758 675340 603786
rect 675404 603772 675432 603894
rect 675128 603294 675156 603758
rect 675116 603288 675168 603294
rect 675116 603230 675168 603236
rect 675128 603146 675418 603174
rect 675128 602993 675156 603146
rect 675114 602984 675170 602993
rect 675114 602919 675170 602928
rect 675390 600944 675446 600953
rect 675390 600879 675446 600888
rect 675404 600644 675432 600879
rect 675114 600400 675170 600409
rect 675114 600335 675170 600344
rect 675128 598278 675156 600335
rect 675496 599865 675524 600100
rect 675482 599856 675538 599865
rect 675482 599791 675538 599800
rect 675312 599474 675418 599502
rect 675312 599010 675340 599474
rect 675300 599004 675352 599010
rect 675300 598946 675352 598952
rect 675496 598641 675524 598808
rect 675482 598632 675538 598641
rect 675482 598567 675538 598576
rect 675128 598250 675418 598278
rect 675114 598088 675170 598097
rect 675114 598023 675170 598032
rect 675128 596442 675156 598023
rect 675404 597417 675432 597652
rect 675390 597408 675446 597417
rect 675390 597343 675446 597352
rect 675128 596414 675418 596442
rect 675404 595377 675432 595816
rect 675390 595368 675446 595377
rect 675390 595303 675446 595312
rect 675496 594833 675524 595136
rect 675482 594824 675538 594833
rect 675482 594759 675538 594768
rect 675404 593473 675432 593980
rect 675390 593464 675446 593473
rect 675390 593399 675446 593408
rect 675482 593192 675538 593201
rect 674944 593150 675248 593178
rect 675022 591560 675078 591569
rect 674840 591524 674892 591530
rect 675022 591495 675078 591504
rect 674840 591466 674892 591472
rect 674656 588600 674708 588606
rect 674656 588542 674708 588548
rect 674208 586486 674420 586514
rect 674208 560294 674236 586486
rect 674380 579760 674432 579766
rect 674378 579728 674380 579737
rect 674432 579728 674434 579737
rect 674378 579663 674434 579672
rect 674472 578468 674524 578474
rect 674472 578410 674524 578416
rect 674484 578241 674512 578410
rect 674470 578232 674526 578241
rect 674470 578167 674526 578176
rect 674380 577584 674432 577590
rect 674378 577552 674380 577561
rect 674432 577552 674434 577561
rect 674378 577487 674434 577496
rect 674562 574832 674618 574841
rect 674562 574767 674618 574776
rect 674380 574116 674432 574122
rect 674380 574058 674432 574064
rect 674392 573889 674420 574058
rect 674378 573880 674434 573889
rect 674378 573815 674434 573824
rect 674576 571606 674604 574767
rect 674564 571600 674616 571606
rect 674564 571542 674616 571548
rect 674380 571464 674432 571470
rect 674378 571432 674380 571441
rect 674432 571432 674434 571441
rect 674378 571367 674434 571376
rect 674838 571160 674894 571169
rect 674838 571095 674894 571104
rect 674852 570518 674880 571095
rect 674840 570512 674892 570518
rect 674840 570454 674892 570460
rect 675036 567194 675064 591495
rect 675220 586265 675248 593150
rect 675482 593127 675538 593136
rect 675206 586256 675262 586265
rect 675206 586191 675262 586200
rect 675496 570518 675524 593127
rect 683396 592680 683448 592686
rect 683396 592622 683448 592628
rect 679624 591524 679676 591530
rect 679624 591466 679676 591472
rect 676218 580544 676274 580553
rect 676218 580479 676274 580488
rect 676232 579766 676260 580479
rect 676220 579760 676272 579766
rect 676220 579702 676272 579708
rect 676218 579320 676274 579329
rect 676218 579255 676274 579264
rect 676232 578474 676260 579255
rect 676220 578468 676272 578474
rect 676220 578410 676272 578416
rect 676218 578096 676274 578105
rect 676218 578031 676274 578040
rect 676232 577590 676260 578031
rect 676220 577584 676272 577590
rect 676220 577526 676272 577532
rect 679636 576473 679664 591466
rect 682382 591424 682438 591433
rect 682382 591359 682438 591368
rect 679622 576464 679678 576473
rect 679622 576399 679678 576408
rect 682396 575657 682424 591359
rect 682382 575648 682438 575657
rect 682382 575583 682438 575592
rect 676218 574832 676274 574841
rect 676218 574767 676274 574776
rect 676232 574122 676260 574767
rect 676220 574116 676272 574122
rect 676220 574058 676272 574064
rect 683408 573209 683436 592622
rect 684222 591152 684278 591161
rect 684222 591087 684278 591096
rect 684040 588600 684092 588606
rect 684040 588542 684092 588548
rect 683394 573200 683450 573209
rect 683394 573135 683450 573144
rect 676218 572384 676274 572393
rect 676218 572319 676274 572328
rect 676036 571600 676088 571606
rect 676036 571542 676088 571548
rect 676048 571305 676076 571542
rect 676232 571470 676260 572319
rect 684052 571985 684080 588542
rect 684236 576065 684264 591087
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 684222 576056 684278 576065
rect 684222 575991 684278 576000
rect 684038 571976 684094 571985
rect 684038 571911 684094 571920
rect 676220 571464 676272 571470
rect 676220 571406 676272 571412
rect 676034 571296 676090 571305
rect 676034 571231 676090 571240
rect 675484 570512 675536 570518
rect 675484 570454 675536 570460
rect 683120 570512 683172 570518
rect 683120 570454 683172 570460
rect 683132 570353 683160 570454
rect 683118 570344 683174 570353
rect 683118 570279 683174 570288
rect 674944 567166 675064 567194
rect 674944 563054 674972 567166
rect 675390 565856 675446 565865
rect 675390 565791 675446 565800
rect 675114 564496 675170 564505
rect 675114 564431 675170 564440
rect 674852 563026 674972 563054
rect 674852 560294 674880 563026
rect 675128 562918 675156 564431
rect 675404 563448 675432 565791
rect 675312 562958 675432 562986
rect 675312 562918 675340 562958
rect 675128 562890 675340 562918
rect 675404 562904 675432 562958
rect 675114 562320 675170 562329
rect 675170 562278 675418 562306
rect 675114 562255 675170 562264
rect 675390 561912 675446 561921
rect 675390 561847 675446 561856
rect 675404 561612 675432 561847
rect 674208 560266 674420 560294
rect 674392 558914 674420 560266
rect 674300 558886 674420 558914
rect 674484 560266 674880 560294
rect 674102 554160 674158 554169
rect 674102 554095 674158 554104
rect 674300 553466 674328 558886
rect 674116 553438 674328 553466
rect 674116 553024 674144 553438
rect 674024 552996 674144 553024
rect 674024 550746 674052 552996
rect 674484 552974 674512 560266
rect 675312 559830 675432 559858
rect 675312 559790 675340 559830
rect 674944 559762 675340 559790
rect 675404 559776 675432 559830
rect 674656 553512 674708 553518
rect 674656 553454 674708 553460
rect 674472 552968 674524 552974
rect 674286 552936 674342 552945
rect 674472 552910 674524 552916
rect 674286 552871 674342 552880
rect 674024 550718 674144 550746
rect 673840 550606 674052 550634
rect 673734 550488 673790 550497
rect 673734 550423 673790 550432
rect 674024 548026 674052 550606
rect 674116 549254 674144 550718
rect 674116 549226 674236 549254
rect 674208 548570 674236 549226
rect 673932 547998 674052 548026
rect 674116 548542 674236 548570
rect 673472 539022 673776 539050
rect 673552 536172 673604 536178
rect 673552 536114 673604 536120
rect 673564 531314 673592 536114
rect 673748 531314 673776 539022
rect 673932 536178 673960 547998
rect 674116 537169 674144 548542
rect 674300 547398 674328 552871
rect 674472 552084 674524 552090
rect 674472 552026 674524 552032
rect 674288 547392 674340 547398
rect 674288 547334 674340 547340
rect 674102 537160 674158 537169
rect 674102 537095 674158 537104
rect 673920 536172 673972 536178
rect 673920 536114 673972 536120
rect 674012 535968 674064 535974
rect 674064 535916 674328 535922
rect 674012 535910 674328 535916
rect 674024 535906 674328 535910
rect 674024 535900 674340 535906
rect 674024 535894 674288 535900
rect 674288 535842 674340 535848
rect 674288 535696 674340 535702
rect 674024 535644 674288 535650
rect 674024 535638 674340 535644
rect 674024 535622 674328 535638
rect 674024 535498 674052 535622
rect 674012 535492 674064 535498
rect 674012 535434 674064 535440
rect 674012 535016 674064 535022
rect 674064 534964 674328 534970
rect 674012 534958 674328 534964
rect 674024 534954 674328 534958
rect 674024 534948 674340 534954
rect 674024 534942 674288 534948
rect 674288 534890 674340 534896
rect 674012 534744 674064 534750
rect 674064 534692 674328 534698
rect 674012 534686 674328 534692
rect 674024 534682 674328 534686
rect 674024 534676 674340 534682
rect 674024 534670 674288 534676
rect 674288 534618 674340 534624
rect 674288 534540 674340 534546
rect 674024 534488 674288 534494
rect 674024 534482 674340 534488
rect 674024 534466 674328 534482
rect 674024 534138 674052 534466
rect 674484 534154 674512 552026
rect 674012 534132 674064 534138
rect 674012 534074 674064 534080
rect 674392 534126 674512 534154
rect 674392 533882 674420 534126
rect 674392 533854 674512 533882
rect 674012 533316 674064 533322
rect 674064 533264 674328 533270
rect 674012 533258 674328 533264
rect 674024 533254 674328 533258
rect 674024 533248 674340 533254
rect 674024 533242 674288 533248
rect 674288 533190 674340 533196
rect 674288 532840 674340 532846
rect 674024 532788 674288 532794
rect 674024 532782 674340 532788
rect 674024 532778 674328 532782
rect 674012 532772 674328 532778
rect 674064 532766 674328 532772
rect 674012 532714 674064 532720
rect 674012 532568 674064 532574
rect 674064 532516 674328 532522
rect 674012 532510 674328 532516
rect 674024 532506 674328 532510
rect 674024 532500 674340 532506
rect 674024 532494 674288 532500
rect 674288 532442 674340 532448
rect 674024 532030 674328 532046
rect 674012 532024 674340 532030
rect 674064 532018 674288 532024
rect 674012 531966 674064 531972
rect 674288 531966 674340 531972
rect 674012 531888 674064 531894
rect 674064 531836 674328 531842
rect 674012 531830 674328 531836
rect 674024 531826 674328 531830
rect 674024 531820 674340 531826
rect 674024 531814 674288 531820
rect 674288 531762 674340 531768
rect 673472 531286 673592 531314
rect 673656 531286 673776 531314
rect 673472 518894 673500 531286
rect 673656 526425 673684 531286
rect 674012 530936 674064 530942
rect 674064 530884 674328 530890
rect 674012 530878 674328 530884
rect 674024 530874 674328 530878
rect 674024 530868 674340 530874
rect 674024 530862 674288 530868
rect 674288 530810 674340 530816
rect 674012 529984 674064 529990
rect 674288 529984 674340 529990
rect 674064 529932 674288 529938
rect 674012 529926 674340 529932
rect 674024 529910 674328 529926
rect 674012 529440 674064 529446
rect 674064 529388 674328 529394
rect 674012 529382 674328 529388
rect 674024 529378 674328 529382
rect 674024 529372 674340 529378
rect 674024 529366 674288 529372
rect 674288 529314 674340 529320
rect 674288 529236 674340 529242
rect 674024 529184 674288 529190
rect 674024 529178 674340 529184
rect 674024 529174 674328 529178
rect 674012 529168 674328 529174
rect 674064 529162 674328 529168
rect 674012 529110 674064 529116
rect 674012 528896 674064 528902
rect 674064 528844 674328 528850
rect 674012 528838 674328 528844
rect 674024 528834 674328 528838
rect 674024 528828 674340 528834
rect 674024 528822 674288 528828
rect 674288 528770 674340 528776
rect 674012 528080 674064 528086
rect 674064 528028 674328 528034
rect 674012 528022 674328 528028
rect 674024 528018 674328 528022
rect 674024 528012 674340 528018
rect 674024 528006 674288 528012
rect 674288 527954 674340 527960
rect 673642 526416 673698 526425
rect 673642 526351 673698 526360
rect 674024 524618 674328 524634
rect 674012 524612 674340 524618
rect 674064 524606 674288 524612
rect 674012 524554 674064 524560
rect 674288 524554 674340 524560
rect 673472 518866 673960 518894
rect 673932 499574 673960 518866
rect 673656 499546 673960 499574
rect 673656 484401 673684 499546
rect 673826 492144 673882 492153
rect 673826 492079 673882 492088
rect 673840 491502 673868 492079
rect 674288 491700 674340 491706
rect 674288 491642 674340 491648
rect 674012 491632 674064 491638
rect 674300 491586 674328 491642
rect 674064 491580 674328 491586
rect 674012 491574 674328 491580
rect 674024 491558 674328 491574
rect 673828 491496 673880 491502
rect 673828 491438 673880 491444
rect 674012 491360 674064 491366
rect 674010 491328 674012 491337
rect 674064 491328 674066 491337
rect 674010 491263 674066 491272
rect 674012 490952 674064 490958
rect 674010 490920 674012 490929
rect 674064 490920 674066 490929
rect 674010 490855 674066 490864
rect 674010 489696 674066 489705
rect 674010 489631 674012 489640
rect 674064 489631 674066 489640
rect 674012 489602 674064 489608
rect 674012 489320 674064 489326
rect 674010 489288 674012 489297
rect 674064 489288 674066 489297
rect 674010 489223 674066 489232
rect 674012 488504 674064 488510
rect 674010 488472 674012 488481
rect 674064 488472 674066 488481
rect 674010 488407 674066 488416
rect 674012 486056 674064 486062
rect 674010 486024 674012 486033
rect 674064 486024 674066 486033
rect 674010 485959 674066 485968
rect 674288 485920 674340 485926
rect 674024 485868 674288 485874
rect 674024 485862 674340 485868
rect 674024 485858 674328 485862
rect 674012 485852 674328 485858
rect 674064 485846 674328 485852
rect 674012 485794 674064 485800
rect 674288 485172 674340 485178
rect 674288 485114 674340 485120
rect 674300 485058 674328 485114
rect 674024 485030 674328 485058
rect 674024 484430 674052 485030
rect 674012 484424 674064 484430
rect 673642 484392 673698 484401
rect 674012 484366 674064 484372
rect 673642 484327 673698 484336
rect 674484 484022 674512 533854
rect 674472 484016 674524 484022
rect 674472 483958 674524 483964
rect 674012 483200 674064 483206
rect 674010 483168 674012 483177
rect 674064 483168 674066 483177
rect 674010 483103 674066 483112
rect 674668 482390 674696 553454
rect 674944 553432 674972 559762
rect 675128 559218 675418 559246
rect 675128 559065 675156 559218
rect 675114 559056 675170 559065
rect 675114 558991 675170 559000
rect 675404 558385 675432 558620
rect 675390 558376 675446 558385
rect 675390 558311 675446 558320
rect 675128 557926 675418 557954
rect 675128 557569 675156 557926
rect 675114 557560 675170 557569
rect 675114 557495 675170 557504
rect 675404 555257 675432 555492
rect 675390 555248 675446 555257
rect 675390 555183 675446 555192
rect 675206 554840 675262 554849
rect 674760 553404 674972 553432
rect 675036 554798 675206 554826
rect 674760 548570 674788 553404
rect 675036 553093 675064 554798
rect 675206 554775 675262 554784
rect 675772 554713 675800 554919
rect 675758 554704 675814 554713
rect 675758 554639 675814 554648
rect 675772 553897 675800 554268
rect 675758 553888 675814 553897
rect 675758 553823 675814 553832
rect 675404 553602 675432 553656
rect 675312 553574 675432 553602
rect 675312 553518 675340 553574
rect 675300 553512 675352 553518
rect 675300 553454 675352 553460
rect 675036 553065 675418 553093
rect 674932 553036 674984 553042
rect 674932 552978 674984 552984
rect 674944 552922 674972 552978
rect 674852 552894 674972 552922
rect 674852 550634 674880 552894
rect 675128 552418 675418 552446
rect 675128 552090 675156 552418
rect 675298 552256 675354 552265
rect 675298 552191 675354 552200
rect 675116 552084 675168 552090
rect 675116 552026 675168 552032
rect 675312 551253 675340 552191
rect 675312 551225 675418 551253
rect 674852 550606 674972 550634
rect 674944 548894 674972 550606
rect 675128 550582 675418 550610
rect 674932 548888 674984 548894
rect 674932 548830 674984 548836
rect 675128 548774 675156 550582
rect 675496 549681 675524 549951
rect 675482 549672 675538 549681
rect 675482 549607 675538 549616
rect 675300 548888 675352 548894
rect 675300 548830 675352 548836
rect 675128 548746 675248 548774
rect 674760 548542 675064 548570
rect 674838 548448 674894 548457
rect 674838 548383 674894 548392
rect 674852 500954 674880 548383
rect 675036 546394 675064 548542
rect 675220 546650 675248 548746
rect 675312 548026 675340 548830
rect 675772 548321 675800 548760
rect 675758 548312 675814 548321
rect 675758 548247 675814 548256
rect 675312 547998 675432 548026
rect 675208 546644 675260 546650
rect 675208 546586 675260 546592
rect 675404 546514 675432 547998
rect 675574 547904 675630 547913
rect 675574 547839 675630 547848
rect 675588 547194 675616 547839
rect 677414 547632 677470 547641
rect 677414 547567 677470 547576
rect 675576 547188 675628 547194
rect 675576 547130 675628 547136
rect 675576 546644 675628 546650
rect 675576 546586 675628 546592
rect 675392 546508 675444 546514
rect 675392 546450 675444 546456
rect 675036 546366 675340 546394
rect 675116 541000 675168 541006
rect 675116 540942 675168 540948
rect 675128 503674 675156 540942
rect 675116 503668 675168 503674
rect 675116 503610 675168 503616
rect 675312 503538 675340 546366
rect 675588 541006 675616 546586
rect 675576 541000 675628 541006
rect 675576 540942 675628 540948
rect 675482 537160 675538 537169
rect 675482 537095 675538 537104
rect 675496 533390 675524 537095
rect 676218 535936 676274 535945
rect 676036 535900 676088 535906
rect 676218 535871 676274 535880
rect 676036 535842 676088 535848
rect 676048 535741 676076 535842
rect 676034 535732 676090 535741
rect 676232 535702 676260 535871
rect 676034 535667 676090 535676
rect 676220 535696 676272 535702
rect 676220 535638 676272 535644
rect 676218 535120 676274 535129
rect 676218 535055 676274 535064
rect 676036 534948 676088 534954
rect 676034 534916 676036 534925
rect 676088 534916 676090 534925
rect 676034 534851 676090 534860
rect 676232 534546 676260 535055
rect 676496 534676 676548 534682
rect 676496 534618 676548 534624
rect 676220 534540 676272 534546
rect 676220 534482 676272 534488
rect 676508 534313 676536 534618
rect 676494 534304 676550 534313
rect 676494 534239 676550 534248
rect 675484 533384 675536 533390
rect 675484 533326 675536 533332
rect 676034 533284 676090 533293
rect 676034 533219 676036 533228
rect 676088 533219 676090 533228
rect 676036 533190 676088 533196
rect 676034 532876 676090 532885
rect 676034 532811 676036 532820
rect 676088 532811 676090 532820
rect 676036 532782 676088 532788
rect 676036 532500 676088 532506
rect 676034 532468 676036 532477
rect 676088 532468 676090 532477
rect 676034 532403 676090 532412
rect 676034 532060 676090 532069
rect 676034 531995 676036 532004
rect 676088 531995 676090 532004
rect 676036 531966 676088 531972
rect 676218 531856 676274 531865
rect 676218 531791 676220 531800
rect 676272 531791 676274 531800
rect 676220 531762 676272 531768
rect 676036 530868 676088 530874
rect 676034 530836 676036 530845
rect 676088 530836 676090 530845
rect 676034 530771 676090 530780
rect 676034 530020 676090 530029
rect 676034 529955 676036 529964
rect 676088 529955 676090 529964
rect 676036 529926 676088 529932
rect 676218 529408 676274 529417
rect 676036 529372 676088 529378
rect 676218 529343 676274 529352
rect 676036 529314 676088 529320
rect 676048 529213 676076 529314
rect 676232 529242 676260 529343
rect 676220 529236 676272 529242
rect 676034 529204 676090 529213
rect 676220 529178 676272 529184
rect 676034 529139 676090 529148
rect 676036 528828 676088 528834
rect 676034 528796 676036 528805
rect 676088 528796 676090 528805
rect 676034 528731 676090 528740
rect 676036 528012 676088 528018
rect 676034 527980 676036 527989
rect 676088 527980 676090 527989
rect 676034 527915 676090 527924
rect 675484 520260 675536 520266
rect 675484 520202 675536 520208
rect 675300 503532 675352 503538
rect 675300 503474 675352 503480
rect 674840 500948 674892 500954
rect 674840 500890 674892 500896
rect 674656 482384 674708 482390
rect 674656 482326 674708 482332
rect 674024 480418 674328 480434
rect 674012 480412 674340 480418
rect 674064 480406 674288 480412
rect 674012 480354 674064 480360
rect 674288 480354 674340 480360
rect 673368 455864 673420 455870
rect 673368 455806 673420 455812
rect 673274 455424 673330 455433
rect 673274 455359 673276 455368
rect 673328 455359 673330 455368
rect 673276 455330 673328 455336
rect 673386 455288 673442 455297
rect 673386 455223 673388 455232
rect 673440 455223 673442 455232
rect 673506 455252 673558 455258
rect 673388 455194 673440 455200
rect 673506 455194 673558 455200
rect 673274 455152 673330 455161
rect 673518 455138 673546 455194
rect 673330 455110 673546 455138
rect 673274 455087 673330 455096
rect 674288 454912 674340 454918
rect 672814 454880 672870 454889
rect 672814 454815 672870 454824
rect 674286 454880 674288 454889
rect 674340 454880 674342 454889
rect 674286 454815 674342 454824
rect 672828 454510 672856 454815
rect 675496 454646 675524 520202
rect 675668 518832 675720 518838
rect 675668 518774 675720 518780
rect 673046 454640 673098 454646
rect 673044 454608 673046 454617
rect 674288 454640 674340 454646
rect 673098 454608 673100 454617
rect 673044 454543 673100 454552
rect 674286 454608 674288 454617
rect 675484 454640 675536 454646
rect 674340 454608 674342 454617
rect 675484 454582 675536 454588
rect 674286 454543 674342 454552
rect 672816 454504 672868 454510
rect 672816 454446 672868 454452
rect 675680 454374 675708 518774
rect 676034 491736 676090 491745
rect 676034 491671 676036 491680
rect 676088 491671 676090 491680
rect 676036 491642 676088 491648
rect 676034 486840 676090 486849
rect 676034 486775 676090 486784
rect 676048 485926 676076 486775
rect 676036 485920 676088 485926
rect 676036 485862 676088 485868
rect 676034 485208 676090 485217
rect 676034 485143 676036 485152
rect 676088 485143 676090 485152
rect 676036 485114 676088 485120
rect 676036 484016 676088 484022
rect 676034 483984 676036 483993
rect 676088 483984 676090 483993
rect 676034 483919 676090 483928
rect 677428 483002 677456 547567
rect 683212 547392 683264 547398
rect 683212 547334 683264 547340
rect 682382 546816 682438 546825
rect 682382 546751 682438 546760
rect 681004 546508 681056 546514
rect 681004 546450 681056 546456
rect 681016 531457 681044 546450
rect 681002 531448 681058 531457
rect 681002 531383 681058 531392
rect 682396 530641 682424 546751
rect 682382 530632 682438 530641
rect 682382 530567 682438 530576
rect 683224 528601 683252 547334
rect 683396 547188 683448 547194
rect 683396 547130 683448 547136
rect 683210 528592 683266 528601
rect 683210 528527 683266 528536
rect 683408 526969 683436 547130
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683580 533384 683632 533390
rect 683580 533326 683632 533332
rect 683592 527785 683620 533326
rect 683578 527776 683634 527785
rect 683578 527711 683634 527720
rect 683394 526960 683450 526969
rect 683394 526895 683450 526904
rect 677874 525736 677930 525745
rect 677874 525671 677930 525680
rect 677888 518838 677916 525671
rect 683118 524920 683174 524929
rect 683118 524855 683174 524864
rect 683132 524618 683160 524855
rect 683120 524612 683172 524618
rect 683120 524554 683172 524560
rect 680358 524512 680414 524521
rect 680358 524447 680414 524456
rect 680372 520266 680400 524447
rect 680360 520260 680412 520266
rect 680360 520202 680412 520208
rect 677876 518832 677928 518838
rect 677876 518774 677928 518780
rect 683210 503704 683266 503713
rect 679624 503668 679676 503674
rect 683210 503639 683266 503648
rect 679624 503610 679676 503616
rect 679636 487257 679664 503610
rect 681004 503532 681056 503538
rect 681004 503474 681056 503480
rect 679622 487248 679678 487257
rect 679622 487183 679678 487192
rect 681016 486441 681044 503474
rect 681188 500948 681240 500954
rect 681188 500890 681240 500896
rect 681200 487665 681228 500890
rect 681186 487656 681242 487665
rect 681186 487591 681242 487600
rect 681002 486432 681058 486441
rect 681002 486367 681058 486376
rect 683224 485625 683252 503639
rect 683394 500984 683450 500993
rect 683394 500919 683450 500928
rect 683210 485616 683266 485625
rect 683210 485551 683266 485560
rect 683408 483585 683436 500919
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683394 483576 683450 483585
rect 683394 483511 683450 483520
rect 676220 482996 676272 483002
rect 676220 482938 676272 482944
rect 677416 482996 677468 483002
rect 677416 482938 677468 482944
rect 676034 482760 676090 482769
rect 676232 482746 676260 482938
rect 676090 482718 676260 482746
rect 676034 482695 676090 482704
rect 676036 482384 676088 482390
rect 676034 482352 676036 482361
rect 676088 482352 676090 482361
rect 676034 482287 676090 482296
rect 680358 481944 680414 481953
rect 680358 481879 680414 481888
rect 675850 480720 675906 480729
rect 675850 480655 675906 480664
rect 675864 454918 675892 480655
rect 680372 475182 680400 481879
rect 683118 481128 683174 481137
rect 683118 481063 683174 481072
rect 683132 480418 683160 481063
rect 683120 480412 683172 480418
rect 683120 480354 683172 480360
rect 676036 475176 676088 475182
rect 676036 475118 676088 475124
rect 680360 475176 680412 475182
rect 680360 475118 680412 475124
rect 675852 454912 675904 454918
rect 675852 454854 675904 454860
rect 672954 454368 673006 454374
rect 672952 454336 672954 454345
rect 674288 454368 674340 454374
rect 673006 454336 673008 454345
rect 672952 454271 673008 454280
rect 674286 454336 674288 454345
rect 675668 454368 675720 454374
rect 674340 454336 674342 454345
rect 675668 454310 675720 454316
rect 674286 454271 674342 454280
rect 676048 453966 676076 475118
rect 674288 453960 674340 453966
rect 674286 453928 674288 453937
rect 676036 453960 676088 453966
rect 674340 453928 674342 453937
rect 676036 453902 676088 453908
rect 674286 453863 674342 453872
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 676218 403336 676274 403345
rect 674564 403300 674616 403306
rect 676218 403271 676220 403280
rect 674564 403242 674616 403248
rect 676272 403271 676274 403280
rect 676220 403242 676272 403248
rect 672630 402520 672686 402529
rect 672630 402455 672686 402464
rect 672446 401976 672502 401985
rect 672446 401911 672502 401920
rect 673182 401704 673238 401713
rect 673182 401639 673238 401648
rect 672814 399664 672870 399673
rect 672814 399599 672870 399608
rect 672630 393952 672686 393961
rect 672630 393887 672686 393896
rect 671894 393680 671950 393689
rect 671894 393615 671950 393624
rect 671710 348936 671766 348945
rect 671710 348871 671766 348880
rect 671724 329769 671752 348871
rect 671710 329760 671766 329769
rect 671710 329695 671766 329704
rect 671526 302288 671582 302297
rect 671526 302223 671582 302232
rect 671344 278724 671396 278730
rect 671344 278666 671396 278672
rect 670974 262168 671030 262177
rect 670974 262103 671030 262112
rect 670698 257272 670754 257281
rect 670698 257207 670754 257216
rect 670514 223952 670570 223961
rect 670514 223887 670570 223896
rect 670422 223680 670478 223689
rect 670422 223615 670424 223624
rect 670476 223615 670478 223624
rect 670424 223586 670476 223592
rect 670068 222822 670464 222850
rect 669884 222166 670280 222194
rect 669780 221400 669832 221406
rect 669780 221342 669832 221348
rect 669780 221128 669832 221134
rect 669700 221076 669780 221082
rect 669700 221070 669832 221076
rect 669700 221054 669820 221070
rect 669412 220924 669464 220930
rect 669412 220866 669464 220872
rect 669412 220788 669464 220794
rect 669412 220730 669464 220736
rect 669240 220646 669360 220674
rect 669056 220510 669268 220538
rect 668950 199200 669006 199209
rect 668950 199135 669006 199144
rect 669042 191720 669098 191729
rect 669042 191655 669098 191664
rect 668766 163296 668822 163305
rect 668766 163231 668822 163240
rect 668858 162344 668914 162353
rect 668858 162279 668914 162288
rect 668872 161474 668900 162279
rect 668872 161446 668992 161474
rect 668766 159080 668822 159089
rect 668766 159015 668822 159024
rect 668780 158409 668808 159015
rect 668766 158400 668822 158409
rect 668766 158335 668822 158344
rect 668964 151814 668992 161446
rect 668872 151786 668992 151814
rect 668872 148617 668900 151786
rect 668858 148608 668914 148617
rect 668858 148543 668914 148552
rect 668768 146056 668820 146062
rect 668768 145998 668820 146004
rect 668780 145353 668808 145998
rect 668766 145344 668822 145353
rect 668766 145279 668822 145288
rect 668582 138816 668638 138825
rect 668582 138751 668638 138760
rect 669056 135561 669084 191655
rect 669240 189417 669268 220510
rect 669332 219434 669360 220646
rect 669424 220538 669452 220730
rect 669424 220510 669544 220538
rect 669516 219434 669544 220510
rect 669700 219434 669728 221054
rect 670054 220824 670110 220833
rect 669872 220788 669924 220794
rect 670252 220794 670280 222166
rect 670054 220759 670110 220768
rect 670240 220788 670292 220794
rect 669872 220730 669924 220736
rect 669884 219434 669912 220730
rect 669332 219406 669452 219434
rect 669516 219406 669636 219434
rect 669700 219406 669820 219434
rect 669884 219406 670004 219434
rect 669424 217297 669452 219406
rect 669410 217288 669466 217297
rect 669410 217223 669466 217232
rect 669410 214840 669466 214849
rect 669410 214775 669466 214784
rect 669424 202881 669452 214775
rect 669410 202872 669466 202881
rect 669410 202807 669466 202816
rect 669226 189408 669282 189417
rect 669226 189343 669282 189352
rect 669228 184884 669280 184890
rect 669228 184826 669280 184832
rect 669042 135552 669098 135561
rect 669042 135487 669098 135496
rect 667202 134600 667258 134609
rect 667202 134535 667258 134544
rect 667940 133816 667992 133822
rect 667938 133784 667940 133793
rect 667992 133784 667994 133793
rect 667938 133719 667994 133728
rect 667018 132696 667074 132705
rect 667018 132631 667074 132640
rect 668858 131200 668914 131209
rect 668858 131135 668914 131144
rect 668676 130688 668728 130694
rect 668674 130656 668676 130665
rect 668728 130656 668730 130665
rect 668674 130591 668730 130600
rect 667940 129600 667992 129606
rect 667940 129542 667992 129548
rect 667952 129033 667980 129542
rect 667938 129024 667994 129033
rect 667938 128959 667994 128968
rect 668582 127800 668638 127809
rect 668582 127735 668638 127744
rect 668398 126984 668454 126993
rect 668398 126919 668454 126928
rect 668412 120873 668440 126919
rect 668398 120864 668454 120873
rect 668398 120799 668454 120808
rect 668124 112940 668176 112946
rect 668124 112882 668176 112888
rect 668136 112713 668164 112882
rect 668122 112704 668178 112713
rect 668122 112639 668178 112648
rect 668400 108044 668452 108050
rect 668400 107986 668452 107992
rect 668412 107817 668440 107986
rect 668398 107808 668454 107817
rect 668398 107743 668454 107752
rect 667940 104576 667992 104582
rect 667938 104544 667940 104553
rect 667992 104544 667994 104553
rect 667938 104479 667994 104488
rect 668596 102921 668624 127735
rect 668872 122834 668900 131135
rect 669240 125769 669268 184826
rect 669608 174758 669636 219406
rect 669596 174752 669648 174758
rect 669596 174694 669648 174700
rect 669594 171184 669650 171193
rect 669594 171119 669650 171128
rect 669608 154465 669636 171119
rect 669792 169726 669820 219406
rect 669780 169720 669832 169726
rect 669780 169662 669832 169668
rect 669778 169552 669834 169561
rect 669778 169487 669834 169496
rect 669594 154456 669650 154465
rect 669594 154391 669650 154400
rect 669792 150385 669820 169487
rect 669778 150376 669834 150385
rect 669778 150311 669834 150320
rect 669976 133822 670004 219406
rect 670068 216186 670096 220759
rect 670240 220730 670292 220736
rect 670436 220674 670464 222822
rect 670160 220646 670464 220674
rect 670160 216458 670188 220646
rect 670330 220416 670386 220425
rect 670330 220351 670386 220360
rect 670344 218113 670372 220351
rect 670330 218104 670386 218113
rect 670330 218039 670386 218048
rect 670514 216608 670570 216617
rect 670514 216543 670570 216552
rect 670330 216472 670386 216481
rect 670160 216430 670330 216458
rect 670330 216407 670386 216416
rect 670068 216158 670372 216186
rect 670146 211168 670202 211177
rect 670146 211103 670202 211112
rect 669964 133816 670016 133822
rect 669964 133758 670016 133764
rect 670160 129606 670188 211103
rect 670344 164966 670372 216158
rect 670528 198257 670556 216543
rect 670514 198248 670570 198257
rect 670514 198183 670570 198192
rect 670712 184890 670740 257207
rect 670988 236201 671016 262103
rect 671252 236904 671304 236910
rect 671252 236846 671304 236852
rect 670974 236192 671030 236201
rect 670974 236127 671030 236136
rect 671068 235952 671120 235958
rect 671068 235894 671120 235900
rect 670882 234016 670938 234025
rect 670882 233951 670884 233960
rect 670936 233951 670938 233960
rect 670884 233922 670936 233928
rect 670884 233232 670936 233238
rect 670884 233174 670936 233180
rect 670896 186314 670924 233174
rect 670896 186286 671016 186314
rect 670700 184884 670752 184890
rect 670700 184826 670752 184832
rect 670792 178016 670844 178022
rect 670790 177984 670792 177993
rect 670844 177984 670846 177993
rect 670790 177919 670846 177928
rect 670988 176654 671016 186286
rect 670896 176626 671016 176654
rect 670606 170368 670662 170377
rect 670606 170303 670662 170312
rect 670332 164960 670384 164966
rect 670332 164902 670384 164908
rect 670620 147665 670648 170303
rect 670896 166994 670924 176626
rect 670804 166966 670924 166994
rect 670804 160070 670832 166966
rect 670792 160064 670844 160070
rect 670792 160006 670844 160012
rect 671080 157334 671108 235894
rect 671264 186314 671292 236846
rect 671372 233776 671424 233782
rect 671356 233724 671372 233730
rect 671356 233718 671424 233724
rect 671356 233702 671412 233718
rect 671356 220814 671384 233702
rect 671540 224369 671568 302223
rect 671710 278624 671766 278633
rect 671710 278559 671712 278568
rect 671764 278559 671766 278568
rect 671712 278530 671764 278536
rect 671710 260536 671766 260545
rect 671710 260471 671766 260480
rect 671724 240281 671752 260471
rect 671710 240272 671766 240281
rect 671710 240207 671766 240216
rect 671712 236496 671764 236502
rect 671712 236438 671764 236444
rect 671526 224360 671582 224369
rect 671526 224295 671582 224304
rect 671724 224210 671752 236438
rect 671908 231985 671936 393615
rect 672644 376281 672672 393887
rect 672630 376272 672686 376281
rect 672630 376207 672686 376216
rect 672538 356280 672594 356289
rect 672538 356215 672594 356224
rect 672354 355464 672410 355473
rect 672354 355399 672410 355408
rect 672170 353424 672226 353433
rect 672170 353359 672226 353368
rect 672184 338065 672212 353359
rect 672170 338056 672226 338065
rect 672170 337991 672226 338000
rect 672368 310865 672396 355399
rect 672552 311681 672580 356215
rect 672828 355065 672856 399599
rect 672998 395040 673054 395049
rect 672998 394975 673054 394984
rect 673012 381041 673040 394975
rect 672998 381032 673054 381041
rect 672998 380967 673054 380976
rect 673196 357513 673224 401639
rect 673918 401432 673974 401441
rect 673918 401367 673974 401376
rect 673366 400480 673422 400489
rect 673366 400415 673422 400424
rect 673182 357504 673238 357513
rect 673182 357439 673238 357448
rect 673182 357096 673238 357105
rect 673182 357031 673238 357040
rect 672814 355056 672870 355065
rect 672814 354991 672870 355000
rect 672998 349752 673054 349761
rect 672998 349687 673054 349696
rect 672722 348528 672778 348537
rect 672722 348463 672778 348472
rect 672538 311672 672594 311681
rect 672538 311607 672594 311616
rect 672354 310856 672410 310865
rect 672354 310791 672410 310800
rect 672172 288448 672224 288454
rect 672172 288390 672224 288396
rect 672184 246265 672212 288390
rect 672736 287054 672764 348463
rect 673012 335617 673040 349687
rect 672998 335608 673054 335617
rect 672998 335543 673054 335552
rect 672906 325000 672962 325009
rect 672906 324935 672962 324944
rect 672644 287026 672764 287054
rect 672356 284368 672408 284374
rect 672356 284310 672408 284316
rect 672368 277394 672396 284310
rect 672644 277394 672672 287026
rect 672920 278633 672948 324935
rect 673196 312497 673224 357031
rect 673380 355881 673408 400415
rect 673734 395720 673790 395729
rect 673734 395655 673790 395664
rect 673748 375465 673776 395655
rect 673734 375456 673790 375465
rect 673734 375391 673790 375400
rect 673932 356561 673960 401367
rect 674576 396681 674604 403242
rect 676586 402928 676642 402937
rect 676586 402863 676642 402872
rect 674838 402248 674894 402257
rect 674838 402183 674894 402192
rect 674852 401713 674880 402183
rect 674838 401704 674894 401713
rect 674838 401639 674894 401648
rect 676600 400897 676628 402863
rect 676586 400888 676642 400897
rect 676586 400823 676642 400832
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 676048 398886 676076 399327
rect 674932 398880 674984 398886
rect 674932 398822 674984 398828
rect 676036 398880 676088 398886
rect 676036 398822 676088 398828
rect 674746 397352 674802 397361
rect 674746 397287 674802 397296
rect 674562 396672 674618 396681
rect 674562 396607 674618 396616
rect 674564 396092 674616 396098
rect 674564 396034 674616 396040
rect 674380 394324 674432 394330
rect 674380 394266 674432 394272
rect 674392 393938 674420 394266
rect 674208 393910 674420 393938
rect 674208 380746 674236 393910
rect 674576 393314 674604 396034
rect 674760 393314 674788 397287
rect 674944 393314 674972 398822
rect 679622 398440 679678 398449
rect 679622 398375 679678 398384
rect 676218 398032 676274 398041
rect 676218 397967 676274 397976
rect 676034 396128 676090 396137
rect 676034 396063 676036 396072
rect 676088 396063 676090 396072
rect 676036 396034 676088 396040
rect 676232 395758 676260 397967
rect 678242 397624 678298 397633
rect 678242 397559 678298 397568
rect 675208 395752 675260 395758
rect 675208 395694 675260 395700
rect 676220 395752 676272 395758
rect 676220 395694 676272 395700
rect 674392 393286 674604 393314
rect 674668 393286 674788 393314
rect 674852 393286 674972 393314
rect 674392 382226 674420 393286
rect 674380 382220 674432 382226
rect 674380 382162 674432 382168
rect 674208 380718 674420 380746
rect 674392 378146 674420 380718
rect 674380 378140 674432 378146
rect 674380 378082 674432 378088
rect 674668 372570 674696 393286
rect 674852 384810 674880 393286
rect 675220 386458 675248 395694
rect 676218 394360 676274 394369
rect 676218 394295 676220 394304
rect 676272 394295 676274 394304
rect 676220 394266 676272 394272
rect 678256 387705 678284 397559
rect 678242 387696 678298 387705
rect 678242 387631 678298 387640
rect 679636 386782 679664 398375
rect 679624 386776 679676 386782
rect 679624 386718 679676 386724
rect 675036 386430 675248 386458
rect 674840 384804 674892 384810
rect 674840 384746 674892 384752
rect 675036 384690 675064 386430
rect 674944 384662 675064 384690
rect 675128 386261 675418 386289
rect 674944 382582 674972 384662
rect 675128 382945 675156 386261
rect 675484 386028 675536 386034
rect 675484 385970 675536 385976
rect 675496 385696 675524 385970
rect 675772 384985 675800 385084
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675392 384804 675444 384810
rect 675392 384746 675444 384752
rect 675404 384435 675432 384746
rect 675114 382936 675170 382945
rect 675114 382871 675170 382880
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 674944 382554 675340 382582
rect 675404 382568 675432 382622
rect 675758 382256 675814 382265
rect 675116 382220 675168 382226
rect 675758 382191 675814 382200
rect 675116 382162 675168 382168
rect 675128 381426 675156 382162
rect 675772 382024 675800 382191
rect 675128 381398 675418 381426
rect 675390 381032 675446 381041
rect 675390 380967 675446 380976
rect 675404 380732 675432 380967
rect 675666 378584 675722 378593
rect 675666 378519 675722 378528
rect 675680 378284 675708 378519
rect 675116 378140 675168 378146
rect 675116 378082 675168 378088
rect 675128 377754 675156 378082
rect 675128 377726 675340 377754
rect 675312 377618 675340 377726
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675758 377496 675814 377505
rect 675758 377431 675814 377440
rect 675772 377060 675800 377431
rect 675404 376281 675432 376448
rect 675390 376272 675446 376281
rect 675390 376207 675446 376216
rect 675114 375456 675170 375465
rect 675114 375391 675170 375400
rect 675128 375238 675156 375391
rect 675128 375210 675418 375238
rect 675758 373688 675814 373697
rect 675758 373623 675814 373632
rect 675772 373388 675800 373623
rect 675114 372872 675170 372881
rect 675114 372807 675170 372816
rect 675128 372722 675156 372807
rect 675404 372722 675432 372776
rect 675036 372694 675432 372722
rect 674656 372564 674708 372570
rect 674656 372506 674708 372512
rect 675036 371249 675064 372694
rect 675300 372564 675352 372570
rect 675300 372506 675352 372512
rect 675312 372042 675340 372506
rect 675312 372014 675432 372042
rect 675404 371552 675432 372014
rect 675022 371240 675078 371249
rect 675022 371175 675078 371184
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 674102 358320 674158 358329
rect 674102 358255 674158 358264
rect 673918 356552 673974 356561
rect 673918 356487 673974 356496
rect 673366 355872 673422 355881
rect 673366 355807 673422 355816
rect 673918 354648 673974 354657
rect 673918 354583 673974 354592
rect 673550 350568 673606 350577
rect 673550 350503 673606 350512
rect 673366 350160 673422 350169
rect 673366 350095 673422 350104
rect 673380 335889 673408 350095
rect 673366 335880 673422 335889
rect 673366 335815 673422 335824
rect 673564 331129 673592 350503
rect 673734 349344 673790 349353
rect 673734 349279 673790 349288
rect 673748 332761 673776 349279
rect 673734 332752 673790 332761
rect 673734 332687 673790 332696
rect 673550 331120 673606 331129
rect 673550 331055 673606 331064
rect 673932 325694 673960 354583
rect 674116 351121 674144 358255
rect 675942 357912 675998 357921
rect 675942 357847 675998 357856
rect 675956 356833 675984 357847
rect 675942 356824 675998 356833
rect 675942 356759 675998 356768
rect 674470 352608 674526 352617
rect 674470 352543 674526 352552
rect 674286 351384 674342 351393
rect 674286 351319 674342 351328
rect 674102 351112 674158 351121
rect 674102 351047 674158 351056
rect 674300 337793 674328 351319
rect 674286 337784 674342 337793
rect 674286 337719 674342 337728
rect 674484 333946 674512 352543
rect 674654 352200 674710 352209
rect 674654 352135 674710 352144
rect 674472 333940 674524 333946
rect 674472 333882 674524 333888
rect 674668 326913 674696 352135
rect 676034 350976 676090 350985
rect 676034 350911 676090 350920
rect 676048 346633 676076 350911
rect 676034 346624 676090 346633
rect 676034 346559 676090 346568
rect 674944 341074 675418 341102
rect 674944 338745 674972 341074
rect 675128 340530 675340 340558
rect 674930 338736 674986 338745
rect 674930 338671 674986 338680
rect 675128 338065 675156 340530
rect 675312 340490 675340 340530
rect 675404 340490 675432 340544
rect 675312 340462 675432 340490
rect 675758 340232 675814 340241
rect 675758 340167 675814 340176
rect 675772 339864 675800 340167
rect 675482 339416 675538 339425
rect 675482 339351 675538 339360
rect 675496 339252 675524 339351
rect 675114 338056 675170 338065
rect 675114 337991 675170 338000
rect 675758 337920 675814 337929
rect 675758 337855 675814 337864
rect 675114 337784 675170 337793
rect 675114 337719 675170 337728
rect 675128 336857 675156 337719
rect 675772 337416 675800 337855
rect 675128 336829 675418 336857
rect 675758 336560 675814 336569
rect 675758 336495 675814 336504
rect 675772 336192 675800 336495
rect 674930 335880 674986 335889
rect 674930 335815 674986 335824
rect 674944 331889 674972 335815
rect 675114 335608 675170 335617
rect 675170 335566 675340 335594
rect 675114 335543 675170 335552
rect 675312 335458 675340 335566
rect 675404 335458 675432 335580
rect 675312 335430 675432 335458
rect 675116 333940 675168 333946
rect 675116 333882 675168 333888
rect 675128 333078 675156 333882
rect 675128 333050 675418 333078
rect 675114 332752 675170 332761
rect 675114 332687 675170 332696
rect 675128 332534 675156 332687
rect 675128 332506 675418 332534
rect 674944 331861 675418 331889
rect 675128 331214 675418 331242
rect 675128 329769 675156 331214
rect 675298 331120 675354 331129
rect 675298 331055 675354 331064
rect 675312 330049 675340 331055
rect 675312 330021 675418 330049
rect 675114 329760 675170 329769
rect 675114 329695 675170 329704
rect 675312 328222 675432 328250
rect 675312 328182 675340 328222
rect 675220 328154 675340 328182
rect 675404 328168 675432 328222
rect 675022 327992 675078 328001
rect 675022 327927 675078 327936
rect 674654 326904 674710 326913
rect 674654 326839 674710 326848
rect 673932 325666 674420 325694
rect 673366 312760 673422 312769
rect 673366 312695 673422 312704
rect 673182 312488 673238 312497
rect 673182 312423 673238 312432
rect 673182 311264 673238 311273
rect 673182 311199 673238 311208
rect 673196 305402 673224 311199
rect 673196 305374 673316 305402
rect 673090 304328 673146 304337
rect 673090 304263 673146 304272
rect 673104 287881 673132 304263
rect 673288 304178 673316 305374
rect 673196 304150 673316 304178
rect 673196 302234 673224 304150
rect 673196 302206 673316 302234
rect 673090 287872 673146 287881
rect 673090 287807 673146 287816
rect 672906 278624 672962 278633
rect 672906 278559 672962 278568
rect 673288 277394 673316 302206
rect 672368 277366 672580 277394
rect 672644 277366 672764 277394
rect 672354 265432 672410 265441
rect 672354 265367 672410 265376
rect 672368 263594 672396 265367
rect 672552 263594 672580 277366
rect 672736 263594 672764 277366
rect 673196 277366 673316 277394
rect 673196 266665 673224 277366
rect 673380 267481 673408 312695
rect 674194 310448 674250 310457
rect 674194 310383 674250 310392
rect 673918 305144 673974 305153
rect 673918 305079 673974 305088
rect 673734 303920 673790 303929
rect 673734 303855 673790 303864
rect 673748 292574 673776 303855
rect 673564 292546 673776 292574
rect 673564 286521 673592 292546
rect 673734 290456 673790 290465
rect 673734 290391 673790 290400
rect 673550 286512 673606 286521
rect 673550 286447 673606 286456
rect 673748 267889 673776 290391
rect 673932 286929 673960 305079
rect 673918 286920 673974 286929
rect 673918 286855 673974 286864
rect 673918 283520 673974 283529
rect 673918 283455 673974 283464
rect 673932 268297 673960 283455
rect 674208 277394 674236 310383
rect 674392 310049 674420 325666
rect 675036 325009 675064 327927
rect 675220 325689 675248 328154
rect 675390 327992 675446 328001
rect 675390 327927 675446 327936
rect 675404 327556 675432 327927
rect 675390 326904 675446 326913
rect 675390 326839 675446 326848
rect 675404 326332 675432 326839
rect 675206 325680 675262 325689
rect 675206 325615 675262 325624
rect 675022 325000 675078 325009
rect 675022 324935 675078 324944
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676218 313984 676274 313993
rect 676218 313919 676274 313928
rect 674654 313032 674710 313041
rect 674654 312967 674710 312976
rect 674668 311953 674696 312967
rect 674838 312760 674894 312769
rect 674838 312695 674894 312704
rect 674852 312089 674880 312695
rect 674838 312080 674894 312089
rect 674838 312015 674894 312024
rect 674654 311944 674710 311953
rect 674654 311879 674710 311888
rect 674378 310040 674434 310049
rect 674378 309975 674434 309984
rect 674654 309632 674710 309641
rect 674654 309567 674710 309576
rect 674470 305552 674526 305561
rect 674470 305487 674526 305496
rect 674484 285666 674512 305487
rect 674668 287054 674696 309567
rect 675850 309360 675906 309369
rect 676232 309346 676260 313919
rect 675906 309318 676260 309346
rect 675850 309295 675906 309304
rect 675850 309088 675906 309097
rect 675850 309023 675906 309032
rect 675022 308000 675078 308009
rect 675022 307935 675078 307944
rect 674838 306368 674894 306377
rect 674838 306303 674894 306312
rect 674852 295610 674880 306303
rect 675036 302234 675064 307935
rect 675390 307592 675446 307601
rect 675390 307527 675446 307536
rect 675206 302968 675262 302977
rect 675206 302903 675262 302912
rect 675036 302206 675156 302234
rect 675128 299474 675156 302206
rect 675036 299446 675156 299474
rect 675220 299474 675248 302903
rect 675404 299474 675432 307527
rect 675864 306649 675892 309023
rect 676034 308408 676090 308417
rect 676090 308366 676444 308394
rect 676034 308343 676090 308352
rect 676034 307184 676090 307193
rect 676090 307142 676260 307170
rect 676034 307119 676090 307128
rect 675850 306640 675906 306649
rect 675850 306575 675906 306584
rect 676232 306406 676260 307142
rect 676220 306400 676272 306406
rect 676220 306342 676272 306348
rect 676034 305960 676090 305969
rect 676090 305918 676260 305946
rect 676034 305895 676090 305904
rect 675852 304972 675904 304978
rect 675852 304914 675904 304920
rect 675864 302977 675892 304914
rect 676034 303512 676090 303521
rect 676034 303447 676090 303456
rect 675850 302968 675906 302977
rect 675850 302903 675906 302912
rect 676048 302025 676076 303447
rect 676034 302016 676090 302025
rect 676034 301951 676090 301960
rect 676232 301617 676260 305918
rect 676416 304978 676444 308366
rect 679622 306776 679678 306785
rect 679622 306711 679678 306720
rect 676864 306400 676916 306406
rect 676864 306342 676916 306348
rect 676404 304972 676456 304978
rect 676404 304914 676456 304920
rect 676218 301608 676274 301617
rect 676218 301543 676274 301552
rect 675220 299446 675340 299474
rect 675404 299446 675524 299474
rect 675036 296562 675064 299446
rect 675036 296534 675156 296562
rect 674852 295582 675064 295610
rect 674838 294536 674894 294545
rect 674838 294471 674894 294480
rect 674852 288062 674880 294471
rect 675036 291870 675064 295582
rect 675128 292414 675156 296534
rect 675312 295905 675340 299446
rect 675496 296721 675524 299446
rect 676876 297401 676904 306342
rect 676862 297392 676918 297401
rect 676862 297327 676918 297336
rect 679636 297090 679664 306711
rect 675852 297084 675904 297090
rect 675852 297026 675904 297032
rect 679624 297084 679676 297090
rect 679624 297026 679676 297032
rect 675482 296712 675538 296721
rect 675482 296647 675538 296656
rect 675864 296562 675892 297026
rect 675496 296534 675892 296562
rect 675496 296410 675524 296534
rect 675484 296404 675536 296410
rect 675484 296346 675536 296352
rect 675666 296304 675722 296313
rect 675666 296239 675722 296248
rect 675680 296072 675708 296239
rect 675298 295896 675354 295905
rect 675298 295831 675354 295840
rect 675666 295896 675722 295905
rect 675666 295831 675722 295840
rect 675680 295528 675708 295831
rect 675484 295248 675536 295254
rect 675484 295190 675536 295196
rect 675496 294879 675524 295190
rect 675758 294536 675814 294545
rect 675758 294471 675814 294480
rect 675772 294236 675800 294471
rect 675128 292386 675418 292414
rect 675036 291842 675418 291870
rect 675758 291544 675814 291553
rect 675758 291479 675814 291488
rect 675772 291176 675800 291479
rect 675758 291000 675814 291009
rect 675758 290935 675814 290944
rect 675772 290564 675800 290935
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 674852 288034 675340 288062
rect 675404 288048 675432 288102
rect 675114 287872 675170 287881
rect 675114 287807 675170 287816
rect 675128 287518 675156 287807
rect 675128 287490 675418 287518
rect 674668 287026 674788 287054
rect 674472 285660 674524 285666
rect 674472 285602 674524 285608
rect 674208 277366 674604 277394
rect 673918 268288 673974 268297
rect 673918 268223 673974 268232
rect 673734 267880 673790 267889
rect 673734 267815 673790 267824
rect 673366 267472 673422 267481
rect 673366 267407 673422 267416
rect 673918 267064 673974 267073
rect 673918 266999 673974 267008
rect 673182 266656 673238 266665
rect 673182 266591 673238 266600
rect 673550 264616 673606 264625
rect 673550 264551 673606 264560
rect 672368 263566 672488 263594
rect 672552 263566 672672 263594
rect 672736 263566 672856 263594
rect 672170 246256 672226 246265
rect 672170 246191 672226 246200
rect 672264 237040 672316 237046
rect 672262 237008 672264 237017
rect 672316 237008 672318 237017
rect 672262 236943 672318 236952
rect 672080 235748 672132 235754
rect 672080 235690 672132 235696
rect 672092 233238 672120 235690
rect 672264 233300 672316 233306
rect 672264 233242 672316 233248
rect 672080 233232 672132 233238
rect 672080 233174 672132 233180
rect 671894 231976 671950 231985
rect 671894 231911 671950 231920
rect 672080 230648 672132 230654
rect 672080 230590 672132 230596
rect 672092 229770 672120 230590
rect 672080 229764 672132 229770
rect 672080 229706 672132 229712
rect 672276 225978 672304 233242
rect 672460 226930 672488 263566
rect 672644 227089 672672 263566
rect 672630 227080 672686 227089
rect 672828 227050 672856 263566
rect 673182 263392 673238 263401
rect 673182 263327 673238 263336
rect 672998 259720 673054 259729
rect 672998 259655 673054 259664
rect 673012 253934 673040 259655
rect 673196 259026 673224 263327
rect 672920 253906 673040 253934
rect 673104 258998 673224 259026
rect 672920 246213 672948 253906
rect 673104 250753 673132 258998
rect 673274 258904 673330 258913
rect 673274 258839 673330 258848
rect 673090 250744 673146 250753
rect 673090 250679 673146 250688
rect 673090 250064 673146 250073
rect 673090 249999 673146 250008
rect 673104 246213 673132 249999
rect 672920 246185 673040 246213
rect 673104 246185 673224 246213
rect 673012 245721 673040 246185
rect 672998 245712 673054 245721
rect 672998 245647 673054 245656
rect 672998 245440 673054 245449
rect 673196 245426 673224 246185
rect 673054 245398 673224 245426
rect 672998 245375 673054 245384
rect 673288 241505 673316 258839
rect 673564 241777 673592 264551
rect 673734 260944 673790 260953
rect 673734 260879 673790 260888
rect 673748 246673 673776 260879
rect 673734 246664 673790 246673
rect 673734 246599 673790 246608
rect 673550 241768 673606 241777
rect 673550 241703 673606 241712
rect 673274 241496 673330 241505
rect 673274 241431 673330 241440
rect 673734 237008 673790 237017
rect 673734 236943 673790 236952
rect 672954 236700 673006 236706
rect 672954 236642 673006 236648
rect 672966 236473 672994 236642
rect 673748 236586 673776 236943
rect 673748 236558 673868 236586
rect 673184 236496 673236 236502
rect 672952 236464 673008 236473
rect 673236 236444 673776 236450
rect 673184 236438 673776 236444
rect 673196 236422 673776 236438
rect 672952 236399 673008 236408
rect 673414 235884 673466 235890
rect 673414 235826 673466 235832
rect 673426 235770 673454 235826
rect 673426 235742 673684 235770
rect 673184 235544 673236 235550
rect 673184 235486 673236 235492
rect 673000 235068 673052 235074
rect 673000 235010 673052 235016
rect 673012 233102 673040 235010
rect 673196 233306 673224 235486
rect 673460 234864 673512 234870
rect 673460 234806 673512 234812
rect 673184 233300 673236 233306
rect 673184 233242 673236 233248
rect 673472 233238 673500 234806
rect 673460 233232 673512 233238
rect 673460 233174 673512 233180
rect 673000 233096 673052 233102
rect 673656 233050 673684 235742
rect 673000 233038 673052 233044
rect 673564 233022 673684 233050
rect 673564 232529 673592 233022
rect 673550 232520 673606 232529
rect 673550 232455 673606 232464
rect 673276 230444 673328 230450
rect 673276 230386 673328 230392
rect 673288 230217 673316 230386
rect 673460 230240 673512 230246
rect 673274 230208 673330 230217
rect 673460 230182 673512 230188
rect 673274 230143 673330 230152
rect 673472 229809 673500 230182
rect 673458 229800 673514 229809
rect 673458 229735 673514 229744
rect 673368 229628 673420 229634
rect 673368 229570 673420 229576
rect 672630 227015 672686 227024
rect 672816 227044 672868 227050
rect 672816 226986 672868 226992
rect 672460 226902 672948 226930
rect 672724 226432 672776 226438
rect 672722 226400 672724 226409
rect 672776 226400 672778 226409
rect 672722 226335 672778 226344
rect 672604 226160 672656 226166
rect 672602 226128 672604 226137
rect 672656 226128 672658 226137
rect 672602 226063 672658 226072
rect 672092 225950 672304 225978
rect 672494 225956 672546 225962
rect 672092 225570 672120 225950
rect 672494 225898 672546 225904
rect 672262 225856 672318 225865
rect 672262 225791 672318 225800
rect 672276 225690 672304 225791
rect 672380 225752 672432 225758
rect 672378 225720 672380 225729
rect 672432 225720 672434 225729
rect 672264 225684 672316 225690
rect 672378 225655 672434 225664
rect 672264 225626 672316 225632
rect 672506 225570 672534 225898
rect 672092 225542 672304 225570
rect 672154 225448 672210 225457
rect 672154 225383 672156 225392
rect 672208 225383 672210 225392
rect 672156 225354 672208 225360
rect 672032 225312 672088 225321
rect 672032 225247 672034 225256
rect 672086 225247 672088 225256
rect 672034 225218 672086 225224
rect 671818 224768 671874 224777
rect 671818 224703 671820 224712
rect 671872 224703 671874 224712
rect 671820 224674 671872 224680
rect 671724 224182 671936 224210
rect 671482 224120 671534 224126
rect 671482 224062 671534 224068
rect 671494 223961 671522 224062
rect 671908 223972 671936 224182
rect 671480 223952 671536 223961
rect 671480 223887 671536 223896
rect 671724 223944 671936 223972
rect 672078 223952 672134 223961
rect 671526 223680 671582 223689
rect 671526 223615 671582 223624
rect 671356 220786 671476 220814
rect 671448 190454 671476 220786
rect 671172 186286 671292 186314
rect 671356 190426 671476 190454
rect 671172 176654 671200 186286
rect 671356 177993 671384 190426
rect 671342 177984 671398 177993
rect 671342 177919 671398 177928
rect 671172 176626 671292 176654
rect 670988 157306 671108 157334
rect 670988 155258 671016 157306
rect 670804 155230 671016 155258
rect 670804 155174 670832 155230
rect 670792 155168 670844 155174
rect 670792 155110 670844 155116
rect 671264 151814 671292 176626
rect 670804 151786 671292 151814
rect 670606 147656 670662 147665
rect 670606 147591 670662 147600
rect 670804 146062 670832 151786
rect 670792 146056 670844 146062
rect 670792 145998 670844 146004
rect 671540 138014 671568 223615
rect 671724 150113 671752 223944
rect 672078 223887 672134 223896
rect 671894 221776 671950 221785
rect 671894 221711 671950 221720
rect 671908 218657 671936 221711
rect 671894 218648 671950 218657
rect 671894 218583 671950 218592
rect 672092 217569 672120 223887
rect 672078 217560 672134 217569
rect 672078 217495 672134 217504
rect 671894 216200 671950 216209
rect 671894 216135 671950 216144
rect 672078 216200 672134 216209
rect 672078 216135 672134 216144
rect 671908 215393 671936 216135
rect 671894 215384 671950 215393
rect 671894 215319 671950 215328
rect 672092 201385 672120 216135
rect 672078 201376 672134 201385
rect 672078 201311 672134 201320
rect 671894 172000 671950 172009
rect 671894 171935 671950 171944
rect 671908 166994 671936 171935
rect 672078 169144 672134 169153
rect 672078 169079 672134 169088
rect 672092 168042 672120 169079
rect 672276 168201 672304 225542
rect 672460 225542 672534 225570
rect 672460 225049 672488 225542
rect 672446 225040 672502 225049
rect 672446 224975 672502 224984
rect 672630 223680 672686 223689
rect 672630 223615 672686 223624
rect 672644 222194 672672 223615
rect 672460 222166 672672 222194
rect 672460 213217 672488 222166
rect 672920 220697 672948 226902
rect 673092 226568 673144 226574
rect 673092 226510 673144 226516
rect 673104 222873 673132 226510
rect 673380 223689 673408 229570
rect 673552 229152 673604 229158
rect 673552 229094 673604 229100
rect 673564 226817 673592 229094
rect 673550 226808 673606 226817
rect 673550 226743 673606 226752
rect 673550 224768 673606 224777
rect 673550 224703 673606 224712
rect 673366 223680 673422 223689
rect 673366 223615 673422 223624
rect 673090 222864 673146 222873
rect 673090 222799 673146 222808
rect 673182 221096 673238 221105
rect 673182 221031 673238 221040
rect 672906 220688 672962 220697
rect 672906 220623 672962 220632
rect 672998 217424 673054 217433
rect 672998 217359 673054 217368
rect 673012 216617 673040 217359
rect 672998 216608 673054 216617
rect 672998 216543 673054 216552
rect 673196 215294 673224 221031
rect 673366 220280 673422 220289
rect 673366 220215 673422 220224
rect 673196 215266 673316 215294
rect 673090 214160 673146 214169
rect 673090 214095 673146 214104
rect 672630 213344 672686 213353
rect 672630 213279 672686 213288
rect 672446 213208 672502 213217
rect 672446 213143 672502 213152
rect 672446 212120 672502 212129
rect 672446 212055 672502 212064
rect 672460 201113 672488 212055
rect 672644 205634 672672 213279
rect 672644 205606 672948 205634
rect 672920 202874 672948 205606
rect 672736 202846 672948 202874
rect 672446 201104 672502 201113
rect 672446 201039 672502 201048
rect 672538 200832 672594 200841
rect 672538 200767 672594 200776
rect 672552 181665 672580 200767
rect 672538 181656 672594 181665
rect 672538 181591 672594 181600
rect 672538 168328 672594 168337
rect 672538 168263 672594 168272
rect 672262 168192 672318 168201
rect 672262 168127 672318 168136
rect 672092 168014 672396 168042
rect 671908 166966 672028 166994
rect 671710 150104 671766 150113
rect 671710 150039 671766 150048
rect 672000 144945 672028 166966
rect 672170 166968 672226 166977
rect 672170 166903 672226 166912
rect 671986 144936 672042 144945
rect 671986 144871 672042 144880
rect 670804 137986 671568 138014
rect 670804 130694 670832 137986
rect 671342 130928 671398 130937
rect 671342 130863 671398 130872
rect 670792 130688 670844 130694
rect 670792 130630 670844 130636
rect 670148 129600 670200 129606
rect 670148 129542 670200 129548
rect 669962 129296 670018 129305
rect 669962 129231 670018 129240
rect 669226 125760 669282 125769
rect 669226 125695 669282 125704
rect 668780 122806 668900 122834
rect 668780 119241 668808 122806
rect 668950 120728 669006 120737
rect 668950 120663 669006 120672
rect 668766 119232 668822 119241
rect 668766 119167 668822 119176
rect 668964 111081 668992 120663
rect 668950 111072 669006 111081
rect 668950 111007 669006 111016
rect 669976 104582 670004 129231
rect 670146 122768 670202 122777
rect 670146 122703 670202 122712
rect 670160 112946 670188 122703
rect 670148 112940 670200 112946
rect 670148 112882 670200 112888
rect 671356 109034 671384 130863
rect 671986 126576 672042 126585
rect 671986 126511 672042 126520
rect 670804 109006 671384 109034
rect 670804 108050 670832 109006
rect 670792 108044 670844 108050
rect 670792 107986 670844 107992
rect 669964 104576 670016 104582
rect 669964 104518 670016 104524
rect 668582 102912 668638 102921
rect 668582 102847 668638 102856
rect 595272 100014 595608 100042
rect 596192 100014 596344 100042
rect 596468 100014 597080 100042
rect 597664 100014 597816 100042
rect 597940 100014 598552 100042
rect 599136 100014 599288 100042
rect 599688 100014 600024 100042
rect 600332 100014 600760 100042
rect 600884 100014 601496 100042
rect 601712 100014 602232 100042
rect 602356 100014 602968 100042
rect 603092 100014 603704 100042
rect 595272 99142 595300 100014
rect 595260 99136 595312 99142
rect 595260 99078 595312 99084
rect 595272 93854 595300 99078
rect 595272 93826 595484 93854
rect 595456 80714 595484 93826
rect 595444 80708 595496 80714
rect 595444 80650 595496 80656
rect 596192 54398 596220 100014
rect 596468 55214 596496 100014
rect 596456 55208 596508 55214
rect 596456 55150 596508 55156
rect 597664 55078 597692 100014
rect 597652 55072 597704 55078
rect 597652 55014 597704 55020
rect 597940 54942 597968 100014
rect 598940 96960 598992 96966
rect 598940 96902 598992 96908
rect 598952 56030 598980 96902
rect 598940 56024 598992 56030
rect 598940 55966 598992 55972
rect 597928 54936 597980 54942
rect 597928 54878 597980 54884
rect 599136 54806 599164 100014
rect 599688 96966 599716 100014
rect 599676 96960 599728 96966
rect 599676 96902 599728 96908
rect 600332 55894 600360 100014
rect 600884 84194 600912 100014
rect 600516 84166 600912 84194
rect 600516 57254 600544 84166
rect 601712 72486 601740 100014
rect 602356 84194 602384 100014
rect 601896 84166 602384 84194
rect 601700 72480 601752 72486
rect 601700 72422 601752 72428
rect 601896 58682 601924 84166
rect 603092 60042 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 606984 100042
rect 607384 100014 607720 100042
rect 608120 100014 608548 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 604426 99742 604500 99770
rect 604472 68338 604500 99742
rect 605484 97306 605512 100014
rect 605472 97300 605524 97306
rect 605472 97242 605524 97248
rect 606220 96966 606248 100014
rect 606208 96960 606260 96966
rect 606208 96902 606260 96908
rect 606956 92886 606984 100014
rect 607128 96960 607180 96966
rect 607128 96902 607180 96908
rect 606944 92880 606996 92886
rect 606944 92822 606996 92828
rect 607140 75206 607168 96902
rect 607692 95946 607720 100014
rect 607680 95940 607732 95946
rect 607680 95882 607732 95888
rect 608520 84182 608548 100014
rect 609164 94518 609192 100014
rect 609152 94512 609204 94518
rect 609152 94454 609204 94460
rect 609900 85406 609928 100014
rect 610636 96762 610664 100014
rect 611050 99770 611078 100028
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 613272 100014 613792 100042
rect 611050 99742 611124 99770
rect 610624 96756 610676 96762
rect 610624 96698 610676 96704
rect 611096 96082 611124 99742
rect 611912 97300 611964 97306
rect 611912 97242 611964 97248
rect 611268 96756 611320 96762
rect 611268 96698 611320 96704
rect 611084 96076 611136 96082
rect 611084 96018 611136 96024
rect 611280 93158 611308 96698
rect 611924 93854 611952 97242
rect 612108 96898 612136 100014
rect 612660 97442 612688 100014
rect 612648 97436 612700 97442
rect 612648 97378 612700 97384
rect 612096 96892 612148 96898
rect 612096 96834 612148 96840
rect 612648 96892 612700 96898
rect 612648 96834 612700 96840
rect 611924 93826 612044 93854
rect 611268 93152 611320 93158
rect 611268 93094 611320 93100
rect 610072 92880 610124 92886
rect 610072 92822 610124 92828
rect 610084 88330 610112 92822
rect 610072 88324 610124 88330
rect 610072 88266 610124 88272
rect 609888 85400 609940 85406
rect 609888 85342 609940 85348
rect 608508 84176 608560 84182
rect 608508 84118 608560 84124
rect 612016 76566 612044 93826
rect 612660 80850 612688 96834
rect 612648 80844 612700 80850
rect 612648 80786 612700 80792
rect 613764 79490 613792 100014
rect 613994 99770 614022 100028
rect 614744 100014 615264 100042
rect 615480 100014 615816 100042
rect 616216 100014 616552 100042
rect 616952 100014 617288 100042
rect 617688 100014 618024 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620232 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 613948 99742 614022 99770
rect 613752 79484 613804 79490
rect 613752 79426 613804 79432
rect 613948 79354 613976 99742
rect 615236 93854 615264 100014
rect 615788 96966 615816 100014
rect 615776 96960 615828 96966
rect 615776 96902 615828 96908
rect 616524 95062 616552 100014
rect 616788 96960 616840 96966
rect 616788 96902 616840 96908
rect 616512 95056 616564 95062
rect 616512 94998 616564 95004
rect 615236 93826 615448 93854
rect 613936 79348 613988 79354
rect 613936 79290 613988 79296
rect 612004 76560 612056 76566
rect 612004 76502 612056 76508
rect 615420 75342 615448 93826
rect 616800 76702 616828 96902
rect 617260 96898 617288 100014
rect 617248 96892 617300 96898
rect 617248 96834 617300 96840
rect 617996 92478 618024 100014
rect 618732 97850 618760 100014
rect 618720 97844 618772 97850
rect 618720 97786 618772 97792
rect 618904 97436 618956 97442
rect 618904 97378 618956 97384
rect 618168 96892 618220 96898
rect 618168 96834 618220 96840
rect 617984 92472 618036 92478
rect 617984 92414 618036 92420
rect 618180 91050 618208 96834
rect 618168 91044 618220 91050
rect 618168 90986 618220 90992
rect 616788 76696 616840 76702
rect 616788 76638 616840 76644
rect 618916 75478 618944 97378
rect 619560 93838 619588 100014
rect 620204 97986 620232 100014
rect 620192 97980 620244 97986
rect 620192 97922 620244 97928
rect 620940 95198 620968 100014
rect 621676 97578 621704 100014
rect 622320 99346 622348 100014
rect 622308 99340 622360 99346
rect 622308 99282 622360 99288
rect 621664 97572 621716 97578
rect 621664 97514 621716 97520
rect 623148 97442 623176 100014
rect 623700 99210 623728 100014
rect 623688 99204 623740 99210
rect 623688 99146 623740 99152
rect 623136 97436 623188 97442
rect 623136 97378 623188 97384
rect 624620 97034 624648 100014
rect 625034 99770 625062 100028
rect 625784 100014 626120 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628328 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 632008 100042
rect 632408 100014 632744 100042
rect 633144 100014 633296 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635596 100042
rect 625034 99742 625108 99770
rect 625080 99074 625108 99742
rect 625068 99068 625120 99074
rect 625068 99010 625120 99016
rect 625804 97844 625856 97850
rect 625804 97786 625856 97792
rect 624608 97028 624660 97034
rect 624608 96970 624660 96976
rect 622124 96076 622176 96082
rect 622124 96018 622176 96024
rect 620928 95192 620980 95198
rect 620928 95134 620980 95140
rect 620284 94512 620336 94518
rect 620284 94454 620336 94460
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 619272 93152 619324 93158
rect 619272 93094 619324 93100
rect 619284 86358 619312 93094
rect 619272 86352 619324 86358
rect 619272 86294 619324 86300
rect 620296 85542 620324 94454
rect 622136 88194 622164 96018
rect 624976 95940 625028 95946
rect 624976 95882 625028 95888
rect 623044 95056 623096 95062
rect 623044 94998 623096 95004
rect 623056 89690 623084 94998
rect 623044 89684 623096 89690
rect 623044 89626 623096 89632
rect 624988 88369 625016 95882
rect 625816 92041 625844 97786
rect 626092 97306 626120 100014
rect 626264 97980 626316 97986
rect 626264 97922 626316 97928
rect 626080 97300 626132 97306
rect 626080 97242 626132 97248
rect 626276 93673 626304 97922
rect 626828 97170 626856 100014
rect 627564 97850 627592 100014
rect 628300 98938 628328 100014
rect 628288 98932 628340 98938
rect 628288 98874 628340 98880
rect 629036 98802 629064 100014
rect 629024 98796 629076 98802
rect 629024 98738 629076 98744
rect 629772 97986 629800 100014
rect 630508 98530 630536 100014
rect 630772 99340 630824 99346
rect 630772 99282 630824 99288
rect 630496 98524 630548 98530
rect 630496 98466 630548 98472
rect 629760 97980 629812 97986
rect 629760 97922 629812 97928
rect 627552 97844 627604 97850
rect 627552 97786 627604 97792
rect 629300 97572 629352 97578
rect 629300 97514 629352 97520
rect 626816 97164 626868 97170
rect 626816 97106 626868 97112
rect 629312 95826 629340 97514
rect 630784 95826 630812 99282
rect 631048 98252 631100 98258
rect 631048 98194 631100 98200
rect 631060 97850 631088 98194
rect 631048 97844 631100 97850
rect 631048 97786 631100 97792
rect 631244 96354 631272 100014
rect 631980 97578 632008 100014
rect 631968 97572 632020 97578
rect 631968 97514 632020 97520
rect 632060 97436 632112 97442
rect 632060 97378 632112 97384
rect 631232 96348 631284 96354
rect 631232 96290 631284 96296
rect 629280 95798 629340 95826
rect 630752 95798 630812 95826
rect 632072 95826 632100 97378
rect 632716 96898 632744 100014
rect 633268 97442 633296 100014
rect 633440 99204 633492 99210
rect 633440 99146 633492 99152
rect 633256 97436 633308 97442
rect 633256 97378 633308 97384
rect 632704 96892 632756 96898
rect 632704 96834 632756 96840
rect 633452 95826 633480 99146
rect 634188 97850 634216 100014
rect 634176 97844 634228 97850
rect 634176 97786 634228 97792
rect 634740 97714 634768 100014
rect 634728 97708 634780 97714
rect 634728 97650 634780 97656
rect 635568 97034 635596 100014
rect 635752 100014 636088 100042
rect 636824 100014 637068 100042
rect 635004 97028 635056 97034
rect 635004 96970 635056 96976
rect 635556 97028 635608 97034
rect 635556 96970 635608 96976
rect 635016 95826 635044 96970
rect 632072 95798 632224 95826
rect 633452 95798 633696 95826
rect 635016 95798 635168 95826
rect 635752 95441 635780 100014
rect 636292 99068 636344 99074
rect 636292 99010 636344 99016
rect 636304 95826 636332 99010
rect 637040 96937 637068 100014
rect 637546 99770 637574 100028
rect 638296 100014 638632 100042
rect 637546 99742 637620 99770
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 96218 637620 99742
rect 637764 97300 637816 97306
rect 637764 97242 637816 97248
rect 637580 96212 637632 96218
rect 637580 96154 637632 96160
rect 637776 95826 637804 97242
rect 636304 95798 636640 95826
rect 637776 95798 638112 95826
rect 638604 95742 638632 100014
rect 639018 99770 639046 100028
rect 639768 100014 640104 100042
rect 639018 99742 639092 99770
rect 639064 96490 639092 99742
rect 639236 97164 639288 97170
rect 639236 97106 639288 97112
rect 639052 96484 639104 96490
rect 639052 96426 639104 96432
rect 639248 95826 639276 97106
rect 639248 95798 639584 95826
rect 638592 95736 638644 95742
rect 638592 95678 638644 95684
rect 640076 95606 640104 100014
rect 640490 99770 640518 100028
rect 641240 100014 641576 100042
rect 640490 99742 640564 99770
rect 640536 96626 640564 99742
rect 640708 98184 640760 98190
rect 640708 98126 640760 98132
rect 640524 96620 640576 96626
rect 640524 96562 640576 96568
rect 640720 95826 640748 98126
rect 640720 95798 641056 95826
rect 640064 95600 640116 95606
rect 640064 95542 640116 95548
rect 641548 95470 641576 100014
rect 641962 99770 641990 100028
rect 642712 100014 643048 100042
rect 641962 99742 642036 99770
rect 642008 96529 642036 99742
rect 642180 98932 642232 98938
rect 642180 98874 642232 98880
rect 641994 96520 642050 96529
rect 641994 96455 642050 96464
rect 642192 95826 642220 98874
rect 643020 97170 643048 100014
rect 643434 99770 643462 100028
rect 644184 100014 644336 100042
rect 643434 99742 643508 99770
rect 643008 97164 643060 97170
rect 643008 97106 643060 97112
rect 643480 95878 643508 99742
rect 643652 98796 643704 98802
rect 643652 98738 643704 98744
rect 643468 95872 643520 95878
rect 642192 95798 642528 95826
rect 643468 95814 643520 95820
rect 643664 95826 643692 98738
rect 644308 97306 644336 100014
rect 644906 99770 644934 100028
rect 645656 100014 645808 100042
rect 644906 99742 644980 99770
rect 644296 97300 644348 97306
rect 644296 97242 644348 97248
rect 644952 96014 644980 99742
rect 645308 98048 645360 98054
rect 645308 97990 645360 97996
rect 645124 96484 645176 96490
rect 645124 96426 645176 96432
rect 644940 96008 644992 96014
rect 644940 95950 644992 95956
rect 643664 95798 644000 95826
rect 645136 95470 645164 96426
rect 645320 95826 645348 97990
rect 645780 96626 645808 100014
rect 646378 99770 646406 100028
rect 647114 99770 647142 100028
rect 647864 100014 648476 100042
rect 648600 100014 648936 100042
rect 649336 100014 649764 100042
rect 650072 100014 650408 100042
rect 650808 100014 651328 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 655224 100014 655468 100042
rect 646378 99742 646452 99770
rect 647114 99742 647188 99770
rect 645768 96620 645820 96626
rect 645768 96562 645820 96568
rect 646424 96490 646452 99742
rect 647160 98666 647188 99742
rect 647148 98660 647200 98666
rect 647148 98602 647200 98608
rect 646596 98524 646648 98530
rect 646596 98466 646648 98472
rect 646412 96484 646464 96490
rect 646412 96426 646464 96432
rect 646608 95826 646636 98466
rect 647516 97572 647568 97578
rect 647516 97514 647568 97520
rect 647148 96348 647200 96354
rect 647148 96290 647200 96296
rect 645320 95798 645472 95826
rect 646608 95798 646944 95826
rect 641536 95464 641588 95470
rect 635738 95432 635794 95441
rect 641536 95406 641588 95412
rect 645124 95464 645176 95470
rect 645124 95406 645176 95412
rect 635738 95367 635794 95376
rect 626448 95192 626500 95198
rect 626448 95134 626500 95140
rect 626460 94489 626488 95134
rect 647160 95033 647188 96290
rect 647332 95736 647384 95742
rect 647332 95678 647384 95684
rect 647146 95024 647202 95033
rect 647146 94959 647202 94968
rect 626446 94480 626502 94489
rect 626446 94415 626502 94424
rect 626448 93832 626500 93838
rect 626448 93774 626500 93780
rect 626262 93664 626318 93673
rect 626262 93599 626318 93608
rect 626460 92857 626488 93774
rect 626446 92848 626502 92857
rect 626446 92783 626502 92792
rect 626448 92472 626500 92478
rect 626448 92414 626500 92420
rect 625802 92032 625858 92041
rect 625802 91967 625858 91976
rect 626460 91225 626488 92414
rect 647344 92410 647372 95678
rect 647528 92449 647556 97514
rect 647700 97028 647752 97034
rect 647700 96970 647752 96976
rect 647712 95198 647740 96970
rect 648252 96892 648304 96898
rect 648252 96834 648304 96840
rect 647884 96756 647936 96762
rect 647884 96698 647936 96704
rect 647896 95742 647924 96698
rect 647884 95736 647936 95742
rect 647884 95678 647936 95684
rect 647884 95600 647936 95606
rect 647884 95542 647936 95548
rect 647700 95192 647752 95198
rect 647700 95134 647752 95140
rect 647514 92440 647570 92449
rect 647332 92404 647384 92410
rect 647514 92375 647570 92384
rect 647332 92346 647384 92352
rect 626446 91216 626502 91225
rect 626446 91151 626502 91160
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90409 626488 90986
rect 626446 90400 626502 90409
rect 626446 90335 626502 90344
rect 626448 89616 626500 89622
rect 626446 89584 626448 89593
rect 626500 89584 626502 89593
rect 626446 89519 626502 89528
rect 624974 88360 625030 88369
rect 624974 88295 625030 88304
rect 626448 88324 626500 88330
rect 626448 88266 626500 88272
rect 622124 88188 622176 88194
rect 622124 88130 622176 88136
rect 626264 88188 626316 88194
rect 626264 88130 626316 88136
rect 626276 87145 626304 88130
rect 626460 87961 626488 88266
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 626262 87136 626318 87145
rect 626262 87071 626318 87080
rect 647896 86630 647924 95542
rect 648264 89593 648292 96834
rect 648250 89584 648306 89593
rect 648250 89519 648306 89528
rect 648448 87038 648476 100014
rect 648620 97436 648672 97442
rect 648620 97378 648672 97384
rect 648632 92546 648660 97378
rect 648908 96354 648936 100014
rect 648896 96348 648948 96354
rect 648896 96290 648948 96296
rect 649080 96008 649132 96014
rect 649080 95950 649132 95956
rect 648804 95192 648856 95198
rect 648804 95134 648856 95140
rect 648620 92540 648672 92546
rect 648620 92482 648672 92488
rect 648436 87032 648488 87038
rect 648436 86974 648488 86980
rect 647884 86624 647936 86630
rect 647884 86566 647936 86572
rect 626448 86352 626500 86358
rect 626446 86320 626448 86329
rect 626500 86320 626502 86329
rect 626446 86255 626502 86264
rect 620284 85536 620336 85542
rect 626448 85536 626500 85542
rect 620284 85478 620336 85484
rect 625342 85504 625398 85513
rect 626448 85478 626500 85484
rect 625342 85439 625398 85448
rect 625356 85338 625384 85439
rect 625344 85332 625396 85338
rect 625344 85274 625396 85280
rect 626460 84697 626488 85478
rect 626446 84688 626502 84697
rect 626446 84623 626502 84632
rect 625804 84176 625856 84182
rect 625804 84118 625856 84124
rect 625816 83881 625844 84118
rect 625802 83872 625858 83881
rect 625802 83807 625858 83816
rect 628746 83328 628802 83337
rect 628746 83263 628802 83272
rect 628760 80986 628788 83263
rect 629206 81696 629262 81705
rect 629206 81631 629262 81640
rect 628748 80980 628800 80986
rect 628748 80922 628800 80928
rect 629220 80034 629248 81631
rect 632808 80974 633144 81002
rect 642456 80980 642508 80986
rect 629208 80028 629260 80034
rect 629208 79970 629260 79976
rect 631048 77988 631100 77994
rect 631048 77930 631100 77936
rect 628472 77784 628524 77790
rect 628472 77726 628524 77732
rect 624422 77344 624478 77353
rect 624422 77279 624478 77288
rect 625804 77308 625856 77314
rect 618904 75472 618956 75478
rect 618904 75414 618956 75420
rect 615408 75336 615460 75342
rect 615408 75278 615460 75284
rect 607128 75200 607180 75206
rect 607128 75142 607180 75148
rect 604460 68332 604512 68338
rect 604460 68274 604512 68280
rect 603080 60036 603132 60042
rect 603080 59978 603132 59984
rect 601884 58676 601936 58682
rect 601884 58618 601936 58624
rect 600504 57248 600556 57254
rect 600504 57190 600556 57196
rect 600320 55888 600372 55894
rect 600320 55830 600372 55836
rect 599124 54800 599176 54806
rect 599124 54742 599176 54748
rect 624436 54670 624464 77279
rect 625804 77250 625856 77256
rect 624424 54664 624476 54670
rect 624424 54606 624476 54612
rect 625816 54534 625844 77250
rect 628484 75290 628512 77726
rect 631060 77314 631088 77930
rect 632808 77790 632836 80974
rect 643080 80974 643140 81002
rect 642456 80922 642508 80928
rect 636752 80708 636804 80714
rect 636752 80650 636804 80656
rect 633440 80028 633492 80034
rect 633440 79970 633492 79976
rect 633452 78130 633480 79970
rect 633898 78568 633954 78577
rect 633898 78503 633954 78512
rect 633440 78124 633492 78130
rect 633440 78066 633492 78072
rect 632796 77784 632848 77790
rect 632796 77726 632848 77732
rect 633912 77353 633940 78503
rect 633898 77344 633954 77353
rect 631048 77308 631100 77314
rect 633898 77279 633954 77288
rect 631048 77250 631100 77256
rect 631060 75290 631088 77250
rect 633912 75290 633940 77279
rect 636764 75290 636792 80650
rect 639602 78160 639658 78169
rect 639602 78095 639658 78104
rect 639616 75290 639644 78095
rect 642468 75290 642496 80922
rect 643112 77994 643140 80974
rect 647424 80844 647476 80850
rect 647424 80786 647476 80792
rect 645952 79484 646004 79490
rect 645952 79426 646004 79432
rect 645308 78124 645360 78130
rect 645308 78066 645360 78072
rect 643100 77988 643152 77994
rect 643100 77930 643152 77936
rect 645320 75290 645348 78066
rect 628176 75262 628512 75290
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 636732 75262 636792 75290
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 645964 64874 645992 79426
rect 646504 79348 646556 79354
rect 646504 79290 646556 79296
rect 646320 76696 646372 76702
rect 646320 76638 646372 76644
rect 646136 75200 646188 75206
rect 646136 75142 646188 75148
rect 646148 74225 646176 75142
rect 646134 74216 646190 74225
rect 646134 74151 646190 74160
rect 646332 71777 646360 76638
rect 646318 71768 646374 71777
rect 646318 71703 646374 71712
rect 646516 67153 646544 79290
rect 646872 75336 646924 75342
rect 646872 75278 646924 75284
rect 646884 74534 646912 75278
rect 646884 74506 647280 74534
rect 647252 68921 647280 74506
rect 647238 68912 647294 68921
rect 647238 68847 647294 68856
rect 646502 67144 646558 67153
rect 646502 67079 646558 67088
rect 647436 64874 647464 80786
rect 648620 75472 648672 75478
rect 648620 75414 648672 75420
rect 645964 64846 646176 64874
rect 646148 64433 646176 64846
rect 647252 64846 647464 64874
rect 646134 64424 646190 64433
rect 646134 64359 646190 64368
rect 647252 59265 647280 64846
rect 648632 62121 648660 75414
rect 648618 62112 648674 62121
rect 648618 62047 648674 62056
rect 647238 59256 647294 59265
rect 647238 59191 647294 59200
rect 648816 57361 648844 95134
rect 649092 93294 649120 95950
rect 649264 95872 649316 95878
rect 649264 95814 649316 95820
rect 649080 93288 649132 93294
rect 649080 93230 649132 93236
rect 649276 86766 649304 95814
rect 649736 88806 649764 100014
rect 650184 97708 650236 97714
rect 650184 97650 650236 97656
rect 649908 96076 649960 96082
rect 649908 96018 649960 96024
rect 649920 95334 649948 96018
rect 649908 95328 649960 95334
rect 649908 95270 649960 95276
rect 650196 93854 650224 97650
rect 650380 97510 650408 100014
rect 650552 97844 650604 97850
rect 650552 97786 650604 97792
rect 650368 97504 650420 97510
rect 650368 97446 650420 97452
rect 650196 93826 650408 93854
rect 650000 92540 650052 92546
rect 650000 92482 650052 92488
rect 649724 88800 649776 88806
rect 649724 88742 649776 88748
rect 650012 87145 650040 92482
rect 649998 87136 650054 87145
rect 649998 87071 650054 87080
rect 649264 86760 649316 86766
rect 649264 86702 649316 86708
rect 650380 82249 650408 93826
rect 650564 84697 650592 97786
rect 651300 93566 651328 100014
rect 651852 97714 651880 100014
rect 651840 97708 651892 97714
rect 651840 97650 651892 97656
rect 652588 96490 652616 100014
rect 652024 96484 652076 96490
rect 652024 96426 652076 96432
rect 652576 96484 652628 96490
rect 652576 96426 652628 96432
rect 651840 95464 651892 95470
rect 651840 95406 651892 95412
rect 651288 93560 651340 93566
rect 651288 93502 651340 93508
rect 651852 90710 651880 95406
rect 651840 90704 651892 90710
rect 651840 90646 651892 90652
rect 652036 86358 652064 96426
rect 653324 95674 653352 100014
rect 653968 96898 653996 100014
rect 654796 96898 654824 100014
rect 655440 97850 655468 100014
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655428 97844 655480 97850
rect 655428 97786 655480 97792
rect 653956 96892 654008 96898
rect 653956 96834 654008 96840
rect 654600 96892 654652 96898
rect 654600 96834 654652 96840
rect 654784 96892 654836 96898
rect 654784 96834 654836 96840
rect 655428 96892 655480 96898
rect 655428 96834 655480 96840
rect 653312 95668 653364 95674
rect 653312 95610 653364 95616
rect 654612 94217 654640 96834
rect 654598 94208 654654 94217
rect 654598 94143 654654 94152
rect 655440 93854 655468 96834
rect 655256 93826 655468 93854
rect 654324 92404 654376 92410
rect 654324 92346 654376 92352
rect 654336 91497 654364 92346
rect 654322 91488 654378 91497
rect 654322 91423 654378 91432
rect 655256 88330 655284 93826
rect 655428 93560 655480 93566
rect 655428 93502 655480 93508
rect 655440 93401 655468 93502
rect 655426 93392 655482 93401
rect 655426 93327 655482 93336
rect 655428 90704 655480 90710
rect 655426 90672 655428 90681
rect 655480 90672 655482 90681
rect 655426 90607 655482 90616
rect 655808 89865 655836 100014
rect 656820 97238 656848 100014
rect 656808 97232 656860 97238
rect 656808 97174 656860 97180
rect 656716 96960 656768 96966
rect 656716 96902 656768 96908
rect 656348 96620 656400 96626
rect 656348 96562 656400 96568
rect 656164 93288 656216 93294
rect 656164 93230 656216 93236
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 655244 88324 655296 88330
rect 655244 88266 655296 88272
rect 656176 86494 656204 93230
rect 656360 88670 656388 96562
rect 656348 88664 656400 88670
rect 656348 88606 656400 88612
rect 656728 86902 656756 96902
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 658108 99742 658182 99770
rect 658108 97374 658136 99742
rect 659212 97986 659240 100014
rect 659200 97980 659252 97986
rect 659200 97922 659252 97928
rect 659948 97850 659976 100014
rect 660132 100014 660376 100042
rect 659936 97844 659988 97850
rect 659936 97786 659988 97792
rect 659568 97708 659620 97714
rect 659568 97650 659620 97656
rect 658280 97504 658332 97510
rect 658280 97446 658332 97452
rect 658096 97368 658148 97374
rect 658096 97310 658148 97316
rect 658292 95132 658320 97446
rect 658832 97096 658884 97102
rect 658832 97038 658884 97044
rect 658844 95132 658872 97038
rect 659580 95132 659608 97650
rect 660132 96966 660160 100014
rect 672000 99385 672028 126511
rect 672184 115841 672212 166903
rect 672368 152697 672396 168014
rect 672354 152688 672410 152697
rect 672354 152623 672410 152632
rect 672552 138014 672580 168263
rect 672368 137986 672580 138014
rect 672368 131209 672396 137986
rect 672538 133376 672594 133385
rect 672538 133311 672594 133320
rect 672552 132705 672580 133311
rect 672538 132696 672594 132705
rect 672538 132631 672594 132640
rect 672538 131744 672594 131753
rect 672538 131679 672594 131688
rect 672354 131200 672410 131209
rect 672354 131135 672410 131144
rect 672552 118694 672580 131679
rect 672736 124137 672764 202846
rect 672906 200696 672962 200705
rect 672906 200631 672962 200640
rect 672920 126993 672948 200631
rect 673104 199753 673132 214095
rect 673090 199744 673146 199753
rect 673090 199679 673146 199688
rect 673288 199594 673316 215266
rect 673196 199566 673316 199594
rect 673196 197849 673224 199566
rect 673182 197840 673238 197849
rect 673182 197775 673238 197784
rect 673380 175681 673408 220215
rect 673564 216889 673592 224703
rect 673550 216880 673606 216889
rect 673550 216815 673606 216824
rect 673550 216608 673606 216617
rect 673550 216543 673606 216552
rect 673564 215937 673592 216543
rect 673550 215928 673606 215937
rect 673550 215863 673606 215872
rect 673748 213738 673776 236422
rect 673564 213710 673776 213738
rect 673564 213246 673592 213710
rect 673840 213330 673868 236558
rect 673932 224954 673960 266999
rect 674378 266248 674434 266257
rect 674378 266183 674434 266192
rect 674392 263594 674420 266183
rect 674576 265849 674604 277366
rect 674562 265840 674618 265849
rect 674562 265775 674618 265784
rect 674760 265033 674788 287026
rect 675114 286920 675170 286929
rect 675170 286878 675340 286906
rect 675114 286855 675170 286864
rect 675312 286770 675340 286878
rect 675404 286770 675432 286892
rect 675312 286742 675432 286770
rect 675390 286512 675446 286521
rect 675390 286447 675446 286456
rect 675404 286212 675432 286447
rect 675116 285660 675168 285666
rect 675116 285602 675168 285608
rect 675128 285070 675156 285602
rect 675128 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675666 282704 675722 282713
rect 675666 282639 675722 282648
rect 675680 282554 675708 282639
rect 675128 282540 675708 282554
rect 675128 282526 675694 282540
rect 675128 278361 675156 282526
rect 675666 281616 675722 281625
rect 675666 281551 675722 281560
rect 675680 281355 675708 281551
rect 675114 278352 675170 278361
rect 675114 278287 675170 278296
rect 675482 278080 675538 278089
rect 675482 278015 675538 278024
rect 674930 276720 674986 276729
rect 674930 276655 674986 276664
rect 674944 273873 674972 276655
rect 674930 273864 674986 273873
rect 674930 273799 674986 273808
rect 674746 265024 674802 265033
rect 674746 264959 674802 264968
rect 675114 264208 675170 264217
rect 675114 264143 675170 264152
rect 674392 263566 674696 263594
rect 674470 262576 674526 262585
rect 674470 262511 674526 262520
rect 674484 260250 674512 262511
rect 674484 260222 674604 260250
rect 674378 260128 674434 260137
rect 674378 260063 674434 260072
rect 674102 259312 674158 259321
rect 674102 259247 674158 259256
rect 674116 242729 674144 259247
rect 674102 242720 674158 242729
rect 674102 242655 674158 242664
rect 674392 242185 674420 260063
rect 674576 253934 674604 260222
rect 674484 253906 674604 253934
rect 674484 243085 674512 253906
rect 674668 244274 674696 263566
rect 674930 254960 674986 254969
rect 674930 254895 674986 254904
rect 674944 249762 674972 254895
rect 674932 249756 674984 249762
rect 674932 249698 674984 249704
rect 675128 249642 675156 264143
rect 675496 258097 675524 278015
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 676402 264072 676458 264081
rect 676402 264007 676458 264016
rect 676218 262848 676274 262857
rect 676218 262783 676274 262792
rect 676232 259570 676260 262783
rect 675680 259542 676260 259570
rect 675482 258088 675538 258097
rect 675482 258023 675538 258032
rect 675680 253934 675708 259542
rect 676416 258806 676444 264007
rect 675852 258800 675904 258806
rect 675852 258742 675904 258748
rect 676404 258800 676456 258806
rect 676404 258742 676456 258748
rect 675864 254969 675892 258742
rect 675850 254960 675906 254969
rect 675850 254895 675906 254904
rect 674760 249614 675156 249642
rect 675220 253906 675708 253934
rect 674760 246213 674788 249614
rect 674930 249520 674986 249529
rect 674930 249455 674986 249464
rect 674944 249218 674972 249455
rect 674932 249212 674984 249218
rect 674932 249154 674984 249160
rect 674932 249076 674984 249082
rect 674932 249018 674984 249024
rect 674944 248962 674972 249018
rect 674852 248934 674972 248962
rect 674852 246378 674880 248934
rect 675220 248690 675248 253906
rect 675128 248662 675248 248690
rect 675312 251110 675432 251138
rect 675128 248010 675156 248662
rect 675312 248169 675340 251110
rect 675404 251056 675432 251110
rect 675482 250744 675538 250753
rect 675482 250679 675538 250688
rect 675496 250512 675524 250679
rect 675758 250336 675814 250345
rect 675758 250271 675814 250280
rect 675772 249900 675800 250271
rect 675484 249756 675536 249762
rect 675484 249698 675536 249704
rect 675496 249220 675524 249698
rect 675298 248160 675354 248169
rect 675298 248095 675354 248104
rect 675128 247982 675340 248010
rect 675312 247398 675340 247982
rect 675312 247370 675418 247398
rect 675772 246673 675800 246840
rect 675298 246664 675354 246673
rect 675298 246599 675354 246608
rect 675758 246664 675814 246673
rect 675758 246599 675814 246608
rect 674852 246350 675156 246378
rect 675128 246265 675156 246350
rect 675114 246256 675170 246265
rect 674760 246185 674880 246213
rect 675114 246191 675170 246200
rect 675312 246213 675340 246599
rect 675312 246185 675418 246213
rect 674852 245478 674880 246185
rect 675298 245712 675354 245721
rect 675298 245647 675354 245656
rect 675312 245562 675340 245647
rect 675312 245534 675418 245562
rect 674840 245472 674892 245478
rect 675208 245472 675260 245478
rect 674840 245414 674892 245420
rect 675022 245440 675078 245449
rect 675208 245414 675260 245420
rect 675022 245375 675078 245384
rect 674668 244246 674788 244274
rect 674484 243057 674604 243085
rect 674576 243001 674604 243057
rect 674562 242992 674618 243001
rect 674562 242927 674618 242936
rect 674760 242842 674788 244246
rect 674760 242814 674880 242842
rect 674378 242176 674434 242185
rect 674378 242111 674434 242120
rect 674654 236464 674710 236473
rect 674654 236399 674710 236408
rect 674088 234728 674140 234734
rect 674088 234670 674140 234676
rect 674100 234614 674128 234670
rect 674100 234586 674144 234614
rect 674116 233782 674144 234586
rect 674104 233776 674156 233782
rect 674104 233718 674156 233724
rect 674288 233232 674340 233238
rect 674288 233174 674340 233180
rect 674104 232688 674156 232694
rect 674102 232656 674104 232665
rect 674156 232656 674158 232665
rect 674102 232591 674158 232600
rect 674104 232416 674156 232422
rect 674102 232384 674104 232393
rect 674156 232384 674158 232393
rect 674102 232319 674158 232328
rect 674102 230480 674158 230489
rect 674102 230415 674158 230424
rect 674116 230042 674144 230415
rect 674104 230036 674156 230042
rect 674104 229978 674156 229984
rect 674104 229832 674156 229838
rect 674102 229800 674104 229809
rect 674156 229800 674158 229809
rect 674102 229735 674158 229744
rect 674104 229356 674156 229362
rect 674104 229298 674156 229304
rect 674116 227089 674144 229298
rect 674102 227080 674158 227089
rect 674300 227066 674328 233174
rect 674102 227015 674158 227024
rect 674254 227038 674328 227066
rect 674254 226930 674282 227038
rect 674208 226902 674282 226930
rect 673932 224926 674052 224954
rect 674024 222329 674052 224926
rect 674010 222320 674066 222329
rect 674010 222255 674066 222264
rect 674010 217968 674066 217977
rect 674010 217903 674066 217912
rect 674024 215294 674052 217903
rect 674208 215294 674236 226902
rect 674668 226794 674696 236399
rect 674852 234614 674880 242814
rect 675036 237289 675064 245375
rect 675022 237280 675078 237289
rect 675022 237215 675078 237224
rect 675220 234614 675248 245414
rect 675390 243264 675446 243273
rect 675390 243199 675446 243208
rect 675404 243071 675432 243199
rect 675482 242720 675538 242729
rect 675482 242655 675538 242664
rect 675496 242519 675524 242655
rect 675482 242176 675538 242185
rect 675482 242111 675538 242120
rect 675496 241876 675524 242111
rect 675482 241496 675538 241505
rect 675482 241431 675538 241440
rect 675496 241231 675524 241431
rect 675482 240272 675538 240281
rect 675482 240207 675538 240216
rect 675496 240040 675524 240207
rect 675482 238640 675538 238649
rect 675482 238575 675538 238584
rect 675496 238204 675524 238575
rect 675496 237289 675524 237524
rect 675482 237280 675538 237289
rect 675482 237215 675538 237224
rect 675496 236201 675524 236368
rect 675482 236192 675538 236201
rect 675482 236127 675538 236136
rect 675482 235512 675538 235521
rect 675482 235447 675538 235456
rect 674852 234586 675064 234614
rect 675220 234586 675340 234614
rect 674840 231600 674892 231606
rect 674840 231542 674892 231548
rect 674852 230858 674880 231542
rect 674840 230852 674892 230858
rect 674840 230794 674892 230800
rect 673748 213314 673868 213330
rect 673736 213308 673868 213314
rect 673788 213302 673868 213308
rect 673932 215266 674052 215294
rect 674116 215266 674236 215294
rect 674300 226766 674696 226794
rect 673736 213250 673788 213256
rect 673552 213240 673604 213246
rect 673552 213182 673604 213188
rect 673552 213104 673604 213110
rect 673552 213046 673604 213052
rect 673564 211154 673592 213046
rect 673736 212968 673788 212974
rect 673736 212910 673788 212916
rect 673564 211126 673684 211154
rect 673366 175672 673422 175681
rect 673366 175607 673422 175616
rect 673274 174448 673330 174457
rect 673274 174383 673330 174392
rect 673288 168858 673316 174383
rect 673656 173894 673684 211126
rect 673564 173866 673684 173894
rect 673748 173894 673776 212910
rect 673932 177313 673960 215266
rect 673918 177304 673974 177313
rect 673918 177239 673974 177248
rect 673918 176896 673974 176905
rect 673918 176831 673974 176840
rect 673748 173866 673868 173894
rect 673564 172281 673592 173866
rect 673550 172272 673606 172281
rect 673550 172207 673606 172216
rect 673458 171592 673514 171601
rect 673458 171527 673514 171536
rect 673288 168830 673408 168858
rect 673182 168736 673238 168745
rect 673182 168671 673238 168680
rect 673196 151337 673224 168671
rect 673182 151328 673238 151337
rect 673182 151263 673238 151272
rect 673380 129713 673408 168830
rect 673472 166994 673500 171527
rect 673472 166966 673592 166994
rect 673564 160041 673592 166966
rect 673840 164234 673868 173866
rect 673932 167090 673960 176831
rect 674116 172961 674144 215266
rect 674102 172952 674158 172961
rect 674102 172887 674158 172896
rect 674102 172272 674158 172281
rect 674102 172207 674158 172216
rect 673932 167062 674052 167090
rect 674024 164234 674052 167062
rect 673748 164206 673868 164234
rect 673932 164206 674052 164234
rect 673748 162602 673776 164206
rect 673656 162574 673776 162602
rect 673656 160154 673684 162574
rect 673656 160126 673776 160154
rect 673550 160032 673606 160041
rect 673550 159967 673606 159976
rect 673748 159089 673776 160126
rect 673734 159080 673790 159089
rect 673734 159015 673790 159024
rect 673932 132161 673960 164206
rect 674116 162353 674144 172207
rect 674102 162344 674158 162353
rect 674102 162279 674158 162288
rect 674102 162072 674158 162081
rect 674102 162007 674158 162016
rect 673918 132152 673974 132161
rect 673918 132087 673974 132096
rect 673366 129704 673422 129713
rect 673366 129639 673422 129648
rect 673182 128480 673238 128489
rect 673182 128415 673238 128424
rect 673196 128354 673224 128415
rect 673196 128326 673408 128354
rect 672906 126984 672962 126993
rect 672906 126919 672962 126928
rect 672722 124128 672778 124137
rect 672722 124063 672778 124072
rect 672722 123856 672778 123865
rect 672722 123791 672778 123800
rect 672368 118666 672580 118694
rect 672170 115832 672226 115841
rect 672170 115767 672226 115776
rect 672368 106185 672396 118666
rect 672736 106321 672764 123791
rect 672906 123176 672962 123185
rect 672906 123111 672962 123120
rect 672920 114345 672948 123111
rect 672906 114336 672962 114345
rect 672906 114271 672962 114280
rect 672722 106312 672778 106321
rect 672722 106247 672778 106256
rect 672354 106176 672410 106185
rect 672354 106111 672410 106120
rect 673380 103465 673408 128326
rect 673918 124808 673974 124817
rect 673918 124743 673974 124752
rect 673932 107001 673960 124743
rect 674116 117473 674144 162007
rect 674300 153241 674328 226766
rect 674838 226128 674894 226137
rect 674838 226063 674894 226072
rect 674852 221513 674880 226063
rect 675036 221513 675064 234586
rect 675312 222194 675340 234586
rect 675496 228585 675524 235447
rect 675852 234048 675904 234054
rect 675850 234016 675852 234025
rect 678244 234048 678296 234054
rect 675904 234016 675906 234025
rect 678244 233990 678296 233996
rect 675850 233951 675906 233960
rect 675852 232688 675904 232694
rect 675850 232656 675852 232665
rect 675904 232656 675906 232665
rect 675850 232591 675906 232600
rect 676036 232552 676088 232558
rect 676036 232494 676088 232500
rect 676048 232393 676076 232494
rect 676034 232384 676090 232393
rect 676034 232319 676090 232328
rect 676586 230208 676642 230217
rect 676586 230143 676642 230152
rect 675482 228576 675538 228585
rect 675482 228511 675538 228520
rect 676402 227080 676458 227089
rect 676402 227015 676458 227024
rect 676036 226840 676088 226846
rect 676036 226782 676088 226788
rect 675482 225720 675538 225729
rect 675482 225655 675538 225664
rect 675220 222166 675340 222194
rect 674838 221504 674894 221513
rect 674838 221439 674894 221448
rect 675022 221504 675078 221513
rect 675022 221439 675078 221448
rect 674838 219056 674894 219065
rect 674838 218991 674894 219000
rect 674470 214976 674526 214985
rect 674470 214911 674526 214920
rect 674484 197169 674512 214911
rect 674654 213752 674710 213761
rect 674654 213687 674710 213696
rect 674668 205634 674696 213687
rect 674576 205606 674696 205634
rect 674576 202874 674604 205606
rect 674852 205170 674880 218991
rect 675022 218240 675078 218249
rect 675022 218175 675078 218184
rect 675036 205337 675064 218175
rect 675220 217410 675248 222166
rect 675496 219881 675524 225655
rect 675850 225448 675906 225457
rect 675850 225383 675906 225392
rect 675864 224954 675892 225383
rect 675680 224926 675892 224954
rect 675680 221785 675708 224926
rect 676048 223145 676076 226782
rect 676416 224954 676444 227015
rect 676232 224926 676444 224954
rect 676034 223136 676090 223145
rect 676034 223071 676090 223080
rect 676034 221912 676090 221921
rect 676034 221847 676090 221856
rect 675666 221776 675722 221785
rect 675666 221711 675722 221720
rect 675482 219872 675538 219881
rect 675482 219807 675538 219816
rect 676048 217977 676076 221847
rect 676034 217968 676090 217977
rect 676034 217903 676090 217912
rect 676232 217682 676260 224926
rect 676048 217654 676260 217682
rect 675220 217382 675340 217410
rect 675312 212537 675340 217382
rect 676048 215937 676076 217654
rect 676034 215928 676090 215937
rect 676034 215863 676090 215872
rect 675852 215416 675904 215422
rect 675666 215384 675722 215393
rect 675722 215364 675852 215370
rect 675722 215358 675904 215364
rect 675722 215342 675892 215358
rect 675666 215319 675722 215328
rect 676600 215294 676628 230143
rect 678256 226846 678284 233990
rect 683212 232688 683264 232694
rect 683212 232630 683264 232636
rect 683224 227089 683252 232630
rect 683396 232552 683448 232558
rect 683396 232494 683448 232500
rect 683210 227080 683266 227089
rect 683210 227015 683266 227024
rect 678244 226840 678296 226846
rect 676954 226808 677010 226817
rect 678244 226782 678296 226788
rect 676954 226743 677010 226752
rect 676968 215422 676996 226743
rect 683408 222737 683436 232494
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 683394 222728 683450 222737
rect 683394 222663 683450 222672
rect 676956 215416 677008 215422
rect 676956 215358 677008 215364
rect 676232 215266 676628 215294
rect 675758 214432 675814 214441
rect 676232 214418 676260 215266
rect 675814 214390 676260 214418
rect 675758 214367 675814 214376
rect 675298 212528 675354 212537
rect 675298 212463 675354 212472
rect 675206 206952 675262 206961
rect 675206 206887 675262 206896
rect 675220 205889 675248 206887
rect 675220 205861 675418 205889
rect 675036 205309 675418 205337
rect 674852 205142 675156 205170
rect 674930 204232 674986 204241
rect 674930 204167 674986 204176
rect 674944 202881 674972 204167
rect 675128 204049 675156 205142
rect 675404 204241 675432 204680
rect 675390 204232 675446 204241
rect 675390 204167 675446 204176
rect 675128 204021 675418 204049
rect 674576 202846 674788 202874
rect 674470 197160 674526 197169
rect 674470 197095 674526 197104
rect 674760 196058 674788 202846
rect 674930 202872 674986 202881
rect 674930 202807 674986 202816
rect 675758 202736 675814 202745
rect 675758 202671 675814 202680
rect 675772 202195 675800 202671
rect 675496 201385 675524 201620
rect 675482 201376 675538 201385
rect 675482 201311 675538 201320
rect 675128 200994 675418 201022
rect 674930 199744 674986 199753
rect 674930 199679 674986 199688
rect 674944 197350 674972 199679
rect 675128 198529 675156 200994
rect 675772 200025 675800 200328
rect 675758 200016 675814 200025
rect 675758 199951 675814 199960
rect 675114 198520 675170 198529
rect 675114 198455 675170 198464
rect 675482 198248 675538 198257
rect 675482 198183 675538 198192
rect 675496 197880 675524 198183
rect 674944 197322 675248 197350
rect 675220 197282 675248 197322
rect 675404 197282 675432 197336
rect 675220 197254 675432 197282
rect 675390 197160 675446 197169
rect 675390 197095 675446 197104
rect 675404 196656 675432 197095
rect 674760 196030 675418 196058
rect 675772 194585 675800 194820
rect 675758 194576 675814 194585
rect 675758 194511 675814 194520
rect 675758 193216 675814 193225
rect 675758 193151 675814 193160
rect 675772 192984 675800 193151
rect 675666 192808 675722 192817
rect 675666 192743 675722 192752
rect 675680 192372 675708 192743
rect 675128 191134 675418 191162
rect 675128 188873 675156 191134
rect 676126 189136 676182 189145
rect 676126 189071 676182 189080
rect 675114 188864 675170 188873
rect 675114 188799 675170 188808
rect 675298 181384 675354 181393
rect 675298 181319 675354 181328
rect 675312 179081 675340 181319
rect 675482 179480 675538 179489
rect 675482 179415 675538 179424
rect 675298 179072 675354 179081
rect 675298 179007 675354 179016
rect 675496 178129 675524 179415
rect 675666 178800 675722 178809
rect 675666 178735 675722 178744
rect 675482 178120 675538 178129
rect 675482 178055 675538 178064
rect 675680 177721 675708 178735
rect 675666 177712 675722 177721
rect 675666 177647 675722 177656
rect 676140 176654 676168 189071
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 675864 176626 676168 176654
rect 674654 176080 674710 176089
rect 674654 176015 674710 176024
rect 674470 175264 674526 175273
rect 674470 175199 674526 175208
rect 674286 153232 674342 153241
rect 674286 153167 674342 153176
rect 674484 130529 674512 175199
rect 674668 131345 674696 176015
rect 675864 167521 675892 176626
rect 676034 174040 676090 174049
rect 676090 173998 676260 174026
rect 676034 173975 676090 173984
rect 676232 169810 676260 173998
rect 679622 173224 679678 173233
rect 679622 173159 679678 173168
rect 676048 169782 676260 169810
rect 675850 167512 675906 167521
rect 675850 167447 675906 167456
rect 676048 166994 676076 169782
rect 676402 169552 676458 169561
rect 676402 169487 676458 169496
rect 675220 166966 676076 166994
rect 675022 161392 675078 161401
rect 675022 161327 675078 161336
rect 675036 157334 675064 161327
rect 675220 159066 675248 166966
rect 676416 166433 676444 169487
rect 676402 166424 676458 166433
rect 676402 166359 676458 166368
rect 679636 163266 679664 173159
rect 681002 172816 681058 172825
rect 681002 172751 681058 172760
rect 675852 163260 675904 163266
rect 675852 163202 675904 163208
rect 679624 163260 679676 163266
rect 679624 163202 679676 163208
rect 675864 161786 675892 163202
rect 681016 162790 681044 172751
rect 683118 167920 683174 167929
rect 683118 167855 683174 167864
rect 676036 162784 676088 162790
rect 676036 162726 676088 162732
rect 681004 162784 681056 162790
rect 681004 162726 681056 162732
rect 675312 161758 675892 161786
rect 675312 160290 675340 161758
rect 676048 161401 676076 162726
rect 683132 162081 683160 167855
rect 683118 162072 683174 162081
rect 683118 162007 683174 162016
rect 676034 161392 676090 161401
rect 676034 161327 676090 161336
rect 675482 161120 675538 161129
rect 675482 161055 675538 161064
rect 675496 160888 675524 161055
rect 675404 160290 675432 160344
rect 675312 160262 675432 160290
rect 675390 160032 675446 160041
rect 675390 159967 675446 159976
rect 675404 159664 675432 159967
rect 675220 159038 675340 159066
rect 675312 158930 675340 159038
rect 675404 158930 675432 159052
rect 675312 158902 675432 158930
rect 675036 157306 675248 157334
rect 675220 157230 675248 157306
rect 675220 157202 675340 157230
rect 675312 157162 675340 157202
rect 675404 157162 675432 157216
rect 675312 157134 675432 157162
rect 675128 156629 675418 156657
rect 675128 154465 675156 156629
rect 675404 155553 675432 155992
rect 675758 155816 675814 155825
rect 675758 155751 675814 155760
rect 675390 155544 675446 155553
rect 675390 155479 675446 155488
rect 675772 155380 675800 155751
rect 675114 154456 675170 154465
rect 675114 154391 675170 154400
rect 674944 152850 675418 152878
rect 674944 150385 674972 152850
rect 675114 152688 675170 152697
rect 675114 152623 675170 152632
rect 675128 152334 675156 152623
rect 675128 152306 675418 152334
rect 675772 151473 675800 151675
rect 675758 151464 675814 151473
rect 675758 151399 675814 151408
rect 675114 151328 675170 151337
rect 675114 151263 675170 151272
rect 675128 151042 675156 151263
rect 675128 151014 675418 151042
rect 674930 150376 674986 150385
rect 674930 150311 674986 150320
rect 675128 149821 675418 149849
rect 675128 147665 675156 149821
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675114 147656 675170 147665
rect 675114 147591 675170 147600
rect 675390 147656 675446 147665
rect 675390 147591 675446 147600
rect 675404 147356 675432 147591
rect 675312 146254 675432 146282
rect 675312 146146 675340 146254
rect 675128 146118 675340 146146
rect 675404 146132 675432 146254
rect 675128 144945 675156 146118
rect 675114 144936 675170 144945
rect 675114 144871 675170 144880
rect 676034 134600 676090 134609
rect 676034 134535 676090 134544
rect 676048 132569 676076 134535
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 676034 132560 676090 132569
rect 676034 132495 676090 132504
rect 674654 131336 674710 131345
rect 674654 131271 674710 131280
rect 674470 130520 674526 130529
rect 674470 130455 674526 130464
rect 676218 130248 676274 130257
rect 676218 130183 676274 130192
rect 675850 128888 675906 128897
rect 675850 128823 675906 128832
rect 675864 128354 675892 128823
rect 674852 128326 675892 128354
rect 674378 125216 674434 125225
rect 674378 125151 674434 125160
rect 674102 117464 674158 117473
rect 674102 117399 674158 117408
rect 673918 106992 673974 107001
rect 673918 106927 673974 106936
rect 674392 104666 674420 125151
rect 674654 123584 674710 123593
rect 674654 123519 674710 123528
rect 674668 105822 674696 123519
rect 674852 113846 674880 128326
rect 676232 127809 676260 130183
rect 676218 127800 676274 127809
rect 676218 127735 676274 127744
rect 676402 127800 676458 127809
rect 676402 127735 676458 127744
rect 676416 120086 676444 127735
rect 682382 126168 682438 126177
rect 682382 126103 682438 126112
rect 681002 125352 681058 125361
rect 681002 125287 681058 125296
rect 675852 120080 675904 120086
rect 675852 120022 675904 120028
rect 676404 120080 676456 120086
rect 676404 120022 676456 120028
rect 675864 118694 675892 120022
rect 675220 118666 675892 118694
rect 675220 115934 675248 118666
rect 681016 117337 681044 125287
rect 681002 117328 681058 117337
rect 681002 117263 681058 117272
rect 682396 116113 682424 126103
rect 683302 125760 683358 125769
rect 683302 125695 683358 125704
rect 683316 120057 683344 125695
rect 683302 120048 683358 120057
rect 683302 119983 683358 119992
rect 682382 116104 682438 116113
rect 682382 116039 682438 116048
rect 675128 115906 675248 115934
rect 675128 115682 675156 115906
rect 675298 115832 675354 115841
rect 675298 115767 675354 115776
rect 675036 115654 675156 115682
rect 675036 115297 675064 115654
rect 675312 115410 675340 115767
rect 675220 115382 675340 115410
rect 675022 115288 675078 115297
rect 675022 115223 675078 115232
rect 675220 114493 675248 115382
rect 675772 115297 675800 115668
rect 675390 115288 675446 115297
rect 675390 115223 675446 115232
rect 675758 115288 675814 115297
rect 675758 115223 675814 115232
rect 675404 115124 675432 115223
rect 675220 114465 675418 114493
rect 674852 113818 675418 113846
rect 675758 112432 675814 112441
rect 675758 112367 675814 112376
rect 675772 111996 675800 112367
rect 675758 111752 675814 111761
rect 675758 111687 675814 111696
rect 675772 111452 675800 111687
rect 675758 111344 675814 111353
rect 675758 111279 675814 111288
rect 675772 110772 675800 111279
rect 675758 110392 675814 110401
rect 675758 110327 675814 110336
rect 675772 110160 675800 110327
rect 675758 108216 675814 108225
rect 675758 108151 675814 108160
rect 675772 107644 675800 108151
rect 675312 107222 675432 107250
rect 675312 107114 675340 107222
rect 675128 107086 675340 107114
rect 675404 107100 675432 107222
rect 675128 106321 675156 107086
rect 675390 106992 675446 107001
rect 675390 106927 675446 106936
rect 675404 106488 675432 106927
rect 675114 106312 675170 106321
rect 675114 106247 675170 106256
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 674668 105794 675340 105822
rect 675404 105808 675432 105862
rect 674392 104638 675340 104666
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 673366 103456 673422 103465
rect 673366 103391 673422 103400
rect 675114 103456 675170 103465
rect 675114 103391 675170 103400
rect 675128 102830 675156 103391
rect 675128 102802 675340 102830
rect 675312 102762 675340 102802
rect 675404 102762 675432 102816
rect 675312 102734 675432 102762
rect 675404 101969 675432 102136
rect 675390 101960 675446 101969
rect 675390 101895 675446 101904
rect 675404 100450 675432 100980
rect 675312 100422 675432 100450
rect 675312 99385 675340 100422
rect 671986 99376 672042 99385
rect 671986 99311 672042 99320
rect 675298 99376 675354 99385
rect 675298 99311 675354 99320
rect 661960 98660 662012 98666
rect 661960 98602 662012 98608
rect 661408 97232 661460 97238
rect 661408 97174 661460 97180
rect 660120 96960 660172 96966
rect 660120 96902 660172 96908
rect 660120 96824 660172 96830
rect 660120 96766 660172 96772
rect 660132 95132 660160 96766
rect 660672 96212 660724 96218
rect 660672 96154 660724 96160
rect 660684 95132 660712 96154
rect 661420 95132 661448 97174
rect 661972 95132 662000 98602
rect 663892 97980 663944 97986
rect 663892 97922 663944 97928
rect 662512 97708 662564 97714
rect 662512 97650 662564 97656
rect 662524 95132 662552 97650
rect 663064 97368 663116 97374
rect 663064 97310 663116 97316
rect 663076 95132 663104 97310
rect 663708 96076 663760 96082
rect 663708 96018 663760 96024
rect 663720 95962 663748 96018
rect 663720 95934 663840 95962
rect 663812 92970 663840 95934
rect 663720 92942 663840 92970
rect 663720 92857 663748 92942
rect 663706 92848 663762 92857
rect 663706 92783 663762 92792
rect 663904 88806 663932 97922
rect 665180 97844 665232 97850
rect 665180 97786 665232 97792
rect 664168 96348 664220 96354
rect 664168 96290 664220 96296
rect 664180 89865 664208 96290
rect 664352 95668 664404 95674
rect 664352 95610 664404 95616
rect 664166 89856 664222 89865
rect 664166 89791 664222 89800
rect 664364 89049 664392 95610
rect 665192 93401 665220 97786
rect 665548 96484 665600 96490
rect 665548 96426 665600 96432
rect 665364 95940 665416 95946
rect 665364 95882 665416 95888
rect 665178 93392 665234 93401
rect 665178 93327 665234 93336
rect 665376 91769 665404 95882
rect 665362 91760 665418 91769
rect 665362 91695 665418 91704
rect 665560 90681 665588 96426
rect 665546 90672 665602 90681
rect 665546 90607 665602 90616
rect 664350 89040 664406 89049
rect 664350 88975 664406 88984
rect 658556 88800 658608 88806
rect 662328 88800 662380 88806
rect 658608 88748 658858 88754
rect 658556 88742 658858 88748
rect 658568 88726 658858 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 663892 88800 663944 88806
rect 663892 88742 663944 88748
rect 661986 88726 662368 88742
rect 657452 88664 657504 88670
rect 657504 88612 657754 88618
rect 657452 88606 657754 88612
rect 657464 88590 657754 88606
rect 658306 88330 658504 88346
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 658464 88266 658516 88272
rect 656716 86896 656768 86902
rect 656716 86838 656768 86844
rect 656164 86488 656216 86494
rect 656164 86430 656216 86436
rect 657188 86358 657216 88196
rect 659580 86902 659608 88196
rect 659568 86896 659620 86902
rect 659568 86838 659620 86844
rect 660132 86630 660160 88196
rect 660120 86624 660172 86630
rect 660120 86566 660172 86572
rect 660684 86494 660712 88196
rect 661420 86766 661448 88196
rect 662524 87038 662552 88196
rect 662512 87032 662564 87038
rect 662512 86974 662564 86980
rect 661408 86760 661460 86766
rect 661408 86702 661460 86708
rect 660672 86488 660724 86494
rect 660672 86430 660724 86436
rect 652024 86352 652076 86358
rect 652024 86294 652076 86300
rect 657176 86352 657228 86358
rect 657176 86294 657228 86300
rect 650550 84688 650606 84697
rect 650550 84623 650606 84632
rect 650366 82240 650422 82249
rect 650366 82175 650422 82184
rect 662420 76560 662472 76566
rect 662420 76502 662472 76508
rect 648802 57352 648858 57361
rect 648802 57287 648858 57296
rect 625804 54528 625856 54534
rect 625804 54470 625856 54476
rect 596180 54392 596232 54398
rect 596180 54334 596232 54340
rect 592684 51740 592736 51746
rect 592684 51682 592736 51688
rect 661590 48510 661646 48519
rect 661590 48445 661646 48454
rect 553674 48104 553730 48113
rect 553674 48039 553730 48048
rect 552018 47832 552074 47841
rect 552018 47767 552074 47776
rect 547878 47560 547934 47569
rect 547878 47495 547934 47504
rect 545670 47288 545726 47297
rect 545670 47223 545726 47232
rect 465262 46744 465318 46753
rect 465262 46679 465318 46688
rect 661604 45554 661632 48445
rect 662432 47433 662460 76502
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 661420 45526 661632 45554
rect 464710 44296 464766 44305
rect 464710 44231 464766 44240
rect 471058 43480 471114 43489
rect 471058 43415 471114 43424
rect 465814 43208 465870 43217
rect 465814 43143 465870 43152
rect 464160 42764 464212 42770
rect 464160 42706 464212 42712
rect 463056 42492 463108 42498
rect 463988 42486 464050 42514
rect 463056 42434 463108 42440
rect 460938 42392 460994 42401
rect 460938 42327 460994 42336
rect 464022 42228 464050 42486
rect 465828 42364 465856 43143
rect 471072 42106 471100 43415
rect 518806 42800 518862 42809
rect 518806 42735 518862 42744
rect 518820 42228 518848 42735
rect 661420 42187 661448 45526
rect 661408 42181 661460 42187
rect 515402 42120 515458 42129
rect 459940 42078 460368 42106
rect 471072 42078 471408 42106
rect 515154 42078 515402 42106
rect 520922 42120 520978 42129
rect 520674 42078 520922 42106
rect 515402 42055 515458 42064
rect 522026 42120 522082 42129
rect 521870 42078 522026 42106
rect 520922 42055 520978 42064
rect 526442 42120 526498 42129
rect 526194 42078 526442 42106
rect 522026 42055 522082 42064
rect 529570 42120 529626 42129
rect 661408 42123 661460 42129
rect 529322 42078 529570 42106
rect 526442 42055 526498 42064
rect 529570 42055 529626 42064
rect 404452 41472 404504 41478
rect 404452 41414 404504 41420
rect 420736 41472 420788 41478
rect 420736 41414 420788 41420
rect 426900 41472 426952 41478
rect 426900 41414 426952 41420
rect 459192 41472 459244 41478
rect 459192 41414 459244 41420
rect 141698 40352 141754 40361
rect 141698 40287 141754 40296
rect 141712 39984 141740 40287
<< via2 >>
rect 676034 897116 676090 897152
rect 676034 897096 676036 897116
rect 676036 897096 676088 897116
rect 676088 897096 676090 897116
rect 651470 868536 651526 868592
rect 675850 896688 675906 896744
rect 676034 896280 676090 896336
rect 652022 867584 652078 867640
rect 651470 866224 651526 866280
rect 651378 865172 651380 865192
rect 651380 865172 651432 865192
rect 651432 865172 651434 865192
rect 651378 865136 651434 865172
rect 651470 863812 651472 863832
rect 651472 863812 651524 863832
rect 651524 863812 651526 863832
rect 651470 863776 651526 863812
rect 651470 862280 651526 862336
rect 35622 817944 35678 818000
rect 35806 817264 35862 817320
rect 35438 816856 35494 816912
rect 35806 816040 35862 816096
rect 35622 815224 35678 815280
rect 35806 814408 35862 814464
rect 41326 813592 41382 813648
rect 40958 812776 41014 812832
rect 32402 811552 32458 811608
rect 31022 809920 31078 809976
rect 41142 812368 41198 812424
rect 34518 811144 34574 811200
rect 33782 809512 33838 809568
rect 40958 808696 41014 808752
rect 41970 810736 42026 810792
rect 41786 809104 41842 809160
rect 41142 807880 41198 807936
rect 41142 806656 41198 806712
rect 41326 806248 41382 806304
rect 40958 805160 41014 805216
rect 42154 810328 42210 810384
rect 41970 805568 42026 805624
rect 42154 804888 42210 804944
rect 41602 804616 41658 804672
rect 40682 800536 40738 800592
rect 41786 800264 41842 800320
rect 41786 799856 41842 799912
rect 41786 794416 41842 794472
rect 42430 793464 42486 793520
rect 42246 791968 42302 792024
rect 42522 789520 42578 789576
rect 42246 788840 42302 788896
rect 41878 788568 41934 788624
rect 42614 789248 42670 789304
rect 43258 808288 43314 808344
rect 43810 807472 43866 807528
rect 35806 774696 35862 774752
rect 35346 773880 35402 773936
rect 35530 773472 35586 773528
rect 35806 773472 35862 773528
rect 41694 773472 41750 773528
rect 35806 773100 35808 773120
rect 35808 773100 35860 773120
rect 35860 773100 35862 773120
rect 35806 773064 35862 773100
rect 40774 773100 40776 773120
rect 40776 773100 40828 773120
rect 40828 773100 40830 773120
rect 40774 773064 40830 773100
rect 35806 772248 35862 772304
rect 35622 771840 35678 771896
rect 42982 773064 43038 773120
rect 40222 771860 40278 771896
rect 40222 771840 40224 771860
rect 40224 771840 40276 771860
rect 40276 771840 40278 771860
rect 42798 771840 42854 771896
rect 35806 771452 35862 771488
rect 35806 771432 35808 771452
rect 35808 771432 35860 771452
rect 35860 771432 35862 771452
rect 41050 771432 41106 771488
rect 35806 771024 35862 771080
rect 41510 771024 41566 771080
rect 35622 770616 35678 770672
rect 35806 770208 35862 770264
rect 39854 770208 39910 770264
rect 35806 769392 35862 769448
rect 35530 768984 35586 769040
rect 35806 768984 35862 769040
rect 35162 768168 35218 768224
rect 32402 767760 32458 767816
rect 33782 766944 33838 767000
rect 35806 767372 35862 767408
rect 35806 767352 35808 767372
rect 35808 767352 35860 767372
rect 35860 767352 35862 767372
rect 35806 766536 35862 766592
rect 35806 765720 35862 765776
rect 35806 764532 35808 764552
rect 35808 764532 35860 764552
rect 35860 764532 35862 764552
rect 35806 764496 35862 764532
rect 35622 764088 35678 764144
rect 35806 763680 35862 763736
rect 35806 762864 35862 762920
rect 39762 765720 39818 765776
rect 41234 767352 41290 767408
rect 39394 764496 39450 764552
rect 41694 763680 41750 763736
rect 40958 763272 41014 763328
rect 41694 762864 41750 762920
rect 36542 757696 36598 757752
rect 39210 757288 39266 757344
rect 41786 757016 41842 757072
rect 41878 756608 41934 756664
rect 42430 762864 42486 762920
rect 42338 755792 42394 755848
rect 42062 754024 42118 754080
rect 42154 752936 42210 752992
rect 42062 751712 42118 751768
rect 42154 751168 42210 751224
rect 42154 750896 42210 750952
rect 42062 749128 42118 749184
rect 41786 746816 41842 746872
rect 42798 754976 42854 755032
rect 42062 746000 42118 746056
rect 42706 746000 42762 746056
rect 42430 745320 42486 745376
rect 42246 744776 42302 744832
rect 42614 745048 42670 745104
rect 42246 730496 42302 730552
rect 40958 729680 41014 729736
rect 43442 771432 43498 771488
rect 43258 763272 43314 763328
rect 42982 730088 43038 730144
rect 41142 729272 41198 729328
rect 42890 728864 42946 728920
rect 40866 728626 40922 728682
rect 41326 727402 41382 727458
rect 41142 726824 41198 726880
rect 40958 726178 41014 726234
rect 40774 725600 40830 725656
rect 32402 725192 32458 725248
rect 31666 723968 31722 724024
rect 35162 724784 35218 724840
rect 37278 724376 37334 724432
rect 39302 723152 39358 723208
rect 37278 716896 37334 716952
rect 41326 726232 41382 726234
rect 41326 726180 41328 726232
rect 41328 726180 41380 726232
rect 41380 726180 41382 726232
rect 41326 726178 41382 726180
rect 41786 725736 41842 725792
rect 41786 723016 41842 723072
rect 41786 722336 41842 722392
rect 40774 719208 40830 719264
rect 41970 721928 42026 721984
rect 41786 718528 41842 718584
rect 41970 718256 42026 718312
rect 40406 714856 40462 714912
rect 38014 714448 38070 714504
rect 42706 719208 42762 719264
rect 42154 714856 42210 714912
rect 42154 714176 42210 714232
rect 41786 713904 41842 713960
rect 42154 713496 42210 713552
rect 42706 714812 42762 714868
rect 42246 710368 42302 710424
rect 42246 709144 42302 709200
rect 42062 708872 42118 708928
rect 42062 708328 42118 708384
rect 41970 707376 42026 707432
rect 42706 709960 42762 710016
rect 42430 706152 42486 706208
rect 41970 704248 42026 704304
rect 42246 701800 42302 701856
rect 41786 700440 41842 700496
rect 42522 701528 42578 701584
rect 41142 686840 41198 686896
rect 40958 686432 41014 686488
rect 40774 685854 40830 685910
rect 41326 685854 41382 685910
rect 35162 681944 35218 682000
rect 33046 681536 33102 681592
rect 33782 681128 33838 681184
rect 36542 680720 36598 680776
rect 33782 672696 33838 672752
rect 42982 684120 43038 684176
rect 41326 683460 41382 683462
rect 41326 683408 41328 683460
rect 41328 683408 41380 683460
rect 41380 683408 41382 683460
rect 41326 683406 41382 683408
rect 40958 682760 41014 682816
rect 42614 682352 42670 682408
rect 41786 678816 41842 678872
rect 41694 678580 41696 678600
rect 41696 678580 41748 678600
rect 41748 678580 41750 678600
rect 41694 678544 41750 678580
rect 41786 678272 41842 678328
rect 40774 677748 40830 677750
rect 40774 677696 40776 677748
rect 40776 677696 40828 677748
rect 40828 677696 40830 677748
rect 40774 677694 40830 677696
rect 41602 671064 41658 671120
rect 40498 670964 40500 670984
rect 40500 670964 40552 670984
rect 40552 670964 40554 670984
rect 40498 670928 40554 670964
rect 41418 670928 41474 670984
rect 41786 670248 41842 670304
rect 42430 677048 42486 677104
rect 42798 679904 42854 679960
rect 42798 671472 42854 671528
rect 42798 671064 42854 671120
rect 42338 667392 42394 667448
rect 42154 666576 42210 666632
rect 42062 665352 42118 665408
rect 41786 665080 41842 665136
rect 42062 664536 42118 664592
rect 41786 658280 41842 658336
rect 41786 657192 41842 657248
rect 42522 658552 42578 658608
rect 35806 644680 35862 644736
rect 38566 644272 38622 644328
rect 35346 643864 35402 643920
rect 35530 643456 35586 643512
rect 35806 643492 35808 643512
rect 35808 643492 35860 643512
rect 35860 643492 35862 643512
rect 35806 643456 35862 643492
rect 35438 642640 35494 642696
rect 35806 642640 35862 642696
rect 35622 642232 35678 642288
rect 39946 642232 40002 642288
rect 35346 641416 35402 641472
rect 40130 641416 40186 641472
rect 35530 641008 35586 641064
rect 35806 641008 35862 641064
rect 39946 640192 40002 640248
rect 40590 641008 40646 641064
rect 34426 639784 34482 639840
rect 40314 639784 40370 639840
rect 35806 639376 35862 639432
rect 35806 638988 35862 639024
rect 35806 638968 35808 638988
rect 35808 638968 35860 638988
rect 35860 638968 35862 638988
rect 35622 638560 35678 638616
rect 32402 637744 32458 637800
rect 35162 637336 35218 637392
rect 32402 629856 32458 629912
rect 35806 638152 35862 638208
rect 35806 636928 35862 636984
rect 35530 636520 35586 636576
rect 35806 636520 35862 636576
rect 35806 635704 35862 635760
rect 35806 634480 35862 634536
rect 35806 633664 35862 633720
rect 39118 636148 39120 636168
rect 39120 636148 39172 636168
rect 39172 636148 39174 636168
rect 39118 636112 39174 636148
rect 39762 633700 39764 633720
rect 39764 633700 39816 633720
rect 39816 633700 39818 633720
rect 39762 633664 39818 633700
rect 40498 635704 40554 635760
rect 40314 634480 40370 634536
rect 41510 633256 41566 633312
rect 40866 632304 40922 632360
rect 42706 634480 42762 634536
rect 42062 633256 42118 633312
rect 40498 630536 40554 630592
rect 40038 630264 40094 630320
rect 39302 629176 39358 629232
rect 40498 628360 40554 628416
rect 42522 630264 42578 630320
rect 42338 628360 42394 628416
rect 41786 627408 41842 627464
rect 41786 627136 41842 627192
rect 41786 621968 41842 622024
rect 41786 620744 41842 620800
rect 43074 632304 43130 632360
rect 42890 630536 42946 630592
rect 41878 615984 41934 616040
rect 42062 615848 42118 615904
rect 42706 615848 42762 615904
rect 42614 615440 42670 615496
rect 41878 613400 41934 613456
rect 42246 612348 42248 612368
rect 42248 612348 42300 612368
rect 42300 612348 42302 612368
rect 42246 612312 42302 612348
rect 43626 752936 43682 752992
rect 43626 731312 43682 731368
rect 43442 723560 43498 723616
rect 43626 720296 43682 720352
rect 43626 707376 43682 707432
rect 43442 688064 43498 688120
rect 43442 687248 43498 687304
rect 43626 680312 43682 680368
rect 43442 677864 43498 677920
rect 43626 633664 43682 633720
rect 43258 612176 43314 612232
rect 46202 773472 46258 773528
rect 44454 771024 44510 771080
rect 44270 770208 44326 770264
rect 43994 751168 44050 751224
rect 44178 728048 44234 728104
rect 45006 765720 45062 765776
rect 45190 764496 45246 764552
rect 44730 754024 44786 754080
rect 44822 751712 44878 751768
rect 45374 763680 45430 763736
rect 45190 750896 45246 750952
rect 46202 730904 46258 730960
rect 44546 727640 44602 727696
rect 44178 721520 44234 721576
rect 44178 708872 44234 708928
rect 43994 708328 44050 708384
rect 44362 685208 44418 685264
rect 44362 684800 44418 684856
rect 44178 679496 44234 679552
rect 43994 679088 44050 679144
rect 44178 664536 44234 664592
rect 45282 722744 45338 722800
rect 44914 721112 44970 721168
rect 44638 684392 44694 684448
rect 44546 641008 44602 641064
rect 44362 636112 44418 636168
rect 43994 635704 44050 635760
rect 43873 612176 43929 612232
rect 44270 611668 44272 611688
rect 44272 611668 44324 611688
rect 44324 611668 44326 611688
rect 44270 611632 44326 611668
rect 44086 611360 44142 611416
rect 40314 601976 40370 602032
rect 35806 601724 35862 601760
rect 35806 601704 35808 601724
rect 35808 601704 35860 601724
rect 35860 601704 35862 601724
rect 35162 595754 35218 595810
rect 33046 595176 33102 595232
rect 31022 594360 31078 594416
rect 33782 593544 33838 593600
rect 35622 591912 35678 591968
rect 35806 591504 35862 591560
rect 39946 601296 40002 601352
rect 37922 594768 37978 594824
rect 36542 589600 36598 589656
rect 40130 600888 40186 600944
rect 45466 687656 45522 687712
rect 45282 678544 45338 678600
rect 45282 642232 45338 642288
rect 46202 641416 46258 641472
rect 45282 640192 45338 640248
rect 45098 639784 45154 639840
rect 44546 600480 44602 600536
rect 44638 600072 44694 600128
rect 43074 597624 43130 597680
rect 42798 596944 42854 597000
rect 42430 596808 42486 596864
rect 40958 596162 41014 596218
rect 41326 595754 41382 595810
rect 41694 595756 41696 595776
rect 41696 595756 41748 595776
rect 41748 595756 41750 595776
rect 41694 595720 41750 595756
rect 41786 594224 41842 594280
rect 41694 592048 41750 592104
rect 39670 589328 39726 589384
rect 39394 586084 39450 586120
rect 39394 586064 39396 586084
rect 39396 586064 39448 586084
rect 39448 586064 39450 586084
rect 37922 585112 37978 585168
rect 39210 584840 39266 584896
rect 40406 585656 40462 585712
rect 39762 584568 39818 584624
rect 42706 586064 42762 586120
rect 41786 580216 41842 580272
rect 42246 580216 42302 580272
rect 42430 579944 42486 580000
rect 42430 579400 42486 579456
rect 42338 579128 42394 579184
rect 42338 578312 42394 578368
rect 42062 578040 42118 578096
rect 41786 577768 41842 577824
rect 41786 574640 41842 574696
rect 42614 573960 42670 574016
rect 41786 573416 41842 573472
rect 42154 573416 42210 573472
rect 42062 572600 42118 572656
rect 42062 571512 42118 571568
rect 42430 571376 42486 571432
rect 41786 570152 41842 570208
rect 40958 558048 41014 558104
rect 37922 553352 37978 553408
rect 29642 551928 29698 551984
rect 42798 555600 42854 555656
rect 44362 593136 44418 593192
rect 43442 589328 43498 589384
rect 43074 554784 43130 554840
rect 43166 554376 43222 554432
rect 40774 549888 40830 549944
rect 41326 553352 41382 553408
rect 41326 552336 41382 552392
rect 41694 551792 41750 551848
rect 42982 551112 43038 551168
rect 42154 550160 42210 550216
rect 42798 549072 42854 549128
rect 41326 548256 41382 548312
rect 41694 547712 41750 547768
rect 41142 545808 41198 545864
rect 40774 545536 40830 545592
rect 42338 545808 42394 545864
rect 37922 542272 37978 542328
rect 42614 539552 42670 539608
rect 42430 538192 42486 538248
rect 42062 537376 42118 537432
rect 42062 536968 42118 537024
rect 42614 536968 42670 537024
rect 42062 535608 42118 535664
rect 41786 535200 41842 535256
rect 42706 536696 42762 536752
rect 42706 535608 42762 535664
rect 42430 533840 42486 533896
rect 42246 533296 42302 533352
rect 42706 532752 42762 532808
rect 42430 531664 42486 531720
rect 42614 530712 42670 530768
rect 42798 529760 42854 529816
rect 42430 528944 42486 529000
rect 42614 526768 42670 526824
rect 35806 430072 35862 430128
rect 35806 428440 35862 428496
rect 43166 427352 43222 427408
rect 42154 427080 42210 427136
rect 41142 426400 41198 426456
rect 41970 426400 42026 426456
rect 42798 426400 42854 426456
rect 40958 425992 41014 426048
rect 39302 425584 39358 425640
rect 32034 424768 32090 424824
rect 34518 424360 34574 424416
rect 33782 423952 33838 424008
rect 41142 423544 41198 423600
rect 41786 423544 41842 423600
rect 41786 422320 41842 422376
rect 41786 421912 41842 421968
rect 41786 421504 41842 421560
rect 41602 418648 41658 418704
rect 41786 418376 41842 418432
rect 39302 415248 39358 415304
rect 33782 414568 33838 414624
rect 42062 408040 42118 408096
rect 42430 407224 42486 407280
rect 41786 406952 41842 407008
rect 41786 406680 41842 406736
rect 42430 404912 42486 404968
rect 42246 404504 42302 404560
rect 42338 402872 42394 402928
rect 42246 402464 42302 402520
rect 41786 400016 41842 400072
rect 41786 399336 41842 399392
rect 41970 398792 42026 398848
rect 42154 395664 42210 395720
rect 41326 387096 41382 387152
rect 41142 386688 41198 386744
rect 40958 385872 41014 385928
rect 41142 385872 41198 385928
rect 41142 383016 41198 383072
rect 40038 382200 40094 382256
rect 40958 382200 41014 382256
rect 35438 381792 35494 381848
rect 33966 380976 34022 381032
rect 39302 381384 39358 381440
rect 35806 379344 35862 379400
rect 35806 378156 35808 378176
rect 35808 378156 35860 378176
rect 35860 378156 35862 378176
rect 35806 378120 35862 378156
rect 35806 376488 35862 376544
rect 35806 376080 35862 376136
rect 35438 374584 35494 374640
rect 41326 382608 41382 382664
rect 41142 381792 41198 381848
rect 41326 379772 41382 379808
rect 41326 379752 41328 379772
rect 41328 379752 41380 379772
rect 41380 379752 41382 379772
rect 41510 379772 41566 379808
rect 41510 379752 41512 379772
rect 41512 379752 41564 379772
rect 41564 379752 41566 379772
rect 40038 379344 40094 379400
rect 42982 425176 43038 425232
rect 43166 422728 43222 422784
rect 42798 385600 42854 385656
rect 43258 385192 43314 385248
rect 41878 381520 41934 381576
rect 42890 380704 42946 380760
rect 41694 378156 41696 378176
rect 41696 378156 41748 378176
rect 41748 378156 41750 378176
rect 41694 378120 41750 378156
rect 40406 376896 40462 376952
rect 41786 364792 41842 364848
rect 41786 364112 41842 364168
rect 42154 363568 42210 363624
rect 42706 363024 42762 363080
rect 42706 362208 42762 362264
rect 41786 360032 41842 360088
rect 42154 359896 42210 359952
rect 42430 358944 42486 359000
rect 41878 358672 41934 358728
rect 41786 356904 41842 356960
rect 43074 376896 43130 376952
rect 42430 355952 42486 356008
rect 41878 355680 41934 355736
rect 44362 578040 44418 578096
rect 45098 599664 45154 599720
rect 44914 599256 44970 599312
rect 44638 558728 44694 558784
rect 46202 611632 46258 611688
rect 45466 598848 45522 598904
rect 45282 598032 45338 598088
rect 45098 580216 45154 580272
rect 45098 556824 45154 556880
rect 44914 556416 44970 556472
rect 44638 556008 44694 556064
rect 44362 555192 44418 555248
rect 43994 551792 44050 551848
rect 43810 550704 43866 550760
rect 43626 547712 43682 547768
rect 43442 354728 43498 354784
rect 44178 548664 44234 548720
rect 44178 536832 44234 536888
rect 43994 533840 44050 533896
rect 43810 532752 43866 532808
rect 44822 550432 44878 550488
rect 45282 551520 45338 551576
rect 44822 539552 44878 539608
rect 44822 537376 44878 537432
rect 45282 529760 45338 529816
rect 45190 527176 45246 527232
rect 45282 430888 45338 430944
rect 45006 429664 45062 429720
rect 45098 429256 45154 429312
rect 44638 428848 44694 428904
rect 44362 428032 44418 428088
rect 44362 427624 44418 427680
rect 44178 426808 44234 426864
rect 43810 422320 43866 422376
rect 43994 421096 44050 421152
rect 43994 408040 44050 408096
rect 43810 402464 43866 402520
rect 44546 423136 44602 423192
rect 44730 407224 44786 407280
rect 45466 420688 45522 420744
rect 44546 402872 44602 402928
rect 45098 386416 45154 386472
rect 44362 384784 44418 384840
rect 45190 384376 45246 384432
rect 44178 383968 44234 384024
rect 45098 383560 45154 383616
rect 44914 382200 44970 382256
rect 44638 380296 44694 380352
rect 43810 379752 43866 379808
rect 43994 378120 44050 378176
rect 44270 377440 44326 377496
rect 43994 363568 44050 363624
rect 43810 359896 43866 359952
rect 43626 354048 43682 354104
rect 44638 363024 44694 363080
rect 44454 358944 44510 359000
rect 44638 355952 44694 356008
rect 44454 354728 44510 354784
rect 44638 354492 44640 354512
rect 44640 354492 44692 354512
rect 44692 354492 44694 354512
rect 44638 354456 44694 354492
rect 44178 353096 44234 353152
rect 40222 345480 40278 345536
rect 43258 345480 43314 345536
rect 35530 344256 35586 344312
rect 35806 344256 35862 344312
rect 40038 344256 40094 344312
rect 33046 343440 33102 343496
rect 35806 342252 35808 342272
rect 35808 342252 35860 342272
rect 35860 342252 35862 342272
rect 35806 342216 35862 342252
rect 44914 343304 44970 343360
rect 40038 341808 40094 341864
rect 35622 341400 35678 341456
rect 40222 341420 40278 341456
rect 40222 341400 40224 341420
rect 40224 341400 40276 341420
rect 40276 341400 40278 341420
rect 35806 340992 35862 341048
rect 39854 340992 39910 341048
rect 45466 354320 45522 354376
rect 45466 354084 45468 354104
rect 45468 354084 45520 354104
rect 45520 354084 45522 354104
rect 45466 354048 45522 354084
rect 45466 353368 45522 353424
rect 45420 353132 45422 353152
rect 45422 353132 45474 353152
rect 45474 353132 45476 353152
rect 45420 353096 45476 353132
rect 40222 340992 40278 341048
rect 45098 340992 45154 341048
rect 45466 341420 45522 341456
rect 45466 341400 45468 341420
rect 45468 341400 45520 341420
rect 45520 341400 45522 341420
rect 40038 340584 40094 340640
rect 45282 340584 45338 340640
rect 35530 339768 35586 339824
rect 35806 339768 35862 339824
rect 39854 339768 39910 339824
rect 35162 338544 35218 338600
rect 35806 336096 35862 336152
rect 35622 334872 35678 334928
rect 35806 334464 35862 334520
rect 45650 338408 45706 338464
rect 45466 336776 45522 336832
rect 38842 336504 38898 336560
rect 43994 334600 44050 334656
rect 40222 334464 40278 334520
rect 43166 334464 43222 334520
rect 36542 332832 36598 332888
rect 39394 332424 39450 332480
rect 42798 332424 42854 332480
rect 35162 331744 35218 331800
rect 41786 324808 41842 324864
rect 42246 324264 42302 324320
rect 41786 321136 41842 321192
rect 42062 321136 42118 321192
rect 42430 320728 42486 320784
rect 42982 321136 43038 321192
rect 42614 319368 42670 319424
rect 42430 319096 42486 319152
rect 41786 317328 41842 317384
rect 41786 315968 41842 316024
rect 41786 315560 41842 315616
rect 42430 314608 42486 314664
rect 41786 313656 41842 313712
rect 42430 312704 42486 312760
rect 42062 310392 42118 310448
rect 42430 310120 42486 310176
rect 41142 300464 41198 300520
rect 42890 299648 42946 299704
rect 41970 297336 42026 297392
rect 41326 296384 41382 296440
rect 40958 295976 41014 296032
rect 39302 295568 39358 295624
rect 33782 294752 33838 294808
rect 37922 294344 37978 294400
rect 41142 295160 41198 295216
rect 42706 292712 42762 292768
rect 41786 292168 41842 292224
rect 41234 291488 41290 291544
rect 41970 291216 42026 291272
rect 41786 290264 41842 290320
rect 41786 289176 41842 289232
rect 37922 284280 37978 284336
rect 42522 284824 42578 284880
rect 41786 282240 41842 282296
rect 42154 281696 42210 281752
rect 42154 280200 42210 280256
rect 42154 279656 42210 279712
rect 42062 278432 42118 278488
rect 42154 277888 42210 277944
rect 41786 277072 41842 277128
rect 41786 274216 41842 274272
rect 42154 272992 42210 273048
rect 43166 293936 43222 293992
rect 42798 277888 42854 277944
rect 42798 275848 42854 275904
rect 43442 293120 43498 293176
rect 41786 270408 41842 270464
rect 41786 269728 41842 269784
rect 41970 269048 42026 269104
rect 42154 266192 42210 266248
rect 43626 291216 43682 291272
rect 43442 279656 43498 279712
rect 43626 278432 43682 278488
rect 43442 273808 43498 273864
rect 35622 257080 35678 257136
rect 39486 257080 39542 257136
rect 42798 257080 42854 257136
rect 35806 256672 35862 256728
rect 35806 256264 35862 256320
rect 35622 253408 35678 253464
rect 40222 253408 40278 253464
rect 42798 253408 42854 253464
rect 35806 253000 35862 253056
rect 35806 252184 35862 252240
rect 35622 250552 35678 250608
rect 35806 250144 35862 250200
rect 35806 247696 35862 247752
rect 34426 246880 34482 246936
rect 40130 245656 40186 245712
rect 39854 244024 39910 244080
rect 40682 240896 40738 240952
rect 42062 240080 42118 240136
rect 42522 238040 42578 238096
rect 41786 236544 41842 236600
rect 42430 235864 42486 235920
rect 41786 234640 41842 234696
rect 42430 234504 42486 234560
rect 42430 232192 42486 232248
rect 42430 231784 42486 231840
rect 42430 229336 42486 229392
rect 41970 228928 42026 228984
rect 42154 226616 42210 226672
rect 42430 225664 42486 225720
rect 41694 224440 41750 224496
rect 35530 217912 35586 217968
rect 35530 214648 35586 214704
rect 35806 214648 35862 214704
rect 42154 223488 42210 223544
rect 43626 245656 43682 245712
rect 43074 240896 43130 240952
rect 43442 244024 43498 244080
rect 44822 334056 44878 334112
rect 44270 298016 44326 298072
rect 44546 297064 44602 297120
rect 44270 255176 44326 255232
rect 44178 254768 44234 254824
rect 43994 230968 44050 231024
rect 43626 229336 43682 229392
rect 35806 213424 35862 213480
rect 39578 213424 39634 213480
rect 42798 213424 42854 213480
rect 35806 210160 35862 210216
rect 35622 209344 35678 209400
rect 40130 209344 40186 209400
rect 42982 209344 43038 209400
rect 35806 208936 35862 208992
rect 40038 208120 40094 208176
rect 35806 207712 35862 207768
rect 39762 207712 39818 207768
rect 40130 206896 40186 206952
rect 42798 206896 42854 206952
rect 35806 206080 35862 206136
rect 35622 204856 35678 204912
rect 40222 204856 40278 204912
rect 35806 204468 35862 204504
rect 35806 204448 35808 204468
rect 35808 204448 35860 204468
rect 35860 204448 35862 204468
rect 41694 204040 41750 204096
rect 35806 203632 35862 203688
rect 41510 203632 41566 203688
rect 37922 198736 37978 198792
rect 42430 197240 42486 197296
rect 41970 195744 42026 195800
rect 41786 195200 41842 195256
rect 42246 194928 42302 194984
rect 41786 193432 41842 193488
rect 42062 191528 42118 191584
rect 42430 190440 42486 190496
rect 42430 187584 42486 187640
rect 42430 186768 42486 186824
rect 41786 186360 41842 186416
rect 41786 185952 41842 186008
rect 43258 204856 43314 204912
rect 42430 182960 42486 183016
rect 42062 179288 42118 179344
rect 44546 254360 44602 254416
rect 44546 251096 44602 251152
rect 44362 249056 44418 249112
rect 44362 231784 44418 231840
rect 44546 226616 44602 226672
rect 44178 212064 44234 212120
rect 44362 208392 44418 208448
rect 43810 207712 43866 207768
rect 43626 203632 43682 203688
rect 44178 207168 44234 207224
rect 43994 204040 44050 204096
rect 43994 191528 44050 191584
rect 44546 205536 44602 205592
rect 44362 197240 44418 197296
rect 44546 190440 44602 190496
rect 44178 186768 44234 186824
rect 43810 182960 43866 183016
rect 45650 319096 45706 319152
rect 45466 314608 45522 314664
rect 45006 298832 45062 298888
rect 45190 293528 45246 293584
rect 45190 272992 45246 273048
rect 46938 579128 46994 579184
rect 47582 558456 47638 558512
rect 46386 547440 46442 547496
rect 47766 430480 47822 430536
rect 47582 419872 47638 419928
rect 46386 376080 46442 376136
rect 46938 339224 46994 339280
rect 47122 338000 47178 338056
rect 47122 324264 47178 324320
rect 46938 310120 46994 310176
rect 47766 387640 47822 387696
rect 47582 290672 47638 290728
rect 46386 258032 46442 258088
rect 45006 255992 45062 256048
rect 45650 255584 45706 255640
rect 45006 248648 45062 248704
rect 45006 234504 45062 234560
rect 46202 253952 46258 254008
rect 45926 252728 45982 252784
rect 45926 225664 45982 225720
rect 45650 212880 45706 212936
rect 46938 251912 46994 251968
rect 46386 248240 46442 248296
rect 46386 235864 46442 235920
rect 47122 251504 47178 251560
rect 47122 240080 47178 240136
rect 46938 232192 46994 232248
rect 46202 211248 46258 211304
rect 46938 208800 46994 208856
rect 46202 204312 46258 204368
rect 46938 187584 46994 187640
rect 47766 179288 47822 179344
rect 49146 290944 49202 291000
rect 62210 790472 62266 790528
rect 62118 789148 62120 789168
rect 62120 789148 62172 789168
rect 62172 789148 62174 789168
rect 62118 789112 62174 789148
rect 62118 787344 62174 787400
rect 61382 786120 61438 786176
rect 62118 784896 62174 784952
rect 51722 538192 51778 538248
rect 51446 404912 51502 404968
rect 51078 395664 51134 395720
rect 51078 362208 51134 362264
rect 51722 354320 51778 354376
rect 51078 310392 51134 310448
rect 50526 278704 50582 278760
rect 62118 746136 62174 746192
rect 62118 744096 62174 744152
rect 62118 743724 62120 743744
rect 62120 743724 62172 743744
rect 62172 743724 62174 743744
rect 62118 743688 62174 743724
rect 62118 742364 62120 742384
rect 62120 742364 62172 742384
rect 62172 742364 62174 742384
rect 62118 742328 62174 742364
rect 53286 301280 53342 301336
rect 53102 276664 53158 276720
rect 51906 266192 51962 266248
rect 50526 247424 50582 247480
rect 51722 223488 51778 223544
rect 62118 704384 62174 704440
rect 62118 703296 62174 703352
rect 61382 699624 61438 699680
rect 62210 697992 62266 698048
rect 57242 275848 57298 275904
rect 55862 264152 55918 264208
rect 62118 660900 62120 660920
rect 62120 660900 62172 660920
rect 62172 660900 62174 660920
rect 62118 660864 62174 660900
rect 62118 659540 62120 659560
rect 62120 659540 62172 659560
rect 62172 659540 62174 659560
rect 62118 659504 62174 659540
rect 62118 658280 62174 658336
rect 61382 656512 61438 656568
rect 62118 655288 62174 655344
rect 62118 616528 62174 616584
rect 62118 614624 62174 614680
rect 61382 613808 61438 613864
rect 62118 612584 62174 612640
rect 60370 319368 60426 319424
rect 60186 278704 60242 278760
rect 60002 278024 60058 278080
rect 60370 256672 60426 256728
rect 62486 594088 62542 594144
rect 62302 590008 62358 590064
rect 62118 574776 62174 574832
rect 62118 573552 62174 573608
rect 62302 569880 62358 569936
rect 62486 568520 62542 568576
rect 62486 550160 62542 550216
rect 62118 531120 62174 531176
rect 62302 530576 62358 530632
rect 62118 528572 62120 528592
rect 62120 528572 62172 528592
rect 62172 528572 62174 528592
rect 62118 528536 62174 528572
rect 62118 527076 62120 527096
rect 62120 527076 62172 527096
rect 62172 527076 62174 527096
rect 62118 527040 62174 527076
rect 62486 525680 62542 525736
rect 62118 404096 62174 404152
rect 62118 402600 62174 402656
rect 62118 400696 62174 400752
rect 62118 399336 62174 399392
rect 62118 398248 62174 398304
rect 62486 381520 62542 381576
rect 62118 360848 62174 360904
rect 62118 359760 62174 359816
rect 62118 357720 62174 357776
rect 62118 355988 62120 356008
rect 62120 355988 62172 356008
rect 62172 355988 62174 356008
rect 62118 355952 62174 355988
rect 62486 354456 62542 354512
rect 62394 341672 62450 341728
rect 62486 332560 62542 332616
rect 62026 320728 62082 320784
rect 62026 317328 62082 317384
rect 62118 315988 62174 316024
rect 62118 315968 62120 315988
rect 62120 315968 62172 315988
rect 62172 315968 62174 315988
rect 62118 314764 62174 314800
rect 62118 314744 62120 314764
rect 62120 314744 62172 314764
rect 62172 314744 62174 314764
rect 62302 314064 62358 314120
rect 62394 312976 62450 313032
rect 62394 297336 62450 297392
rect 62118 295704 62174 295760
rect 62118 294092 62174 294128
rect 62118 294072 62120 294092
rect 62120 294072 62172 294092
rect 62172 294072 62174 294092
rect 62118 292712 62174 292768
rect 62394 292440 62450 292496
rect 62118 290944 62174 291000
rect 62394 288496 62450 288552
rect 62302 287136 62358 287192
rect 62118 284436 62174 284472
rect 62118 284416 62120 284436
rect 62120 284416 62172 284436
rect 62172 284416 62174 284436
rect 62118 283192 62174 283248
rect 62118 282104 62174 282160
rect 62118 280336 62174 280392
rect 62210 273808 62266 273864
rect 62946 787072 63002 787128
rect 651470 778368 651526 778424
rect 652022 777008 652078 777064
rect 651470 776056 651526 776112
rect 651378 775276 651380 775296
rect 651380 775276 651432 775296
rect 651432 775276 651434 775296
rect 651378 775240 651434 775276
rect 651470 774172 651526 774208
rect 651470 774152 651472 774172
rect 651472 774152 651524 774172
rect 651524 774152 651526 774172
rect 651470 773336 651526 773392
rect 62946 747632 63002 747688
rect 63038 741784 63094 741840
rect 651470 734168 651526 734224
rect 652666 732808 652722 732864
rect 651470 731720 651526 731776
rect 651378 731076 651380 731096
rect 651380 731076 651432 731096
rect 651432 731076 651434 731096
rect 651378 731040 651434 731076
rect 651470 729816 651526 729872
rect 651470 728492 651472 728512
rect 651472 728492 651524 728512
rect 651524 728492 651526 728512
rect 651470 728456 651526 728492
rect 62946 701256 63002 701312
rect 63130 700848 63186 700904
rect 651470 689424 651526 689480
rect 651654 688744 651710 688800
rect 651470 687384 651526 687440
rect 651470 686704 651526 686760
rect 651470 685208 651526 685264
rect 652574 684392 652630 684448
rect 62946 657600 63002 657656
rect 651470 643184 651526 643240
rect 652022 641824 652078 641880
rect 651470 640736 651526 640792
rect 651378 640092 651380 640112
rect 651380 640092 651432 640112
rect 651432 640092 651434 640112
rect 651378 640056 651434 640092
rect 651470 638560 651526 638616
rect 651654 638152 651710 638208
rect 63130 618024 63186 618080
rect 62946 612040 63002 612096
rect 64142 611360 64198 611416
rect 63406 595720 63462 595776
rect 63038 590688 63094 590744
rect 62854 585656 62910 585712
rect 58806 217912 58862 217968
rect 62670 224168 62726 224224
rect 63406 571104 63462 571160
rect 63222 556688 63278 556744
rect 63222 527992 63278 528048
rect 63314 427080 63370 427136
rect 63314 400152 63370 400208
rect 63222 385872 63278 385928
rect 63222 357312 63278 357368
rect 63314 341400 63370 341456
rect 63314 311752 63370 311808
rect 63314 299512 63370 299568
rect 63314 289720 63370 289776
rect 63038 285912 63094 285968
rect 63222 280880 63278 280936
rect 62854 223488 62910 223544
rect 651470 597896 651526 597952
rect 651470 596672 651526 596728
rect 651470 595312 651526 595368
rect 651654 595040 651710 595096
rect 651470 594088 651526 594144
rect 651470 592864 651526 592920
rect 651470 553424 651526 553480
rect 651654 552064 651710 552120
rect 651470 551112 651526 551168
rect 651378 550332 651380 550352
rect 651380 550332 651432 550352
rect 651432 550332 651434 550352
rect 651378 550296 651434 550332
rect 651470 549228 651526 549264
rect 651470 549208 651472 549228
rect 651472 549208 651524 549228
rect 651524 549208 651526 549228
rect 651470 548392 651526 548448
rect 64326 353368 64382 353424
rect 461030 272856 461086 272912
rect 460846 272584 460902 272640
rect 461858 272620 461860 272640
rect 461860 272620 461912 272640
rect 461912 272620 461914 272640
rect 461858 272584 461914 272620
rect 464710 272448 464766 272504
rect 466274 272856 466330 272912
rect 470690 272484 470692 272504
rect 470692 272484 470744 272504
rect 470744 272484 470746 272504
rect 470690 272448 470746 272484
rect 470598 271904 470654 271960
rect 478050 271904 478106 271960
rect 479522 272040 479578 272096
rect 480534 272076 480536 272096
rect 480536 272076 480588 272096
rect 480588 272076 480590 272096
rect 480534 272040 480590 272076
rect 501602 271904 501658 271960
rect 504546 271940 504548 271960
rect 504548 271940 504600 271960
rect 504600 271940 504602 271960
rect 504546 271904 504602 271940
rect 509238 269864 509294 269920
rect 509146 269456 509202 269512
rect 509882 269492 509884 269512
rect 509884 269492 509936 269512
rect 509936 269492 509938 269512
rect 509882 269456 509938 269492
rect 516598 269864 516654 269920
rect 530398 270136 530454 270192
rect 534078 270136 534134 270192
rect 536562 272448 536618 272504
rect 539322 273944 539378 274000
rect 538034 269728 538090 269784
rect 545946 273964 546002 274000
rect 545946 273944 545948 273964
rect 545948 273944 546000 273964
rect 546000 273944 546002 273964
rect 541346 269764 541348 269784
rect 541348 269764 541400 269784
rect 541400 269764 541402 269784
rect 541346 269728 541402 269764
rect 547694 272448 547750 272504
rect 547510 272076 547512 272096
rect 547512 272076 547564 272096
rect 547564 272076 547566 272096
rect 547510 272040 547566 272076
rect 547878 272040 547934 272096
rect 554410 262112 554466 262168
rect 554318 259936 554374 259992
rect 553950 257760 554006 257816
rect 554502 255604 554558 255640
rect 554502 255584 554504 255604
rect 554504 255584 554556 255604
rect 554556 255584 554558 255604
rect 554410 253408 554466 253464
rect 554134 251252 554190 251288
rect 554134 251232 554136 251252
rect 554136 251232 554188 251252
rect 554188 251232 554190 251252
rect 554042 249056 554098 249112
rect 553858 246880 553914 246936
rect 553490 244704 553546 244760
rect 553674 242528 553730 242584
rect 553766 236000 553822 236056
rect 63222 224440 63278 224496
rect 140042 229064 140098 229120
rect 136638 227860 136694 227896
rect 136638 227840 136640 227860
rect 136640 227840 136692 227860
rect 136692 227840 136694 227860
rect 137282 223896 137338 223952
rect 138294 221604 138350 221640
rect 138294 221584 138296 221604
rect 138296 221584 138348 221604
rect 138348 221584 138350 221604
rect 140778 221992 140834 222048
rect 141514 227860 141570 227896
rect 141514 227840 141516 227860
rect 141516 227840 141568 227860
rect 141568 227840 141570 227860
rect 143538 229064 143594 229120
rect 141606 226500 141662 226536
rect 141606 226480 141608 226500
rect 141608 226480 141660 226500
rect 141660 226480 141662 226500
rect 142250 226500 142306 226536
rect 142250 226480 142252 226500
rect 142252 226480 142304 226500
rect 142304 226480 142306 226500
rect 141330 221584 141386 221640
rect 142112 225564 142114 225584
rect 142114 225564 142166 225584
rect 142166 225564 142168 225584
rect 142112 225528 142168 225564
rect 142250 223896 142306 223952
rect 142434 223896 142490 223952
rect 141974 222844 141976 222864
rect 141976 222844 142028 222864
rect 142028 222844 142030 222864
rect 141974 222808 142030 222844
rect 142158 222844 142160 222864
rect 142160 222844 142212 222864
rect 142212 222844 142214 222864
rect 142158 222808 142214 222844
rect 141974 221992 142030 222048
rect 142112 220924 142168 220960
rect 142112 220904 142114 220924
rect 142114 220904 142166 220924
rect 142166 220904 142168 220924
rect 144642 230424 144698 230480
rect 144458 229764 144514 229800
rect 144458 229744 144460 229764
rect 144460 229744 144512 229764
rect 144512 229744 144514 229764
rect 145838 229356 145894 229392
rect 145838 229336 145840 229356
rect 145840 229336 145892 229356
rect 145892 229336 145894 229356
rect 146206 227976 146262 228032
rect 145562 221176 145618 221232
rect 145654 220380 145710 220416
rect 145654 220360 145656 220380
rect 145656 220360 145708 220380
rect 145708 220360 145710 220380
rect 147126 227976 147182 228032
rect 147954 229336 148010 229392
rect 147770 225528 147826 225584
rect 146390 221176 146446 221232
rect 148874 225936 148930 225992
rect 148322 220360 148378 220416
rect 150346 230152 150402 230208
rect 151082 230424 151138 230480
rect 151910 230152 151966 230208
rect 150530 229744 150586 229800
rect 151634 229200 151690 229256
rect 151910 225972 151912 225992
rect 151912 225972 151964 225992
rect 151964 225972 151966 225992
rect 151910 225936 151966 225972
rect 151174 220904 151230 220960
rect 151726 225700 151728 225720
rect 151728 225700 151780 225720
rect 151780 225700 151782 225720
rect 151726 225664 151782 225700
rect 151634 224440 151690 224496
rect 151634 223896 151690 223952
rect 154026 229764 154082 229800
rect 154026 229744 154028 229764
rect 154028 229744 154080 229764
rect 154080 229744 154082 229764
rect 153658 229200 153714 229256
rect 153106 228384 153162 228440
rect 152370 224440 152426 224496
rect 154394 228404 154450 228440
rect 154394 228384 154396 228404
rect 154396 228384 154448 228404
rect 154448 228384 154450 228404
rect 155866 227024 155922 227080
rect 157522 225664 157578 225720
rect 158350 220904 158406 220960
rect 160006 228384 160062 228440
rect 160834 229744 160890 229800
rect 161294 229336 161350 229392
rect 161754 229336 161810 229392
rect 161432 228812 161488 228848
rect 161432 228792 161434 228812
rect 161434 228792 161486 228812
rect 161486 228792 161488 228812
rect 161570 228384 161626 228440
rect 161432 227316 161488 227352
rect 161432 227296 161434 227316
rect 161434 227296 161486 227316
rect 161486 227296 161488 227316
rect 161570 227024 161626 227080
rect 161432 221740 161488 221776
rect 161432 221720 161434 221740
rect 161434 221720 161486 221740
rect 161486 221720 161488 221740
rect 161570 220924 161626 220960
rect 161570 220904 161572 220924
rect 161572 220904 161624 220924
rect 161624 220904 161626 220924
rect 164238 228792 164294 228848
rect 166906 227296 166962 227352
rect 166998 221720 167054 221776
rect 169574 227160 169630 227216
rect 168930 219428 168986 219464
rect 170770 227452 170826 227488
rect 170770 227432 170772 227452
rect 170772 227432 170824 227452
rect 170824 227432 170826 227452
rect 168930 219408 168932 219428
rect 168932 219408 168984 219428
rect 168984 219408 168986 219428
rect 169758 219428 169814 219464
rect 169758 219408 169760 219428
rect 169760 219408 169812 219428
rect 169812 219408 169814 219428
rect 171690 227432 171746 227488
rect 171092 227160 171148 227216
rect 171414 221448 171470 221504
rect 171966 221468 172022 221504
rect 171966 221448 171968 221468
rect 171968 221448 172020 221468
rect 172020 221448 172022 221468
rect 173162 228792 173218 228848
rect 175370 227588 175426 227624
rect 175370 227568 175372 227588
rect 175372 227568 175424 227588
rect 175424 227568 175426 227588
rect 171414 218320 171470 218376
rect 171966 218320 172022 218376
rect 176106 228812 176162 228848
rect 176106 228792 176108 228812
rect 176108 228792 176160 228812
rect 176160 228792 176162 228812
rect 175922 227296 175978 227352
rect 176290 221876 176346 221912
rect 176290 221856 176292 221876
rect 176292 221856 176344 221876
rect 176344 221856 176346 221876
rect 177210 227568 177266 227624
rect 176750 227316 176806 227352
rect 176750 227296 176752 227316
rect 176752 227296 176804 227316
rect 176804 227296 176806 227316
rect 179326 224848 179382 224904
rect 177394 221856 177450 221912
rect 177210 220788 177266 220824
rect 177210 220768 177212 220788
rect 177212 220768 177264 220788
rect 177264 220768 177266 220788
rect 181994 224884 181996 224904
rect 181996 224884 182048 224904
rect 182048 224884 182050 224904
rect 181994 224848 182050 224884
rect 180522 218748 180578 218784
rect 180522 218728 180524 218748
rect 180524 218728 180576 218748
rect 180576 218728 180578 218748
rect 182270 218728 182326 218784
rect 185398 229880 185454 229936
rect 186042 229880 186098 229936
rect 185122 220768 185178 220824
rect 185950 220768 186006 220824
rect 193034 228928 193090 228984
rect 190550 220788 190606 220824
rect 190550 220768 190552 220788
rect 190552 220768 190604 220788
rect 190604 220768 190606 220788
rect 195426 228948 195482 228984
rect 195426 228928 195428 228948
rect 195428 228928 195480 228948
rect 195480 228928 195482 228948
rect 194874 219292 194930 219328
rect 194874 219272 194876 219292
rect 194876 219272 194928 219292
rect 194928 219272 194930 219292
rect 197818 219272 197874 219328
rect 486974 220224 487030 220280
rect 487802 218048 487858 218104
rect 488814 217096 488870 217152
rect 492954 219680 493010 219736
rect 493690 219680 493746 219736
rect 494702 218320 494758 218376
rect 495162 217096 495218 217152
rect 502246 217232 502302 217288
rect 510986 217504 511042 217560
rect 513562 221448 513618 221504
rect 515770 221176 515826 221232
rect 515126 219952 515182 220008
rect 520186 219408 520242 219464
rect 520002 217504 520058 217560
rect 522670 220904 522726 220960
rect 531502 217504 531558 217560
rect 533250 221992 533306 222048
rect 532514 217504 532570 217560
rect 535734 221720 535790 221776
rect 538494 221992 538550 222048
rect 538678 221720 538734 221776
rect 543738 224440 543794 224496
rect 544290 224476 544292 224496
rect 544292 224476 544344 224496
rect 544344 224476 544346 224496
rect 544290 224440 544346 224476
rect 545762 221720 545818 221776
rect 549258 221740 549314 221776
rect 549258 221720 549260 221740
rect 549260 221720 549312 221740
rect 549312 221720 549314 221740
rect 554502 240352 554558 240408
rect 554318 238176 554374 238232
rect 554410 233824 554466 233880
rect 554870 224440 554926 224496
rect 556066 224440 556122 224496
rect 553306 221720 553362 221776
rect 556802 221992 556858 222048
rect 557630 224712 557686 224768
rect 557630 224440 557686 224496
rect 557538 221992 557594 222048
rect 557170 221720 557226 221776
rect 559378 222028 559380 222048
rect 559380 222028 559432 222048
rect 559432 222028 559434 222048
rect 559378 221992 559434 222028
rect 561954 224712 562010 224768
rect 562138 224748 562140 224768
rect 562140 224748 562192 224768
rect 562192 224748 562194 224768
rect 562138 224712 562194 224748
rect 563702 224712 563758 224768
rect 561494 221992 561550 222048
rect 561310 217776 561366 217832
rect 560758 217504 560814 217560
rect 560942 217504 560998 217560
rect 561770 220496 561826 220552
rect 562046 219136 562102 219192
rect 561770 218728 561826 218784
rect 563702 221720 563758 221776
rect 563058 220652 563114 220688
rect 563058 220632 563060 220652
rect 563060 220632 563112 220652
rect 563112 220632 563114 220652
rect 562598 219136 562654 219192
rect 563058 218592 563114 218648
rect 563334 217504 563390 217560
rect 565634 220496 565690 220552
rect 564806 219000 564862 219056
rect 564162 218612 564218 218648
rect 564162 218592 564164 218612
rect 564164 218592 564216 218612
rect 564216 218592 564218 218612
rect 566462 218728 566518 218784
rect 571982 217504 572038 217560
rect 572626 221720 572682 221776
rect 574742 220496 574798 220552
rect 572672 219020 572728 219056
rect 572672 219000 572674 219020
rect 572674 219000 572726 219020
rect 572726 219000 572728 219020
rect 572350 218592 572406 218648
rect 574374 218592 574430 218648
rect 574190 217504 574246 217560
rect 52458 215056 52514 215112
rect 53286 215056 53342 215112
rect 574742 217776 574798 217832
rect 575478 216688 575534 216744
rect 52458 214240 52514 214296
rect 591486 224168 591542 224224
rect 582378 220632 582434 220688
rect 587530 220652 587586 220688
rect 587530 220632 587532 220652
rect 587532 220632 587584 220652
rect 587584 220632 587586 220652
rect 578882 213968 578938 214024
rect 578514 211656 578570 211712
rect 579526 209788 579528 209808
rect 579528 209788 579580 209808
rect 579580 209788 579582 209808
rect 579526 209752 579582 209788
rect 579526 207440 579582 207496
rect 579526 205828 579582 205864
rect 579526 205808 579528 205828
rect 579528 205808 579580 205828
rect 579580 205808 579582 205828
rect 578330 203224 578386 203280
rect 578790 200776 578846 200832
rect 579526 198872 579582 198928
rect 578514 196424 578570 196480
rect 579526 194928 579582 194984
rect 579526 192208 579582 192264
rect 579526 190712 579582 190768
rect 579526 187992 579582 188048
rect 579526 186260 579528 186280
rect 579528 186260 579580 186280
rect 579580 186260 579582 186280
rect 579526 186224 579582 186260
rect 579526 184320 579582 184376
rect 579526 181872 579582 181928
rect 578790 180104 578846 180160
rect 579526 177656 579582 177712
rect 578790 175072 578846 175128
rect 578422 173440 578478 173496
rect 578238 170992 578294 171048
rect 578698 169224 578754 169280
rect 578238 166912 578294 166968
rect 579526 164464 579582 164520
rect 579342 162696 579398 162752
rect 578238 159840 578294 159896
rect 578422 158344 578478 158400
rect 578882 155896 578938 155952
rect 578330 153584 578386 153640
rect 578238 151680 578294 151736
rect 578882 149640 578938 149696
rect 579526 147464 579582 147520
rect 578606 140528 578662 140584
rect 578606 138760 578662 138816
rect 579250 144644 579252 144664
rect 579252 144644 579304 144664
rect 579304 144644 579306 144664
rect 579250 144608 579306 144644
rect 579526 142976 579582 143032
rect 578882 136584 578938 136640
rect 579526 134408 579582 134464
rect 579066 132232 579122 132288
rect 578882 129648 578938 129704
rect 579526 127880 579582 127936
rect 578330 125296 578386 125352
rect 578422 123564 578424 123584
rect 578424 123564 578476 123584
rect 578476 123564 578478 123584
rect 578422 123528 578478 123564
rect 578882 121352 578938 121408
rect 578514 118396 578516 118416
rect 578516 118396 578568 118416
rect 578568 118396 578570 118416
rect 578514 118360 578570 118396
rect 578330 108296 578386 108352
rect 578606 99220 578608 99240
rect 578608 99220 578660 99240
rect 578660 99220 578662 99240
rect 578606 99184 578662 99220
rect 578330 97416 578386 97472
rect 578514 93064 578570 93120
rect 579526 116900 579528 116920
rect 579528 116900 579580 116920
rect 579580 116900 579582 116920
rect 579526 116864 579582 116900
rect 579250 114452 579252 114472
rect 579252 114452 579304 114472
rect 579304 114452 579306 114472
rect 579250 114416 579306 114452
rect 579526 112512 579582 112568
rect 579342 110100 579344 110120
rect 579344 110100 579396 110120
rect 579396 110100 579398 110120
rect 579342 110064 579398 110100
rect 579066 105848 579122 105904
rect 579526 103264 579582 103320
rect 579526 101632 579582 101688
rect 579526 95004 579528 95024
rect 579528 95004 579580 95024
rect 579580 95004 579582 95024
rect 579526 94968 579582 95004
rect 579066 90888 579122 90944
rect 579526 88068 579528 88088
rect 579528 88068 579580 88088
rect 579580 88068 579582 88088
rect 579526 88032 579582 88068
rect 579342 86400 579398 86456
rect 579158 83952 579214 84008
rect 579066 82184 579122 82240
rect 578882 80008 578938 80064
rect 578238 75520 578294 75576
rect 579526 77832 579582 77888
rect 589462 207984 589518 208040
rect 589462 206352 589518 206408
rect 589462 204720 589518 204776
rect 589462 203088 589518 203144
rect 589462 201456 589518 201512
rect 589462 199824 589518 199880
rect 590382 198192 590438 198248
rect 589462 196560 589518 196616
rect 589278 194928 589334 194984
rect 589462 193296 589518 193352
rect 589462 191664 589518 191720
rect 590566 190032 590622 190088
rect 589646 188400 589702 188456
rect 589462 186768 589518 186824
rect 589462 185136 589518 185192
rect 589462 183504 589518 183560
rect 590566 181872 590622 181928
rect 589646 180240 589702 180296
rect 589462 178608 589518 178664
rect 589646 176976 589702 177032
rect 589462 175364 589518 175400
rect 589462 175344 589464 175364
rect 589464 175344 589516 175364
rect 589516 175344 589518 175364
rect 589462 173712 589518 173768
rect 589462 172080 589518 172136
rect 589646 170448 589702 170504
rect 589462 168816 589518 168872
rect 589462 167184 589518 167240
rect 589462 165552 589518 165608
rect 589462 163920 589518 163976
rect 589462 162288 589518 162344
rect 589462 160656 589518 160712
rect 589462 159024 589518 159080
rect 589278 157412 589334 157448
rect 589278 157392 589280 157412
rect 589280 157392 589332 157412
rect 589332 157392 589334 157412
rect 589462 155760 589518 155816
rect 589462 154128 589518 154184
rect 589462 152496 589518 152552
rect 590014 150864 590070 150920
rect 589462 149232 589518 149288
rect 588542 147600 588598 147656
rect 589462 145968 589518 146024
rect 589462 144336 589518 144392
rect 589830 142704 589886 142760
rect 589462 141072 589518 141128
rect 589462 139460 589518 139496
rect 589462 139440 589464 139460
rect 589464 139440 589516 139460
rect 589516 139440 589518 139460
rect 589462 137808 589518 137864
rect 589462 136176 589518 136232
rect 590382 134544 590438 134600
rect 589462 132912 589518 132968
rect 589462 131300 589518 131336
rect 589462 131280 589464 131300
rect 589464 131280 589516 131300
rect 589516 131280 589518 131300
rect 588542 129648 588598 129704
rect 581642 77832 581698 77888
rect 579066 73072 579122 73128
rect 576122 54984 576178 55040
rect 579066 71168 579122 71224
rect 580262 54712 580318 54768
rect 578882 54440 578938 54496
rect 589462 128016 589518 128072
rect 589922 126384 589978 126440
rect 589462 124752 589518 124808
rect 589462 123120 589518 123176
rect 590014 121488 590070 121544
rect 589646 119856 589702 119912
rect 589462 116592 589518 116648
rect 590106 118224 590162 118280
rect 589462 113328 589518 113384
rect 590290 114960 590346 115016
rect 589462 111696 589518 111752
rect 589278 110064 589334 110120
rect 589462 108432 589518 108488
rect 589830 106800 589886 106856
rect 589462 105168 589518 105224
rect 588726 103536 588782 103592
rect 589462 101904 589518 101960
rect 577502 54168 577558 54224
rect 459834 53624 459890 53680
rect 460754 53624 460810 53680
rect 461674 53624 461730 53680
rect 462594 53624 462650 53680
rect 460386 53352 460442 53408
rect 465446 53352 465502 53408
rect 130382 44240 130438 44296
rect 458178 46960 458234 47016
rect 522946 47776 523002 47832
rect 458362 46688 458418 46744
rect 132774 44252 132776 44296
rect 132776 44252 132828 44296
rect 132828 44252 132830 44296
rect 132774 44240 132830 44252
rect 142618 44240 142674 44296
rect 255870 44104 255926 44160
rect 419722 43832 419778 43888
rect 440238 43852 440294 43888
rect 440238 43832 440240 43852
rect 440240 43832 440292 43852
rect 440292 43832 440294 43852
rect 441066 43852 441122 43888
rect 441066 43832 441068 43852
rect 441068 43832 441120 43852
rect 441120 43832 441122 43852
rect 361946 41792 362002 41848
rect 365166 41792 365222 41848
rect 416686 42200 416742 42256
rect 415582 42064 415638 42120
rect 446218 42200 446274 42256
rect 446218 41520 446274 41576
rect 460110 44104 460166 44160
rect 460754 43424 460810 43480
rect 461950 44240 462006 44296
rect 462870 43968 462926 44024
rect 462686 43152 462742 43208
rect 461766 42880 461822 42936
rect 463698 44240 463754 44296
rect 463974 42880 464030 42936
rect 465078 46960 465134 47016
rect 549994 48864 550050 48920
rect 591486 101632 591542 101688
rect 599490 221448 599546 221504
rect 595166 217232 595222 217288
rect 595718 216960 595774 217016
rect 599030 215600 599086 215656
rect 600870 221176 600926 221232
rect 611634 220224 611690 220280
rect 612738 219680 612794 219736
rect 618258 220904 618314 220960
rect 617154 219952 617210 220008
rect 617798 215872 617854 215928
rect 618442 219408 618498 219464
rect 621110 215328 621166 215384
rect 623962 218048 624018 218104
rect 630678 218320 630734 218376
rect 667662 698264 667718 698320
rect 667478 645768 667534 645824
rect 667294 600888 667350 600944
rect 668398 689424 668454 689480
rect 668214 687792 668270 687848
rect 668858 730088 668914 730144
rect 669410 728728 669466 728784
rect 669042 690512 669098 690568
rect 668398 593408 668454 593464
rect 671250 733760 671306 733816
rect 670882 694864 670938 694920
rect 669778 683848 669834 683904
rect 669042 594768 669098 594824
rect 668766 562264 668822 562320
rect 669594 644272 669650 644328
rect 670606 684936 670662 684992
rect 669594 552200 669650 552256
rect 675850 895464 675906 895520
rect 676034 894648 676090 894704
rect 675850 893832 675906 893888
rect 671526 668072 671582 668128
rect 671342 638696 671398 638752
rect 671710 647808 671766 647864
rect 670422 549616 670478 549672
rect 669778 455368 669834 455424
rect 671158 608504 671214 608560
rect 670974 578176 671030 578232
rect 670974 533976 671030 534032
rect 676034 893036 676090 893072
rect 676034 893016 676036 893036
rect 676036 893016 676088 893036
rect 676088 893016 676090 893036
rect 676034 892608 676090 892664
rect 676034 891384 676090 891440
rect 675206 890976 675262 891032
rect 676034 890160 676090 890216
rect 676034 889344 676090 889400
rect 676034 888956 676090 888992
rect 676034 888936 676036 888956
rect 676036 888936 676088 888956
rect 676088 888936 676090 888956
rect 676034 888548 676090 888584
rect 676034 888528 676036 888548
rect 676036 888528 676088 888548
rect 676088 888528 676090 888548
rect 676034 887324 676090 887360
rect 676034 887304 676036 887324
rect 676036 887304 676088 887324
rect 676088 887304 676090 887324
rect 676034 886916 676090 886952
rect 676034 886896 676036 886916
rect 676036 886896 676088 886916
rect 676088 886896 676090 886916
rect 676034 885692 676090 885728
rect 676034 885672 676036 885692
rect 676036 885672 676088 885692
rect 676088 885672 676090 885692
rect 675758 878464 675814 878520
rect 679622 891792 679678 891848
rect 678242 889752 678298 889808
rect 681002 890568 681058 890624
rect 683118 888120 683174 888176
rect 681002 880640 681058 880696
rect 683118 880368 683174 880424
rect 679622 878464 679678 878520
rect 675390 877920 675446 877976
rect 675574 874112 675630 874168
rect 675758 872752 675814 872808
rect 675758 869760 675814 869816
rect 675298 865680 675354 865736
rect 675758 865408 675814 865464
rect 675666 864864 675722 864920
rect 675758 788024 675814 788080
rect 675114 786664 675170 786720
rect 675390 786664 675446 786720
rect 673274 777416 673330 777472
rect 673090 714040 673146 714096
rect 672906 712816 672962 712872
rect 672722 711592 672778 711648
rect 673458 734168 673514 734224
rect 673274 708328 673330 708384
rect 673182 696904 673238 696960
rect 672998 688780 673000 688800
rect 673000 688780 673052 688800
rect 673052 688780 673054 688800
rect 672998 688744 673054 688780
rect 672814 685616 672870 685672
rect 672630 669840 672686 669896
rect 672170 652432 672226 652488
rect 672630 649168 672686 649224
rect 672998 648760 673054 648816
rect 672814 621424 672870 621480
rect 672538 620644 672540 620664
rect 672540 620644 672592 620664
rect 672592 620644 672594 620664
rect 672538 620608 672594 620644
rect 672170 609048 672226 609104
rect 670606 455096 670662 455152
rect 657542 403280 657598 403336
rect 652022 400832 652078 400888
rect 651470 373224 651526 373280
rect 652206 396616 652262 396672
rect 654782 382880 654838 382936
rect 652206 373904 652262 373960
rect 652022 372136 652078 372192
rect 670514 392536 670570 392592
rect 668582 371184 668638 371240
rect 651470 370640 651526 370696
rect 654782 358536 654838 358592
rect 652022 356632 652078 356688
rect 651378 328072 651434 328128
rect 652390 351056 652446 351112
rect 653402 338680 653458 338736
rect 652390 329704 652446 329760
rect 652022 326848 652078 326904
rect 651378 325644 651434 325680
rect 669410 347248 669466 347304
rect 651378 325624 651380 325644
rect 651380 325624 651432 325644
rect 651432 325624 651434 325644
rect 653402 313248 653458 313304
rect 652298 309848 652354 309904
rect 651378 303320 651434 303376
rect 660302 311888 660358 311944
rect 652298 302096 652354 302152
rect 651470 300600 651526 300656
rect 652574 298560 652630 298616
rect 652114 297472 652170 297528
rect 651930 296812 651986 296848
rect 651930 296792 651932 296812
rect 651932 296792 651984 296812
rect 651984 296792 651986 296812
rect 651654 295296 651710 295352
rect 651470 294208 651526 294264
rect 651470 291624 651526 291680
rect 651378 290420 651434 290456
rect 651378 290400 651380 290420
rect 651380 290400 651432 290420
rect 651432 290400 651434 290420
rect 651654 290400 651710 290456
rect 651470 288632 651526 288688
rect 651470 287408 651526 287464
rect 651470 285912 651526 285968
rect 651470 284688 651526 284744
rect 652850 293800 652906 293856
rect 652390 292712 652446 292768
rect 652206 289176 652262 289232
rect 652022 283464 652078 283520
rect 651470 283192 651526 283248
rect 652022 282104 652078 282160
rect 651470 280880 651526 280936
rect 649814 221448 649870 221504
rect 646042 219816 646098 219872
rect 648526 218592 648582 218648
rect 651102 217232 651158 217288
rect 651470 221720 651526 221776
rect 652574 280336 652630 280392
rect 652206 228520 652262 228576
rect 665822 268504 665878 268560
rect 664442 247968 664498 248024
rect 666558 245656 666614 245712
rect 663890 229744 663946 229800
rect 652574 226888 652630 226944
rect 653586 226344 653642 226400
rect 653402 222808 653458 222864
rect 659106 225528 659162 225584
rect 654782 224984 654838 225040
rect 654138 220768 654194 220824
rect 653770 217504 653826 217560
rect 656162 223896 656218 223952
rect 657542 223624 657598 223680
rect 656714 218864 656770 218920
rect 658922 222264 658978 222320
rect 657910 215328 657966 215384
rect 658738 213424 658794 213480
rect 660394 214512 660450 214568
rect 661498 213152 661554 213208
rect 662418 215600 662474 215656
rect 664442 225800 664498 225856
rect 665822 230424 665878 230480
rect 666006 230152 666062 230208
rect 667018 223624 667074 223680
rect 667018 222264 667074 222320
rect 666650 218864 666706 218920
rect 666650 217776 666706 217832
rect 666834 215600 666890 215656
rect 666834 198464 666890 198520
rect 666650 188808 666706 188864
rect 667754 224168 667810 224224
rect 667754 220768 667810 220824
rect 667754 219408 667810 219464
rect 667570 181328 667626 181384
rect 667386 178744 667442 178800
rect 668674 232464 668730 232520
rect 668306 231104 668362 231160
rect 669962 301960 670018 302016
rect 670330 263744 670386 263800
rect 670146 258440 670202 258496
rect 670330 238584 670386 238640
rect 668490 221720 668546 221776
rect 668306 204040 668362 204096
rect 668398 198736 668454 198792
rect 668122 194248 668178 194304
rect 667938 184456 667994 184512
rect 668214 177964 668216 177984
rect 668216 177964 668268 177984
rect 668268 177964 668270 177984
rect 668214 177928 668270 177964
rect 667754 174936 667810 174992
rect 667938 174700 667940 174720
rect 667940 174700 667992 174720
rect 667992 174700 667994 174720
rect 667938 174664 667994 174700
rect 667938 169668 667940 169688
rect 667940 169668 667992 169688
rect 667992 169668 667994 169688
rect 667938 169632 667994 169668
rect 668030 164908 668032 164928
rect 668032 164908 668084 164928
rect 668084 164908 668086 164928
rect 668030 164872 668086 164908
rect 668214 160012 668216 160032
rect 668216 160012 668268 160032
rect 668268 160012 668270 160032
rect 668214 159976 668270 160012
rect 668214 155116 668216 155136
rect 668216 155116 668268 155136
rect 668268 155116 668270 155136
rect 668214 155080 668270 155116
rect 668398 143656 668454 143712
rect 670330 224576 670386 224632
rect 670974 296248 671030 296304
rect 670974 293800 671030 293856
rect 671802 557504 671858 557560
rect 672354 604288 672410 604344
rect 672538 597352 672594 597408
rect 672722 573552 672778 573608
rect 674378 779320 674434 779376
rect 674010 734984 674066 735040
rect 674562 778776 674618 778832
rect 674930 777008 674986 777064
rect 674930 775668 674986 775704
rect 674930 775648 674932 775668
rect 674932 775648 674984 775668
rect 674984 775648 674986 775668
rect 675482 779320 675538 779376
rect 675482 778776 675538 778832
rect 675390 777416 675446 777472
rect 675482 777008 675538 777064
rect 675390 775648 675446 775704
rect 675114 743280 675170 743336
rect 675114 738112 675170 738168
rect 675482 734984 675538 735040
rect 675482 734168 675538 734224
rect 675482 733760 675538 733816
rect 675298 730768 675354 730824
rect 675114 729816 675170 729872
rect 675482 730088 675538 730144
rect 675482 728728 675538 728784
rect 682382 726552 682438 726608
rect 674010 721656 674066 721712
rect 674930 721656 674986 721712
rect 674010 719752 674066 719808
rect 674010 715708 674012 715728
rect 674012 715708 674064 715728
rect 674064 715708 674066 715728
rect 674010 715672 674066 715708
rect 674010 715300 674012 715320
rect 674012 715300 674064 715320
rect 674064 715300 674066 715320
rect 674010 715264 674066 715300
rect 674010 714484 674012 714504
rect 674012 714484 674064 714504
rect 674064 714484 674066 714504
rect 674010 714448 674066 714484
rect 674010 713668 674012 713688
rect 674012 713668 674064 713688
rect 674064 713668 674066 713688
rect 674010 713632 674066 713668
rect 674010 713244 674066 713280
rect 674010 713224 674012 713244
rect 674012 713224 674064 713244
rect 674064 713224 674066 713244
rect 674010 712428 674066 712464
rect 674010 712408 674012 712428
rect 674012 712408 674064 712428
rect 674064 712408 674066 712428
rect 674010 709996 674012 710016
rect 674012 709996 674064 710016
rect 674064 709996 674066 710016
rect 674010 709960 674066 709996
rect 674010 709180 674012 709200
rect 674012 709180 674064 709200
rect 674064 709180 674066 709200
rect 674010 709144 674066 709180
rect 673734 707512 673790 707568
rect 676034 716508 676090 716544
rect 676034 716488 676036 716508
rect 676036 716488 676088 716508
rect 676088 716488 676090 716508
rect 676034 716080 676090 716136
rect 676034 714892 676036 714912
rect 676036 714892 676088 714912
rect 676088 714892 676090 714912
rect 676034 714856 676090 714892
rect 675298 712000 675354 712056
rect 682382 711184 682438 711240
rect 681002 710776 681058 710832
rect 676034 710368 676090 710424
rect 676034 708756 676090 708792
rect 676034 708736 676036 708756
rect 676036 708736 676088 708756
rect 676088 708736 676090 708756
rect 676034 707140 676036 707160
rect 676036 707140 676088 707160
rect 676088 707140 676090 707160
rect 676034 707104 676090 707140
rect 684222 726280 684278 726336
rect 684222 709552 684278 709608
rect 684038 707920 684094 707976
rect 683394 706696 683450 706752
rect 675850 706288 675906 706344
rect 683118 705472 683174 705528
rect 676034 705064 676090 705120
rect 673734 701156 673736 701176
rect 673736 701156 673788 701176
rect 673788 701156 673790 701176
rect 673734 701120 673790 701156
rect 673458 682352 673514 682408
rect 675114 701120 675170 701176
rect 675114 698264 675170 698320
rect 675114 696904 675170 696960
rect 675482 696768 675538 696824
rect 674010 692960 674066 693016
rect 673458 682080 673514 682136
rect 673550 671356 673606 671392
rect 673550 671336 673552 671356
rect 673552 671336 673604 671356
rect 673604 671336 673606 671356
rect 673550 670928 673606 670984
rect 673550 670520 673606 670576
rect 673366 670112 673422 670168
rect 673366 669432 673422 669488
rect 673550 668888 673606 668944
rect 673550 668516 673552 668536
rect 673552 668516 673604 668536
rect 673604 668516 673606 668536
rect 673550 668480 673606 668516
rect 673550 668108 673552 668128
rect 673552 668108 673604 668128
rect 673604 668108 673606 668128
rect 673550 668072 673606 668108
rect 673550 667664 673606 667720
rect 673550 666712 673606 666768
rect 673550 665252 673552 665272
rect 673552 665252 673604 665272
rect 673604 665252 673606 665272
rect 673550 665216 673606 665252
rect 673550 664420 673606 664456
rect 673550 664400 673552 664420
rect 673552 664400 673604 664420
rect 673604 664400 673606 664420
rect 673366 663992 673422 664048
rect 673550 663720 673606 663776
rect 673550 661952 673606 662008
rect 673366 659640 673422 659696
rect 673182 619384 673238 619440
rect 673182 608232 673238 608288
rect 673182 598032 673238 598088
rect 673182 581052 673238 581088
rect 673182 581032 673184 581052
rect 673184 581032 673236 581052
rect 673236 581032 673238 581052
rect 673182 580252 673184 580272
rect 673184 580252 673236 580272
rect 673236 580252 673238 580272
rect 673182 580216 673238 580252
rect 673182 579980 673184 580000
rect 673184 579980 673236 580000
rect 673236 579980 673238 580000
rect 673182 579944 673238 579980
rect 673182 579692 673238 579728
rect 673182 579672 673184 579692
rect 673184 579672 673236 579692
rect 673236 579672 673238 579692
rect 673182 578892 673184 578912
rect 673184 578892 673236 578912
rect 673236 578892 673238 578912
rect 673182 578856 673238 578892
rect 673182 577904 673238 577960
rect 673182 577652 673238 577688
rect 673182 577632 673184 577652
rect 673184 577632 673236 577652
rect 673236 577632 673238 577652
rect 673182 577396 673184 577416
rect 673184 577396 673236 577416
rect 673236 577396 673238 577416
rect 673182 577360 673238 577396
rect 673182 577124 673184 577144
rect 673184 577124 673236 577144
rect 673236 577124 673238 577144
rect 673182 577088 673238 577124
rect 673182 576852 673184 576872
rect 673184 576852 673236 576872
rect 673236 576852 673238 576872
rect 673182 576816 673238 576852
rect 672998 572736 673054 572792
rect 673090 559000 673146 559056
rect 672906 555192 672962 555248
rect 672722 554804 672778 554840
rect 672722 554784 672724 554804
rect 672724 554784 672776 554804
rect 672776 554784 672778 554804
rect 672722 533568 672778 533624
rect 672906 490456 672962 490512
rect 672722 490048 672778 490104
rect 672262 453908 672264 453928
rect 672264 453908 672316 453928
rect 672316 453908 672318 453928
rect 672262 453872 672318 453908
rect 673090 484744 673146 484800
rect 673550 625948 673552 625968
rect 673552 625948 673604 625968
rect 673604 625948 673606 625968
rect 673550 625912 673606 625948
rect 674010 690260 674066 690296
rect 674010 690240 674012 690260
rect 674012 690240 674064 690260
rect 674064 690240 674066 690260
rect 675114 694864 675170 694920
rect 675114 694592 675170 694648
rect 675482 692960 675538 693016
rect 675114 690512 675170 690568
rect 674930 690240 674986 690296
rect 673918 663176 673974 663232
rect 673918 661580 673920 661600
rect 673920 661580 673972 661600
rect 673972 661580 673974 661600
rect 673918 661544 673974 661580
rect 673918 661156 673974 661192
rect 673918 661136 673920 661156
rect 673920 661136 673972 661156
rect 673972 661136 673974 661156
rect 673918 660084 673920 660104
rect 673920 660084 673972 660104
rect 673972 660084 673974 660104
rect 673918 660048 673974 660084
rect 673918 655580 673974 655616
rect 673918 655560 673920 655580
rect 673920 655560 673972 655580
rect 673972 655560 673974 655580
rect 675114 689424 675170 689480
rect 674930 688744 674986 688800
rect 675114 687792 675170 687848
rect 675298 686160 675354 686216
rect 675022 685888 675078 685944
rect 674746 682388 674748 682408
rect 674748 682388 674800 682408
rect 674800 682388 674802 682408
rect 674746 682352 674802 682388
rect 675022 676368 675078 676424
rect 674010 645496 674066 645552
rect 674010 643456 674066 643512
rect 674010 643084 674012 643104
rect 674012 643084 674064 643104
rect 674064 643084 674066 643104
rect 674010 643048 674066 643084
rect 673918 641688 673974 641744
rect 673642 620200 673698 620256
rect 673642 619828 673644 619848
rect 673644 619828 673696 619848
rect 673696 619828 673698 619848
rect 673642 619792 673698 619828
rect 673642 619112 673698 619168
rect 673642 618160 673698 618216
rect 673642 617752 673698 617808
rect 673642 615476 673644 615496
rect 673644 615476 673696 615496
rect 673696 615476 673698 615496
rect 673642 615440 673698 615476
rect 673642 614916 673698 614952
rect 673642 614896 673644 614916
rect 673644 614896 673696 614916
rect 673696 614896 673698 614916
rect 673642 611380 673698 611416
rect 673642 611360 673644 611380
rect 673644 611360 673696 611380
rect 673696 611360 673698 611380
rect 674838 669840 674894 669896
rect 674838 667392 674894 667448
rect 675482 685616 675538 685672
rect 675482 684936 675538 684992
rect 675482 683848 675538 683904
rect 684130 682624 684186 682680
rect 675482 682080 675538 682136
rect 676494 669468 676496 669488
rect 676496 669468 676548 669488
rect 676548 669468 676550 669488
rect 676494 669432 676550 669468
rect 676494 667020 676496 667040
rect 676496 667020 676548 667040
rect 676548 667020 676550 667040
rect 676494 666984 676550 667020
rect 675298 666440 675354 666496
rect 676034 664808 676090 664864
rect 674838 663756 674840 663776
rect 674840 663756 674892 663776
rect 674892 663756 674894 663776
rect 674838 663720 674894 663756
rect 683210 663720 683266 663776
rect 684130 666168 684186 666224
rect 683486 662904 683542 662960
rect 674838 660048 674894 660104
rect 683118 660048 683174 660104
rect 675114 655560 675170 655616
rect 675390 652840 675446 652896
rect 675114 652432 675170 652488
rect 675390 649168 675446 649224
rect 675114 648760 675170 648816
rect 675390 647808 675446 647864
rect 675022 646040 675078 646096
rect 675114 645768 675170 645824
rect 675114 645496 675170 645552
rect 675298 644272 675354 644328
rect 675298 643456 675354 643512
rect 675114 643048 675170 643104
rect 674838 640212 674894 640248
rect 674838 640192 674840 640212
rect 674840 640192 674892 640212
rect 674892 640192 674894 640212
rect 675298 641688 675354 641744
rect 674010 626320 674066 626376
rect 674010 625504 674066 625560
rect 674010 624996 674012 625016
rect 674012 624996 674064 625016
rect 674064 624996 674066 625016
rect 674010 624960 674066 624996
rect 674010 624708 674066 624744
rect 674010 624688 674012 624708
rect 674012 624688 674064 624708
rect 674064 624688 674066 624708
rect 674010 624316 674012 624336
rect 674012 624316 674064 624336
rect 674064 624316 674066 624336
rect 674010 624280 674066 624316
rect 674010 623892 674066 623928
rect 674010 623872 674012 623892
rect 674012 623872 674064 623892
rect 674064 623872 674066 623892
rect 674010 623500 674012 623520
rect 674012 623500 674064 623520
rect 674064 623500 674066 623520
rect 674010 623464 674066 623500
rect 674010 623076 674066 623112
rect 674010 623056 674012 623076
rect 674012 623056 674064 623076
rect 674064 623056 674066 623076
rect 674010 622684 674012 622704
rect 674012 622684 674064 622704
rect 674064 622684 674066 622704
rect 674010 622648 674066 622684
rect 674010 622260 674066 622296
rect 674010 622240 674012 622260
rect 674012 622240 674064 622260
rect 674064 622240 674066 622260
rect 674010 621152 674066 621208
rect 674746 625912 674802 625968
rect 674286 619112 674342 619168
rect 674286 615476 674288 615496
rect 674288 615476 674340 615496
rect 674340 615476 674342 615496
rect 674286 615440 674342 615476
rect 674286 609048 674342 609104
rect 673826 600616 673882 600672
rect 673826 600380 673828 600400
rect 673828 600380 673880 600400
rect 673880 600380 673882 600400
rect 673826 600344 673882 600380
rect 673734 599800 673790 599856
rect 673550 598576 673606 598632
rect 675482 638696 675538 638752
rect 679622 637472 679678 637528
rect 675482 631352 675538 631408
rect 675666 631352 675722 631408
rect 676494 625676 676496 625696
rect 676496 625676 676548 625696
rect 676548 625676 676550 625696
rect 676494 625640 676550 625676
rect 679622 621968 679678 622024
rect 683210 618704 683266 618760
rect 676218 617516 676220 617536
rect 676220 617516 676272 617536
rect 676272 617516 676274 617536
rect 676218 617480 676274 617516
rect 675298 617072 675354 617128
rect 683578 617072 683634 617128
rect 683394 616664 683450 616720
rect 683118 615476 683120 615496
rect 683120 615476 683172 615496
rect 683172 615476 683174 615496
rect 683118 615440 683174 615476
rect 675298 611360 675354 611416
rect 675022 608504 675078 608560
rect 674930 608232 674986 608288
rect 674286 600616 674342 600672
rect 673918 574776 673974 574832
rect 673918 574540 673920 574560
rect 673920 574540 673972 574560
rect 673972 574540 673974 574560
rect 673918 574504 673974 574540
rect 673918 574096 673974 574152
rect 673918 573860 673920 573880
rect 673920 573860 673972 573880
rect 673972 573860 673974 573880
rect 673918 573824 673974 573860
rect 673918 572056 673974 572112
rect 673918 571396 673974 571432
rect 673918 571376 673920 571396
rect 673920 571376 673972 571396
rect 673972 571376 673974 571396
rect 673918 571124 673974 571160
rect 673918 571104 673920 571124
rect 673920 571104 673972 571124
rect 673972 571104 673974 571124
rect 673918 570832 673974 570888
rect 673918 569608 673974 569664
rect 673918 565836 673920 565856
rect 673920 565836 673972 565856
rect 673972 565836 673974 565856
rect 673918 565800 673974 565836
rect 673918 564460 673974 564496
rect 673918 564440 673920 564460
rect 673920 564440 673972 564460
rect 673972 564440 673974 564460
rect 673918 558320 673974 558376
rect 675114 604288 675170 604344
rect 675114 602928 675170 602984
rect 675390 600888 675446 600944
rect 675114 600344 675170 600400
rect 675482 599800 675538 599856
rect 675482 598576 675538 598632
rect 675114 598032 675170 598088
rect 675390 597352 675446 597408
rect 675390 595312 675446 595368
rect 675482 594768 675538 594824
rect 675390 593408 675446 593464
rect 675022 591504 675078 591560
rect 674378 579708 674380 579728
rect 674380 579708 674432 579728
rect 674432 579708 674434 579728
rect 674378 579672 674434 579708
rect 674470 578176 674526 578232
rect 674378 577532 674380 577552
rect 674380 577532 674432 577552
rect 674432 577532 674434 577552
rect 674378 577496 674434 577532
rect 674562 574776 674618 574832
rect 674378 573824 674434 573880
rect 674378 571412 674380 571432
rect 674380 571412 674432 571432
rect 674432 571412 674434 571432
rect 674378 571376 674434 571412
rect 674838 571104 674894 571160
rect 675482 593136 675538 593192
rect 675206 586200 675262 586256
rect 676218 580488 676274 580544
rect 676218 579264 676274 579320
rect 676218 578040 676274 578096
rect 682382 591368 682438 591424
rect 679622 576408 679678 576464
rect 682382 575592 682438 575648
rect 676218 574776 676274 574832
rect 684222 591096 684278 591152
rect 683394 573144 683450 573200
rect 676218 572328 676274 572384
rect 684222 576000 684278 576056
rect 684038 571920 684094 571976
rect 676034 571240 676090 571296
rect 683118 570288 683174 570344
rect 675390 565800 675446 565856
rect 675114 564440 675170 564496
rect 675114 562264 675170 562320
rect 675390 561856 675446 561912
rect 674102 554104 674158 554160
rect 674286 552880 674342 552936
rect 673734 550432 673790 550488
rect 674102 537104 674158 537160
rect 673642 526360 673698 526416
rect 673826 492088 673882 492144
rect 674010 491308 674012 491328
rect 674012 491308 674064 491328
rect 674064 491308 674066 491328
rect 674010 491272 674066 491308
rect 674010 490900 674012 490920
rect 674012 490900 674064 490920
rect 674064 490900 674066 490920
rect 674010 490864 674066 490900
rect 674010 489660 674066 489696
rect 674010 489640 674012 489660
rect 674012 489640 674064 489660
rect 674064 489640 674066 489660
rect 674010 489268 674012 489288
rect 674012 489268 674064 489288
rect 674064 489268 674066 489288
rect 674010 489232 674066 489268
rect 674010 488452 674012 488472
rect 674012 488452 674064 488472
rect 674064 488452 674066 488472
rect 674010 488416 674066 488452
rect 674010 486004 674012 486024
rect 674012 486004 674064 486024
rect 674064 486004 674066 486024
rect 674010 485968 674066 486004
rect 673642 484336 673698 484392
rect 674010 483148 674012 483168
rect 674012 483148 674064 483168
rect 674064 483148 674066 483168
rect 674010 483112 674066 483148
rect 675114 559000 675170 559056
rect 675390 558320 675446 558376
rect 675114 557504 675170 557560
rect 675390 555192 675446 555248
rect 675206 554784 675262 554840
rect 675758 554648 675814 554704
rect 675758 553832 675814 553888
rect 675298 552200 675354 552256
rect 675482 549616 675538 549672
rect 674838 548392 674894 548448
rect 675758 548256 675814 548312
rect 675574 547848 675630 547904
rect 677414 547576 677470 547632
rect 675482 537104 675538 537160
rect 676218 535880 676274 535936
rect 676034 535676 676090 535732
rect 676218 535064 676274 535120
rect 676034 534896 676036 534916
rect 676036 534896 676088 534916
rect 676088 534896 676090 534916
rect 676034 534860 676090 534896
rect 676494 534248 676550 534304
rect 676034 533248 676090 533284
rect 676034 533228 676036 533248
rect 676036 533228 676088 533248
rect 676088 533228 676090 533248
rect 676034 532840 676090 532876
rect 676034 532820 676036 532840
rect 676036 532820 676088 532840
rect 676088 532820 676090 532840
rect 676034 532448 676036 532468
rect 676036 532448 676088 532468
rect 676088 532448 676090 532468
rect 676034 532412 676090 532448
rect 676034 532024 676090 532060
rect 676034 532004 676036 532024
rect 676036 532004 676088 532024
rect 676088 532004 676090 532024
rect 676218 531820 676274 531856
rect 676218 531800 676220 531820
rect 676220 531800 676272 531820
rect 676272 531800 676274 531820
rect 676034 530816 676036 530836
rect 676036 530816 676088 530836
rect 676088 530816 676090 530836
rect 676034 530780 676090 530816
rect 676034 529984 676090 530020
rect 676034 529964 676036 529984
rect 676036 529964 676088 529984
rect 676088 529964 676090 529984
rect 676218 529352 676274 529408
rect 676034 529148 676090 529204
rect 676034 528776 676036 528796
rect 676036 528776 676088 528796
rect 676088 528776 676090 528796
rect 676034 528740 676090 528776
rect 676034 527960 676036 527980
rect 676036 527960 676088 527980
rect 676088 527960 676090 527980
rect 676034 527924 676090 527960
rect 673274 455388 673330 455424
rect 673274 455368 673276 455388
rect 673276 455368 673328 455388
rect 673328 455368 673330 455388
rect 673386 455252 673442 455288
rect 673386 455232 673388 455252
rect 673388 455232 673440 455252
rect 673440 455232 673442 455252
rect 673274 455096 673330 455152
rect 672814 454824 672870 454880
rect 674286 454860 674288 454880
rect 674288 454860 674340 454880
rect 674340 454860 674342 454880
rect 674286 454824 674342 454860
rect 673044 454588 673046 454608
rect 673046 454588 673098 454608
rect 673098 454588 673100 454608
rect 673044 454552 673100 454588
rect 674286 454588 674288 454608
rect 674288 454588 674340 454608
rect 674340 454588 674342 454608
rect 674286 454552 674342 454588
rect 676034 491700 676090 491736
rect 676034 491680 676036 491700
rect 676036 491680 676088 491700
rect 676088 491680 676090 491700
rect 676034 486784 676090 486840
rect 676034 485172 676090 485208
rect 676034 485152 676036 485172
rect 676036 485152 676088 485172
rect 676088 485152 676090 485172
rect 676034 483964 676036 483984
rect 676036 483964 676088 483984
rect 676088 483964 676090 483984
rect 676034 483928 676090 483964
rect 682382 546760 682438 546816
rect 681002 531392 681058 531448
rect 682382 530576 682438 530632
rect 683210 528536 683266 528592
rect 683578 527720 683634 527776
rect 683394 526904 683450 526960
rect 677874 525680 677930 525736
rect 683118 524864 683174 524920
rect 680358 524456 680414 524512
rect 683210 503648 683266 503704
rect 679622 487192 679678 487248
rect 681186 487600 681242 487656
rect 681002 486376 681058 486432
rect 683394 500928 683450 500984
rect 683210 485560 683266 485616
rect 683394 483520 683450 483576
rect 676034 482704 676090 482760
rect 676034 482332 676036 482352
rect 676036 482332 676088 482352
rect 676088 482332 676090 482352
rect 676034 482296 676090 482332
rect 680358 481888 680414 481944
rect 675850 480664 675906 480720
rect 683118 481072 683174 481128
rect 672952 454316 672954 454336
rect 672954 454316 673006 454336
rect 673006 454316 673008 454336
rect 672952 454280 673008 454316
rect 674286 454316 674288 454336
rect 674288 454316 674340 454336
rect 674340 454316 674342 454336
rect 674286 454280 674342 454316
rect 674286 453908 674288 453928
rect 674288 453908 674340 453928
rect 674340 453908 674342 453928
rect 674286 453872 674342 453908
rect 676218 403300 676274 403336
rect 676218 403280 676220 403300
rect 676220 403280 676272 403300
rect 676272 403280 676274 403300
rect 672630 402464 672686 402520
rect 672446 401920 672502 401976
rect 673182 401648 673238 401704
rect 672814 399608 672870 399664
rect 672630 393896 672686 393952
rect 671894 393624 671950 393680
rect 671710 348880 671766 348936
rect 671710 329704 671766 329760
rect 671526 302232 671582 302288
rect 670974 262112 671030 262168
rect 670698 257216 670754 257272
rect 670514 223896 670570 223952
rect 670422 223644 670478 223680
rect 670422 223624 670424 223644
rect 670424 223624 670476 223644
rect 670476 223624 670478 223644
rect 668950 199144 669006 199200
rect 669042 191664 669098 191720
rect 668766 163240 668822 163296
rect 668858 162288 668914 162344
rect 668766 159024 668822 159080
rect 668766 158344 668822 158400
rect 668858 148552 668914 148608
rect 668766 145288 668822 145344
rect 668582 138760 668638 138816
rect 670054 220768 670110 220824
rect 669410 217232 669466 217288
rect 669410 214784 669466 214840
rect 669410 202816 669466 202872
rect 669226 189352 669282 189408
rect 669042 135496 669098 135552
rect 667202 134544 667258 134600
rect 667938 133764 667940 133784
rect 667940 133764 667992 133784
rect 667992 133764 667994 133784
rect 667938 133728 667994 133764
rect 667018 132640 667074 132696
rect 668858 131144 668914 131200
rect 668674 130636 668676 130656
rect 668676 130636 668728 130656
rect 668728 130636 668730 130656
rect 668674 130600 668730 130636
rect 667938 128968 667994 129024
rect 668582 127744 668638 127800
rect 668398 126928 668454 126984
rect 668398 120808 668454 120864
rect 668122 112648 668178 112704
rect 668398 107752 668454 107808
rect 667938 104524 667940 104544
rect 667940 104524 667992 104544
rect 667992 104524 667994 104544
rect 667938 104488 667994 104524
rect 669594 171128 669650 171184
rect 669778 169496 669834 169552
rect 669594 154400 669650 154456
rect 669778 150320 669834 150376
rect 670330 220360 670386 220416
rect 670330 218048 670386 218104
rect 670514 216552 670570 216608
rect 670330 216416 670386 216472
rect 670146 211112 670202 211168
rect 670514 198192 670570 198248
rect 670974 236136 671030 236192
rect 670882 233980 670938 234016
rect 670882 233960 670884 233980
rect 670884 233960 670936 233980
rect 670936 233960 670938 233980
rect 670790 177964 670792 177984
rect 670792 177964 670844 177984
rect 670844 177964 670846 177984
rect 670790 177928 670846 177964
rect 670606 170312 670662 170368
rect 671710 278588 671766 278624
rect 671710 278568 671712 278588
rect 671712 278568 671764 278588
rect 671764 278568 671766 278588
rect 671710 260480 671766 260536
rect 671710 240216 671766 240272
rect 671526 224304 671582 224360
rect 672630 376216 672686 376272
rect 672538 356224 672594 356280
rect 672354 355408 672410 355464
rect 672170 353368 672226 353424
rect 672170 338000 672226 338056
rect 672998 394984 673054 395040
rect 672998 380976 673054 381032
rect 673918 401376 673974 401432
rect 673366 400424 673422 400480
rect 673182 357448 673238 357504
rect 673182 357040 673238 357096
rect 672814 355000 672870 355056
rect 672998 349696 673054 349752
rect 672722 348472 672778 348528
rect 672538 311616 672594 311672
rect 672354 310800 672410 310856
rect 672998 335552 673054 335608
rect 672906 324944 672962 325000
rect 673734 395664 673790 395720
rect 673734 375400 673790 375456
rect 676586 402872 676642 402928
rect 674838 402192 674894 402248
rect 674838 401648 674894 401704
rect 676586 400832 676642 400888
rect 676034 399336 676090 399392
rect 674746 397296 674802 397352
rect 674562 396616 674618 396672
rect 679622 398384 679678 398440
rect 676218 397976 676274 398032
rect 676034 396092 676090 396128
rect 676034 396072 676036 396092
rect 676036 396072 676088 396092
rect 676088 396072 676090 396092
rect 678242 397568 678298 397624
rect 676218 394324 676274 394360
rect 676218 394304 676220 394324
rect 676220 394304 676272 394324
rect 676272 394304 676274 394324
rect 678242 387640 678298 387696
rect 675758 384920 675814 384976
rect 675114 382880 675170 382936
rect 675758 382200 675814 382256
rect 675390 380976 675446 381032
rect 675666 378528 675722 378584
rect 675758 377440 675814 377496
rect 675390 376216 675446 376272
rect 675114 375400 675170 375456
rect 675758 373632 675814 373688
rect 675114 372816 675170 372872
rect 675022 371184 675078 371240
rect 674102 358264 674158 358320
rect 673918 356496 673974 356552
rect 673366 355816 673422 355872
rect 673918 354592 673974 354648
rect 673550 350512 673606 350568
rect 673366 350104 673422 350160
rect 673366 335824 673422 335880
rect 673734 349288 673790 349344
rect 673734 332696 673790 332752
rect 673550 331064 673606 331120
rect 675942 357856 675998 357912
rect 675942 356768 675998 356824
rect 674470 352552 674526 352608
rect 674286 351328 674342 351384
rect 674102 351056 674158 351112
rect 674286 337728 674342 337784
rect 674654 352144 674710 352200
rect 676034 350920 676090 350976
rect 676034 346568 676090 346624
rect 674930 338680 674986 338736
rect 675758 340176 675814 340232
rect 675482 339360 675538 339416
rect 675114 338000 675170 338056
rect 675758 337864 675814 337920
rect 675114 337728 675170 337784
rect 675758 336504 675814 336560
rect 674930 335824 674986 335880
rect 675114 335552 675170 335608
rect 675114 332696 675170 332752
rect 675298 331064 675354 331120
rect 675114 329704 675170 329760
rect 675022 327936 675078 327992
rect 674654 326848 674710 326904
rect 673366 312704 673422 312760
rect 673182 312432 673238 312488
rect 673182 311208 673238 311264
rect 673090 304272 673146 304328
rect 673090 287816 673146 287872
rect 672906 278568 672962 278624
rect 672354 265376 672410 265432
rect 674194 310392 674250 310448
rect 673918 305088 673974 305144
rect 673734 303864 673790 303920
rect 673734 290400 673790 290456
rect 673550 286456 673606 286512
rect 673918 286864 673974 286920
rect 673918 283464 673974 283520
rect 675390 327936 675446 327992
rect 675390 326848 675446 326904
rect 675206 325624 675262 325680
rect 675022 324944 675078 325000
rect 676218 313928 676274 313984
rect 674654 312976 674710 313032
rect 674838 312704 674894 312760
rect 674838 312024 674894 312080
rect 674654 311888 674710 311944
rect 674378 309984 674434 310040
rect 674654 309576 674710 309632
rect 674470 305496 674526 305552
rect 675850 309304 675906 309360
rect 675850 309032 675906 309088
rect 675022 307944 675078 308000
rect 674838 306312 674894 306368
rect 675390 307536 675446 307592
rect 675206 302912 675262 302968
rect 676034 308352 676090 308408
rect 676034 307128 676090 307184
rect 675850 306584 675906 306640
rect 676034 305904 676090 305960
rect 676034 303456 676090 303512
rect 675850 302912 675906 302968
rect 676034 301960 676090 302016
rect 679622 306720 679678 306776
rect 676218 301552 676274 301608
rect 674838 294480 674894 294536
rect 676862 297336 676918 297392
rect 675482 296656 675538 296712
rect 675666 296248 675722 296304
rect 675298 295840 675354 295896
rect 675666 295840 675722 295896
rect 675758 294480 675814 294536
rect 675758 291488 675814 291544
rect 675758 290944 675814 291000
rect 675114 287816 675170 287872
rect 673918 268232 673974 268288
rect 673734 267824 673790 267880
rect 673366 267416 673422 267472
rect 673918 267008 673974 267064
rect 673182 266600 673238 266656
rect 673550 264560 673606 264616
rect 672170 246200 672226 246256
rect 672262 236988 672264 237008
rect 672264 236988 672316 237008
rect 672316 236988 672318 237008
rect 672262 236952 672318 236988
rect 671894 231920 671950 231976
rect 672630 227024 672686 227080
rect 673182 263336 673238 263392
rect 672998 259664 673054 259720
rect 673274 258848 673330 258904
rect 673090 250688 673146 250744
rect 673090 250008 673146 250064
rect 672998 245656 673054 245712
rect 672998 245384 673054 245440
rect 673734 260888 673790 260944
rect 673734 246608 673790 246664
rect 673550 241712 673606 241768
rect 673274 241440 673330 241496
rect 673734 236952 673790 237008
rect 672952 236408 673008 236464
rect 673550 232464 673606 232520
rect 673274 230152 673330 230208
rect 673458 229744 673514 229800
rect 672722 226380 672724 226400
rect 672724 226380 672776 226400
rect 672776 226380 672778 226400
rect 672722 226344 672778 226380
rect 672602 226108 672604 226128
rect 672604 226108 672656 226128
rect 672656 226108 672658 226128
rect 672602 226072 672658 226108
rect 672262 225800 672318 225856
rect 672378 225700 672380 225720
rect 672380 225700 672432 225720
rect 672432 225700 672434 225720
rect 672378 225664 672434 225700
rect 672154 225412 672210 225448
rect 672154 225392 672156 225412
rect 672156 225392 672208 225412
rect 672208 225392 672210 225412
rect 672032 225276 672088 225312
rect 672032 225256 672034 225276
rect 672034 225256 672086 225276
rect 672086 225256 672088 225276
rect 671818 224732 671874 224768
rect 671818 224712 671820 224732
rect 671820 224712 671872 224732
rect 671872 224712 671874 224732
rect 671480 223896 671536 223952
rect 671526 223624 671582 223680
rect 671342 177928 671398 177984
rect 670606 147600 670662 147656
rect 672078 223896 672134 223952
rect 671894 221720 671950 221776
rect 671894 218592 671950 218648
rect 672078 217504 672134 217560
rect 671894 216144 671950 216200
rect 672078 216144 672134 216200
rect 671894 215328 671950 215384
rect 672078 201320 672134 201376
rect 671894 171944 671950 172000
rect 672078 169088 672134 169144
rect 672446 224984 672502 225040
rect 672630 223624 672686 223680
rect 673550 226752 673606 226808
rect 673550 224712 673606 224768
rect 673366 223624 673422 223680
rect 673090 222808 673146 222864
rect 673182 221040 673238 221096
rect 672906 220632 672962 220688
rect 672998 217368 673054 217424
rect 672998 216552 673054 216608
rect 673366 220224 673422 220280
rect 673090 214104 673146 214160
rect 672630 213288 672686 213344
rect 672446 213152 672502 213208
rect 672446 212064 672502 212120
rect 672446 201048 672502 201104
rect 672538 200776 672594 200832
rect 672538 181600 672594 181656
rect 672538 168272 672594 168328
rect 672262 168136 672318 168192
rect 671710 150048 671766 150104
rect 672170 166912 672226 166968
rect 671986 144880 672042 144936
rect 671342 130872 671398 130928
rect 669962 129240 670018 129296
rect 669226 125704 669282 125760
rect 668950 120672 669006 120728
rect 668766 119176 668822 119232
rect 668950 111016 669006 111072
rect 670146 122712 670202 122768
rect 671986 126520 672042 126576
rect 668582 102856 668638 102912
rect 637026 96872 637082 96928
rect 641994 96464 642050 96520
rect 635738 95376 635794 95432
rect 647146 94968 647202 95024
rect 626446 94424 626502 94480
rect 626262 93608 626318 93664
rect 626446 92792 626502 92848
rect 625802 91976 625858 92032
rect 647514 92384 647570 92440
rect 626446 91160 626502 91216
rect 626446 90344 626502 90400
rect 626446 89564 626448 89584
rect 626448 89564 626500 89584
rect 626500 89564 626502 89584
rect 626446 89528 626502 89564
rect 624974 88304 625030 88360
rect 626446 87896 626502 87952
rect 626262 87080 626318 87136
rect 648250 89528 648306 89584
rect 626446 86300 626448 86320
rect 626448 86300 626500 86320
rect 626500 86300 626502 86320
rect 626446 86264 626502 86300
rect 625342 85448 625398 85504
rect 626446 84632 626502 84688
rect 625802 83816 625858 83872
rect 628746 83272 628802 83328
rect 629206 81640 629262 81696
rect 624422 77288 624478 77344
rect 633898 78512 633954 78568
rect 633898 77288 633954 77344
rect 639602 78104 639658 78160
rect 646134 74160 646190 74216
rect 646318 71712 646374 71768
rect 647238 68856 647294 68912
rect 646502 67088 646558 67144
rect 646134 64368 646190 64424
rect 648618 62056 648674 62112
rect 647238 59200 647294 59256
rect 649998 87080 650054 87136
rect 654598 94152 654654 94208
rect 654322 91432 654378 91488
rect 655426 93336 655482 93392
rect 655426 90652 655428 90672
rect 655428 90652 655480 90672
rect 655480 90652 655482 90672
rect 655426 90616 655482 90652
rect 655794 89800 655850 89856
rect 672354 152632 672410 152688
rect 672538 133320 672594 133376
rect 672538 132640 672594 132696
rect 672538 131688 672594 131744
rect 672354 131144 672410 131200
rect 672906 200640 672962 200696
rect 673090 199688 673146 199744
rect 673182 197784 673238 197840
rect 673550 216824 673606 216880
rect 673550 216552 673606 216608
rect 673550 215872 673606 215928
rect 674378 266192 674434 266248
rect 674562 265784 674618 265840
rect 675114 286864 675170 286920
rect 675390 286456 675446 286512
rect 675758 283600 675814 283656
rect 675666 282648 675722 282704
rect 675666 281560 675722 281616
rect 675114 278296 675170 278352
rect 675482 278024 675538 278080
rect 674930 276664 674986 276720
rect 674930 273808 674986 273864
rect 674746 264968 674802 265024
rect 675114 264152 675170 264208
rect 674470 262520 674526 262576
rect 674378 260072 674434 260128
rect 674102 259256 674158 259312
rect 674102 242664 674158 242720
rect 674930 254904 674986 254960
rect 676402 264016 676458 264072
rect 676218 262792 676274 262848
rect 675482 258032 675538 258088
rect 675850 254904 675906 254960
rect 674930 249464 674986 249520
rect 675482 250688 675538 250744
rect 675758 250280 675814 250336
rect 675298 248104 675354 248160
rect 675298 246608 675354 246664
rect 675758 246608 675814 246664
rect 675114 246200 675170 246256
rect 675298 245656 675354 245712
rect 675022 245384 675078 245440
rect 674562 242936 674618 242992
rect 674378 242120 674434 242176
rect 674654 236408 674710 236464
rect 674102 232636 674104 232656
rect 674104 232636 674156 232656
rect 674156 232636 674158 232656
rect 674102 232600 674158 232636
rect 674102 232364 674104 232384
rect 674104 232364 674156 232384
rect 674156 232364 674158 232384
rect 674102 232328 674158 232364
rect 674102 230424 674158 230480
rect 674102 229780 674104 229800
rect 674104 229780 674156 229800
rect 674156 229780 674158 229800
rect 674102 229744 674158 229780
rect 674102 227024 674158 227080
rect 674010 222264 674066 222320
rect 674010 217912 674066 217968
rect 675022 237224 675078 237280
rect 675390 243208 675446 243264
rect 675482 242664 675538 242720
rect 675482 242120 675538 242176
rect 675482 241440 675538 241496
rect 675482 240216 675538 240272
rect 675482 238584 675538 238640
rect 675482 237224 675538 237280
rect 675482 236136 675538 236192
rect 675482 235456 675538 235512
rect 673366 175616 673422 175672
rect 673274 174392 673330 174448
rect 673918 177248 673974 177304
rect 673918 176840 673974 176896
rect 673550 172216 673606 172272
rect 673458 171536 673514 171592
rect 673182 168680 673238 168736
rect 673182 151272 673238 151328
rect 674102 172896 674158 172952
rect 674102 172216 674158 172272
rect 673550 159976 673606 160032
rect 673734 159024 673790 159080
rect 674102 162288 674158 162344
rect 674102 162016 674158 162072
rect 673918 132096 673974 132152
rect 673366 129648 673422 129704
rect 673182 128424 673238 128480
rect 672906 126928 672962 126984
rect 672722 124072 672778 124128
rect 672722 123800 672778 123856
rect 672170 115776 672226 115832
rect 672906 123120 672962 123176
rect 672906 114280 672962 114336
rect 672722 106256 672778 106312
rect 672354 106120 672410 106176
rect 673918 124752 673974 124808
rect 674838 226072 674894 226128
rect 675850 233996 675852 234016
rect 675852 233996 675904 234016
rect 675904 233996 675906 234016
rect 675850 233960 675906 233996
rect 675850 232636 675852 232656
rect 675852 232636 675904 232656
rect 675904 232636 675906 232656
rect 675850 232600 675906 232636
rect 676034 232328 676090 232384
rect 676586 230152 676642 230208
rect 675482 228520 675538 228576
rect 676402 227024 676458 227080
rect 675482 225664 675538 225720
rect 674838 221448 674894 221504
rect 675022 221448 675078 221504
rect 674838 219000 674894 219056
rect 674470 214920 674526 214976
rect 674654 213696 674710 213752
rect 675022 218184 675078 218240
rect 675850 225392 675906 225448
rect 676034 223080 676090 223136
rect 676034 221856 676090 221912
rect 675666 221720 675722 221776
rect 675482 219816 675538 219872
rect 676034 217912 676090 217968
rect 676034 215872 676090 215928
rect 675666 215328 675722 215384
rect 683210 227024 683266 227080
rect 676954 226752 677010 226808
rect 683394 222672 683450 222728
rect 675758 214376 675814 214432
rect 675298 212472 675354 212528
rect 675206 206896 675262 206952
rect 674930 204176 674986 204232
rect 675390 204176 675446 204232
rect 674470 197104 674526 197160
rect 674930 202816 674986 202872
rect 675758 202680 675814 202736
rect 675482 201320 675538 201376
rect 674930 199688 674986 199744
rect 675758 199960 675814 200016
rect 675114 198464 675170 198520
rect 675482 198192 675538 198248
rect 675390 197104 675446 197160
rect 675758 194520 675814 194576
rect 675758 193160 675814 193216
rect 675666 192752 675722 192808
rect 676126 189080 676182 189136
rect 675114 188808 675170 188864
rect 675298 181328 675354 181384
rect 675482 179424 675538 179480
rect 675298 179016 675354 179072
rect 675666 178744 675722 178800
rect 675482 178064 675538 178120
rect 675666 177656 675722 177712
rect 674654 176024 674710 176080
rect 674470 175208 674526 175264
rect 674286 153176 674342 153232
rect 676034 173984 676090 174040
rect 679622 173168 679678 173224
rect 675850 167456 675906 167512
rect 676402 169496 676458 169552
rect 675022 161336 675078 161392
rect 676402 166368 676458 166424
rect 681002 172760 681058 172816
rect 683118 167864 683174 167920
rect 683118 162016 683174 162072
rect 676034 161336 676090 161392
rect 675482 161064 675538 161120
rect 675390 159976 675446 160032
rect 675758 155760 675814 155816
rect 675390 155488 675446 155544
rect 675114 154400 675170 154456
rect 675114 152632 675170 152688
rect 675758 151408 675814 151464
rect 675114 151272 675170 151328
rect 674930 150320 674986 150376
rect 675758 148416 675814 148472
rect 675114 147600 675170 147656
rect 675390 147600 675446 147656
rect 675114 144880 675170 144936
rect 676034 134544 676090 134600
rect 676034 132504 676090 132560
rect 674654 131280 674710 131336
rect 674470 130464 674526 130520
rect 676218 130192 676274 130248
rect 675850 128832 675906 128888
rect 674378 125160 674434 125216
rect 674102 117408 674158 117464
rect 673918 106936 673974 106992
rect 674654 123528 674710 123584
rect 676218 127744 676274 127800
rect 676402 127744 676458 127800
rect 682382 126112 682438 126168
rect 681002 125296 681058 125352
rect 681002 117272 681058 117328
rect 683302 125704 683358 125760
rect 683302 119992 683358 120048
rect 682382 116048 682438 116104
rect 675298 115776 675354 115832
rect 675022 115232 675078 115288
rect 675390 115232 675446 115288
rect 675758 115232 675814 115288
rect 675758 112376 675814 112432
rect 675758 111696 675814 111752
rect 675758 111288 675814 111344
rect 675758 110336 675814 110392
rect 675758 108160 675814 108216
rect 675390 106936 675446 106992
rect 675114 106256 675170 106312
rect 673366 103400 673422 103456
rect 675114 103400 675170 103456
rect 675390 101904 675446 101960
rect 671986 99320 672042 99376
rect 675298 99320 675354 99376
rect 663706 92792 663762 92848
rect 664166 89800 664222 89856
rect 665178 93336 665234 93392
rect 665362 91704 665418 91760
rect 665546 90616 665602 90672
rect 664350 88984 664406 89040
rect 650550 84632 650606 84688
rect 650366 82184 650422 82240
rect 648802 57296 648858 57352
rect 661590 48454 661646 48510
rect 553674 48048 553730 48104
rect 552018 47776 552074 47832
rect 547878 47504 547934 47560
rect 545670 47232 545726 47288
rect 465262 46688 465318 46744
rect 662418 47368 662474 47424
rect 464710 44240 464766 44296
rect 471058 43424 471114 43480
rect 465814 43152 465870 43208
rect 460938 42336 460994 42392
rect 518806 42744 518862 42800
rect 515402 42064 515458 42120
rect 520922 42064 520978 42120
rect 522026 42064 522082 42120
rect 526442 42064 526498 42120
rect 529570 42064 529626 42120
rect 141698 40296 141754 40352
<< metal3 >>
rect 676029 897154 676095 897157
rect 676029 897152 676292 897154
rect 676029 897096 676034 897152
rect 676090 897096 676292 897152
rect 676029 897094 676292 897096
rect 676029 897091 676095 897094
rect 675845 896746 675911 896749
rect 675845 896744 676292 896746
rect 675845 896688 675850 896744
rect 675906 896688 676292 896744
rect 675845 896686 676292 896688
rect 675845 896683 675911 896686
rect 676029 896338 676095 896341
rect 676029 896336 676292 896338
rect 676029 896280 676034 896336
rect 676090 896280 676292 896336
rect 676029 896278 676292 896280
rect 676029 896275 676095 896278
rect 675845 895522 675911 895525
rect 675845 895520 676292 895522
rect 675845 895464 675850 895520
rect 675906 895464 676292 895520
rect 675845 895462 676292 895464
rect 675845 895459 675911 895462
rect 676029 894706 676095 894709
rect 676029 894704 676292 894706
rect 676029 894648 676034 894704
rect 676090 894648 676292 894704
rect 676029 894646 676292 894648
rect 676029 894643 676095 894646
rect 675845 893890 675911 893893
rect 675845 893888 676292 893890
rect 675845 893832 675850 893888
rect 675906 893832 676292 893888
rect 675845 893830 676292 893832
rect 675845 893827 675911 893830
rect 676029 893074 676095 893077
rect 676029 893072 676292 893074
rect 676029 893016 676034 893072
rect 676090 893016 676292 893072
rect 676029 893014 676292 893016
rect 676029 893011 676095 893014
rect 676029 892666 676095 892669
rect 676029 892664 676292 892666
rect 676029 892608 676034 892664
rect 676090 892608 676292 892664
rect 676029 892606 676292 892608
rect 676029 892603 676095 892606
rect 675886 892196 675892 892260
rect 675956 892258 675962 892260
rect 675956 892198 676292 892258
rect 675956 892196 675962 892198
rect 679617 891850 679683 891853
rect 679604 891848 679683 891850
rect 679604 891792 679622 891848
rect 679678 891792 679683 891848
rect 679604 891790 679683 891792
rect 679617 891787 679683 891790
rect 676029 891442 676095 891445
rect 676029 891440 676292 891442
rect 676029 891384 676034 891440
rect 676090 891384 676292 891440
rect 676029 891382 676292 891384
rect 676029 891379 676095 891382
rect 675201 891034 675267 891037
rect 675201 891032 676292 891034
rect 675201 890976 675206 891032
rect 675262 890976 676292 891032
rect 675201 890974 676292 890976
rect 675201 890971 675267 890974
rect 680997 890626 681063 890629
rect 680997 890624 681076 890626
rect 680997 890568 681002 890624
rect 681058 890568 681076 890624
rect 680997 890566 681076 890568
rect 680997 890563 681063 890566
rect 676029 890218 676095 890221
rect 676029 890216 676292 890218
rect 676029 890160 676034 890216
rect 676090 890160 676292 890216
rect 676029 890158 676292 890160
rect 676029 890155 676095 890158
rect 678237 889810 678303 889813
rect 678237 889808 678316 889810
rect 678237 889752 678242 889808
rect 678298 889752 678316 889808
rect 678237 889750 678316 889752
rect 678237 889747 678303 889750
rect 676029 889402 676095 889405
rect 676029 889400 676292 889402
rect 676029 889344 676034 889400
rect 676090 889344 676292 889400
rect 676029 889342 676292 889344
rect 676029 889339 676095 889342
rect 676029 888994 676095 888997
rect 676029 888992 676292 888994
rect 676029 888936 676034 888992
rect 676090 888936 676292 888992
rect 676029 888934 676292 888936
rect 676029 888931 676095 888934
rect 676029 888586 676095 888589
rect 676029 888584 676292 888586
rect 676029 888528 676034 888584
rect 676090 888528 676292 888584
rect 676029 888526 676292 888528
rect 676029 888523 676095 888526
rect 683113 888178 683179 888181
rect 683100 888176 683179 888178
rect 683100 888120 683118 888176
rect 683174 888120 683179 888176
rect 683100 888118 683179 888120
rect 683113 888115 683179 888118
rect 675886 887708 675892 887772
rect 675956 887770 675962 887772
rect 675956 887710 676292 887770
rect 675956 887708 675962 887710
rect 676029 887362 676095 887365
rect 676029 887360 676292 887362
rect 676029 887304 676034 887360
rect 676090 887304 676292 887360
rect 676029 887302 676292 887304
rect 676029 887299 676095 887302
rect 676029 886954 676095 886957
rect 676029 886952 676292 886954
rect 676029 886896 676034 886952
rect 676090 886896 676292 886952
rect 676029 886894 676292 886896
rect 676029 886891 676095 886894
rect 683070 886138 683130 886516
rect 675894 886108 683130 886138
rect 675894 886078 683100 886108
rect 675702 885804 675708 885868
rect 675772 885866 675778 885868
rect 675894 885866 675954 886078
rect 675772 885806 675954 885866
rect 675772 885804 675778 885806
rect 676029 885730 676095 885733
rect 676029 885728 676292 885730
rect 676029 885672 676034 885728
rect 676090 885672 676292 885728
rect 676029 885670 676292 885672
rect 676029 885667 676095 885670
rect 675518 880636 675524 880700
rect 675588 880698 675594 880700
rect 680997 880698 681063 880701
rect 675588 880696 681063 880698
rect 675588 880640 681002 880696
rect 681058 880640 681063 880696
rect 675588 880638 681063 880640
rect 675588 880636 675594 880638
rect 680997 880635 681063 880638
rect 676438 880364 676444 880428
rect 676508 880426 676514 880428
rect 683113 880426 683179 880429
rect 676508 880424 683179 880426
rect 676508 880368 683118 880424
rect 683174 880368 683179 880424
rect 676508 880366 683179 880368
rect 676508 880364 676514 880366
rect 683113 880363 683179 880366
rect 675334 878460 675340 878524
rect 675404 878522 675410 878524
rect 675753 878522 675819 878525
rect 679617 878522 679683 878525
rect 675404 878520 675819 878522
rect 675404 878464 675758 878520
rect 675814 878464 675819 878520
rect 675404 878462 675819 878464
rect 675404 878460 675410 878462
rect 675753 878459 675819 878462
rect 676032 878520 679683 878522
rect 676032 878464 679622 878520
rect 679678 878464 679683 878520
rect 676032 878462 679683 878464
rect 675385 877978 675451 877981
rect 676032 877978 676092 878462
rect 679617 878459 679683 878462
rect 675385 877976 676092 877978
rect 675385 877920 675390 877976
rect 675446 877920 676092 877976
rect 675385 877918 676092 877920
rect 675385 877915 675451 877918
rect 675334 874108 675340 874172
rect 675404 874170 675410 874172
rect 675569 874170 675635 874173
rect 675404 874168 675635 874170
rect 675404 874112 675574 874168
rect 675630 874112 675635 874168
rect 675404 874110 675635 874112
rect 675404 874108 675410 874110
rect 675569 874107 675635 874110
rect 675753 872810 675819 872813
rect 676438 872810 676444 872812
rect 675753 872808 676444 872810
rect 675753 872752 675758 872808
rect 675814 872752 676444 872808
rect 675753 872750 676444 872752
rect 675753 872747 675819 872750
rect 676438 872748 676444 872750
rect 676508 872748 676514 872812
rect 675753 869818 675819 869821
rect 676254 869818 676260 869820
rect 675753 869816 676260 869818
rect 675753 869760 675758 869816
rect 675814 869760 676260 869816
rect 675753 869758 676260 869760
rect 675753 869755 675819 869758
rect 676254 869756 676260 869758
rect 676324 869756 676330 869820
rect 651465 868594 651531 868597
rect 649950 868592 651531 868594
rect 649950 868536 651470 868592
rect 651526 868536 651531 868592
rect 649950 868534 651531 868536
rect 649950 868246 650010 868534
rect 651465 868531 651531 868534
rect 652017 867642 652083 867645
rect 649950 867640 652083 867642
rect 649950 867584 652022 867640
rect 652078 867584 652083 867640
rect 649950 867582 652083 867584
rect 649950 867064 650010 867582
rect 652017 867579 652083 867582
rect 651465 866282 651531 866285
rect 649950 866280 651531 866282
rect 649950 866224 651470 866280
rect 651526 866224 651531 866280
rect 649950 866222 651531 866224
rect 649950 865882 650010 866222
rect 651465 866219 651531 866222
rect 675293 865738 675359 865741
rect 675702 865738 675708 865740
rect 675293 865736 675708 865738
rect 675293 865680 675298 865736
rect 675354 865680 675708 865736
rect 675293 865678 675708 865680
rect 675293 865675 675359 865678
rect 675702 865676 675708 865678
rect 675772 865676 675778 865740
rect 675753 865466 675819 865469
rect 676070 865466 676076 865468
rect 675753 865464 676076 865466
rect 675753 865408 675758 865464
rect 675814 865408 676076 865464
rect 675753 865406 676076 865408
rect 675753 865403 675819 865406
rect 676070 865404 676076 865406
rect 676140 865404 676146 865468
rect 651373 865194 651439 865197
rect 649950 865192 651439 865194
rect 649950 865136 651378 865192
rect 651434 865136 651439 865192
rect 649950 865134 651439 865136
rect 649950 864700 650010 865134
rect 651373 865131 651439 865134
rect 675661 864922 675727 864925
rect 675886 864922 675892 864924
rect 675661 864920 675892 864922
rect 675661 864864 675666 864920
rect 675722 864864 675892 864920
rect 675661 864862 675892 864864
rect 675661 864859 675727 864862
rect 675886 864860 675892 864862
rect 675956 864860 675962 864924
rect 651465 863834 651531 863837
rect 649766 863832 651531 863834
rect 649766 863776 651470 863832
rect 651526 863776 651531 863832
rect 649766 863774 651531 863776
rect 649766 863518 649826 863774
rect 651465 863771 651531 863774
rect 651465 862338 651531 862341
rect 649766 862336 651531 862338
rect 649766 862280 651470 862336
rect 651526 862280 651531 862336
rect 649766 862278 651531 862280
rect 651465 862275 651531 862278
rect 35617 818002 35683 818005
rect 35574 818000 35683 818002
rect 35574 817944 35622 818000
rect 35678 817944 35683 818000
rect 35574 817939 35683 817944
rect 35574 817700 35634 817939
rect 35801 817322 35867 817325
rect 35788 817320 35867 817322
rect 35788 817264 35806 817320
rect 35862 817264 35867 817320
rect 35788 817262 35867 817264
rect 35801 817259 35867 817262
rect 35433 816914 35499 816917
rect 35420 816912 35499 816914
rect 35420 816856 35438 816912
rect 35494 816856 35499 816912
rect 35420 816854 35499 816856
rect 35433 816851 35499 816854
rect 35801 816098 35867 816101
rect 35788 816096 35867 816098
rect 35788 816040 35806 816096
rect 35862 816040 35867 816096
rect 35788 816038 35867 816040
rect 35801 816035 35867 816038
rect 35617 815282 35683 815285
rect 35604 815280 35683 815282
rect 35604 815224 35622 815280
rect 35678 815224 35683 815280
rect 35604 815222 35683 815224
rect 35617 815219 35683 815222
rect 35801 814466 35867 814469
rect 35788 814464 35867 814466
rect 35788 814408 35806 814464
rect 35862 814408 35867 814464
rect 35788 814406 35867 814408
rect 35801 814403 35867 814406
rect 41321 813650 41387 813653
rect 41308 813648 41387 813650
rect 41308 813592 41326 813648
rect 41382 813592 41387 813648
rect 41308 813590 41387 813592
rect 41321 813587 41387 813590
rect 41822 813242 41828 813244
rect 41492 813182 41828 813242
rect 41822 813180 41828 813182
rect 41892 813180 41898 813244
rect 40953 812834 41019 812837
rect 40940 812832 41019 812834
rect 40940 812776 40958 812832
rect 41014 812776 41019 812832
rect 40940 812774 41019 812776
rect 40953 812771 41019 812774
rect 41137 812426 41203 812429
rect 41124 812424 41203 812426
rect 41124 812368 41142 812424
rect 41198 812368 41203 812424
rect 41124 812366 41203 812368
rect 41137 812363 41203 812366
rect 42006 812018 42012 812020
rect 41492 811958 42012 812018
rect 42006 811956 42012 811958
rect 42076 811956 42082 812020
rect 32397 811610 32463 811613
rect 32397 811608 32476 811610
rect 32397 811552 32402 811608
rect 32458 811552 32476 811608
rect 32397 811550 32476 811552
rect 32397 811547 32463 811550
rect 34513 811202 34579 811205
rect 34500 811200 34579 811202
rect 34500 811144 34518 811200
rect 34574 811144 34579 811200
rect 34500 811142 34579 811144
rect 34513 811139 34579 811142
rect 41965 810794 42031 810797
rect 41492 810792 42031 810794
rect 41492 810736 41970 810792
rect 42026 810736 42031 810792
rect 41492 810734 42031 810736
rect 41965 810731 42031 810734
rect 42149 810386 42215 810389
rect 41492 810384 42215 810386
rect 41492 810328 42154 810384
rect 42210 810328 42215 810384
rect 41492 810326 42215 810328
rect 42149 810323 42215 810326
rect 31017 809978 31083 809981
rect 31004 809976 31083 809978
rect 31004 809920 31022 809976
rect 31078 809920 31083 809976
rect 31004 809918 31083 809920
rect 31017 809915 31083 809918
rect 33777 809570 33843 809573
rect 33764 809568 33843 809570
rect 33764 809512 33782 809568
rect 33838 809512 33843 809568
rect 33764 809510 33843 809512
rect 33777 809507 33843 809510
rect 41781 809162 41847 809165
rect 41492 809160 41847 809162
rect 41492 809104 41786 809160
rect 41842 809104 41847 809160
rect 41492 809102 41847 809104
rect 41781 809099 41847 809102
rect 40953 808754 41019 808757
rect 40940 808752 41019 808754
rect 40940 808696 40958 808752
rect 41014 808696 41019 808752
rect 40940 808694 41019 808696
rect 40953 808691 41019 808694
rect 43253 808346 43319 808349
rect 41492 808344 43319 808346
rect 41492 808288 43258 808344
rect 43314 808288 43319 808344
rect 41492 808286 43319 808288
rect 43253 808283 43319 808286
rect 41137 807938 41203 807941
rect 41124 807936 41203 807938
rect 41124 807880 41142 807936
rect 41198 807880 41203 807936
rect 41124 807878 41203 807880
rect 41137 807875 41203 807878
rect 43805 807530 43871 807533
rect 41492 807528 43871 807530
rect 41492 807472 43810 807528
rect 43866 807472 43871 807528
rect 41492 807470 43871 807472
rect 43805 807467 43871 807470
rect 41094 806717 41154 807092
rect 41094 806712 41203 806717
rect 41094 806684 41142 806712
rect 41124 806656 41142 806684
rect 41198 806656 41203 806712
rect 41124 806654 41203 806656
rect 41137 806651 41203 806654
rect 41321 806306 41387 806309
rect 41308 806304 41387 806306
rect 41308 806248 41326 806304
rect 41382 806248 41387 806304
rect 41308 806246 41387 806248
rect 41321 806243 41387 806246
rect 40534 805564 40540 805628
rect 40604 805626 40610 805628
rect 41965 805626 42031 805629
rect 40604 805624 42031 805626
rect 40604 805568 41970 805624
rect 42026 805568 42031 805624
rect 40604 805566 42031 805568
rect 40604 805564 40610 805566
rect 41965 805563 42031 805566
rect 40953 805220 41019 805221
rect 40902 805218 40908 805220
rect 40862 805158 40908 805218
rect 40972 805216 41019 805220
rect 41014 805160 41019 805216
rect 40902 805156 40908 805158
rect 40972 805156 41019 805160
rect 40953 805155 41019 805156
rect 40718 804884 40724 804948
rect 40788 804946 40794 804948
rect 42149 804946 42215 804949
rect 40788 804944 42215 804946
rect 40788 804888 42154 804944
rect 42210 804888 42215 804944
rect 40788 804886 42215 804888
rect 40788 804884 40794 804886
rect 42149 804883 42215 804886
rect 41597 804676 41663 804677
rect 41597 804674 41644 804676
rect 41552 804672 41644 804674
rect 41552 804616 41602 804672
rect 41552 804614 41644 804616
rect 41597 804612 41644 804614
rect 41708 804612 41714 804676
rect 41597 804611 41663 804612
rect 40677 800594 40743 800597
rect 41086 800594 41092 800596
rect 40677 800592 41092 800594
rect 40677 800536 40682 800592
rect 40738 800536 41092 800592
rect 40677 800534 41092 800536
rect 40677 800531 40743 800534
rect 41086 800532 41092 800534
rect 41156 800532 41162 800596
rect 41781 800322 41847 800325
rect 41781 800320 41890 800322
rect 41781 800264 41786 800320
rect 41842 800264 41890 800320
rect 41781 800259 41890 800264
rect 41830 799917 41890 800259
rect 41781 799912 41890 799917
rect 41781 799856 41786 799912
rect 41842 799856 41890 799912
rect 41781 799854 41890 799856
rect 41781 799851 41847 799854
rect 41086 794412 41092 794476
rect 41156 794474 41162 794476
rect 41781 794474 41847 794477
rect 41156 794472 41847 794474
rect 41156 794416 41786 794472
rect 41842 794416 41847 794472
rect 41156 794414 41847 794416
rect 41156 794412 41162 794414
rect 41781 794411 41847 794414
rect 40902 793460 40908 793524
rect 40972 793522 40978 793524
rect 42425 793522 42491 793525
rect 40972 793520 42491 793522
rect 40972 793464 42430 793520
rect 42486 793464 42491 793520
rect 40972 793462 42491 793464
rect 40972 793460 40978 793462
rect 42425 793459 42491 793462
rect 40718 791964 40724 792028
rect 40788 792026 40794 792028
rect 42241 792026 42307 792029
rect 40788 792024 42307 792026
rect 40788 791968 42246 792024
rect 42302 791968 42307 792024
rect 40788 791966 42307 791968
rect 40788 791964 40794 791966
rect 42241 791963 42307 791966
rect 62205 790530 62271 790533
rect 62205 790528 64706 790530
rect 62205 790472 62210 790528
rect 62266 790472 64706 790528
rect 62205 790470 64706 790472
rect 62205 790467 62271 790470
rect 64646 790304 64706 790470
rect 40534 789516 40540 789580
rect 40604 789578 40610 789580
rect 42517 789578 42583 789581
rect 40604 789576 42583 789578
rect 40604 789520 42522 789576
rect 42578 789520 42583 789576
rect 40604 789518 42583 789520
rect 40604 789516 40610 789518
rect 42517 789515 42583 789518
rect 41638 789244 41644 789308
rect 41708 789306 41714 789308
rect 42609 789306 42675 789309
rect 41708 789304 42675 789306
rect 41708 789248 42614 789304
rect 42670 789248 42675 789304
rect 41708 789246 42675 789248
rect 41708 789244 41714 789246
rect 42609 789243 42675 789246
rect 62113 789170 62179 789173
rect 62113 789168 64706 789170
rect 62113 789112 62118 789168
rect 62174 789112 64706 789168
rect 62113 789110 64706 789112
rect 62113 789107 62179 789110
rect 41454 788836 41460 788900
rect 41524 788898 41530 788900
rect 42241 788898 42307 788901
rect 41524 788896 42307 788898
rect 41524 788840 42246 788896
rect 42302 788840 42307 788896
rect 41524 788838 42307 788840
rect 41524 788836 41530 788838
rect 42241 788835 42307 788838
rect 41873 788628 41939 788629
rect 41822 788626 41828 788628
rect 41782 788566 41828 788626
rect 41892 788624 41939 788628
rect 41934 788568 41939 788624
rect 41822 788564 41828 788566
rect 41892 788564 41939 788568
rect 41873 788563 41939 788564
rect 675753 788082 675819 788085
rect 676070 788082 676076 788084
rect 675753 788080 676076 788082
rect 675753 788024 675758 788080
rect 675814 788024 676076 788080
rect 675753 788022 676076 788024
rect 675753 788019 675819 788022
rect 676070 788020 676076 788022
rect 676140 788020 676146 788084
rect 62113 787402 62179 787405
rect 64646 787402 64706 787940
rect 62113 787400 64706 787402
rect 62113 787344 62118 787400
rect 62174 787344 64706 787400
rect 62113 787342 64706 787344
rect 62113 787339 62179 787342
rect 62941 787130 63007 787133
rect 62941 787128 64706 787130
rect 62941 787072 62946 787128
rect 63002 787072 64706 787128
rect 62941 787070 64706 787072
rect 62941 787067 63007 787070
rect 64646 786758 64706 787070
rect 674414 786660 674420 786724
rect 674484 786722 674490 786724
rect 675109 786722 675175 786725
rect 675385 786724 675451 786725
rect 675334 786722 675340 786724
rect 674484 786720 675175 786722
rect 674484 786664 675114 786720
rect 675170 786664 675175 786720
rect 674484 786662 675175 786664
rect 675294 786662 675340 786722
rect 675404 786720 675451 786724
rect 675446 786664 675451 786720
rect 674484 786660 674490 786662
rect 675109 786659 675175 786662
rect 675334 786660 675340 786662
rect 675404 786660 675451 786664
rect 675385 786659 675451 786660
rect 61377 786178 61443 786181
rect 61377 786176 64706 786178
rect 61377 786120 61382 786176
rect 61438 786120 64706 786176
rect 61377 786118 64706 786120
rect 61377 786115 61443 786118
rect 64646 785576 64706 786118
rect 62113 784954 62179 784957
rect 62113 784952 64706 784954
rect 62113 784896 62118 784952
rect 62174 784896 64706 784952
rect 62113 784894 64706 784896
rect 62113 784891 62179 784894
rect 64646 784394 64706 784894
rect 674373 779378 674439 779381
rect 675477 779378 675543 779381
rect 674373 779376 675543 779378
rect 674373 779320 674378 779376
rect 674434 779320 675482 779376
rect 675538 779320 675543 779376
rect 674373 779318 675543 779320
rect 674373 779315 674439 779318
rect 675477 779315 675543 779318
rect 674557 778834 674623 778837
rect 675477 778834 675543 778837
rect 674557 778832 675543 778834
rect 649950 778426 650010 778824
rect 674557 778776 674562 778832
rect 674618 778776 675482 778832
rect 675538 778776 675543 778832
rect 674557 778774 675543 778776
rect 674557 778771 674623 778774
rect 675477 778771 675543 778774
rect 651465 778426 651531 778429
rect 649950 778424 651531 778426
rect 649950 778368 651470 778424
rect 651526 778368 651531 778424
rect 649950 778366 651531 778368
rect 651465 778363 651531 778366
rect 649950 777066 650010 777642
rect 673269 777474 673335 777477
rect 675385 777474 675451 777477
rect 673269 777472 675451 777474
rect 673269 777416 673274 777472
rect 673330 777416 675390 777472
rect 675446 777416 675451 777472
rect 673269 777414 675451 777416
rect 673269 777411 673335 777414
rect 675385 777411 675451 777414
rect 652017 777066 652083 777069
rect 649950 777064 652083 777066
rect 649950 777008 652022 777064
rect 652078 777008 652083 777064
rect 649950 777006 652083 777008
rect 652017 777003 652083 777006
rect 674925 777066 674991 777069
rect 675477 777066 675543 777069
rect 674925 777064 675543 777066
rect 674925 777008 674930 777064
rect 674986 777008 675482 777064
rect 675538 777008 675543 777064
rect 674925 777006 675543 777008
rect 674925 777003 674991 777006
rect 675477 777003 675543 777006
rect 649950 776114 650010 776460
rect 651465 776114 651531 776117
rect 649950 776112 651531 776114
rect 649950 776056 651470 776112
rect 651526 776056 651531 776112
rect 649950 776054 651531 776056
rect 651465 776051 651531 776054
rect 674925 775706 674991 775709
rect 675385 775706 675451 775709
rect 674925 775704 675451 775706
rect 674925 775648 674930 775704
rect 674986 775648 675390 775704
rect 675446 775648 675451 775704
rect 674925 775646 675451 775648
rect 674925 775643 674991 775646
rect 675385 775643 675451 775646
rect 651373 775298 651439 775301
rect 649950 775296 651439 775298
rect 649950 775240 651378 775296
rect 651434 775240 651439 775296
rect 649950 775238 651439 775240
rect 651373 775235 651439 775238
rect 35801 774754 35867 774757
rect 35758 774752 35867 774754
rect 35758 774696 35806 774752
rect 35862 774696 35867 774752
rect 35758 774691 35867 774696
rect 35758 774452 35818 774691
rect 651465 774210 651531 774213
rect 649950 774208 651531 774210
rect 649950 774152 651470 774208
rect 651526 774152 651531 774208
rect 649950 774150 651531 774152
rect 649950 774096 650010 774150
rect 651465 774147 651531 774150
rect 35390 773941 35450 774044
rect 35341 773936 35450 773941
rect 35341 773880 35346 773936
rect 35402 773880 35450 773936
rect 35341 773878 35450 773880
rect 35341 773875 35407 773878
rect 35758 773533 35818 773636
rect 35525 773530 35591 773533
rect 35525 773528 35634 773530
rect 35525 773472 35530 773528
rect 35586 773472 35634 773528
rect 35525 773467 35634 773472
rect 35758 773528 35867 773533
rect 35758 773472 35806 773528
rect 35862 773472 35867 773528
rect 35758 773470 35867 773472
rect 35801 773467 35867 773470
rect 41689 773530 41755 773533
rect 46197 773530 46263 773533
rect 41689 773528 46263 773530
rect 41689 773472 41694 773528
rect 41750 773472 46202 773528
rect 46258 773472 46263 773528
rect 41689 773470 46263 773472
rect 41689 773467 41755 773470
rect 46197 773467 46263 773470
rect 35574 773228 35634 773467
rect 651465 773394 651531 773397
rect 649950 773392 651531 773394
rect 649950 773336 651470 773392
rect 651526 773336 651531 773392
rect 649950 773334 651531 773336
rect 35801 773122 35867 773125
rect 35758 773120 35867 773122
rect 35758 773064 35806 773120
rect 35862 773064 35867 773120
rect 35758 773059 35867 773064
rect 40769 773122 40835 773125
rect 42977 773122 43043 773125
rect 40769 773120 43043 773122
rect 40769 773064 40774 773120
rect 40830 773064 42982 773120
rect 43038 773064 43043 773120
rect 40769 773062 43043 773064
rect 40769 773059 40835 773062
rect 42977 773059 43043 773062
rect 35758 772820 35818 773059
rect 649950 772914 650010 773334
rect 651465 773331 651531 773334
rect 35758 772309 35818 772412
rect 35758 772304 35867 772309
rect 35758 772248 35806 772304
rect 35862 772248 35867 772304
rect 35758 772246 35867 772248
rect 35801 772243 35867 772246
rect 35574 771901 35634 772004
rect 35574 771896 35683 771901
rect 35574 771840 35622 771896
rect 35678 771840 35683 771896
rect 35574 771838 35683 771840
rect 35617 771835 35683 771838
rect 40217 771898 40283 771901
rect 42793 771898 42859 771901
rect 40217 771896 42859 771898
rect 40217 771840 40222 771896
rect 40278 771840 42798 771896
rect 42854 771840 42859 771896
rect 40217 771838 42859 771840
rect 40217 771835 40283 771838
rect 42793 771835 42859 771838
rect 35758 771493 35818 771596
rect 35758 771488 35867 771493
rect 35758 771432 35806 771488
rect 35862 771432 35867 771488
rect 35758 771430 35867 771432
rect 35801 771427 35867 771430
rect 41045 771490 41111 771493
rect 43437 771490 43503 771493
rect 41045 771488 43503 771490
rect 41045 771432 41050 771488
rect 41106 771432 43442 771488
rect 43498 771432 43503 771488
rect 41045 771430 43503 771432
rect 41045 771427 41111 771430
rect 43437 771427 43503 771430
rect 35758 771085 35818 771188
rect 35758 771080 35867 771085
rect 35758 771024 35806 771080
rect 35862 771024 35867 771080
rect 35758 771022 35867 771024
rect 35801 771019 35867 771022
rect 41505 771082 41571 771085
rect 44449 771082 44515 771085
rect 41505 771080 44515 771082
rect 41505 771024 41510 771080
rect 41566 771024 44454 771080
rect 44510 771024 44515 771080
rect 41505 771022 44515 771024
rect 41505 771019 41571 771022
rect 44449 771019 44515 771022
rect 35574 770677 35634 770780
rect 35574 770672 35683 770677
rect 35574 770616 35622 770672
rect 35678 770616 35683 770672
rect 35574 770614 35683 770616
rect 35617 770611 35683 770614
rect 35758 770269 35818 770372
rect 35758 770264 35867 770269
rect 35758 770208 35806 770264
rect 35862 770208 35867 770264
rect 35758 770206 35867 770208
rect 35801 770203 35867 770206
rect 39849 770266 39915 770269
rect 44265 770266 44331 770269
rect 39849 770264 44331 770266
rect 39849 770208 39854 770264
rect 39910 770208 44270 770264
rect 44326 770208 44331 770264
rect 39849 770206 44331 770208
rect 39849 770203 39915 770206
rect 44265 770203 44331 770206
rect 41462 769858 41522 769964
rect 41638 769858 41644 769860
rect 41462 769798 41644 769858
rect 41638 769796 41644 769798
rect 41708 769796 41714 769860
rect 35758 769453 35818 769556
rect 35758 769448 35867 769453
rect 35758 769392 35806 769448
rect 35862 769392 35867 769448
rect 35758 769390 35867 769392
rect 35801 769387 35867 769390
rect 35574 769045 35634 769148
rect 35525 769040 35634 769045
rect 35801 769042 35867 769045
rect 35525 768984 35530 769040
rect 35586 768984 35634 769040
rect 35525 768982 35634 768984
rect 35758 769040 35867 769042
rect 35758 768984 35806 769040
rect 35862 768984 35867 769040
rect 35525 768979 35591 768982
rect 35758 768979 35867 768984
rect 35758 768740 35818 768979
rect 35206 768229 35266 768332
rect 35157 768224 35266 768229
rect 35157 768168 35162 768224
rect 35218 768168 35266 768224
rect 35157 768166 35266 768168
rect 35157 768163 35223 768166
rect 32446 767821 32506 767924
rect 32397 767816 32506 767821
rect 32397 767760 32402 767816
rect 32458 767760 32506 767816
rect 32397 767758 32506 767760
rect 32397 767755 32463 767758
rect 35758 767413 35818 767516
rect 35758 767408 35867 767413
rect 35758 767352 35806 767408
rect 35862 767352 35867 767408
rect 35758 767350 35867 767352
rect 35801 767347 35867 767350
rect 41229 767410 41295 767413
rect 41454 767410 41460 767412
rect 41229 767408 41460 767410
rect 41229 767352 41234 767408
rect 41290 767352 41460 767408
rect 41229 767350 41460 767352
rect 41229 767347 41295 767350
rect 41454 767348 41460 767350
rect 41524 767348 41530 767412
rect 33734 767005 33794 767108
rect 33734 767000 33843 767005
rect 33734 766944 33782 767000
rect 33838 766944 33843 767000
rect 33734 766942 33843 766944
rect 33777 766939 33843 766942
rect 35801 766594 35867 766597
rect 40726 766596 40786 766700
rect 35758 766592 35867 766594
rect 35758 766536 35806 766592
rect 35862 766536 35867 766592
rect 35758 766531 35867 766536
rect 40718 766532 40724 766596
rect 40788 766532 40794 766596
rect 35758 766292 35818 766531
rect 35758 765781 35818 765884
rect 35758 765776 35867 765781
rect 35758 765720 35806 765776
rect 35862 765720 35867 765776
rect 35758 765718 35867 765720
rect 35801 765715 35867 765718
rect 39757 765778 39823 765781
rect 45001 765778 45067 765781
rect 39757 765776 45067 765778
rect 39757 765720 39762 765776
rect 39818 765720 45006 765776
rect 45062 765720 45067 765776
rect 39757 765718 45067 765720
rect 39757 765715 39823 765718
rect 45001 765715 45067 765718
rect 40542 765372 40602 765476
rect 40534 765308 40540 765372
rect 40604 765308 40610 765372
rect 40910 764964 40970 765068
rect 40902 764900 40908 764964
rect 40972 764900 40978 764964
rect 35758 764557 35818 764660
rect 35758 764552 35867 764557
rect 35758 764496 35806 764552
rect 35862 764496 35867 764552
rect 35758 764494 35867 764496
rect 35801 764491 35867 764494
rect 39389 764554 39455 764557
rect 45185 764554 45251 764557
rect 39389 764552 45251 764554
rect 39389 764496 39394 764552
rect 39450 764496 45190 764552
rect 45246 764496 45251 764552
rect 39389 764494 45251 764496
rect 39389 764491 39455 764494
rect 45185 764491 45251 764494
rect 35574 764149 35634 764252
rect 35574 764144 35683 764149
rect 35574 764088 35622 764144
rect 35678 764088 35683 764144
rect 35574 764086 35683 764088
rect 35617 764083 35683 764086
rect 35801 763738 35867 763741
rect 35758 763736 35867 763738
rect 35758 763680 35806 763736
rect 35862 763680 35867 763736
rect 35758 763675 35867 763680
rect 41689 763738 41755 763741
rect 45369 763738 45435 763741
rect 41689 763736 45435 763738
rect 41689 763680 41694 763736
rect 41750 763680 45374 763736
rect 45430 763680 45435 763736
rect 41689 763678 45435 763680
rect 41689 763675 41755 763678
rect 45369 763675 45435 763678
rect 35758 763436 35818 763675
rect 40953 763330 41019 763333
rect 43253 763330 43319 763333
rect 40953 763328 43319 763330
rect 40953 763272 40958 763328
rect 41014 763272 43258 763328
rect 43314 763272 43319 763328
rect 40953 763270 43319 763272
rect 40953 763267 41019 763270
rect 43253 763267 43319 763270
rect 35758 762925 35818 763028
rect 35758 762920 35867 762925
rect 35758 762864 35806 762920
rect 35862 762864 35867 762920
rect 35758 762862 35867 762864
rect 35801 762859 35867 762862
rect 41689 762922 41755 762925
rect 42425 762922 42491 762925
rect 41689 762920 42491 762922
rect 41689 762864 41694 762920
rect 41750 762864 42430 762920
rect 42486 762864 42491 762920
rect 41689 762862 42491 762864
rect 41689 762859 41755 762862
rect 42425 762859 42491 762862
rect 36537 757754 36603 757757
rect 41822 757754 41828 757756
rect 36537 757752 41828 757754
rect 36537 757696 36542 757752
rect 36598 757696 41828 757752
rect 36537 757694 41828 757696
rect 36537 757691 36603 757694
rect 41822 757692 41828 757694
rect 41892 757692 41898 757756
rect 39205 757346 39271 757349
rect 40350 757346 40356 757348
rect 39205 757344 40356 757346
rect 39205 757288 39210 757344
rect 39266 757288 40356 757344
rect 39205 757286 40356 757288
rect 39205 757283 39271 757286
rect 40350 757284 40356 757286
rect 40420 757284 40426 757348
rect 41781 757074 41847 757077
rect 41781 757072 41890 757074
rect 41781 757016 41786 757072
rect 41842 757016 41890 757072
rect 41781 757011 41890 757016
rect 41830 756669 41890 757011
rect 41830 756664 41939 756669
rect 41830 756608 41878 756664
rect 41934 756608 41939 756664
rect 41830 756606 41939 756608
rect 41873 756603 41939 756606
rect 40902 755788 40908 755852
rect 40972 755850 40978 755852
rect 42333 755850 42399 755853
rect 40972 755848 42399 755850
rect 40972 755792 42338 755848
rect 42394 755792 42399 755848
rect 40972 755790 42399 755792
rect 40972 755788 40978 755790
rect 42333 755787 42399 755790
rect 40350 754972 40356 755036
rect 40420 755034 40426 755036
rect 42793 755034 42859 755037
rect 40420 755032 42859 755034
rect 40420 754976 42798 755032
rect 42854 754976 42859 755032
rect 40420 754974 42859 754976
rect 40420 754972 40426 754974
rect 42793 754971 42859 754974
rect 42057 754082 42123 754085
rect 44725 754082 44791 754085
rect 42057 754080 44791 754082
rect 42057 754024 42062 754080
rect 42118 754024 44730 754080
rect 44786 754024 44791 754080
rect 42057 754022 44791 754024
rect 42057 754019 42123 754022
rect 44725 754019 44791 754022
rect 42149 752994 42215 752997
rect 43621 752994 43687 752997
rect 42149 752992 43687 752994
rect 42149 752936 42154 752992
rect 42210 752936 43626 752992
rect 43682 752936 43687 752992
rect 42149 752934 43687 752936
rect 42149 752931 42215 752934
rect 43621 752931 43687 752934
rect 42057 751770 42123 751773
rect 44817 751770 44883 751773
rect 42057 751768 44883 751770
rect 42057 751712 42062 751768
rect 42118 751712 44822 751768
rect 44878 751712 44883 751768
rect 42057 751710 44883 751712
rect 42057 751707 42123 751710
rect 44817 751707 44883 751710
rect 42149 751226 42215 751229
rect 43989 751226 44055 751229
rect 42149 751224 44055 751226
rect 42149 751168 42154 751224
rect 42210 751168 43994 751224
rect 44050 751168 44055 751224
rect 42149 751166 44055 751168
rect 42149 751163 42215 751166
rect 43989 751163 44055 751166
rect 42149 750954 42215 750957
rect 45185 750954 45251 750957
rect 42149 750952 45251 750954
rect 42149 750896 42154 750952
rect 42210 750896 45190 750952
rect 45246 750896 45251 750952
rect 42149 750894 45251 750896
rect 42149 750891 42215 750894
rect 45185 750891 45251 750894
rect 40534 749396 40540 749460
rect 40604 749458 40610 749460
rect 40604 749398 42074 749458
rect 40604 749396 40610 749398
rect 42014 749189 42074 749398
rect 42014 749184 42123 749189
rect 42014 749128 42062 749184
rect 42118 749128 42123 749184
rect 42014 749126 42123 749128
rect 42057 749123 42123 749126
rect 62941 747690 63007 747693
rect 62941 747688 64706 747690
rect 62941 747632 62946 747688
rect 63002 747632 64706 747688
rect 62941 747630 64706 747632
rect 62941 747627 63007 747630
rect 64646 747082 64706 747630
rect 40718 746812 40724 746876
rect 40788 746874 40794 746876
rect 41781 746874 41847 746877
rect 40788 746872 41847 746874
rect 40788 746816 41786 746872
rect 41842 746816 41847 746872
rect 40788 746814 41847 746816
rect 40788 746812 40794 746814
rect 41781 746811 41847 746814
rect 62113 746194 62179 746197
rect 62113 746192 64706 746194
rect 62113 746136 62118 746192
rect 62174 746136 64706 746192
rect 62113 746134 64706 746136
rect 62113 746131 62179 746134
rect 42057 746058 42123 746061
rect 42701 746058 42767 746061
rect 42057 746056 42767 746058
rect 42057 746000 42062 746056
rect 42118 746000 42706 746056
rect 42762 746000 42767 746056
rect 42057 745998 42767 746000
rect 42057 745995 42123 745998
rect 42701 745995 42767 745998
rect 64646 745900 64706 746134
rect 41822 745316 41828 745380
rect 41892 745378 41898 745380
rect 42425 745378 42491 745381
rect 41892 745376 42491 745378
rect 41892 745320 42430 745376
rect 42486 745320 42491 745376
rect 41892 745318 42491 745320
rect 41892 745316 41898 745318
rect 42425 745315 42491 745318
rect 41454 745044 41460 745108
rect 41524 745106 41530 745108
rect 42609 745106 42675 745109
rect 41524 745104 42675 745106
rect 41524 745048 42614 745104
rect 42670 745048 42675 745104
rect 41524 745046 42675 745048
rect 41524 745044 41530 745046
rect 42609 745043 42675 745046
rect 41638 744772 41644 744836
rect 41708 744834 41714 744836
rect 42241 744834 42307 744837
rect 41708 744832 42307 744834
rect 41708 744776 42246 744832
rect 42302 744776 42307 744832
rect 41708 744774 42307 744776
rect 41708 744772 41714 744774
rect 42241 744771 42307 744774
rect 62113 744154 62179 744157
rect 64646 744154 64706 744718
rect 62113 744152 64706 744154
rect 62113 744096 62118 744152
rect 62174 744096 64706 744152
rect 62113 744094 64706 744096
rect 62113 744091 62179 744094
rect 62113 743746 62179 743749
rect 62113 743744 64706 743746
rect 62113 743688 62118 743744
rect 62174 743688 64706 743744
rect 62113 743686 64706 743688
rect 62113 743683 62179 743686
rect 64646 743536 64706 743686
rect 674230 743276 674236 743340
rect 674300 743338 674306 743340
rect 675109 743338 675175 743341
rect 674300 743336 675175 743338
rect 674300 743280 675114 743336
rect 675170 743280 675175 743336
rect 674300 743278 675175 743280
rect 674300 743276 674306 743278
rect 675109 743275 675175 743278
rect 62113 742386 62179 742389
rect 62113 742384 64706 742386
rect 62113 742328 62118 742384
rect 62174 742328 64706 742384
rect 62113 742326 64706 742328
rect 62113 742323 62179 742326
rect 63033 741842 63099 741845
rect 63033 741840 64706 741842
rect 63033 741784 63038 741840
rect 63094 741784 64706 741840
rect 63033 741782 64706 741784
rect 63033 741779 63099 741782
rect 64646 741172 64706 741782
rect 674598 738108 674604 738172
rect 674668 738170 674674 738172
rect 675109 738170 675175 738173
rect 674668 738168 675175 738170
rect 674668 738112 675114 738168
rect 675170 738112 675175 738168
rect 674668 738110 675175 738112
rect 674668 738108 674674 738110
rect 675109 738107 675175 738110
rect 674005 735042 674071 735045
rect 675477 735042 675543 735045
rect 674005 735040 675543 735042
rect 674005 734984 674010 735040
rect 674066 734984 675482 735040
rect 675538 734984 675543 735040
rect 674005 734982 675543 734984
rect 674005 734979 674071 734982
rect 675477 734979 675543 734982
rect 649950 734226 650010 734402
rect 651465 734226 651531 734229
rect 649950 734224 651531 734226
rect 649950 734168 651470 734224
rect 651526 734168 651531 734224
rect 649950 734166 651531 734168
rect 651465 734163 651531 734166
rect 673453 734226 673519 734229
rect 675477 734226 675543 734229
rect 673453 734224 675543 734226
rect 673453 734168 673458 734224
rect 673514 734168 675482 734224
rect 675538 734168 675543 734224
rect 673453 734166 675543 734168
rect 673453 734163 673519 734166
rect 675477 734163 675543 734166
rect 671245 733818 671311 733821
rect 675477 733818 675543 733821
rect 671245 733816 675543 733818
rect 671245 733760 671250 733816
rect 671306 733760 675482 733816
rect 675538 733760 675543 733816
rect 671245 733758 675543 733760
rect 671245 733755 671311 733758
rect 675477 733755 675543 733758
rect 649950 732866 650010 733220
rect 652661 732866 652727 732869
rect 649950 732864 652727 732866
rect 649950 732808 652666 732864
rect 652722 732808 652727 732864
rect 649950 732806 652727 732808
rect 652661 732803 652727 732806
rect 649950 731778 650010 732038
rect 651465 731778 651531 731781
rect 649950 731776 651531 731778
rect 649950 731720 651470 731776
rect 651526 731720 651531 731776
rect 649950 731718 651531 731720
rect 651465 731715 651531 731718
rect 43621 731370 43687 731373
rect 41492 731368 43687 731370
rect 41492 731312 43626 731368
rect 43682 731312 43687 731368
rect 41492 731310 43687 731312
rect 43621 731307 43687 731310
rect 651373 731098 651439 731101
rect 649950 731096 651439 731098
rect 649950 731040 651378 731096
rect 651434 731040 651439 731096
rect 649950 731038 651439 731040
rect 46197 730962 46263 730965
rect 41492 730960 46263 730962
rect 41492 730904 46202 730960
rect 46258 730904 46263 730960
rect 41492 730902 46263 730904
rect 46197 730899 46263 730902
rect 649950 730856 650010 731038
rect 651373 731035 651439 731038
rect 675293 730828 675359 730829
rect 675293 730826 675340 730828
rect 675248 730824 675340 730826
rect 675248 730768 675298 730824
rect 675248 730766 675340 730768
rect 675293 730764 675340 730766
rect 675404 730764 675410 730828
rect 675293 730763 675359 730764
rect 42241 730554 42307 730557
rect 41492 730552 42307 730554
rect 41492 730496 42246 730552
rect 42302 730496 42307 730552
rect 41492 730494 42307 730496
rect 42241 730491 42307 730494
rect 42977 730146 43043 730149
rect 41492 730144 43043 730146
rect 41492 730088 42982 730144
rect 43038 730088 43043 730144
rect 41492 730086 43043 730088
rect 42977 730083 43043 730086
rect 668853 730146 668919 730149
rect 675477 730146 675543 730149
rect 668853 730144 675543 730146
rect 668853 730088 668858 730144
rect 668914 730088 675482 730144
rect 675538 730088 675543 730144
rect 668853 730086 675543 730088
rect 668853 730083 668919 730086
rect 675477 730083 675543 730086
rect 651465 729874 651531 729877
rect 649950 729872 651531 729874
rect 649950 729816 651470 729872
rect 651526 729816 651531 729872
rect 649950 729814 651531 729816
rect 40953 729738 41019 729741
rect 40940 729736 41019 729738
rect 40940 729680 40958 729736
rect 41014 729680 41019 729736
rect 40940 729678 41019 729680
rect 40953 729675 41019 729678
rect 649950 729674 650010 729814
rect 651465 729811 651531 729814
rect 675109 729874 675175 729877
rect 676806 729874 676812 729876
rect 675109 729872 676812 729874
rect 675109 729816 675114 729872
rect 675170 729816 676812 729872
rect 675109 729814 676812 729816
rect 675109 729811 675175 729814
rect 676806 729812 676812 729814
rect 676876 729812 676882 729876
rect 41137 729330 41203 729333
rect 41124 729328 41203 729330
rect 41124 729272 41142 729328
rect 41198 729272 41203 729328
rect 41124 729270 41203 729272
rect 41137 729267 41203 729270
rect 42885 728922 42951 728925
rect 41492 728920 42951 728922
rect 41492 728864 42890 728920
rect 42946 728864 42951 728920
rect 41492 728862 42951 728864
rect 42885 728859 42951 728862
rect 669405 728786 669471 728789
rect 675477 728786 675543 728789
rect 669405 728784 675543 728786
rect 669405 728728 669410 728784
rect 669466 728728 675482 728784
rect 675538 728728 675543 728784
rect 669405 728726 675543 728728
rect 669405 728723 669471 728726
rect 675477 728723 675543 728726
rect 40861 728684 40927 728687
rect 40861 728682 40970 728684
rect 40861 728626 40866 728682
rect 40922 728626 40970 728682
rect 40861 728621 40970 728626
rect 40910 728484 40970 728621
rect 651465 728514 651531 728517
rect 649950 728512 651531 728514
rect 649950 728456 651470 728512
rect 651526 728456 651531 728512
rect 649950 728454 651531 728456
rect 651465 728451 651531 728454
rect 44173 728106 44239 728109
rect 41492 728104 44239 728106
rect 41492 728048 44178 728104
rect 44234 728048 44239 728104
rect 41492 728046 44239 728048
rect 44173 728043 44239 728046
rect 44541 727698 44607 727701
rect 41492 727696 44607 727698
rect 41492 727640 44546 727696
rect 44602 727640 44607 727696
rect 41492 727638 44607 727640
rect 44541 727635 44607 727638
rect 41321 727460 41387 727463
rect 41278 727458 41387 727460
rect 41278 727402 41326 727458
rect 41382 727402 41387 727458
rect 41278 727397 41387 727402
rect 41278 727260 41338 727397
rect 41137 726882 41203 726885
rect 41124 726880 41203 726882
rect 41124 726824 41142 726880
rect 41198 726824 41203 726880
rect 41124 726822 41203 726824
rect 41137 726819 41203 726822
rect 676070 726548 676076 726612
rect 676140 726610 676146 726612
rect 682377 726610 682443 726613
rect 676140 726608 682443 726610
rect 676140 726552 682382 726608
rect 682438 726552 682443 726608
rect 676140 726550 682443 726552
rect 676140 726548 676146 726550
rect 682377 726547 682443 726550
rect 41278 726239 41338 726444
rect 674414 726276 674420 726340
rect 674484 726338 674490 726340
rect 684217 726338 684283 726341
rect 674484 726336 684283 726338
rect 674484 726280 684222 726336
rect 684278 726280 684283 726336
rect 674484 726278 684283 726280
rect 674484 726276 674490 726278
rect 684217 726275 684283 726278
rect 40953 726236 41019 726239
rect 40910 726234 41019 726236
rect 40910 726178 40958 726234
rect 41014 726178 41019 726234
rect 40910 726173 41019 726178
rect 41278 726234 41387 726239
rect 41278 726178 41326 726234
rect 41382 726178 41387 726234
rect 41278 726176 41387 726178
rect 41321 726173 41387 726176
rect 40910 726036 40970 726173
rect 41781 725796 41847 725797
rect 41781 725794 41828 725796
rect 41736 725792 41828 725794
rect 41736 725736 41786 725792
rect 41736 725734 41828 725736
rect 41781 725732 41828 725734
rect 41892 725732 41898 725796
rect 41781 725731 41847 725732
rect 40769 725658 40835 725661
rect 40756 725656 40835 725658
rect 40756 725600 40774 725656
rect 40830 725600 40835 725656
rect 40756 725598 40835 725600
rect 40769 725595 40835 725598
rect 32397 725250 32463 725253
rect 32397 725248 32476 725250
rect 32397 725192 32402 725248
rect 32458 725192 32476 725248
rect 32397 725190 32476 725192
rect 32397 725187 32463 725190
rect 35157 724842 35223 724845
rect 35157 724840 35236 724842
rect 35157 724784 35162 724840
rect 35218 724784 35236 724840
rect 35157 724782 35236 724784
rect 35157 724779 35223 724782
rect 37273 724434 37339 724437
rect 37260 724432 37339 724434
rect 37260 724376 37278 724432
rect 37334 724376 37339 724432
rect 37260 724374 37339 724376
rect 37273 724371 37339 724374
rect 31661 724026 31727 724029
rect 31661 724024 31740 724026
rect 31661 723968 31666 724024
rect 31722 723968 31740 724024
rect 31661 723966 31740 723968
rect 31661 723963 31727 723966
rect 43437 723618 43503 723621
rect 41492 723616 43503 723618
rect 41492 723560 43442 723616
rect 43498 723560 43503 723616
rect 41492 723558 43503 723560
rect 43437 723555 43503 723558
rect 39297 723210 39363 723213
rect 39284 723208 39363 723210
rect 39284 723152 39302 723208
rect 39358 723152 39363 723208
rect 39284 723150 39363 723152
rect 39297 723147 39363 723150
rect 41781 723076 41847 723077
rect 41781 723072 41828 723076
rect 41892 723074 41898 723076
rect 41781 723016 41786 723072
rect 41781 723012 41828 723016
rect 41892 723014 41938 723074
rect 41892 723012 41898 723014
rect 41781 723011 41847 723012
rect 45277 722802 45343 722805
rect 41492 722800 45343 722802
rect 41492 722744 45282 722800
rect 45338 722744 45343 722800
rect 41492 722742 45343 722744
rect 45277 722739 45343 722742
rect 41781 722394 41847 722397
rect 41492 722392 41847 722394
rect 41492 722336 41786 722392
rect 41842 722336 41847 722392
rect 41492 722334 41847 722336
rect 41781 722331 41847 722334
rect 41965 721986 42031 721989
rect 41492 721984 42031 721986
rect 41492 721928 41970 721984
rect 42026 721928 42031 721984
rect 41492 721926 42031 721928
rect 41965 721923 42031 721926
rect 674005 721716 674071 721717
rect 674005 721712 674052 721716
rect 674116 721714 674122 721716
rect 674925 721714 674991 721717
rect 674005 721656 674010 721712
rect 674005 721652 674052 721656
rect 674116 721654 674162 721714
rect 674925 721712 675034 721714
rect 674925 721656 674930 721712
rect 674986 721656 675034 721712
rect 674116 721652 674122 721654
rect 674005 721651 674071 721652
rect 674925 721651 675034 721656
rect 44173 721578 44239 721581
rect 41492 721576 44239 721578
rect 41492 721520 44178 721576
rect 44234 721520 44239 721576
rect 41492 721518 44239 721520
rect 674974 721578 675034 721651
rect 675334 721578 675340 721580
rect 674974 721518 675340 721578
rect 44173 721515 44239 721518
rect 675334 721516 675340 721518
rect 675404 721516 675410 721580
rect 44909 721170 44975 721173
rect 41492 721168 44975 721170
rect 41492 721112 44914 721168
rect 44970 721112 44975 721168
rect 41492 721110 44975 721112
rect 44909 721107 44975 721110
rect 43621 720354 43687 720357
rect 41492 720352 43687 720354
rect 41492 720296 43626 720352
rect 43682 720296 43687 720352
rect 41492 720294 43687 720296
rect 43621 720291 43687 720294
rect 674005 719812 674071 719813
rect 674005 719810 674052 719812
rect 673960 719808 674052 719810
rect 673960 719752 674010 719808
rect 673960 719750 674052 719752
rect 674005 719748 674052 719750
rect 674116 719748 674122 719812
rect 674005 719747 674071 719748
rect 40769 719266 40835 719269
rect 42701 719266 42767 719269
rect 40769 719264 42767 719266
rect 40769 719208 40774 719264
rect 40830 719208 42706 719264
rect 42762 719208 42767 719264
rect 40769 719206 42767 719208
rect 40769 719203 40835 719206
rect 42701 719203 42767 719206
rect 40534 718524 40540 718588
rect 40604 718586 40610 718588
rect 41781 718586 41847 718589
rect 40604 718584 41847 718586
rect 40604 718528 41786 718584
rect 41842 718528 41847 718584
rect 40604 718526 41847 718528
rect 40604 718524 40610 718526
rect 41781 718523 41847 718526
rect 40718 718252 40724 718316
rect 40788 718314 40794 718316
rect 41965 718314 42031 718317
rect 40788 718312 42031 718314
rect 40788 718256 41970 718312
rect 42026 718256 42031 718312
rect 40788 718254 42031 718256
rect 40788 718252 40794 718254
rect 41965 718251 42031 718254
rect 37273 716954 37339 716957
rect 41822 716954 41828 716956
rect 37273 716952 41828 716954
rect 37273 716896 37278 716952
rect 37334 716896 41828 716952
rect 37273 716894 41828 716896
rect 37273 716891 37339 716894
rect 41822 716892 41828 716894
rect 41892 716892 41898 716956
rect 676029 716546 676095 716549
rect 676029 716544 676292 716546
rect 676029 716488 676034 716544
rect 676090 716488 676292 716544
rect 676029 716486 676292 716488
rect 676029 716483 676095 716486
rect 676029 716138 676095 716141
rect 676029 716136 676292 716138
rect 676029 716080 676034 716136
rect 676090 716080 676292 716136
rect 676029 716078 676292 716080
rect 676029 716075 676095 716078
rect 674005 715730 674071 715733
rect 674005 715728 676292 715730
rect 674005 715672 674010 715728
rect 674066 715672 676292 715728
rect 674005 715670 676292 715672
rect 674005 715667 674071 715670
rect 674005 715322 674071 715325
rect 674005 715320 676292 715322
rect 674005 715264 674010 715320
rect 674066 715264 676292 715320
rect 674005 715262 676292 715264
rect 674005 715259 674071 715262
rect 40401 714914 40467 714917
rect 42149 714914 42215 714917
rect 40401 714912 42215 714914
rect 40401 714856 40406 714912
rect 40462 714856 42154 714912
rect 42210 714856 42215 714912
rect 676029 714914 676095 714917
rect 676029 714912 676292 714914
rect 40401 714854 42215 714856
rect 40401 714851 40467 714854
rect 42149 714851 42215 714854
rect 42701 714870 42767 714873
rect 42701 714868 42810 714870
rect 42701 714812 42706 714868
rect 42762 714812 42810 714868
rect 676029 714856 676034 714912
rect 676090 714856 676292 714912
rect 676029 714854 676292 714856
rect 676029 714851 676095 714854
rect 42701 714807 42810 714812
rect 42750 714644 42810 714807
rect 42742 714580 42748 714644
rect 42812 714580 42818 714644
rect 38009 714506 38075 714509
rect 42374 714506 42380 714508
rect 38009 714504 42380 714506
rect 38009 714448 38014 714504
rect 38070 714448 42380 714504
rect 38009 714446 42380 714448
rect 38009 714443 38075 714446
rect 42374 714444 42380 714446
rect 42444 714444 42450 714508
rect 674005 714506 674071 714509
rect 674005 714504 676292 714506
rect 674005 714448 674010 714504
rect 674066 714448 676292 714504
rect 674005 714446 676292 714448
rect 674005 714443 674071 714446
rect 42149 714234 42215 714237
rect 42149 714232 42442 714234
rect 42149 714176 42154 714232
rect 42210 714176 42442 714232
rect 42149 714174 42442 714176
rect 42149 714171 42215 714174
rect 41781 713962 41847 713965
rect 42190 713962 42196 713964
rect 41781 713960 42196 713962
rect 41781 713904 41786 713960
rect 41842 713904 42196 713960
rect 41781 713902 42196 713904
rect 41781 713899 41847 713902
rect 42190 713900 42196 713902
rect 42260 713900 42266 713964
rect 42149 713554 42215 713557
rect 42382 713554 42442 714174
rect 673085 714098 673151 714101
rect 673085 714096 676292 714098
rect 673085 714040 673090 714096
rect 673146 714040 676292 714096
rect 673085 714038 676292 714040
rect 673085 714035 673151 714038
rect 674005 713690 674071 713693
rect 674005 713688 676292 713690
rect 674005 713632 674010 713688
rect 674066 713632 676292 713688
rect 674005 713630 676292 713632
rect 674005 713627 674071 713630
rect 42149 713552 42442 713554
rect 42149 713496 42154 713552
rect 42210 713496 42442 713552
rect 42149 713494 42442 713496
rect 42149 713491 42215 713494
rect 674005 713282 674071 713285
rect 674005 713280 676292 713282
rect 674005 713224 674010 713280
rect 674066 713224 676292 713280
rect 674005 713222 676292 713224
rect 674005 713219 674071 713222
rect 672901 712874 672967 712877
rect 672901 712872 676292 712874
rect 672901 712816 672906 712872
rect 672962 712816 676292 712872
rect 672901 712814 676292 712816
rect 672901 712811 672967 712814
rect 674005 712466 674071 712469
rect 674005 712464 676292 712466
rect 674005 712408 674010 712464
rect 674066 712408 676292 712464
rect 674005 712406 676292 712408
rect 674005 712403 674071 712406
rect 675293 712058 675359 712061
rect 675293 712056 676292 712058
rect 675293 712000 675298 712056
rect 675354 712000 676292 712056
rect 675293 711998 676292 712000
rect 675293 711995 675359 711998
rect 672717 711650 672783 711653
rect 672717 711648 676292 711650
rect 672717 711592 672722 711648
rect 672778 711592 676292 711648
rect 672717 711590 676292 711592
rect 672717 711587 672783 711590
rect 682377 711242 682443 711245
rect 682364 711240 682443 711242
rect 682364 711184 682382 711240
rect 682438 711184 682443 711240
rect 682364 711182 682443 711184
rect 682377 711179 682443 711182
rect 680997 710834 681063 710837
rect 680997 710832 681076 710834
rect 680997 710776 681002 710832
rect 681058 710776 681076 710832
rect 680997 710774 681076 710776
rect 680997 710771 681063 710774
rect 42241 710428 42307 710429
rect 42190 710426 42196 710428
rect 42150 710366 42196 710426
rect 42260 710424 42307 710428
rect 42302 710368 42307 710424
rect 42190 710364 42196 710366
rect 42260 710364 42307 710368
rect 42241 710363 42307 710364
rect 676029 710426 676095 710429
rect 676029 710424 676292 710426
rect 676029 710368 676034 710424
rect 676090 710368 676292 710424
rect 676029 710366 676292 710368
rect 676029 710363 676095 710366
rect 42701 710020 42767 710021
rect 42701 710018 42748 710020
rect 42656 710016 42748 710018
rect 42656 709960 42706 710016
rect 42656 709958 42748 709960
rect 42701 709956 42748 709958
rect 42812 709956 42818 710020
rect 674005 710018 674071 710021
rect 674005 710016 676292 710018
rect 674005 709960 674010 710016
rect 674066 709960 676292 710016
rect 674005 709958 676292 709960
rect 42701 709955 42767 709956
rect 674005 709955 674071 709958
rect 684217 709610 684283 709613
rect 684204 709608 684283 709610
rect 684204 709552 684222 709608
rect 684278 709552 684283 709608
rect 684204 709550 684283 709552
rect 684217 709547 684283 709550
rect 40718 709412 40724 709476
rect 40788 709474 40794 709476
rect 40788 709414 42258 709474
rect 40788 709412 40794 709414
rect 42198 709205 42258 709414
rect 42198 709200 42307 709205
rect 42198 709144 42246 709200
rect 42302 709144 42307 709200
rect 42198 709142 42307 709144
rect 42241 709139 42307 709142
rect 674005 709202 674071 709205
rect 674005 709200 676292 709202
rect 674005 709144 674010 709200
rect 674066 709144 676292 709200
rect 674005 709142 676292 709144
rect 674005 709139 674071 709142
rect 42057 708930 42123 708933
rect 44173 708930 44239 708933
rect 42057 708928 44239 708930
rect 42057 708872 42062 708928
rect 42118 708872 44178 708928
rect 44234 708872 44239 708928
rect 42057 708870 44239 708872
rect 42057 708867 42123 708870
rect 44173 708867 44239 708870
rect 676029 708794 676095 708797
rect 676029 708792 676292 708794
rect 676029 708736 676034 708792
rect 676090 708736 676292 708792
rect 676029 708734 676292 708736
rect 676029 708731 676095 708734
rect 42057 708386 42123 708389
rect 43989 708386 44055 708389
rect 42057 708384 44055 708386
rect 42057 708328 42062 708384
rect 42118 708328 43994 708384
rect 44050 708328 44055 708384
rect 42057 708326 44055 708328
rect 42057 708323 42123 708326
rect 43989 708323 44055 708326
rect 673269 708386 673335 708389
rect 673269 708384 676292 708386
rect 673269 708328 673274 708384
rect 673330 708328 676292 708384
rect 673269 708326 676292 708328
rect 673269 708323 673335 708326
rect 40534 707916 40540 707980
rect 40604 707978 40610 707980
rect 42190 707978 42196 707980
rect 40604 707918 42196 707978
rect 40604 707916 40610 707918
rect 42190 707916 42196 707918
rect 42260 707916 42266 707980
rect 684033 707978 684099 707981
rect 684020 707976 684099 707978
rect 684020 707920 684038 707976
rect 684094 707920 684099 707976
rect 684020 707918 684099 707920
rect 684033 707915 684099 707918
rect 673729 707570 673795 707573
rect 673729 707568 676292 707570
rect 673729 707512 673734 707568
rect 673790 707512 676292 707568
rect 673729 707510 676292 707512
rect 673729 707507 673795 707510
rect 41965 707434 42031 707437
rect 43621 707434 43687 707437
rect 41965 707432 43687 707434
rect 41965 707376 41970 707432
rect 42026 707376 43626 707432
rect 43682 707376 43687 707432
rect 41965 707374 43687 707376
rect 41965 707371 42031 707374
rect 43621 707371 43687 707374
rect 676029 707162 676095 707165
rect 676029 707160 676292 707162
rect 676029 707104 676034 707160
rect 676090 707104 676292 707160
rect 676029 707102 676292 707104
rect 676029 707099 676095 707102
rect 683389 706754 683455 706757
rect 683389 706752 683468 706754
rect 683389 706696 683394 706752
rect 683450 706696 683468 706752
rect 683389 706694 683468 706696
rect 683389 706691 683455 706694
rect 675845 706346 675911 706349
rect 675845 706344 676292 706346
rect 675845 706288 675850 706344
rect 675906 706288 676292 706344
rect 675845 706286 676292 706288
rect 675845 706283 675911 706286
rect 42425 706212 42491 706213
rect 42374 706210 42380 706212
rect 42334 706150 42380 706210
rect 42444 706208 42491 706212
rect 42486 706152 42491 706208
rect 42374 706148 42380 706150
rect 42444 706148 42491 706152
rect 42425 706147 42491 706148
rect 678470 705530 678530 705908
rect 683113 705530 683179 705533
rect 678470 705528 683179 705530
rect 678470 705500 683118 705528
rect 678500 705472 683118 705500
rect 683174 705472 683179 705528
rect 678500 705470 683179 705472
rect 683113 705467 683179 705470
rect 676029 705122 676095 705125
rect 676029 705120 676292 705122
rect 676029 705064 676034 705120
rect 676090 705064 676292 705120
rect 676029 705062 676292 705064
rect 676029 705059 676095 705062
rect 62113 704442 62179 704445
rect 62113 704440 64706 704442
rect 62113 704384 62118 704440
rect 62174 704384 64706 704440
rect 62113 704382 64706 704384
rect 62113 704379 62179 704382
rect 41965 704306 42031 704309
rect 42190 704306 42196 704308
rect 41965 704304 42196 704306
rect 41965 704248 41970 704304
rect 42026 704248 42196 704304
rect 41965 704246 42196 704248
rect 41965 704243 42031 704246
rect 42190 704244 42196 704246
rect 42260 704244 42266 704308
rect 64646 703860 64706 704382
rect 62113 703354 62179 703357
rect 62113 703352 64706 703354
rect 62113 703296 62118 703352
rect 62174 703296 64706 703352
rect 62113 703294 64706 703296
rect 62113 703291 62179 703294
rect 64646 702678 64706 703294
rect 41822 701796 41828 701860
rect 41892 701858 41898 701860
rect 42241 701858 42307 701861
rect 41892 701856 42307 701858
rect 41892 701800 42246 701856
rect 42302 701800 42307 701856
rect 41892 701798 42307 701800
rect 41892 701796 41898 701798
rect 42241 701795 42307 701798
rect 41638 701524 41644 701588
rect 41708 701586 41714 701588
rect 42517 701586 42583 701589
rect 41708 701584 42583 701586
rect 41708 701528 42522 701584
rect 42578 701528 42583 701584
rect 41708 701526 42583 701528
rect 41708 701524 41714 701526
rect 42517 701523 42583 701526
rect 62941 701314 63007 701317
rect 64646 701314 64706 701496
rect 62941 701312 64706 701314
rect 62941 701256 62946 701312
rect 63002 701256 64706 701312
rect 62941 701254 64706 701256
rect 62941 701251 63007 701254
rect 673729 701178 673795 701181
rect 675109 701178 675175 701181
rect 673729 701176 675175 701178
rect 673729 701120 673734 701176
rect 673790 701120 675114 701176
rect 675170 701120 675175 701176
rect 673729 701118 675175 701120
rect 673729 701115 673795 701118
rect 675109 701115 675175 701118
rect 63125 700906 63191 700909
rect 63125 700904 64706 700906
rect 63125 700848 63130 700904
rect 63186 700848 64706 700904
rect 63125 700846 64706 700848
rect 63125 700843 63191 700846
rect 41454 700436 41460 700500
rect 41524 700498 41530 700500
rect 41781 700498 41847 700501
rect 41524 700496 41847 700498
rect 41524 700440 41786 700496
rect 41842 700440 41847 700496
rect 41524 700438 41847 700440
rect 41524 700436 41530 700438
rect 41781 700435 41847 700438
rect 64646 700314 64706 700846
rect 61377 699682 61443 699685
rect 61377 699680 64706 699682
rect 61377 699624 61382 699680
rect 61438 699624 64706 699680
rect 61377 699622 64706 699624
rect 61377 699619 61443 699622
rect 64646 699132 64706 699622
rect 667657 698322 667723 698325
rect 675109 698322 675175 698325
rect 667657 698320 675175 698322
rect 667657 698264 667662 698320
rect 667718 698264 675114 698320
rect 675170 698264 675175 698320
rect 667657 698262 675175 698264
rect 667657 698259 667723 698262
rect 675109 698259 675175 698262
rect 62205 698050 62271 698053
rect 62205 698048 64706 698050
rect 62205 697992 62210 698048
rect 62266 697992 64706 698048
rect 62205 697990 64706 697992
rect 62205 697987 62271 697990
rect 64646 697950 64706 697990
rect 673177 696962 673243 696965
rect 675109 696962 675175 696965
rect 673177 696960 675175 696962
rect 673177 696904 673182 696960
rect 673238 696904 675114 696960
rect 675170 696904 675175 696960
rect 673177 696902 675175 696904
rect 673177 696899 673243 696902
rect 675109 696899 675175 696902
rect 675477 696828 675543 696829
rect 675477 696824 675524 696828
rect 675588 696826 675594 696828
rect 675477 696768 675482 696824
rect 675477 696764 675524 696768
rect 675588 696766 675634 696826
rect 675588 696764 675594 696766
rect 675477 696763 675543 696764
rect 670877 694922 670943 694925
rect 675109 694922 675175 694925
rect 670877 694920 675175 694922
rect 670877 694864 670882 694920
rect 670938 694864 675114 694920
rect 675170 694864 675175 694920
rect 670877 694862 675175 694864
rect 670877 694859 670943 694862
rect 675109 694859 675175 694862
rect 674414 694588 674420 694652
rect 674484 694650 674490 694652
rect 675109 694650 675175 694653
rect 674484 694648 675175 694650
rect 674484 694592 675114 694648
rect 675170 694592 675175 694648
rect 674484 694590 675175 694592
rect 674484 694588 674490 694590
rect 675109 694587 675175 694590
rect 674005 693018 674071 693021
rect 675477 693018 675543 693021
rect 674005 693016 675543 693018
rect 674005 692960 674010 693016
rect 674066 692960 675482 693016
rect 675538 692960 675543 693016
rect 674005 692958 675543 692960
rect 674005 692955 674071 692958
rect 675477 692955 675543 692958
rect 669037 690570 669103 690573
rect 675109 690570 675175 690573
rect 669037 690568 675175 690570
rect 669037 690512 669042 690568
rect 669098 690512 675114 690568
rect 675170 690512 675175 690568
rect 669037 690510 675175 690512
rect 669037 690507 669103 690510
rect 675109 690507 675175 690510
rect 674005 690298 674071 690301
rect 674925 690298 674991 690301
rect 674005 690296 674991 690298
rect 674005 690240 674010 690296
rect 674066 690240 674930 690296
rect 674986 690240 674991 690296
rect 674005 690238 674991 690240
rect 674005 690235 674071 690238
rect 674925 690235 674991 690238
rect 649950 689482 650010 689980
rect 651465 689482 651531 689485
rect 649950 689480 651531 689482
rect 649950 689424 651470 689480
rect 651526 689424 651531 689480
rect 649950 689422 651531 689424
rect 651465 689419 651531 689422
rect 668393 689482 668459 689485
rect 675109 689482 675175 689485
rect 668393 689480 675175 689482
rect 668393 689424 668398 689480
rect 668454 689424 675114 689480
rect 675170 689424 675175 689480
rect 668393 689422 675175 689424
rect 668393 689419 668459 689422
rect 675109 689419 675175 689422
rect 649980 688802 650562 688828
rect 651649 688802 651715 688805
rect 649980 688800 651715 688802
rect 649980 688768 651654 688800
rect 650502 688744 651654 688768
rect 651710 688744 651715 688800
rect 650502 688742 651715 688744
rect 651649 688739 651715 688742
rect 672993 688802 673059 688805
rect 674925 688802 674991 688805
rect 672993 688800 674991 688802
rect 672993 688744 672998 688800
rect 673054 688744 674930 688800
rect 674986 688744 674991 688800
rect 672993 688742 674991 688744
rect 672993 688739 673059 688742
rect 674925 688739 674991 688742
rect 43437 688122 43503 688125
rect 41492 688120 43503 688122
rect 41492 688064 43442 688120
rect 43498 688064 43503 688120
rect 41492 688062 43503 688064
rect 43437 688059 43503 688062
rect 668209 687850 668275 687853
rect 675109 687850 675175 687853
rect 668209 687848 675175 687850
rect 668209 687792 668214 687848
rect 668270 687792 675114 687848
rect 675170 687792 675175 687848
rect 668209 687790 675175 687792
rect 668209 687787 668275 687790
rect 675109 687787 675175 687790
rect 45461 687714 45527 687717
rect 41492 687712 45527 687714
rect 41492 687656 45466 687712
rect 45522 687656 45527 687712
rect 41492 687654 45527 687656
rect 45461 687651 45527 687654
rect 649950 687442 650010 687616
rect 651465 687442 651531 687445
rect 649950 687440 651531 687442
rect 649950 687384 651470 687440
rect 651526 687384 651531 687440
rect 649950 687382 651531 687384
rect 651465 687379 651531 687382
rect 43437 687306 43503 687309
rect 41492 687304 43503 687306
rect 41492 687248 43442 687304
rect 43498 687248 43503 687304
rect 41492 687246 43503 687248
rect 43437 687243 43503 687246
rect 41137 686898 41203 686901
rect 41124 686896 41203 686898
rect 41124 686840 41142 686896
rect 41198 686840 41203 686896
rect 41124 686838 41203 686840
rect 41137 686835 41203 686838
rect 651465 686762 651531 686765
rect 649950 686760 651531 686762
rect 649950 686704 651470 686760
rect 651526 686704 651531 686760
rect 649950 686702 651531 686704
rect 40953 686490 41019 686493
rect 40940 686488 41019 686490
rect 40940 686432 40958 686488
rect 41014 686432 41019 686488
rect 649950 686434 650010 686702
rect 651465 686699 651531 686702
rect 40940 686430 41019 686432
rect 40953 686427 41019 686430
rect 675293 686220 675359 686221
rect 675293 686218 675340 686220
rect 675248 686216 675340 686218
rect 675248 686160 675298 686216
rect 675248 686158 675340 686160
rect 675293 686156 675340 686158
rect 675404 686156 675410 686220
rect 675293 686155 675359 686156
rect 41278 685915 41338 686052
rect 675017 685946 675083 685949
rect 675518 685946 675524 685948
rect 675017 685944 675524 685946
rect 40769 685912 40835 685915
rect 40726 685910 40835 685912
rect 40726 685854 40774 685910
rect 40830 685854 40835 685910
rect 40726 685849 40835 685854
rect 41278 685910 41387 685915
rect 41278 685854 41326 685910
rect 41382 685854 41387 685910
rect 675017 685888 675022 685944
rect 675078 685888 675524 685944
rect 675017 685886 675524 685888
rect 675017 685883 675083 685886
rect 675518 685884 675524 685886
rect 675588 685884 675594 685948
rect 41278 685852 41387 685854
rect 41321 685849 41387 685852
rect 40726 685644 40786 685849
rect 672809 685674 672875 685677
rect 675477 685674 675543 685677
rect 672809 685672 675543 685674
rect 672809 685616 672814 685672
rect 672870 685616 675482 685672
rect 675538 685616 675543 685672
rect 672809 685614 675543 685616
rect 672809 685611 672875 685614
rect 675477 685611 675543 685614
rect 44357 685266 44423 685269
rect 651465 685266 651531 685269
rect 41492 685264 44423 685266
rect 41492 685208 44362 685264
rect 44418 685208 44423 685264
rect 41492 685206 44423 685208
rect 649950 685264 651531 685266
rect 649950 685208 651470 685264
rect 651526 685208 651531 685264
rect 649950 685206 651531 685208
rect 44357 685203 44423 685206
rect 651465 685203 651531 685206
rect 670601 684994 670667 684997
rect 675477 684994 675543 684997
rect 670601 684992 675543 684994
rect 670601 684936 670606 684992
rect 670662 684936 675482 684992
rect 675538 684936 675543 684992
rect 670601 684934 675543 684936
rect 670601 684931 670667 684934
rect 675477 684931 675543 684934
rect 44357 684858 44423 684861
rect 41492 684856 44423 684858
rect 41492 684800 44362 684856
rect 44418 684800 44423 684856
rect 41492 684798 44423 684800
rect 44357 684795 44423 684798
rect 44633 684450 44699 684453
rect 652569 684450 652635 684453
rect 41492 684448 44699 684450
rect 41492 684392 44638 684448
rect 44694 684392 44699 684448
rect 41492 684390 44699 684392
rect 44633 684387 44699 684390
rect 649950 684448 652635 684450
rect 649950 684392 652574 684448
rect 652630 684392 652635 684448
rect 649950 684390 652635 684392
rect 42977 684178 43043 684181
rect 41784 684176 43043 684178
rect 41784 684120 42982 684176
rect 43038 684120 43043 684176
rect 41784 684118 43043 684120
rect 41784 684042 41844 684118
rect 42977 684115 43043 684118
rect 649950 684070 650010 684390
rect 652569 684387 652635 684390
rect 41492 683982 41844 684042
rect 669773 683906 669839 683909
rect 675477 683906 675543 683909
rect 669773 683904 675543 683906
rect 669773 683848 669778 683904
rect 669834 683848 675482 683904
rect 675538 683848 675543 683904
rect 669773 683846 675543 683848
rect 669773 683843 669839 683846
rect 675477 683843 675543 683846
rect 41094 683466 41154 683604
rect 41086 683402 41092 683466
rect 41156 683402 41162 683466
rect 41321 683464 41387 683467
rect 41278 683462 41387 683464
rect 41278 683406 41326 683462
rect 41382 683406 41387 683462
rect 41278 683401 41387 683406
rect 41278 683196 41338 683401
rect 40953 682818 41019 682821
rect 40940 682816 41019 682818
rect 40940 682760 40958 682816
rect 41014 682760 41019 682816
rect 40940 682758 41019 682760
rect 40953 682755 41019 682758
rect 674230 682620 674236 682684
rect 674300 682682 674306 682684
rect 684125 682682 684191 682685
rect 674300 682680 684191 682682
rect 674300 682624 684130 682680
rect 684186 682624 684191 682680
rect 674300 682622 684191 682624
rect 674300 682620 674306 682622
rect 684125 682619 684191 682622
rect 42609 682410 42675 682413
rect 41492 682408 42675 682410
rect 41492 682352 42614 682408
rect 42670 682352 42675 682408
rect 41492 682350 42675 682352
rect 42609 682347 42675 682350
rect 673453 682410 673519 682413
rect 674741 682410 674807 682413
rect 673453 682408 674807 682410
rect 673453 682352 673458 682408
rect 673514 682352 674746 682408
rect 674802 682352 674807 682408
rect 673453 682350 674807 682352
rect 673453 682347 673519 682350
rect 674741 682347 674807 682350
rect 673453 682138 673519 682141
rect 675477 682138 675543 682141
rect 673453 682136 675543 682138
rect 673453 682080 673458 682136
rect 673514 682080 675482 682136
rect 675538 682080 675543 682136
rect 673453 682078 675543 682080
rect 673453 682075 673519 682078
rect 675477 682075 675543 682078
rect 35157 682002 35223 682005
rect 35157 682000 35236 682002
rect 35157 681944 35162 682000
rect 35218 681944 35236 682000
rect 35157 681942 35236 681944
rect 35157 681939 35223 681942
rect 33041 681594 33107 681597
rect 33028 681592 33107 681594
rect 33028 681536 33046 681592
rect 33102 681536 33107 681592
rect 33028 681534 33107 681536
rect 33041 681531 33107 681534
rect 33777 681186 33843 681189
rect 33764 681184 33843 681186
rect 33764 681128 33782 681184
rect 33838 681128 33843 681184
rect 33764 681126 33843 681128
rect 33777 681123 33843 681126
rect 36537 680778 36603 680781
rect 36524 680776 36603 680778
rect 36524 680720 36542 680776
rect 36598 680720 36603 680776
rect 36524 680718 36603 680720
rect 36537 680715 36603 680718
rect 43621 680370 43687 680373
rect 41492 680368 43687 680370
rect 41492 680312 43626 680368
rect 43682 680312 43687 680368
rect 41492 680310 43687 680312
rect 43621 680307 43687 680310
rect 42793 679962 42859 679965
rect 41492 679960 42859 679962
rect 41492 679904 42798 679960
rect 42854 679904 42859 679960
rect 41492 679902 42859 679904
rect 42793 679899 42859 679902
rect 44173 679554 44239 679557
rect 41492 679552 44239 679554
rect 41492 679496 44178 679552
rect 44234 679496 44239 679552
rect 41492 679494 44239 679496
rect 44173 679491 44239 679494
rect 43989 679146 44055 679149
rect 41492 679144 44055 679146
rect 41492 679088 43994 679144
rect 44050 679088 44055 679144
rect 41492 679086 44055 679088
rect 43989 679083 44055 679086
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 40542 678708 40602 678928
rect 41781 678876 41847 678877
rect 41781 678872 41828 678876
rect 41892 678874 41898 678876
rect 41781 678816 41786 678872
rect 41781 678812 41828 678816
rect 41892 678814 41938 678874
rect 41892 678812 41898 678814
rect 41781 678811 41847 678812
rect 41689 678602 41755 678605
rect 45277 678602 45343 678605
rect 41689 678600 45343 678602
rect 41689 678544 41694 678600
rect 41750 678544 45282 678600
rect 45338 678544 45343 678600
rect 41689 678542 45343 678544
rect 41689 678539 41755 678542
rect 45277 678539 45343 678542
rect 41781 678330 41847 678333
rect 41492 678328 41847 678330
rect 41492 678272 41786 678328
rect 41842 678272 41847 678328
rect 41492 678270 41847 678272
rect 41781 678267 41847 678270
rect 43437 677922 43503 677925
rect 41492 677920 43503 677922
rect 41492 677864 43442 677920
rect 43498 677864 43503 677920
rect 41492 677862 43503 677864
rect 43437 677859 43503 677862
rect 40769 677754 40835 677755
rect 40718 677752 40724 677754
rect 40678 677692 40724 677752
rect 40788 677750 40835 677754
rect 40830 677694 40835 677750
rect 40718 677690 40724 677692
rect 40788 677690 40835 677694
rect 40769 677689 40835 677690
rect 42425 677106 42491 677109
rect 41492 677104 42491 677106
rect 41492 677048 42430 677104
rect 42486 677048 42491 677104
rect 41492 677046 42491 677048
rect 42425 677043 42491 677046
rect 675017 676426 675083 676429
rect 676070 676426 676076 676428
rect 675017 676424 676076 676426
rect 675017 676368 675022 676424
rect 675078 676368 676076 676424
rect 675017 676366 676076 676368
rect 675017 676363 675083 676366
rect 676070 676364 676076 676366
rect 676140 676364 676146 676428
rect 33777 672754 33843 672757
rect 41822 672754 41828 672756
rect 33777 672752 41828 672754
rect 33777 672696 33782 672752
rect 33838 672696 41828 672752
rect 33777 672694 41828 672696
rect 33777 672691 33843 672694
rect 41822 672692 41828 672694
rect 41892 672692 41898 672756
rect 42190 671468 42196 671532
rect 42260 671530 42266 671532
rect 42793 671530 42859 671533
rect 42260 671528 42859 671530
rect 42260 671472 42798 671528
rect 42854 671472 42859 671528
rect 42260 671470 42859 671472
rect 42260 671468 42266 671470
rect 42793 671467 42859 671470
rect 673545 671394 673611 671397
rect 673545 671392 676292 671394
rect 673545 671336 673550 671392
rect 673606 671336 676292 671392
rect 673545 671334 676292 671336
rect 673545 671331 673611 671334
rect 41597 671122 41663 671125
rect 42793 671122 42859 671125
rect 41597 671120 42859 671122
rect 41597 671064 41602 671120
rect 41658 671064 42798 671120
rect 42854 671064 42859 671120
rect 41597 671062 42859 671064
rect 41597 671059 41663 671062
rect 42793 671059 42859 671062
rect 40493 670986 40559 670989
rect 40902 670986 40908 670988
rect 40493 670984 40908 670986
rect 40493 670928 40498 670984
rect 40554 670928 40908 670984
rect 40493 670926 40908 670928
rect 40493 670923 40559 670926
rect 40902 670924 40908 670926
rect 40972 670924 40978 670988
rect 41413 670986 41479 670989
rect 673545 670986 673611 670989
rect 41413 670984 41522 670986
rect 41413 670928 41418 670984
rect 41474 670928 41522 670984
rect 41413 670923 41522 670928
rect 673545 670984 676292 670986
rect 673545 670928 673550 670984
rect 673606 670928 676292 670984
rect 673545 670926 676292 670928
rect 673545 670923 673611 670926
rect 41462 670306 41522 670923
rect 673545 670578 673611 670581
rect 673545 670576 676292 670578
rect 673545 670520 673550 670576
rect 673606 670520 676292 670576
rect 673545 670518 676292 670520
rect 673545 670515 673611 670518
rect 41781 670306 41847 670309
rect 41462 670304 41847 670306
rect 41462 670248 41786 670304
rect 41842 670248 41847 670304
rect 41462 670246 41847 670248
rect 41781 670243 41847 670246
rect 673361 670170 673427 670173
rect 673361 670168 676292 670170
rect 673361 670112 673366 670168
rect 673422 670112 676292 670168
rect 673361 670110 676292 670112
rect 673361 670107 673427 670110
rect 672625 669898 672691 669901
rect 674833 669898 674899 669901
rect 672625 669896 674899 669898
rect 672625 669840 672630 669896
rect 672686 669840 674838 669896
rect 674894 669840 674899 669896
rect 672625 669838 674899 669840
rect 672625 669835 672691 669838
rect 674833 669835 674899 669838
rect 673361 669490 673427 669493
rect 676262 669490 676322 669732
rect 676489 669490 676555 669493
rect 673361 669488 676322 669490
rect 673361 669432 673366 669488
rect 673422 669432 676322 669488
rect 673361 669430 676322 669432
rect 676446 669488 676555 669490
rect 676446 669432 676494 669488
rect 676550 669432 676555 669488
rect 673361 669427 673427 669430
rect 676446 669427 676555 669432
rect 676446 669324 676506 669427
rect 673545 668946 673611 668949
rect 673545 668944 676292 668946
rect 673545 668888 673550 668944
rect 673606 668888 676292 668944
rect 673545 668886 676292 668888
rect 673545 668883 673611 668886
rect 673545 668538 673611 668541
rect 673545 668536 676292 668538
rect 673545 668480 673550 668536
rect 673606 668480 676292 668536
rect 673545 668478 676292 668480
rect 673545 668475 673611 668478
rect 671521 668130 671587 668133
rect 673545 668130 673611 668133
rect 671521 668128 672090 668130
rect 671521 668072 671526 668128
rect 671582 668072 672090 668128
rect 671521 668070 672090 668072
rect 671521 668067 671587 668070
rect 672030 667586 672090 668070
rect 673545 668128 676292 668130
rect 673545 668072 673550 668128
rect 673606 668072 676292 668128
rect 673545 668070 676292 668072
rect 673545 668067 673611 668070
rect 673545 667722 673611 667725
rect 673545 667720 676292 667722
rect 673545 667664 673550 667720
rect 673606 667664 676292 667720
rect 673545 667662 676292 667664
rect 673545 667659 673611 667662
rect 672030 667526 673470 667586
rect 40902 667388 40908 667452
rect 40972 667450 40978 667452
rect 42333 667450 42399 667453
rect 40972 667448 42399 667450
rect 40972 667392 42338 667448
rect 42394 667392 42399 667448
rect 40972 667390 42399 667392
rect 673410 667450 673470 667526
rect 674833 667450 674899 667453
rect 673410 667448 674899 667450
rect 673410 667392 674838 667448
rect 674894 667392 674899 667448
rect 673410 667390 674899 667392
rect 40972 667388 40978 667390
rect 42333 667387 42399 667390
rect 674833 667387 674899 667390
rect 676262 667042 676322 667284
rect 676489 667042 676555 667045
rect 675894 666982 676322 667042
rect 676446 667040 676555 667042
rect 676446 666984 676494 667040
rect 676550 666984 676555 667040
rect 673545 666770 673611 666773
rect 675894 666770 675954 666982
rect 676446 666979 676555 666984
rect 676446 666876 676506 666979
rect 673545 666768 675954 666770
rect 673545 666712 673550 666768
rect 673606 666712 675954 666768
rect 673545 666710 675954 666712
rect 673545 666707 673611 666710
rect 42149 666636 42215 666637
rect 42149 666634 42196 666636
rect 42104 666632 42196 666634
rect 42104 666576 42154 666632
rect 42104 666574 42196 666576
rect 42149 666572 42196 666574
rect 42260 666572 42266 666636
rect 42149 666571 42215 666572
rect 675293 666498 675359 666501
rect 675293 666496 676292 666498
rect 675293 666440 675298 666496
rect 675354 666440 676292 666496
rect 675293 666438 676292 666440
rect 675293 666435 675359 666438
rect 684125 666226 684191 666229
rect 684125 666224 684234 666226
rect 684125 666168 684130 666224
rect 684186 666168 684234 666224
rect 684125 666163 684234 666168
rect 684174 666060 684234 666163
rect 676806 665756 676812 665820
rect 676876 665756 676882 665820
rect 676814 665652 676874 665756
rect 40534 665348 40540 665412
rect 40604 665410 40610 665412
rect 42057 665410 42123 665413
rect 40604 665408 42123 665410
rect 40604 665352 42062 665408
rect 42118 665352 42123 665408
rect 40604 665350 42123 665352
rect 40604 665348 40610 665350
rect 42057 665347 42123 665350
rect 673545 665274 673611 665277
rect 673545 665272 676292 665274
rect 673545 665216 673550 665272
rect 673606 665216 676292 665272
rect 673545 665214 676292 665216
rect 673545 665211 673611 665214
rect 40718 665076 40724 665140
rect 40788 665138 40794 665140
rect 41781 665138 41847 665141
rect 40788 665136 41847 665138
rect 40788 665080 41786 665136
rect 41842 665080 41847 665136
rect 40788 665078 41847 665080
rect 40788 665076 40794 665078
rect 41781 665075 41847 665078
rect 676029 664866 676095 664869
rect 676029 664864 676292 664866
rect 676029 664808 676034 664864
rect 676090 664808 676292 664864
rect 676029 664806 676292 664808
rect 676029 664803 676095 664806
rect 42057 664594 42123 664597
rect 44173 664594 44239 664597
rect 42057 664592 44239 664594
rect 42057 664536 42062 664592
rect 42118 664536 44178 664592
rect 44234 664536 44239 664592
rect 42057 664534 44239 664536
rect 42057 664531 42123 664534
rect 44173 664531 44239 664534
rect 673545 664458 673611 664461
rect 673545 664456 676292 664458
rect 673545 664400 673550 664456
rect 673606 664400 676292 664456
rect 673545 664398 676292 664400
rect 673545 664395 673611 664398
rect 673361 664050 673427 664053
rect 673361 664048 676292 664050
rect 673361 663992 673366 664048
rect 673422 663992 676292 664048
rect 673361 663990 676292 663992
rect 673361 663987 673427 663990
rect 673545 663778 673611 663781
rect 674833 663778 674899 663781
rect 673545 663776 674899 663778
rect 673545 663720 673550 663776
rect 673606 663720 674838 663776
rect 674894 663720 674899 663776
rect 673545 663718 674899 663720
rect 673545 663715 673611 663718
rect 674833 663715 674899 663718
rect 683205 663778 683271 663781
rect 683205 663776 683314 663778
rect 683205 663720 683210 663776
rect 683266 663720 683314 663776
rect 683205 663715 683314 663720
rect 683254 663612 683314 663715
rect 673913 663234 673979 663237
rect 673913 663232 676292 663234
rect 673913 663176 673918 663232
rect 673974 663176 676292 663232
rect 673913 663174 676292 663176
rect 673913 663171 673979 663174
rect 683481 662962 683547 662965
rect 683438 662960 683547 662962
rect 683438 662904 683486 662960
rect 683542 662904 683547 662960
rect 683438 662899 683547 662904
rect 683438 662796 683498 662899
rect 674598 662356 674604 662420
rect 674668 662418 674674 662420
rect 674668 662358 676292 662418
rect 674668 662356 674674 662358
rect 673545 662010 673611 662013
rect 673545 662008 676292 662010
rect 673545 661952 673550 662008
rect 673606 661952 676292 662008
rect 673545 661950 676292 661952
rect 673545 661947 673611 661950
rect 673913 661602 673979 661605
rect 673913 661600 676292 661602
rect 673913 661544 673918 661600
rect 673974 661544 676292 661600
rect 673913 661542 676292 661544
rect 673913 661539 673979 661542
rect 673913 661194 673979 661197
rect 673913 661192 676292 661194
rect 673913 661136 673918 661192
rect 673974 661136 676292 661192
rect 673913 661134 676292 661136
rect 673913 661131 673979 661134
rect 62113 660922 62179 660925
rect 62113 660920 64706 660922
rect 62113 660864 62118 660920
rect 62174 660864 64706 660920
rect 62113 660862 64706 660864
rect 62113 660859 62179 660862
rect 64646 660638 64706 660862
rect 683070 660109 683130 660756
rect 673913 660106 673979 660109
rect 674833 660106 674899 660109
rect 673913 660104 674899 660106
rect 673913 660048 673918 660104
rect 673974 660048 674838 660104
rect 674894 660048 674899 660104
rect 673913 660046 674899 660048
rect 683070 660104 683179 660109
rect 683070 660048 683118 660104
rect 683174 660048 683179 660104
rect 683070 660046 683179 660048
rect 673913 660043 673979 660046
rect 674833 660043 674899 660046
rect 683113 660043 683179 660046
rect 673361 659698 673427 659701
rect 676262 659698 676322 659940
rect 673361 659696 676322 659698
rect 673361 659640 673366 659696
rect 673422 659640 676322 659696
rect 673361 659638 676322 659640
rect 673361 659635 673427 659638
rect 62113 659562 62179 659565
rect 62113 659560 64706 659562
rect 62113 659504 62118 659560
rect 62174 659504 64706 659560
rect 62113 659502 64706 659504
rect 62113 659499 62179 659502
rect 64646 659456 64706 659502
rect 41638 658548 41644 658612
rect 41708 658610 41714 658612
rect 42517 658610 42583 658613
rect 41708 658608 42583 658610
rect 41708 658552 42522 658608
rect 42578 658552 42583 658608
rect 41708 658550 42583 658552
rect 41708 658548 41714 658550
rect 42517 658547 42583 658550
rect 41781 658340 41847 658341
rect 41781 658336 41828 658340
rect 41892 658338 41898 658340
rect 62113 658338 62179 658341
rect 41781 658280 41786 658336
rect 41781 658276 41828 658280
rect 41892 658278 41938 658338
rect 62113 658336 64706 658338
rect 62113 658280 62118 658336
rect 62174 658280 64706 658336
rect 62113 658278 64706 658280
rect 41892 658276 41898 658278
rect 41781 658275 41847 658276
rect 62113 658275 62179 658278
rect 64646 658274 64706 658278
rect 62941 657658 63007 657661
rect 62941 657656 64706 657658
rect 62941 657600 62946 657656
rect 63002 657600 64706 657656
rect 62941 657598 64706 657600
rect 62941 657595 63007 657598
rect 41454 657188 41460 657252
rect 41524 657250 41530 657252
rect 41781 657250 41847 657253
rect 41524 657248 41847 657250
rect 41524 657192 41786 657248
rect 41842 657192 41847 657248
rect 41524 657190 41847 657192
rect 41524 657188 41530 657190
rect 41781 657187 41847 657190
rect 64646 657092 64706 657598
rect 61377 656570 61443 656573
rect 61377 656568 64706 656570
rect 61377 656512 61382 656568
rect 61438 656512 64706 656568
rect 61377 656510 64706 656512
rect 61377 656507 61443 656510
rect 64646 655910 64706 656510
rect 673913 655618 673979 655621
rect 675109 655618 675175 655621
rect 673913 655616 675175 655618
rect 673913 655560 673918 655616
rect 673974 655560 675114 655616
rect 675170 655560 675175 655616
rect 673913 655558 675175 655560
rect 673913 655555 673979 655558
rect 675109 655555 675175 655558
rect 62113 655346 62179 655349
rect 62113 655344 64706 655346
rect 62113 655288 62118 655344
rect 62174 655288 64706 655344
rect 62113 655286 64706 655288
rect 62113 655283 62179 655286
rect 64646 654728 64706 655286
rect 674230 652836 674236 652900
rect 674300 652898 674306 652900
rect 675385 652898 675451 652901
rect 674300 652896 675451 652898
rect 674300 652840 675390 652896
rect 675446 652840 675451 652896
rect 674300 652838 675451 652840
rect 674300 652836 674306 652838
rect 675385 652835 675451 652838
rect 672165 652490 672231 652493
rect 675109 652490 675175 652493
rect 672165 652488 675175 652490
rect 672165 652432 672170 652488
rect 672226 652432 675114 652488
rect 675170 652432 675175 652488
rect 672165 652430 675175 652432
rect 672165 652427 672231 652430
rect 675109 652427 675175 652430
rect 672625 649226 672691 649229
rect 675385 649226 675451 649229
rect 672625 649224 675451 649226
rect 672625 649168 672630 649224
rect 672686 649168 675390 649224
rect 675446 649168 675451 649224
rect 672625 649166 675451 649168
rect 672625 649163 672691 649166
rect 675385 649163 675451 649166
rect 672993 648818 673059 648821
rect 675109 648818 675175 648821
rect 672993 648816 675175 648818
rect 672993 648760 672998 648816
rect 673054 648760 675114 648816
rect 675170 648760 675175 648816
rect 672993 648758 675175 648760
rect 672993 648755 673059 648758
rect 675109 648755 675175 648758
rect 671705 647866 671771 647869
rect 675385 647866 675451 647869
rect 671705 647864 675451 647866
rect 671705 647808 671710 647864
rect 671766 647808 675390 647864
rect 675446 647808 675451 647864
rect 671705 647806 675451 647808
rect 671705 647803 671771 647806
rect 675385 647803 675451 647806
rect 674782 646036 674788 646100
rect 674852 646098 674858 646100
rect 675017 646098 675083 646101
rect 674852 646096 675083 646098
rect 674852 646040 675022 646096
rect 675078 646040 675083 646096
rect 674852 646038 675083 646040
rect 674852 646036 674858 646038
rect 675017 646035 675083 646038
rect 667473 645826 667539 645829
rect 675109 645826 675175 645829
rect 667473 645824 675175 645826
rect 667473 645768 667478 645824
rect 667534 645768 675114 645824
rect 675170 645768 675175 645824
rect 667473 645766 675175 645768
rect 667473 645763 667539 645766
rect 675109 645763 675175 645766
rect 674005 645554 674071 645557
rect 675109 645554 675175 645557
rect 674005 645552 675175 645554
rect 674005 645496 674010 645552
rect 674066 645496 675114 645552
rect 675170 645496 675175 645552
rect 674005 645494 675175 645496
rect 674005 645491 674071 645494
rect 675109 645491 675175 645494
rect 35758 644741 35818 644912
rect 35758 644736 35867 644741
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644678 35867 644680
rect 35801 644675 35867 644678
rect 38518 644333 38578 644504
rect 38518 644328 38627 644333
rect 38518 644272 38566 644328
rect 38622 644272 38627 644328
rect 38518 644270 38627 644272
rect 38561 644267 38627 644270
rect 669589 644330 669655 644333
rect 675293 644330 675359 644333
rect 669589 644328 675359 644330
rect 669589 644272 669594 644328
rect 669650 644272 675298 644328
rect 675354 644272 675359 644328
rect 669589 644270 675359 644272
rect 669589 644267 669655 644270
rect 675293 644267 675359 644270
rect 35390 643925 35450 644096
rect 35341 643920 35450 643925
rect 35341 643864 35346 643920
rect 35402 643864 35450 643920
rect 35341 643862 35450 643864
rect 35341 643859 35407 643862
rect 35574 643517 35634 643688
rect 35525 643512 35634 643517
rect 35801 643514 35867 643517
rect 35525 643456 35530 643512
rect 35586 643456 35634 643512
rect 35525 643454 35634 643456
rect 35758 643512 35867 643514
rect 35758 643456 35806 643512
rect 35862 643456 35867 643512
rect 35525 643451 35591 643454
rect 35758 643451 35867 643456
rect 35758 643280 35818 643451
rect 649950 643242 650010 643558
rect 674005 643514 674071 643517
rect 675293 643514 675359 643517
rect 674005 643512 675359 643514
rect 674005 643456 674010 643512
rect 674066 643456 675298 643512
rect 675354 643456 675359 643512
rect 674005 643454 675359 643456
rect 674005 643451 674071 643454
rect 675293 643451 675359 643454
rect 651465 643242 651531 643245
rect 649950 643240 651531 643242
rect 649950 643184 651470 643240
rect 651526 643184 651531 643240
rect 649950 643182 651531 643184
rect 651465 643179 651531 643182
rect 674005 643106 674071 643109
rect 675109 643106 675175 643109
rect 674005 643104 675175 643106
rect 674005 643048 674010 643104
rect 674066 643048 675114 643104
rect 675170 643048 675175 643104
rect 674005 643046 675175 643048
rect 674005 643043 674071 643046
rect 675109 643043 675175 643046
rect 35390 642701 35450 642872
rect 35390 642696 35499 642701
rect 35801 642698 35867 642701
rect 35390 642640 35438 642696
rect 35494 642640 35499 642696
rect 35390 642638 35499 642640
rect 35433 642635 35499 642638
rect 35758 642696 35867 642698
rect 35758 642640 35806 642696
rect 35862 642640 35867 642696
rect 35758 642635 35867 642640
rect 35758 642464 35818 642635
rect 35617 642290 35683 642293
rect 35574 642288 35683 642290
rect 35574 642232 35622 642288
rect 35678 642232 35683 642288
rect 35574 642227 35683 642232
rect 39941 642290 40007 642293
rect 45277 642290 45343 642293
rect 39941 642288 45343 642290
rect 39941 642232 39946 642288
rect 40002 642232 45282 642288
rect 45338 642232 45343 642288
rect 39941 642230 45343 642232
rect 39941 642227 40007 642230
rect 45277 642227 45343 642230
rect 35574 642056 35634 642227
rect 649950 641882 650010 642376
rect 652017 641882 652083 641885
rect 649950 641880 652083 641882
rect 649950 641824 652022 641880
rect 652078 641824 652083 641880
rect 649950 641822 652083 641824
rect 652017 641819 652083 641822
rect 673913 641746 673979 641749
rect 675293 641746 675359 641749
rect 673913 641744 675359 641746
rect 673913 641688 673918 641744
rect 673974 641688 675298 641744
rect 675354 641688 675359 641744
rect 673913 641686 675359 641688
rect 673913 641683 673979 641686
rect 675293 641683 675359 641686
rect 35390 641477 35450 641648
rect 35341 641472 35450 641477
rect 35341 641416 35346 641472
rect 35402 641416 35450 641472
rect 35341 641414 35450 641416
rect 40125 641474 40191 641477
rect 46197 641474 46263 641477
rect 40125 641472 46263 641474
rect 40125 641416 40130 641472
rect 40186 641416 46202 641472
rect 46258 641416 46263 641472
rect 40125 641414 46263 641416
rect 35341 641411 35407 641414
rect 40125 641411 40191 641414
rect 46197 641411 46263 641414
rect 35574 641069 35634 641240
rect 35525 641064 35634 641069
rect 35801 641066 35867 641069
rect 35525 641008 35530 641064
rect 35586 641008 35634 641064
rect 35525 641006 35634 641008
rect 35758 641064 35867 641066
rect 35758 641008 35806 641064
rect 35862 641008 35867 641064
rect 35525 641003 35591 641006
rect 35758 641003 35867 641008
rect 40585 641066 40651 641069
rect 44541 641066 44607 641069
rect 40585 641064 44607 641066
rect 40585 641008 40590 641064
rect 40646 641008 44546 641064
rect 44602 641008 44607 641064
rect 40585 641006 44607 641008
rect 40585 641003 40651 641006
rect 44541 641003 44607 641006
rect 35758 640832 35818 641003
rect 649950 640794 650010 641194
rect 651465 640794 651531 640797
rect 649950 640792 651531 640794
rect 649950 640736 651470 640792
rect 651526 640736 651531 640792
rect 649950 640734 651531 640736
rect 651465 640731 651531 640734
rect 41454 640596 41460 640660
rect 41524 640596 41530 640660
rect 41462 640424 41522 640596
rect 39941 640250 40007 640253
rect 45277 640250 45343 640253
rect 674833 640252 674899 640253
rect 39941 640248 45343 640250
rect 39941 640192 39946 640248
rect 40002 640192 45282 640248
rect 45338 640192 45343 640248
rect 39941 640190 45343 640192
rect 39941 640187 40007 640190
rect 45277 640187 45343 640190
rect 674782 640188 674788 640252
rect 674852 640250 674899 640252
rect 674852 640248 674944 640250
rect 674894 640192 674944 640248
rect 674852 640190 674944 640192
rect 674852 640188 674899 640190
rect 674833 640187 674899 640188
rect 651373 640114 651439 640117
rect 649950 640112 651439 640114
rect 649950 640056 651378 640112
rect 651434 640056 651439 640112
rect 649950 640054 651439 640056
rect 34470 639845 34530 640016
rect 649950 640012 650010 640054
rect 651373 640051 651439 640054
rect 34421 639840 34530 639845
rect 34421 639784 34426 639840
rect 34482 639784 34530 639840
rect 34421 639782 34530 639784
rect 40309 639842 40375 639845
rect 45093 639842 45159 639845
rect 40309 639840 45159 639842
rect 40309 639784 40314 639840
rect 40370 639784 45098 639840
rect 45154 639784 45159 639840
rect 40309 639782 45159 639784
rect 34421 639779 34487 639782
rect 40309 639779 40375 639782
rect 45093 639779 45159 639782
rect 35758 639437 35818 639608
rect 35758 639432 35867 639437
rect 35758 639376 35806 639432
rect 35862 639376 35867 639432
rect 35758 639374 35867 639376
rect 35801 639371 35867 639374
rect 35758 639029 35818 639200
rect 35758 639024 35867 639029
rect 35758 638968 35806 639024
rect 35862 638968 35867 639024
rect 35758 638966 35867 638968
rect 35801 638963 35867 638966
rect 35574 638621 35634 638792
rect 35574 638616 35683 638621
rect 35574 638560 35622 638616
rect 35678 638560 35683 638616
rect 35574 638558 35683 638560
rect 649766 638618 649826 638830
rect 671337 638754 671403 638757
rect 675477 638754 675543 638757
rect 671337 638752 675543 638754
rect 671337 638696 671342 638752
rect 671398 638696 675482 638752
rect 675538 638696 675543 638752
rect 671337 638694 675543 638696
rect 671337 638691 671403 638694
rect 675477 638691 675543 638694
rect 651465 638618 651531 638621
rect 649766 638616 651531 638618
rect 649766 638560 651470 638616
rect 651526 638560 651531 638616
rect 649766 638558 651531 638560
rect 35617 638555 35683 638558
rect 651465 638555 651531 638558
rect 35758 638213 35818 638384
rect 35758 638208 35867 638213
rect 651649 638210 651715 638213
rect 35758 638152 35806 638208
rect 35862 638152 35867 638208
rect 35758 638150 35867 638152
rect 35801 638147 35867 638150
rect 649950 638208 651715 638210
rect 649950 638152 651654 638208
rect 651710 638152 651715 638208
rect 649950 638150 651715 638152
rect 32446 637805 32506 637976
rect 32397 637800 32506 637805
rect 32397 637744 32402 637800
rect 32458 637744 32506 637800
rect 32397 637742 32506 637744
rect 32397 637739 32463 637742
rect 649950 637648 650010 638150
rect 651649 638147 651715 638150
rect 35206 637397 35266 637568
rect 676070 637468 676076 637532
rect 676140 637530 676146 637532
rect 679617 637530 679683 637533
rect 676140 637528 679683 637530
rect 676140 637472 679622 637528
rect 679678 637472 679683 637528
rect 676140 637470 679683 637472
rect 676140 637468 676146 637470
rect 679617 637467 679683 637470
rect 35157 637392 35266 637397
rect 35157 637336 35162 637392
rect 35218 637336 35266 637392
rect 35157 637334 35266 637336
rect 35157 637331 35223 637334
rect 35758 636989 35818 637160
rect 35758 636984 35867 636989
rect 35758 636928 35806 636984
rect 35862 636928 35867 636984
rect 35758 636926 35867 636928
rect 35801 636923 35867 636926
rect 35574 636581 35634 636752
rect 35525 636576 35634 636581
rect 35801 636578 35867 636581
rect 35525 636520 35530 636576
rect 35586 636520 35634 636576
rect 35525 636518 35634 636520
rect 35758 636576 35867 636578
rect 35758 636520 35806 636576
rect 35862 636520 35867 636576
rect 35525 636515 35591 636518
rect 35758 636515 35867 636520
rect 35758 636344 35818 636515
rect 39113 636170 39179 636173
rect 44357 636170 44423 636173
rect 39113 636168 44423 636170
rect 39113 636112 39118 636168
rect 39174 636112 44362 636168
rect 44418 636112 44423 636168
rect 39113 636110 44423 636112
rect 39113 636107 39179 636110
rect 44357 636107 44423 636110
rect 35758 635765 35818 635936
rect 35758 635760 35867 635765
rect 35758 635704 35806 635760
rect 35862 635704 35867 635760
rect 35758 635702 35867 635704
rect 35801 635699 35867 635702
rect 40493 635762 40559 635765
rect 43989 635762 44055 635765
rect 40493 635760 44055 635762
rect 40493 635704 40498 635760
rect 40554 635704 43994 635760
rect 44050 635704 44055 635760
rect 40493 635702 44055 635704
rect 40493 635699 40559 635702
rect 43989 635699 44055 635702
rect 40542 635356 40602 635528
rect 40534 635292 40540 635356
rect 40604 635292 40610 635356
rect 40726 634948 40786 635120
rect 40718 634884 40724 634948
rect 40788 634884 40794 634948
rect 35758 634541 35818 634712
rect 35758 634536 35867 634541
rect 35758 634480 35806 634536
rect 35862 634480 35867 634536
rect 35758 634478 35867 634480
rect 35801 634475 35867 634478
rect 40309 634538 40375 634541
rect 42701 634538 42767 634541
rect 40309 634536 42767 634538
rect 40309 634480 40314 634536
rect 40370 634480 42706 634536
rect 42762 634480 42767 634536
rect 40309 634478 42767 634480
rect 40309 634475 40375 634478
rect 42701 634475 42767 634478
rect 35758 633725 35818 633896
rect 35758 633720 35867 633725
rect 35758 633664 35806 633720
rect 35862 633664 35867 633720
rect 35758 633662 35867 633664
rect 35801 633659 35867 633662
rect 39757 633722 39823 633725
rect 43621 633722 43687 633725
rect 39757 633720 43687 633722
rect 39757 633664 39762 633720
rect 39818 633664 43626 633720
rect 43682 633664 43687 633720
rect 39757 633662 43687 633664
rect 39757 633659 39823 633662
rect 43621 633659 43687 633662
rect 41505 633314 41571 633317
rect 42057 633314 42123 633317
rect 41505 633312 42123 633314
rect 41505 633256 41510 633312
rect 41566 633256 42062 633312
rect 42118 633256 42123 633312
rect 41505 633254 42123 633256
rect 41505 633251 41571 633254
rect 42057 633251 42123 633254
rect 40861 632362 40927 632365
rect 43069 632362 43135 632365
rect 40861 632360 43135 632362
rect 40861 632304 40866 632360
rect 40922 632304 43074 632360
rect 43130 632304 43135 632360
rect 40861 632302 43135 632304
rect 40861 632299 40927 632302
rect 43069 632299 43135 632302
rect 675150 631348 675156 631412
rect 675220 631410 675226 631412
rect 675477 631410 675543 631413
rect 675220 631408 675543 631410
rect 675220 631352 675482 631408
rect 675538 631352 675543 631408
rect 675220 631350 675543 631352
rect 675220 631348 675226 631350
rect 675477 631347 675543 631350
rect 675661 631410 675727 631413
rect 676070 631410 676076 631412
rect 675661 631408 676076 631410
rect 675661 631352 675666 631408
rect 675722 631352 676076 631408
rect 675661 631350 676076 631352
rect 675661 631347 675727 631350
rect 676070 631348 676076 631350
rect 676140 631348 676146 631412
rect 40493 630594 40559 630597
rect 42885 630594 42951 630597
rect 40493 630592 42951 630594
rect 40493 630536 40498 630592
rect 40554 630536 42890 630592
rect 42946 630536 42951 630592
rect 40493 630534 42951 630536
rect 40493 630531 40559 630534
rect 42885 630531 42951 630534
rect 40033 630322 40099 630325
rect 42517 630322 42583 630325
rect 40033 630320 42583 630322
rect 40033 630264 40038 630320
rect 40094 630264 42522 630320
rect 42578 630264 42583 630320
rect 40033 630262 42583 630264
rect 40033 630259 40099 630262
rect 42517 630259 42583 630262
rect 32397 629914 32463 629917
rect 41638 629914 41644 629916
rect 32397 629912 41644 629914
rect 32397 629856 32402 629912
rect 32458 629856 41644 629912
rect 32397 629854 41644 629856
rect 32397 629851 32463 629854
rect 41638 629852 41644 629854
rect 41708 629852 41714 629916
rect 39297 629234 39363 629237
rect 41822 629234 41828 629236
rect 39297 629232 41828 629234
rect 39297 629176 39302 629232
rect 39358 629176 41828 629232
rect 39297 629174 41828 629176
rect 39297 629171 39363 629174
rect 41822 629172 41828 629174
rect 41892 629172 41898 629236
rect 40493 628418 40559 628421
rect 42333 628418 42399 628421
rect 40493 628416 42399 628418
rect 40493 628360 40498 628416
rect 40554 628360 42338 628416
rect 42394 628360 42399 628416
rect 40493 628358 42399 628360
rect 40493 628355 40559 628358
rect 42333 628355 42399 628358
rect 41781 627464 41847 627469
rect 41781 627408 41786 627464
rect 41842 627408 41847 627464
rect 41781 627403 41847 627408
rect 41784 627197 41844 627403
rect 41781 627192 41847 627197
rect 41781 627136 41786 627192
rect 41842 627136 41847 627192
rect 41781 627131 41847 627136
rect 674005 626378 674071 626381
rect 674005 626376 676292 626378
rect 674005 626320 674010 626376
rect 674066 626320 676292 626376
rect 674005 626318 676292 626320
rect 674005 626315 674071 626318
rect 673545 625970 673611 625973
rect 674741 625970 674807 625973
rect 673545 625968 674807 625970
rect 673545 625912 673550 625968
rect 673606 625912 674746 625968
rect 674802 625912 674807 625968
rect 673545 625910 674807 625912
rect 673545 625907 673611 625910
rect 674741 625907 674807 625910
rect 676262 625698 676322 625940
rect 676489 625698 676555 625701
rect 674238 625638 676322 625698
rect 676446 625696 676555 625698
rect 676446 625640 676494 625696
rect 676550 625640 676555 625696
rect 674005 625562 674071 625565
rect 674238 625562 674298 625638
rect 674005 625560 674298 625562
rect 674005 625504 674010 625560
rect 674066 625504 674298 625560
rect 676446 625635 676555 625640
rect 676446 625532 676506 625635
rect 674005 625502 674298 625504
rect 674005 625499 674071 625502
rect 676170 625094 676292 625154
rect 674005 625018 674071 625021
rect 676170 625018 676230 625094
rect 674005 625016 676230 625018
rect 674005 624960 674010 625016
rect 674066 624960 676230 625016
rect 674005 624958 676230 624960
rect 674005 624955 674071 624958
rect 674005 624746 674071 624749
rect 674005 624744 676292 624746
rect 674005 624688 674010 624744
rect 674066 624688 676292 624744
rect 674005 624686 676292 624688
rect 674005 624683 674071 624686
rect 674005 624338 674071 624341
rect 674005 624336 676292 624338
rect 674005 624280 674010 624336
rect 674066 624280 676292 624336
rect 674005 624278 676292 624280
rect 674005 624275 674071 624278
rect 674005 623930 674071 623933
rect 674005 623928 676292 623930
rect 674005 623872 674010 623928
rect 674066 623872 676292 623928
rect 674005 623870 676292 623872
rect 674005 623867 674071 623870
rect 674005 623522 674071 623525
rect 674005 623520 676292 623522
rect 674005 623464 674010 623520
rect 674066 623464 676292 623520
rect 674005 623462 676292 623464
rect 674005 623459 674071 623462
rect 674005 623114 674071 623117
rect 674005 623112 676292 623114
rect 674005 623056 674010 623112
rect 674066 623056 676292 623112
rect 674005 623054 676292 623056
rect 674005 623051 674071 623054
rect 674005 622706 674071 622709
rect 674005 622704 676292 622706
rect 674005 622648 674010 622704
rect 674066 622648 676292 622704
rect 674005 622646 676292 622648
rect 674005 622643 674071 622646
rect 674005 622298 674071 622301
rect 674005 622296 676292 622298
rect 674005 622240 674010 622296
rect 674066 622240 676292 622296
rect 674005 622238 676292 622240
rect 674005 622235 674071 622238
rect 40718 621964 40724 622028
rect 40788 622026 40794 622028
rect 41781 622026 41847 622029
rect 679617 622026 679683 622029
rect 40788 622024 41847 622026
rect 40788 621968 41786 622024
rect 41842 621968 41847 622024
rect 40788 621966 41847 621968
rect 40788 621964 40794 621966
rect 41781 621963 41847 621966
rect 679574 622024 679683 622026
rect 679574 621968 679622 622024
rect 679678 621968 679683 622024
rect 679574 621963 679683 621968
rect 679574 621860 679634 621963
rect 672809 621482 672875 621485
rect 672809 621480 676292 621482
rect 672809 621424 672814 621480
rect 672870 621424 676292 621480
rect 672809 621422 676292 621424
rect 672809 621419 672875 621422
rect 674005 621210 674071 621213
rect 674005 621208 676322 621210
rect 674005 621152 674010 621208
rect 674066 621152 676322 621208
rect 674005 621150 676322 621152
rect 674005 621147 674071 621150
rect 676262 621044 676322 621150
rect 40534 620740 40540 620804
rect 40604 620802 40610 620804
rect 41781 620802 41847 620805
rect 40604 620800 41847 620802
rect 40604 620744 41786 620800
rect 41842 620744 41847 620800
rect 40604 620742 41847 620744
rect 40604 620740 40610 620742
rect 41781 620739 41847 620742
rect 672533 620666 672599 620669
rect 672533 620664 676292 620666
rect 672533 620608 672538 620664
rect 672594 620608 676292 620664
rect 672533 620606 676292 620608
rect 672533 620603 672599 620606
rect 673637 620258 673703 620261
rect 673637 620256 676292 620258
rect 673637 620200 673642 620256
rect 673698 620200 676292 620256
rect 673637 620198 676292 620200
rect 673637 620195 673703 620198
rect 673637 619850 673703 619853
rect 673637 619848 676292 619850
rect 673637 619792 673642 619848
rect 673698 619792 676292 619848
rect 673637 619790 676292 619792
rect 673637 619787 673703 619790
rect 673177 619442 673243 619445
rect 673177 619440 676292 619442
rect 673177 619384 673182 619440
rect 673238 619384 676292 619440
rect 673177 619382 676292 619384
rect 673177 619379 673243 619382
rect 673637 619170 673703 619173
rect 674281 619170 674347 619173
rect 673637 619168 674347 619170
rect 673637 619112 673642 619168
rect 673698 619112 674286 619168
rect 674342 619112 674347 619168
rect 673637 619110 674347 619112
rect 673637 619107 673703 619110
rect 674281 619107 674347 619110
rect 674414 618972 674420 619036
rect 674484 619034 674490 619036
rect 674484 618974 676292 619034
rect 674484 618972 674490 618974
rect 683205 618762 683271 618765
rect 683205 618760 683314 618762
rect 683205 618704 683210 618760
rect 683266 618704 683314 618760
rect 683205 618699 683314 618704
rect 683254 618596 683314 618699
rect 673637 618218 673703 618221
rect 673637 618216 676292 618218
rect 673637 618160 673642 618216
rect 673698 618160 676292 618216
rect 673637 618158 676292 618160
rect 673637 618155 673703 618158
rect 63125 618082 63191 618085
rect 63125 618080 64706 618082
rect 63125 618024 63130 618080
rect 63186 618024 64706 618080
rect 63125 618022 64706 618024
rect 63125 618019 63191 618022
rect 64646 617416 64706 618022
rect 673637 617810 673703 617813
rect 673637 617808 676292 617810
rect 673637 617752 673642 617808
rect 673698 617752 676292 617808
rect 673637 617750 676292 617752
rect 673637 617747 673703 617750
rect 676213 617538 676279 617541
rect 676213 617536 676322 617538
rect 676213 617480 676218 617536
rect 676274 617480 676322 617536
rect 676213 617475 676322 617480
rect 676262 617372 676322 617475
rect 675293 617130 675359 617133
rect 676806 617130 676812 617132
rect 675293 617128 676812 617130
rect 675293 617072 675298 617128
rect 675354 617072 676812 617128
rect 675293 617070 676812 617072
rect 675293 617067 675359 617070
rect 676806 617068 676812 617070
rect 676876 617068 676882 617132
rect 683573 617130 683639 617133
rect 683573 617128 683682 617130
rect 683573 617072 683578 617128
rect 683634 617072 683682 617128
rect 683573 617067 683682 617072
rect 683622 616964 683682 617067
rect 683389 616722 683455 616725
rect 683389 616720 683498 616722
rect 683389 616664 683394 616720
rect 683450 616664 683498 616720
rect 683389 616659 683498 616664
rect 62113 616586 62179 616589
rect 62113 616584 64706 616586
rect 62113 616528 62118 616584
rect 62174 616528 64706 616584
rect 683438 616556 683498 616659
rect 62113 616526 64706 616528
rect 62113 616523 62179 616526
rect 64646 616234 64706 616526
rect 673862 616116 673868 616180
rect 673932 616178 673938 616180
rect 673932 616118 676292 616178
rect 673932 616116 673938 616118
rect 41454 615980 41460 616044
rect 41524 616042 41530 616044
rect 41873 616042 41939 616045
rect 41524 616040 41939 616042
rect 41524 615984 41878 616040
rect 41934 615984 41939 616040
rect 41524 615982 41939 615984
rect 41524 615980 41530 615982
rect 41873 615979 41939 615982
rect 42057 615906 42123 615909
rect 42701 615906 42767 615909
rect 42057 615904 42767 615906
rect 42057 615848 42062 615904
rect 42118 615848 42706 615904
rect 42762 615848 42767 615904
rect 42057 615846 42767 615848
rect 42057 615843 42123 615846
rect 42701 615843 42767 615846
rect 683070 615501 683130 615740
rect 41822 615436 41828 615500
rect 41892 615498 41898 615500
rect 42609 615498 42675 615501
rect 41892 615496 42675 615498
rect 41892 615440 42614 615496
rect 42670 615440 42675 615496
rect 41892 615438 42675 615440
rect 41892 615436 41898 615438
rect 42609 615435 42675 615438
rect 673637 615498 673703 615501
rect 674281 615498 674347 615501
rect 673637 615496 674347 615498
rect 673637 615440 673642 615496
rect 673698 615440 674286 615496
rect 674342 615440 674347 615496
rect 673637 615438 674347 615440
rect 673637 615435 673703 615438
rect 674281 615435 674347 615438
rect 683070 615498 683179 615501
rect 683070 615496 683260 615498
rect 683070 615440 683118 615496
rect 683174 615440 683260 615496
rect 683070 615438 683260 615440
rect 683070 615435 683179 615438
rect 683070 615332 683130 615435
rect 62113 614682 62179 614685
rect 64646 614682 64706 615052
rect 673637 614954 673703 614957
rect 673637 614952 676292 614954
rect 673637 614896 673642 614952
rect 673698 614896 676292 614952
rect 673637 614894 676292 614896
rect 673637 614891 673703 614894
rect 62113 614680 64706 614682
rect 62113 614624 62118 614680
rect 62174 614624 64706 614680
rect 62113 614622 64706 614624
rect 62113 614619 62179 614622
rect 61377 613866 61443 613869
rect 64646 613866 64706 613870
rect 61377 613864 64706 613866
rect 61377 613808 61382 613864
rect 61438 613808 64706 613864
rect 61377 613806 64706 613808
rect 61377 613803 61443 613806
rect 41873 613460 41939 613461
rect 41822 613458 41828 613460
rect 41782 613398 41828 613458
rect 41892 613456 41939 613460
rect 41934 613400 41939 613456
rect 41822 613396 41828 613398
rect 41892 613396 41939 613400
rect 41873 613395 41939 613396
rect 62113 612642 62179 612645
rect 64646 612642 64706 612688
rect 62113 612640 64706 612642
rect 62113 612584 62118 612640
rect 62174 612584 64706 612640
rect 62113 612582 64706 612584
rect 62113 612579 62179 612582
rect 40534 612308 40540 612372
rect 40604 612370 40610 612372
rect 42241 612370 42307 612373
rect 40604 612368 42307 612370
rect 40604 612312 42246 612368
rect 42302 612312 42307 612368
rect 40604 612310 42307 612312
rect 40604 612308 40610 612310
rect 42241 612307 42307 612310
rect 43253 612234 43319 612237
rect 43868 612234 43934 612237
rect 43253 612232 43934 612234
rect 43253 612176 43258 612232
rect 43314 612176 43873 612232
rect 43929 612176 43934 612232
rect 43253 612174 43934 612176
rect 43253 612171 43319 612174
rect 43868 612171 43934 612174
rect 62941 612098 63007 612101
rect 62941 612096 64706 612098
rect 62941 612040 62946 612096
rect 63002 612040 64706 612096
rect 62941 612038 64706 612040
rect 62941 612035 63007 612038
rect 44265 611690 44331 611693
rect 46197 611690 46263 611693
rect 44265 611688 46263 611690
rect 44265 611632 44270 611688
rect 44326 611632 46202 611688
rect 46258 611632 46263 611688
rect 44265 611630 46263 611632
rect 44265 611627 44331 611630
rect 46197 611627 46263 611630
rect 64646 611506 64706 612038
rect 44081 611418 44147 611421
rect 64137 611418 64203 611421
rect 44081 611416 64203 611418
rect 44081 611360 44086 611416
rect 44142 611360 64142 611416
rect 64198 611360 64203 611416
rect 44081 611358 64203 611360
rect 44081 611355 44147 611358
rect 64137 611355 64203 611358
rect 673637 611418 673703 611421
rect 675293 611418 675359 611421
rect 673637 611416 675359 611418
rect 673637 611360 673642 611416
rect 673698 611360 675298 611416
rect 675354 611360 675359 611416
rect 673637 611358 675359 611360
rect 673637 611355 673703 611358
rect 675293 611355 675359 611358
rect 672165 609106 672231 609109
rect 674281 609106 674347 609109
rect 672165 609104 674347 609106
rect 672165 609048 672170 609104
rect 672226 609048 674286 609104
rect 674342 609048 674347 609104
rect 672165 609046 674347 609048
rect 672165 609043 672231 609046
rect 674281 609043 674347 609046
rect 671153 608562 671219 608565
rect 675017 608562 675083 608565
rect 671153 608560 675083 608562
rect 671153 608504 671158 608560
rect 671214 608504 675022 608560
rect 675078 608504 675083 608560
rect 671153 608502 675083 608504
rect 671153 608499 671219 608502
rect 675017 608499 675083 608502
rect 673177 608290 673243 608293
rect 674925 608290 674991 608293
rect 673177 608288 674991 608290
rect 673177 608232 673182 608288
rect 673238 608232 674930 608288
rect 674986 608232 674991 608288
rect 673177 608230 674991 608232
rect 673177 608227 673243 608230
rect 674925 608227 674991 608230
rect 672349 604346 672415 604349
rect 675109 604346 675175 604349
rect 672349 604344 675175 604346
rect 672349 604288 672354 604344
rect 672410 604288 675114 604344
rect 675170 604288 675175 604344
rect 672349 604286 675175 604288
rect 672349 604283 672415 604286
rect 675109 604283 675175 604286
rect 674414 602924 674420 602988
rect 674484 602986 674490 602988
rect 675109 602986 675175 602989
rect 674484 602984 675175 602986
rect 674484 602928 675114 602984
rect 675170 602928 675175 602984
rect 674484 602926 675175 602928
rect 674484 602924 674490 602926
rect 675109 602923 675175 602926
rect 40309 602034 40375 602037
rect 40534 602034 40540 602036
rect 40309 602032 40540 602034
rect 40309 601976 40314 602032
rect 40370 601976 40540 602032
rect 40309 601974 40540 601976
rect 40309 601971 40375 601974
rect 40534 601972 40540 601974
rect 40604 601972 40610 602036
rect 35801 601762 35867 601765
rect 35788 601760 35867 601762
rect 35788 601704 35806 601760
rect 35862 601704 35867 601760
rect 35788 601702 35867 601704
rect 35801 601699 35867 601702
rect 39941 601354 40007 601357
rect 39941 601352 40020 601354
rect 39941 601296 39946 601352
rect 40002 601296 40020 601352
rect 39941 601294 40020 601296
rect 39941 601291 40007 601294
rect 40125 600946 40191 600949
rect 667289 600946 667355 600949
rect 675385 600946 675451 600949
rect 40125 600944 40204 600946
rect 40125 600888 40130 600944
rect 40186 600888 40204 600944
rect 40125 600886 40204 600888
rect 667289 600944 675451 600946
rect 667289 600888 667294 600944
rect 667350 600888 675390 600944
rect 675446 600888 675451 600944
rect 667289 600886 675451 600888
rect 40125 600883 40191 600886
rect 667289 600883 667355 600886
rect 675385 600883 675451 600886
rect 673821 600674 673887 600677
rect 674281 600674 674347 600677
rect 673821 600672 674347 600674
rect 673821 600616 673826 600672
rect 673882 600616 674286 600672
rect 674342 600616 674347 600672
rect 673821 600614 674347 600616
rect 673821 600611 673887 600614
rect 674281 600611 674347 600614
rect 44541 600538 44607 600541
rect 41492 600536 44607 600538
rect 41492 600480 44546 600536
rect 44602 600480 44607 600536
rect 41492 600478 44607 600480
rect 44541 600475 44607 600478
rect 673821 600402 673887 600405
rect 675109 600402 675175 600405
rect 673821 600400 675175 600402
rect 673821 600344 673826 600400
rect 673882 600344 675114 600400
rect 675170 600344 675175 600400
rect 673821 600342 675175 600344
rect 673821 600339 673887 600342
rect 675109 600339 675175 600342
rect 44633 600130 44699 600133
rect 41492 600128 44699 600130
rect 41492 600072 44638 600128
rect 44694 600072 44699 600128
rect 41492 600070 44699 600072
rect 44633 600067 44699 600070
rect 673729 599858 673795 599861
rect 675477 599858 675543 599861
rect 673729 599856 675543 599858
rect 673729 599800 673734 599856
rect 673790 599800 675482 599856
rect 675538 599800 675543 599856
rect 673729 599798 675543 599800
rect 673729 599795 673795 599798
rect 675477 599795 675543 599798
rect 45093 599722 45159 599725
rect 41492 599720 45159 599722
rect 41492 599664 45098 599720
rect 45154 599664 45159 599720
rect 41492 599662 45159 599664
rect 45093 599659 45159 599662
rect 44909 599314 44975 599317
rect 41492 599312 44975 599314
rect 41492 599256 44914 599312
rect 44970 599256 44975 599312
rect 41492 599254 44975 599256
rect 44909 599251 44975 599254
rect 45461 598906 45527 598909
rect 41492 598904 45527 598906
rect 41492 598848 45466 598904
rect 45522 598848 45527 598904
rect 41492 598846 45527 598848
rect 45461 598843 45527 598846
rect 673545 598634 673611 598637
rect 675477 598634 675543 598637
rect 673545 598632 675543 598634
rect 673545 598576 673550 598632
rect 673606 598576 675482 598632
rect 675538 598576 675543 598632
rect 673545 598574 675543 598576
rect 673545 598571 673611 598574
rect 675477 598571 675543 598574
rect 42742 598498 42748 598500
rect 41492 598438 42748 598498
rect 42742 598436 42748 598438
rect 42812 598436 42818 598500
rect 45277 598090 45343 598093
rect 41492 598088 45343 598090
rect 41492 598032 45282 598088
rect 45338 598032 45343 598088
rect 41492 598030 45343 598032
rect 45277 598027 45343 598030
rect 649950 597954 650010 598336
rect 673177 598090 673243 598093
rect 675109 598090 675175 598093
rect 673177 598088 675175 598090
rect 673177 598032 673182 598088
rect 673238 598032 675114 598088
rect 675170 598032 675175 598088
rect 673177 598030 675175 598032
rect 673177 598027 673243 598030
rect 675109 598027 675175 598030
rect 651465 597954 651531 597957
rect 649950 597952 651531 597954
rect 649950 597896 651470 597952
rect 651526 597896 651531 597952
rect 649950 597894 651531 597896
rect 651465 597891 651531 597894
rect 43069 597682 43135 597685
rect 41492 597680 43135 597682
rect 41492 597624 43074 597680
rect 43130 597624 43135 597680
rect 41492 597622 43135 597624
rect 43069 597619 43135 597622
rect 672533 597410 672599 597413
rect 675385 597410 675451 597413
rect 672533 597408 675451 597410
rect 672533 597352 672538 597408
rect 672594 597352 675390 597408
rect 675446 597352 675451 597408
rect 672533 597350 675451 597352
rect 672533 597347 672599 597350
rect 675385 597347 675451 597350
rect 42006 597274 42012 597276
rect 41492 597214 42012 597274
rect 42006 597212 42012 597214
rect 42076 597212 42082 597276
rect 42793 597004 42859 597005
rect 42742 597002 42748 597004
rect 42702 596942 42748 597002
rect 42812 597000 42859 597004
rect 42854 596944 42859 597000
rect 42742 596940 42748 596942
rect 42812 596940 42859 596944
rect 42793 596939 42859 596940
rect 42425 596866 42491 596869
rect 41492 596864 42491 596866
rect 41492 596808 42430 596864
rect 42486 596808 42491 596864
rect 41492 596806 42491 596808
rect 42425 596803 42491 596806
rect 649950 596730 650010 597154
rect 651465 596730 651531 596733
rect 649950 596728 651531 596730
rect 649950 596672 651470 596728
rect 651526 596672 651531 596728
rect 649950 596670 651531 596672
rect 651465 596667 651531 596670
rect 40910 596223 40970 596428
rect 40910 596218 41019 596223
rect 40910 596162 40958 596218
rect 41014 596162 41019 596218
rect 40910 596160 41019 596162
rect 40953 596157 41019 596160
rect 41278 595815 41338 596020
rect 35157 595812 35223 595815
rect 35157 595810 35266 595812
rect 35157 595754 35162 595810
rect 35218 595754 35266 595810
rect 35157 595749 35266 595754
rect 41278 595810 41387 595815
rect 41278 595754 41326 595810
rect 41382 595754 41387 595810
rect 41278 595752 41387 595754
rect 41321 595749 41387 595752
rect 41689 595778 41755 595781
rect 63401 595778 63467 595781
rect 41689 595776 63467 595778
rect 35206 595612 35266 595749
rect 41689 595720 41694 595776
rect 41750 595720 63406 595776
rect 63462 595720 63467 595776
rect 41689 595718 63467 595720
rect 41689 595715 41755 595718
rect 63401 595715 63467 595718
rect 649950 595370 650010 595972
rect 651465 595370 651531 595373
rect 675385 595372 675451 595373
rect 675334 595370 675340 595372
rect 649950 595368 651531 595370
rect 649950 595312 651470 595368
rect 651526 595312 651531 595368
rect 649950 595310 651531 595312
rect 675294 595310 675340 595370
rect 675404 595368 675451 595372
rect 675446 595312 675451 595368
rect 651465 595307 651531 595310
rect 675334 595308 675340 595310
rect 675404 595308 675451 595312
rect 675385 595307 675451 595308
rect 33041 595234 33107 595237
rect 33028 595232 33107 595234
rect 33028 595176 33046 595232
rect 33102 595176 33107 595232
rect 33028 595174 33107 595176
rect 33041 595171 33107 595174
rect 651649 595098 651715 595101
rect 649950 595096 651715 595098
rect 649950 595040 651654 595096
rect 651710 595040 651715 595096
rect 649950 595038 651715 595040
rect 37917 594826 37983 594829
rect 37917 594824 37996 594826
rect 37917 594768 37922 594824
rect 37978 594768 37996 594824
rect 649950 594790 650010 595038
rect 651649 595035 651715 595038
rect 669037 594826 669103 594829
rect 675477 594826 675543 594829
rect 669037 594824 675543 594826
rect 37917 594766 37996 594768
rect 669037 594768 669042 594824
rect 669098 594768 675482 594824
rect 675538 594768 675543 594824
rect 669037 594766 675543 594768
rect 37917 594763 37983 594766
rect 669037 594763 669103 594766
rect 675477 594763 675543 594766
rect 31017 594418 31083 594421
rect 31004 594416 31083 594418
rect 31004 594360 31022 594416
rect 31078 594360 31083 594416
rect 31004 594358 31083 594360
rect 31017 594355 31083 594358
rect 41781 594282 41847 594285
rect 41781 594280 51090 594282
rect 41781 594224 41786 594280
rect 41842 594224 51090 594280
rect 41781 594222 51090 594224
rect 41781 594219 41847 594222
rect 51030 594146 51090 594222
rect 62481 594146 62547 594149
rect 651465 594146 651531 594149
rect 51030 594144 62547 594146
rect 51030 594088 62486 594144
rect 62542 594088 62547 594144
rect 51030 594086 62547 594088
rect 62481 594083 62547 594086
rect 649950 594144 651531 594146
rect 649950 594088 651470 594144
rect 651526 594088 651531 594144
rect 649950 594086 651531 594088
rect 41822 594010 41828 594012
rect 41492 593950 41828 594010
rect 41822 593948 41828 593950
rect 41892 593948 41898 594012
rect 649950 593608 650010 594086
rect 651465 594083 651531 594086
rect 33777 593602 33843 593605
rect 33764 593600 33843 593602
rect 33764 593544 33782 593600
rect 33838 593544 33843 593600
rect 33764 593542 33843 593544
rect 33777 593539 33843 593542
rect 668393 593466 668459 593469
rect 675385 593466 675451 593469
rect 668393 593464 675451 593466
rect 668393 593408 668398 593464
rect 668454 593408 675390 593464
rect 675446 593408 675451 593464
rect 668393 593406 675451 593408
rect 668393 593403 668459 593406
rect 675385 593403 675451 593406
rect 44357 593194 44423 593197
rect 41492 593192 44423 593194
rect 41492 593136 44362 593192
rect 44418 593136 44423 593192
rect 41492 593134 44423 593136
rect 44357 593131 44423 593134
rect 675150 593132 675156 593196
rect 675220 593194 675226 593196
rect 675477 593194 675543 593197
rect 675220 593192 675543 593194
rect 675220 593136 675482 593192
rect 675538 593136 675543 593192
rect 675220 593134 675543 593136
rect 675220 593132 675226 593134
rect 675477 593131 675543 593134
rect 651465 592922 651531 592925
rect 649950 592920 651531 592922
rect 649950 592864 651470 592920
rect 651526 592864 651531 592920
rect 649950 592862 651531 592864
rect 40726 592550 40786 592756
rect 40718 592486 40724 592550
rect 40788 592486 40794 592550
rect 649950 592426 650010 592862
rect 651465 592859 651531 592862
rect 41822 592378 41828 592380
rect 41492 592318 41828 592378
rect 41822 592316 41828 592318
rect 41892 592316 41898 592380
rect 41689 592106 41755 592109
rect 42190 592106 42196 592108
rect 41689 592104 42196 592106
rect 41689 592048 41694 592104
rect 41750 592048 42196 592104
rect 41689 592046 42196 592048
rect 41689 592043 41755 592046
rect 42190 592044 42196 592046
rect 42260 592044 42266 592108
rect 35617 591970 35683 591973
rect 35604 591968 35683 591970
rect 35604 591912 35622 591968
rect 35678 591912 35683 591968
rect 35604 591910 35683 591912
rect 35617 591907 35683 591910
rect 35801 591562 35867 591565
rect 35788 591560 35867 591562
rect 35788 591504 35806 591560
rect 35862 591504 35867 591560
rect 35788 591502 35867 591504
rect 35801 591499 35867 591502
rect 675017 591562 675083 591565
rect 675334 591562 675340 591564
rect 675017 591560 675340 591562
rect 675017 591504 675022 591560
rect 675078 591504 675340 591560
rect 675017 591502 675340 591504
rect 675017 591499 675083 591502
rect 675334 591500 675340 591502
rect 675404 591500 675410 591564
rect 676070 591364 676076 591428
rect 676140 591426 676146 591428
rect 682377 591426 682443 591429
rect 676140 591424 682443 591426
rect 676140 591368 682382 591424
rect 682438 591368 682443 591424
rect 676140 591366 682443 591368
rect 676140 591364 676146 591366
rect 682377 591363 682443 591366
rect 41462 590746 41522 591124
rect 674230 591092 674236 591156
rect 674300 591154 674306 591156
rect 684217 591154 684283 591157
rect 674300 591152 684283 591154
rect 674300 591096 684222 591152
rect 684278 591096 684283 591152
rect 674300 591094 684283 591096
rect 674300 591092 674306 591094
rect 684217 591091 684283 591094
rect 63033 590746 63099 590749
rect 41462 590744 63099 590746
rect 41462 590716 63038 590744
rect 41492 590688 63038 590716
rect 63094 590688 63099 590744
rect 41492 590686 63099 590688
rect 63033 590683 63099 590686
rect 62297 590066 62363 590069
rect 51030 590064 62363 590066
rect 51030 590008 62302 590064
rect 62358 590008 62363 590064
rect 51030 590006 62363 590008
rect 36537 589658 36603 589661
rect 51030 589658 51090 590006
rect 62297 590003 62363 590006
rect 36537 589656 51090 589658
rect 36537 589600 36542 589656
rect 36598 589600 51090 589656
rect 36537 589598 51090 589600
rect 36537 589595 36603 589598
rect 39665 589386 39731 589389
rect 43437 589386 43503 589389
rect 39665 589384 43503 589386
rect 39665 589328 39670 589384
rect 39726 589328 43442 589384
rect 43498 589328 43503 589384
rect 39665 589326 43503 589328
rect 39665 589323 39731 589326
rect 43437 589323 43503 589326
rect 675201 586258 675267 586261
rect 676070 586258 676076 586260
rect 675201 586256 676076 586258
rect 675201 586200 675206 586256
rect 675262 586200 676076 586256
rect 675201 586198 676076 586200
rect 675201 586195 675267 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 39389 586122 39455 586125
rect 42701 586122 42767 586125
rect 39389 586120 42767 586122
rect 39389 586064 39394 586120
rect 39450 586064 42706 586120
rect 42762 586064 42767 586120
rect 39389 586062 42767 586064
rect 39389 586059 39455 586062
rect 42701 586059 42767 586062
rect 40401 585714 40467 585717
rect 62849 585714 62915 585717
rect 40401 585712 62915 585714
rect 40401 585656 40406 585712
rect 40462 585656 62854 585712
rect 62910 585656 62915 585712
rect 40401 585654 62915 585656
rect 40401 585651 40467 585654
rect 62849 585651 62915 585654
rect 37917 585170 37983 585173
rect 41822 585170 41828 585172
rect 37917 585168 41828 585170
rect 37917 585112 37922 585168
rect 37978 585112 41828 585168
rect 37917 585110 41828 585112
rect 37917 585107 37983 585110
rect 41822 585108 41828 585110
rect 41892 585108 41898 585172
rect 39205 584898 39271 584901
rect 41086 584898 41092 584900
rect 39205 584896 41092 584898
rect 39205 584840 39210 584896
rect 39266 584840 41092 584896
rect 39205 584838 41092 584840
rect 39205 584835 39271 584838
rect 41086 584836 41092 584838
rect 41156 584836 41162 584900
rect 39757 584626 39823 584629
rect 40350 584626 40356 584628
rect 39757 584624 40356 584626
rect 39757 584568 39762 584624
rect 39818 584568 40356 584624
rect 39757 584566 40356 584568
rect 39757 584563 39823 584566
rect 40350 584564 40356 584566
rect 40420 584564 40426 584628
rect 673177 581090 673243 581093
rect 673177 581088 676292 581090
rect 673177 581032 673182 581088
rect 673238 581032 676292 581088
rect 673177 581030 676292 581032
rect 673177 581027 673243 581030
rect 676262 580549 676322 580652
rect 676213 580544 676322 580549
rect 676213 580488 676218 580544
rect 676274 580488 676322 580544
rect 676213 580486 676322 580488
rect 676213 580483 676279 580486
rect 40350 580212 40356 580276
rect 40420 580274 40426 580276
rect 41781 580274 41847 580277
rect 40420 580272 41847 580274
rect 40420 580216 41786 580272
rect 41842 580216 41847 580272
rect 40420 580214 41847 580216
rect 40420 580212 40426 580214
rect 41781 580211 41847 580214
rect 42241 580274 42307 580277
rect 45093 580274 45159 580277
rect 42241 580272 45159 580274
rect 42241 580216 42246 580272
rect 42302 580216 45098 580272
rect 45154 580216 45159 580272
rect 42241 580214 45159 580216
rect 42241 580211 42307 580214
rect 45093 580211 45159 580214
rect 673177 580274 673243 580277
rect 673177 580272 676292 580274
rect 673177 580216 673182 580272
rect 673238 580216 676292 580272
rect 673177 580214 676292 580216
rect 673177 580211 673243 580214
rect 41086 579940 41092 580004
rect 41156 580002 41162 580004
rect 42425 580002 42491 580005
rect 41156 580000 42491 580002
rect 41156 579944 42430 580000
rect 42486 579944 42491 580000
rect 41156 579942 42491 579944
rect 41156 579940 41162 579942
rect 42425 579939 42491 579942
rect 673177 580002 673243 580005
rect 673177 580000 676322 580002
rect 673177 579944 673182 580000
rect 673238 579944 676322 580000
rect 673177 579942 676322 579944
rect 673177 579939 673243 579942
rect 676262 579836 676322 579942
rect 673177 579730 673243 579733
rect 674373 579730 674439 579733
rect 673177 579728 674439 579730
rect 673177 579672 673182 579728
rect 673238 579672 674378 579728
rect 674434 579672 674439 579728
rect 673177 579670 674439 579672
rect 673177 579667 673243 579670
rect 674373 579667 674439 579670
rect 42190 579396 42196 579460
rect 42260 579458 42266 579460
rect 42425 579458 42491 579461
rect 42260 579456 42491 579458
rect 42260 579400 42430 579456
rect 42486 579400 42491 579456
rect 42260 579398 42491 579400
rect 42260 579396 42266 579398
rect 42425 579395 42491 579398
rect 676262 579325 676322 579428
rect 676213 579320 676322 579325
rect 676213 579264 676218 579320
rect 676274 579264 676322 579320
rect 676213 579262 676322 579264
rect 676213 579259 676279 579262
rect 42333 579186 42399 579189
rect 46933 579186 46999 579189
rect 42333 579184 46999 579186
rect 42333 579128 42338 579184
rect 42394 579128 46938 579184
rect 46994 579128 46999 579184
rect 42333 579126 46999 579128
rect 42333 579123 42399 579126
rect 46933 579123 46999 579126
rect 673177 578914 673243 578917
rect 676262 578914 676322 579020
rect 673177 578912 676322 578914
rect 673177 578856 673182 578912
rect 673238 578856 676322 578912
rect 673177 578854 676322 578856
rect 673177 578851 673243 578854
rect 673678 578580 673684 578644
rect 673748 578642 673754 578644
rect 673748 578582 676292 578642
rect 673748 578580 673754 578582
rect 42006 578308 42012 578372
rect 42076 578370 42082 578372
rect 42333 578370 42399 578373
rect 42076 578368 42399 578370
rect 42076 578312 42338 578368
rect 42394 578312 42399 578368
rect 42076 578310 42399 578312
rect 42076 578308 42082 578310
rect 42333 578307 42399 578310
rect 670969 578234 671035 578237
rect 674465 578234 674531 578237
rect 670969 578232 674531 578234
rect 670969 578176 670974 578232
rect 671030 578176 674470 578232
rect 674526 578176 674531 578232
rect 670969 578174 674531 578176
rect 670969 578171 671035 578174
rect 674465 578171 674531 578174
rect 676262 578101 676322 578204
rect 42057 578098 42123 578101
rect 44357 578098 44423 578101
rect 42057 578096 44423 578098
rect 42057 578040 42062 578096
rect 42118 578040 44362 578096
rect 44418 578040 44423 578096
rect 42057 578038 44423 578040
rect 42057 578035 42123 578038
rect 44357 578035 44423 578038
rect 676213 578096 676322 578101
rect 676213 578040 676218 578096
rect 676274 578040 676322 578096
rect 676213 578038 676322 578040
rect 676213 578035 676279 578038
rect 673177 577962 673243 577965
rect 673494 577962 673500 577964
rect 673177 577960 673500 577962
rect 673177 577904 673182 577960
rect 673238 577904 673500 577960
rect 673177 577902 673500 577904
rect 673177 577899 673243 577902
rect 673494 577900 673500 577902
rect 673564 577900 673570 577964
rect 40902 577764 40908 577828
rect 40972 577826 40978 577828
rect 41781 577826 41847 577829
rect 40972 577824 41847 577826
rect 40972 577768 41786 577824
rect 41842 577768 41847 577824
rect 40972 577766 41847 577768
rect 40972 577764 40978 577766
rect 41781 577763 41847 577766
rect 673686 577766 676292 577826
rect 673177 577690 673243 577693
rect 673686 577690 673746 577766
rect 673177 577688 673746 577690
rect 673177 577632 673182 577688
rect 673238 577632 673746 577688
rect 673177 577630 673746 577632
rect 673177 577627 673243 577630
rect 674373 577554 674439 577557
rect 673870 577552 674439 577554
rect 673870 577496 674378 577552
rect 674434 577496 674439 577552
rect 673870 577494 674439 577496
rect 673177 577418 673243 577421
rect 673870 577418 673930 577494
rect 674373 577491 674439 577494
rect 673177 577416 673930 577418
rect 673177 577360 673182 577416
rect 673238 577360 673930 577416
rect 673177 577358 673930 577360
rect 673177 577355 673243 577358
rect 676262 577282 676322 577388
rect 674054 577222 676322 577282
rect 673177 577146 673243 577149
rect 674054 577146 674114 577222
rect 673177 577144 674114 577146
rect 673177 577088 673182 577144
rect 673238 577088 674114 577144
rect 673177 577086 674114 577088
rect 673177 577083 673243 577086
rect 673177 576874 673243 576877
rect 676262 576874 676322 576980
rect 673177 576872 676322 576874
rect 673177 576816 673182 576872
rect 673238 576816 676322 576872
rect 673177 576814 676322 576816
rect 673177 576811 673243 576814
rect 676806 576812 676812 576876
rect 676876 576812 676882 576876
rect 676814 576572 676874 576812
rect 679617 576466 679683 576469
rect 679574 576464 679683 576466
rect 679574 576408 679622 576464
rect 679678 576408 679683 576464
rect 679574 576403 679683 576408
rect 679574 576164 679634 576403
rect 684217 576058 684283 576061
rect 684174 576056 684283 576058
rect 684174 576000 684222 576056
rect 684278 576000 684283 576056
rect 684174 575995 684283 576000
rect 684174 575756 684234 575995
rect 682377 575650 682443 575653
rect 682334 575648 682443 575650
rect 682334 575592 682382 575648
rect 682438 575592 682443 575648
rect 682334 575587 682443 575592
rect 682334 575348 682394 575587
rect 676262 574837 676322 574940
rect 62113 574834 62179 574837
rect 673913 574834 673979 574837
rect 674557 574834 674623 574837
rect 62113 574832 64706 574834
rect 62113 574776 62118 574832
rect 62174 574776 64706 574832
rect 62113 574774 64706 574776
rect 62113 574771 62179 574774
rect 40718 574636 40724 574700
rect 40788 574698 40794 574700
rect 41781 574698 41847 574701
rect 40788 574696 41847 574698
rect 40788 574640 41786 574696
rect 41842 574640 41847 574696
rect 40788 574638 41847 574640
rect 40788 574636 40794 574638
rect 41781 574635 41847 574638
rect 64646 574194 64706 574774
rect 673913 574832 674623 574834
rect 673913 574776 673918 574832
rect 673974 574776 674562 574832
rect 674618 574776 674623 574832
rect 673913 574774 674623 574776
rect 673913 574771 673979 574774
rect 674557 574771 674623 574774
rect 676213 574832 676322 574837
rect 676213 574776 676218 574832
rect 676274 574776 676322 574832
rect 676213 574774 676322 574776
rect 676213 574771 676279 574774
rect 673913 574562 673979 574565
rect 673913 574560 676292 574562
rect 673913 574504 673918 574560
rect 673974 574504 676292 574560
rect 673913 574502 676292 574504
rect 673913 574499 673979 574502
rect 673913 574154 673979 574157
rect 673913 574152 676292 574154
rect 673913 574096 673918 574152
rect 673974 574096 676292 574152
rect 673913 574094 676292 574096
rect 673913 574091 673979 574094
rect 41454 573956 41460 574020
rect 41524 574018 41530 574020
rect 42609 574018 42675 574021
rect 41524 574016 42675 574018
rect 41524 573960 42614 574016
rect 42670 573960 42675 574016
rect 41524 573958 42675 573960
rect 41524 573956 41530 573958
rect 42609 573955 42675 573958
rect 673913 573882 673979 573885
rect 674373 573882 674439 573885
rect 673913 573880 674439 573882
rect 673913 573824 673918 573880
rect 673974 573824 674378 573880
rect 674434 573824 674439 573880
rect 673913 573822 674439 573824
rect 673913 573819 673979 573822
rect 674373 573819 674439 573822
rect 62113 573610 62179 573613
rect 672717 573610 672783 573613
rect 676262 573610 676322 573716
rect 62113 573608 64706 573610
rect 62113 573552 62118 573608
rect 62174 573552 64706 573608
rect 62113 573550 64706 573552
rect 62113 573547 62179 573550
rect 40534 573412 40540 573476
rect 40604 573474 40610 573476
rect 41781 573474 41847 573477
rect 42149 573476 42215 573477
rect 42149 573474 42196 573476
rect 40604 573472 41847 573474
rect 40604 573416 41786 573472
rect 41842 573416 41847 573472
rect 40604 573414 41847 573416
rect 42104 573472 42196 573474
rect 42104 573416 42154 573472
rect 42104 573414 42196 573416
rect 40604 573412 40610 573414
rect 41781 573411 41847 573414
rect 42149 573412 42196 573414
rect 42260 573412 42266 573476
rect 42149 573411 42215 573412
rect 64646 573012 64706 573550
rect 672717 573608 676322 573610
rect 672717 573552 672722 573608
rect 672778 573552 676322 573608
rect 672717 573550 676322 573552
rect 672717 573547 672783 573550
rect 676262 573202 676322 573308
rect 673686 573142 676322 573202
rect 683389 573202 683455 573205
rect 683389 573200 683498 573202
rect 683389 573144 683394 573200
rect 683450 573144 683498 573200
rect 672993 572794 673059 572797
rect 673686 572794 673746 573142
rect 683389 573139 683498 573144
rect 683438 572900 683498 573139
rect 672993 572792 673746 572794
rect 672993 572736 672998 572792
rect 673054 572736 673746 572792
rect 672993 572734 673746 572736
rect 672993 572731 673059 572734
rect 42057 572660 42123 572661
rect 42006 572596 42012 572660
rect 42076 572658 42123 572660
rect 42076 572656 42168 572658
rect 42118 572600 42168 572656
rect 42076 572598 42168 572600
rect 42076 572596 42123 572598
rect 42057 572595 42123 572596
rect 676262 572389 676322 572492
rect 676213 572384 676322 572389
rect 676213 572328 676218 572384
rect 676274 572328 676322 572384
rect 676213 572326 676322 572328
rect 676213 572323 676279 572326
rect 673913 572114 673979 572117
rect 673913 572112 676292 572114
rect 673913 572056 673918 572112
rect 673974 572056 676292 572112
rect 673913 572054 676292 572056
rect 673913 572051 673979 572054
rect 684033 571978 684099 571981
rect 683990 571976 684099 571978
rect 683990 571920 684038 571976
rect 684094 571920 684099 571976
rect 683990 571915 684099 571920
rect 41638 571508 41644 571572
rect 41708 571570 41714 571572
rect 42057 571570 42123 571573
rect 41708 571568 42123 571570
rect 41708 571512 42062 571568
rect 42118 571512 42123 571568
rect 41708 571510 42123 571512
rect 41708 571508 41714 571510
rect 42057 571507 42123 571510
rect 42425 571434 42491 571437
rect 64646 571434 64706 571830
rect 683990 571676 684050 571915
rect 42425 571432 64706 571434
rect 42425 571376 42430 571432
rect 42486 571376 64706 571432
rect 42425 571374 64706 571376
rect 673913 571434 673979 571437
rect 674373 571434 674439 571437
rect 673913 571432 674439 571434
rect 673913 571376 673918 571432
rect 673974 571376 674378 571432
rect 674434 571376 674439 571432
rect 673913 571374 674439 571376
rect 42425 571371 42491 571374
rect 673913 571371 673979 571374
rect 674373 571371 674439 571374
rect 676029 571298 676095 571301
rect 676029 571296 676292 571298
rect 676029 571240 676034 571296
rect 676090 571240 676292 571296
rect 676029 571238 676292 571240
rect 676029 571235 676095 571238
rect 63401 571162 63467 571165
rect 673913 571162 673979 571165
rect 674833 571162 674899 571165
rect 63401 571160 64706 571162
rect 63401 571104 63406 571160
rect 63462 571104 64706 571160
rect 63401 571102 64706 571104
rect 63401 571099 63467 571102
rect 64646 570648 64706 571102
rect 673913 571160 674899 571162
rect 673913 571104 673918 571160
rect 673974 571104 674838 571160
rect 674894 571104 674899 571160
rect 673913 571102 674899 571104
rect 673913 571099 673979 571102
rect 674833 571099 674899 571102
rect 673913 570890 673979 570893
rect 673913 570888 676292 570890
rect 673913 570832 673918 570888
rect 673974 570832 676292 570888
rect 673913 570830 676292 570832
rect 673913 570827 673979 570830
rect 682886 570346 682946 570452
rect 683113 570346 683179 570349
rect 682886 570344 683179 570346
rect 682886 570288 683118 570344
rect 683174 570288 683179 570344
rect 682886 570286 683179 570288
rect 41781 570212 41847 570213
rect 41781 570208 41828 570212
rect 41892 570210 41898 570212
rect 41781 570152 41786 570208
rect 41781 570148 41828 570152
rect 41892 570150 41938 570210
rect 41892 570148 41898 570150
rect 41781 570147 41847 570148
rect 682886 570044 682946 570286
rect 683113 570283 683179 570286
rect 62297 569938 62363 569941
rect 62297 569936 64706 569938
rect 62297 569880 62302 569936
rect 62358 569880 64706 569936
rect 62297 569878 64706 569880
rect 62297 569875 62363 569878
rect 64646 569466 64706 569878
rect 673913 569666 673979 569669
rect 673913 569664 676292 569666
rect 673913 569608 673918 569664
rect 673974 569608 676292 569664
rect 673913 569606 676292 569608
rect 673913 569603 673979 569606
rect 62481 568578 62547 568581
rect 62481 568576 64706 568578
rect 62481 568520 62486 568576
rect 62542 568520 64706 568576
rect 62481 568518 64706 568520
rect 62481 568515 62547 568518
rect 64646 568284 64706 568518
rect 673913 565858 673979 565861
rect 675385 565858 675451 565861
rect 673913 565856 675451 565858
rect 673913 565800 673918 565856
rect 673974 565800 675390 565856
rect 675446 565800 675451 565856
rect 673913 565798 675451 565800
rect 673913 565795 673979 565798
rect 675385 565795 675451 565798
rect 673913 564498 673979 564501
rect 675109 564498 675175 564501
rect 673913 564496 675175 564498
rect 673913 564440 673918 564496
rect 673974 564440 675114 564496
rect 675170 564440 675175 564496
rect 673913 564438 675175 564440
rect 673913 564435 673979 564438
rect 675109 564435 675175 564438
rect 668761 562322 668827 562325
rect 675109 562322 675175 562325
rect 668761 562320 675175 562322
rect 668761 562264 668766 562320
rect 668822 562264 675114 562320
rect 675170 562264 675175 562320
rect 668761 562262 675175 562264
rect 668761 562259 668827 562262
rect 675109 562259 675175 562262
rect 675385 561916 675451 561917
rect 675334 561914 675340 561916
rect 675294 561854 675340 561914
rect 675404 561912 675451 561916
rect 675446 561856 675451 561912
rect 675334 561852 675340 561854
rect 675404 561852 675451 561856
rect 675385 561851 675451 561852
rect 673085 559058 673151 559061
rect 675109 559058 675175 559061
rect 673085 559056 675175 559058
rect 673085 559000 673090 559056
rect 673146 559000 675114 559056
rect 675170 559000 675175 559056
rect 673085 558998 675175 559000
rect 673085 558995 673151 558998
rect 675109 558995 675175 558998
rect 41086 558724 41092 558788
rect 41156 558786 41162 558788
rect 44633 558786 44699 558789
rect 41156 558784 44699 558786
rect 41156 558728 44638 558784
rect 44694 558728 44699 558784
rect 41156 558726 44699 558728
rect 41156 558724 41162 558726
rect 44633 558723 44699 558726
rect 47577 558514 47643 558517
rect 41492 558512 47643 558514
rect 41492 558456 47582 558512
rect 47638 558456 47643 558512
rect 41492 558454 47643 558456
rect 47577 558451 47643 558454
rect 673913 558378 673979 558381
rect 675385 558378 675451 558381
rect 673913 558376 675451 558378
rect 673913 558320 673918 558376
rect 673974 558320 675390 558376
rect 675446 558320 675451 558376
rect 673913 558318 675451 558320
rect 673913 558315 673979 558318
rect 675385 558315 675451 558318
rect 40953 558106 41019 558109
rect 40940 558104 41019 558106
rect 40940 558048 40958 558104
rect 41014 558048 41019 558104
rect 40940 558046 41019 558048
rect 40953 558043 41019 558046
rect 41086 557488 41092 557552
rect 41156 557488 41162 557552
rect 41278 557550 41338 557668
rect 671797 557562 671863 557565
rect 675109 557562 675175 557565
rect 671797 557560 675175 557562
rect 41278 557490 41890 557550
rect 671797 557504 671802 557560
rect 671858 557504 675114 557560
rect 675170 557504 675175 557560
rect 671797 557502 675175 557504
rect 671797 557499 671863 557502
rect 675109 557499 675175 557502
rect 41094 557260 41154 557488
rect 41830 557426 41890 557490
rect 41830 557366 51090 557426
rect 45093 556882 45159 556885
rect 41492 556880 45159 556882
rect 41492 556824 45098 556880
rect 45154 556824 45159 556880
rect 41492 556822 45159 556824
rect 45093 556819 45159 556822
rect 51030 556746 51090 557366
rect 63217 556746 63283 556749
rect 51030 556744 63283 556746
rect 51030 556688 63222 556744
rect 63278 556688 63283 556744
rect 51030 556686 63283 556688
rect 63217 556683 63283 556686
rect 44909 556474 44975 556477
rect 41492 556472 44975 556474
rect 41492 556416 44914 556472
rect 44970 556416 44975 556472
rect 41492 556414 44975 556416
rect 44909 556411 44975 556414
rect 44633 556066 44699 556069
rect 41492 556064 44699 556066
rect 41492 556008 44638 556064
rect 44694 556008 44699 556064
rect 41492 556006 44699 556008
rect 44633 556003 44699 556006
rect 42793 555658 42859 555661
rect 41492 555656 42859 555658
rect 41492 555600 42798 555656
rect 42854 555600 42859 555656
rect 41492 555598 42859 555600
rect 42793 555595 42859 555598
rect 44357 555250 44423 555253
rect 41492 555248 44423 555250
rect 41492 555192 44362 555248
rect 44418 555192 44423 555248
rect 41492 555190 44423 555192
rect 44357 555187 44423 555190
rect 672901 555250 672967 555253
rect 675385 555250 675451 555253
rect 672901 555248 675451 555250
rect 672901 555192 672906 555248
rect 672962 555192 675390 555248
rect 675446 555192 675451 555248
rect 672901 555190 675451 555192
rect 672901 555187 672967 555190
rect 675385 555187 675451 555190
rect 43069 554842 43135 554845
rect 41492 554840 43135 554842
rect 41492 554784 43074 554840
rect 43130 554784 43135 554840
rect 41492 554782 43135 554784
rect 43069 554779 43135 554782
rect 672717 554842 672783 554845
rect 675201 554842 675267 554845
rect 672717 554840 675267 554842
rect 672717 554784 672722 554840
rect 672778 554784 675206 554840
rect 675262 554784 675267 554840
rect 672717 554782 675267 554784
rect 672717 554779 672783 554782
rect 675201 554779 675267 554782
rect 675753 554706 675819 554709
rect 676254 554706 676260 554708
rect 675753 554704 676260 554706
rect 675753 554648 675758 554704
rect 675814 554648 676260 554704
rect 675753 554646 676260 554648
rect 675753 554643 675819 554646
rect 676254 554644 676260 554646
rect 676324 554644 676330 554708
rect 43161 554434 43227 554437
rect 41492 554432 43227 554434
rect 41492 554376 43166 554432
rect 43222 554376 43227 554432
rect 41492 554374 43227 554376
rect 43161 554371 43227 554374
rect 674097 554164 674163 554165
rect 674046 554100 674052 554164
rect 674116 554162 674163 554164
rect 674116 554160 674208 554162
rect 674158 554104 674208 554160
rect 674116 554102 674208 554104
rect 674116 554100 674163 554102
rect 674097 554099 674163 554100
rect 41822 554026 41828 554028
rect 41492 553966 41828 554026
rect 41822 553964 41828 553966
rect 41892 553964 41898 554028
rect 41278 553413 41338 553588
rect 649950 553482 650010 553914
rect 675753 553890 675819 553893
rect 676806 553890 676812 553892
rect 675753 553888 676812 553890
rect 675753 553832 675758 553888
rect 675814 553832 676812 553888
rect 675753 553830 676812 553832
rect 675753 553827 675819 553830
rect 676806 553828 676812 553830
rect 676876 553828 676882 553892
rect 651465 553482 651531 553485
rect 649950 553480 651531 553482
rect 649950 553424 651470 553480
rect 651526 553424 651531 553480
rect 649950 553422 651531 553424
rect 651465 553419 651531 553422
rect 37917 553410 37983 553413
rect 37917 553408 38026 553410
rect 37917 553352 37922 553408
rect 37978 553352 38026 553408
rect 37917 553347 38026 553352
rect 41278 553408 41387 553413
rect 41278 553352 41326 553408
rect 41382 553352 41387 553408
rect 41278 553350 41387 553352
rect 41321 553347 41387 553350
rect 37966 553180 38026 553347
rect 674046 552876 674052 552940
rect 674116 552938 674122 552940
rect 674281 552938 674347 552941
rect 674116 552936 674347 552938
rect 674116 552880 674286 552936
rect 674342 552880 674347 552936
rect 674116 552878 674347 552880
rect 674116 552876 674122 552878
rect 674281 552875 674347 552878
rect 41822 552802 41828 552804
rect 41492 552742 41828 552802
rect 41822 552740 41828 552742
rect 41892 552740 41898 552804
rect 41321 552394 41387 552397
rect 41308 552392 41387 552394
rect 41308 552336 41326 552392
rect 41382 552336 41387 552392
rect 41308 552334 41387 552336
rect 41321 552331 41387 552334
rect 649950 552122 650010 552732
rect 669589 552258 669655 552261
rect 675293 552258 675359 552261
rect 669589 552256 675359 552258
rect 669589 552200 669594 552256
rect 669650 552200 675298 552256
rect 675354 552200 675359 552256
rect 669589 552198 675359 552200
rect 669589 552195 669655 552198
rect 675293 552195 675359 552198
rect 651649 552122 651715 552125
rect 649950 552120 651715 552122
rect 649950 552064 651654 552120
rect 651710 552064 651715 552120
rect 649950 552062 651715 552064
rect 651649 552059 651715 552062
rect 29637 551986 29703 551989
rect 29637 551984 29716 551986
rect 29637 551928 29642 551984
rect 29698 551928 29716 551984
rect 29637 551926 29716 551928
rect 29637 551923 29703 551926
rect 41689 551850 41755 551853
rect 43989 551850 44055 551853
rect 41689 551848 44055 551850
rect 41689 551792 41694 551848
rect 41750 551792 43994 551848
rect 44050 551792 44055 551848
rect 41689 551790 44055 551792
rect 41689 551787 41755 551790
rect 43989 551787 44055 551790
rect 45277 551578 45343 551581
rect 41492 551576 45343 551578
rect 41492 551520 45282 551576
rect 45338 551520 45343 551576
rect 41492 551518 45343 551520
rect 45277 551515 45343 551518
rect 42977 551170 43043 551173
rect 41492 551168 43043 551170
rect 41492 551112 42982 551168
rect 43038 551112 43043 551168
rect 41492 551110 43043 551112
rect 649950 551170 650010 551550
rect 651465 551170 651531 551173
rect 649950 551168 651531 551170
rect 649950 551112 651470 551168
rect 651526 551112 651531 551168
rect 649950 551110 651531 551112
rect 42977 551107 43043 551110
rect 651465 551107 651531 551110
rect 43805 550762 43871 550765
rect 41492 550760 43871 550762
rect 41492 550704 43810 550760
rect 43866 550704 43871 550760
rect 41492 550702 43871 550704
rect 43805 550699 43871 550702
rect 44817 550490 44883 550493
rect 41830 550488 44883 550490
rect 41830 550432 44822 550488
rect 44878 550432 44883 550488
rect 41830 550430 44883 550432
rect 41830 550354 41890 550430
rect 44817 550427 44883 550430
rect 673729 550490 673795 550493
rect 674046 550490 674052 550492
rect 673729 550488 674052 550490
rect 673729 550432 673734 550488
rect 673790 550432 674052 550488
rect 673729 550430 674052 550432
rect 673729 550427 673795 550430
rect 674046 550428 674052 550430
rect 674116 550428 674122 550492
rect 41492 550294 41890 550354
rect 649950 550354 650010 550368
rect 651373 550354 651439 550357
rect 649950 550352 651439 550354
rect 649950 550296 651378 550352
rect 651434 550296 651439 550352
rect 649950 550294 651439 550296
rect 651373 550291 651439 550294
rect 42149 550218 42215 550221
rect 62481 550218 62547 550221
rect 42149 550216 62547 550218
rect 42149 550160 42154 550216
rect 42210 550160 62486 550216
rect 62542 550160 62547 550216
rect 42149 550158 62547 550160
rect 42149 550155 42215 550158
rect 62481 550155 62547 550158
rect 40769 549946 40835 549949
rect 40756 549944 40835 549946
rect 40756 549888 40774 549944
rect 40830 549888 40835 549944
rect 40756 549886 40835 549888
rect 40769 549883 40835 549886
rect 670417 549674 670483 549677
rect 675477 549674 675543 549677
rect 670417 549672 675543 549674
rect 670417 549616 670422 549672
rect 670478 549616 675482 549672
rect 675538 549616 675543 549672
rect 670417 549614 675543 549616
rect 670417 549611 670483 549614
rect 675477 549611 675543 549614
rect 42190 549538 42196 549540
rect 41492 549478 42196 549538
rect 42190 549476 42196 549478
rect 42260 549476 42266 549540
rect 651465 549266 651531 549269
rect 649950 549264 651531 549266
rect 649950 549208 651470 549264
rect 651526 549208 651531 549264
rect 649950 549206 651531 549208
rect 649950 549186 650010 549206
rect 651465 549203 651531 549206
rect 42793 549130 42859 549133
rect 41492 549128 42859 549130
rect 41492 549072 42798 549128
rect 42854 549072 42859 549128
rect 41492 549070 42859 549072
rect 42793 549067 42859 549070
rect 44173 548722 44239 548725
rect 41492 548720 44239 548722
rect 41492 548664 44178 548720
rect 44234 548664 44239 548720
rect 41492 548662 44239 548664
rect 44173 548659 44239 548662
rect 651465 548450 651531 548453
rect 649950 548448 651531 548450
rect 649950 548392 651470 548448
rect 651526 548392 651531 548448
rect 649950 548390 651531 548392
rect 41321 548314 41387 548317
rect 41308 548312 41387 548314
rect 41308 548256 41326 548312
rect 41382 548256 41387 548312
rect 41308 548254 41387 548256
rect 41321 548251 41387 548254
rect 649950 548004 650010 548390
rect 651465 548387 651531 548390
rect 674833 548450 674899 548453
rect 675334 548450 675340 548452
rect 674833 548448 675340 548450
rect 674833 548392 674838 548448
rect 674894 548392 675340 548448
rect 674833 548390 675340 548392
rect 674833 548387 674899 548390
rect 675334 548388 675340 548390
rect 675404 548388 675410 548452
rect 675753 548314 675819 548317
rect 676990 548314 676996 548316
rect 675753 548312 676996 548314
rect 675753 548256 675758 548312
rect 675814 548256 676996 548312
rect 675753 548254 676996 548256
rect 675753 548251 675819 548254
rect 676990 548252 676996 548254
rect 677060 548252 677066 548316
rect 41462 547498 41522 547876
rect 674046 547844 674052 547908
rect 674116 547906 674122 547908
rect 675569 547906 675635 547909
rect 674116 547904 675635 547906
rect 674116 547848 675574 547904
rect 675630 547848 675635 547904
rect 674116 547846 675635 547848
rect 674116 547844 674122 547846
rect 675569 547843 675635 547846
rect 41689 547770 41755 547773
rect 43621 547770 43687 547773
rect 41689 547768 43687 547770
rect 41689 547712 41694 547768
rect 41750 547712 43626 547768
rect 43682 547712 43687 547768
rect 41689 547710 43687 547712
rect 41689 547707 41755 547710
rect 43621 547707 43687 547710
rect 676254 547572 676260 547636
rect 676324 547634 676330 547636
rect 677409 547634 677475 547637
rect 676324 547632 677475 547634
rect 676324 547576 677414 547632
rect 677470 547576 677475 547632
rect 676324 547574 677475 547576
rect 676324 547572 676330 547574
rect 677409 547571 677475 547574
rect 46381 547498 46447 547501
rect 41462 547496 46447 547498
rect 41462 547468 46386 547496
rect 41492 547440 46386 547468
rect 46442 547440 46447 547496
rect 41492 547438 46447 547440
rect 46381 547435 46447 547438
rect 676070 546756 676076 546820
rect 676140 546818 676146 546820
rect 682377 546818 682443 546821
rect 676140 546816 682443 546818
rect 676140 546760 682382 546816
rect 682438 546760 682443 546816
rect 676140 546758 682443 546760
rect 676140 546756 676146 546758
rect 682377 546755 682443 546758
rect 41137 545866 41203 545869
rect 42333 545866 42399 545869
rect 41137 545864 42399 545866
rect 41137 545808 41142 545864
rect 41198 545808 42338 545864
rect 42394 545808 42399 545864
rect 41137 545806 42399 545808
rect 41137 545803 41203 545806
rect 42333 545803 42399 545806
rect 40769 545596 40835 545597
rect 40718 545594 40724 545596
rect 40678 545534 40724 545594
rect 40788 545592 40835 545596
rect 40830 545536 40835 545592
rect 40718 545532 40724 545534
rect 40788 545532 40835 545536
rect 40769 545531 40835 545532
rect 40534 545260 40540 545324
rect 40604 545322 40610 545324
rect 42190 545322 42196 545324
rect 40604 545262 42196 545322
rect 40604 545260 40610 545262
rect 42190 545260 42196 545262
rect 42260 545260 42266 545324
rect 37917 542330 37983 542333
rect 41822 542330 41828 542332
rect 37917 542328 41828 542330
rect 37917 542272 37922 542328
rect 37978 542272 41828 542328
rect 37917 542270 41828 542272
rect 37917 542267 37983 542270
rect 41822 542268 41828 542270
rect 41892 542268 41898 542332
rect 42609 539610 42675 539613
rect 44817 539610 44883 539613
rect 42609 539608 44883 539610
rect 42609 539552 42614 539608
rect 42670 539552 44822 539608
rect 44878 539552 44883 539608
rect 42609 539550 44883 539552
rect 42609 539547 42675 539550
rect 44817 539547 44883 539550
rect 42425 538250 42491 538253
rect 51717 538250 51783 538253
rect 42425 538248 51783 538250
rect 42425 538192 42430 538248
rect 42486 538192 51722 538248
rect 51778 538192 51783 538248
rect 42425 538190 51783 538192
rect 42425 538187 42491 538190
rect 51717 538187 51783 538190
rect 42057 537434 42123 537437
rect 44817 537434 44883 537437
rect 42057 537432 44883 537434
rect 42057 537376 42062 537432
rect 42118 537376 44822 537432
rect 44878 537376 44883 537432
rect 42057 537374 44883 537376
rect 42057 537371 42123 537374
rect 44817 537371 44883 537374
rect 674097 537162 674163 537165
rect 675477 537162 675543 537165
rect 674097 537160 675543 537162
rect 674097 537104 674102 537160
rect 674158 537104 675482 537160
rect 675538 537104 675543 537160
rect 674097 537102 675543 537104
rect 674097 537099 674163 537102
rect 675477 537099 675543 537102
rect 42057 537026 42123 537029
rect 42609 537026 42675 537029
rect 42057 537024 42675 537026
rect 42057 536968 42062 537024
rect 42118 536968 42614 537024
rect 42670 536968 42675 537024
rect 42057 536966 42675 536968
rect 42057 536963 42123 536966
rect 42609 536963 42675 536966
rect 44173 536890 44239 536893
rect 42750 536888 44239 536890
rect 42750 536832 44178 536888
rect 44234 536832 44239 536888
rect 42750 536830 44239 536832
rect 42750 536757 42810 536830
rect 44173 536827 44239 536830
rect 42701 536752 42810 536757
rect 42701 536696 42706 536752
rect 42762 536696 42810 536752
rect 42701 536694 42810 536696
rect 42701 536691 42767 536694
rect 676262 535941 676322 536112
rect 676213 535936 676322 535941
rect 676213 535880 676218 535936
rect 676274 535880 676322 535936
rect 676213 535878 676322 535880
rect 676213 535875 676279 535878
rect 676029 535734 676095 535737
rect 676029 535732 676292 535734
rect 676029 535676 676034 535732
rect 676090 535676 676292 535732
rect 676029 535674 676292 535676
rect 676029 535671 676095 535674
rect 42057 535666 42123 535669
rect 42701 535666 42767 535669
rect 42057 535664 42767 535666
rect 42057 535608 42062 535664
rect 42118 535608 42706 535664
rect 42762 535608 42767 535664
rect 42057 535606 42767 535608
rect 42057 535603 42123 535606
rect 42701 535603 42767 535606
rect 40718 535196 40724 535260
rect 40788 535258 40794 535260
rect 41781 535258 41847 535261
rect 40788 535256 41847 535258
rect 40788 535200 41786 535256
rect 41842 535200 41847 535256
rect 40788 535198 41847 535200
rect 40788 535196 40794 535198
rect 41781 535195 41847 535198
rect 676262 535125 676322 535296
rect 676213 535120 676322 535125
rect 676213 535064 676218 535120
rect 676274 535064 676322 535120
rect 676213 535062 676322 535064
rect 676213 535059 676279 535062
rect 676029 534918 676095 534921
rect 676029 534916 676292 534918
rect 676029 534860 676034 534916
rect 676090 534860 676292 534916
rect 676029 534858 676292 534860
rect 676029 534855 676095 534858
rect 676262 534306 676322 534480
rect 676489 534306 676555 534309
rect 675894 534246 676322 534306
rect 676446 534304 676555 534306
rect 676446 534248 676494 534304
rect 676550 534248 676555 534304
rect 670969 534034 671035 534037
rect 675894 534034 675954 534246
rect 676446 534243 676555 534248
rect 676446 534072 676506 534243
rect 670969 534032 675954 534034
rect 670969 533976 670974 534032
rect 671030 533976 675954 534032
rect 670969 533974 675954 533976
rect 670969 533971 671035 533974
rect 42425 533898 42491 533901
rect 43989 533898 44055 533901
rect 42425 533896 44055 533898
rect 42425 533840 42430 533896
rect 42486 533840 43994 533896
rect 44050 533840 44055 533896
rect 42425 533838 44055 533840
rect 42425 533835 42491 533838
rect 43989 533835 44055 533838
rect 672717 533626 672783 533629
rect 676262 533626 676322 533664
rect 672717 533624 676322 533626
rect 672717 533568 672722 533624
rect 672778 533568 676322 533624
rect 672717 533566 676322 533568
rect 672717 533563 672783 533566
rect 40534 533292 40540 533356
rect 40604 533354 40610 533356
rect 42241 533354 42307 533357
rect 40604 533352 42307 533354
rect 40604 533296 42246 533352
rect 42302 533296 42307 533352
rect 40604 533294 42307 533296
rect 40604 533292 40610 533294
rect 42241 533291 42307 533294
rect 676029 533286 676095 533289
rect 676029 533284 676292 533286
rect 676029 533228 676034 533284
rect 676090 533228 676292 533284
rect 676029 533226 676292 533228
rect 676029 533223 676095 533226
rect 676029 532878 676095 532881
rect 676029 532876 676292 532878
rect 676029 532820 676034 532876
rect 676090 532820 676292 532876
rect 676029 532818 676292 532820
rect 676029 532815 676095 532818
rect 42701 532810 42767 532813
rect 43805 532810 43871 532813
rect 42701 532808 43871 532810
rect 42701 532752 42706 532808
rect 42762 532752 43810 532808
rect 43866 532752 43871 532808
rect 42701 532750 43871 532752
rect 42701 532747 42767 532750
rect 43805 532747 43871 532750
rect 676029 532470 676095 532473
rect 676029 532468 676292 532470
rect 676029 532412 676034 532468
rect 676090 532412 676292 532468
rect 676029 532410 676292 532412
rect 676029 532407 676095 532410
rect 676029 532062 676095 532065
rect 676029 532060 676292 532062
rect 676029 532004 676034 532060
rect 676090 532004 676292 532060
rect 676029 532002 676292 532004
rect 676029 531999 676095 532002
rect 676213 531858 676279 531861
rect 676213 531856 676322 531858
rect 676213 531800 676218 531856
rect 676274 531800 676322 531856
rect 676213 531795 676322 531800
rect 41638 531660 41644 531724
rect 41708 531722 41714 531724
rect 42425 531722 42491 531725
rect 41708 531720 42491 531722
rect 41708 531664 42430 531720
rect 42486 531664 42491 531720
rect 41708 531662 42491 531664
rect 41708 531660 41714 531662
rect 42425 531659 42491 531662
rect 676262 531624 676322 531795
rect 680997 531450 681063 531453
rect 680997 531448 681106 531450
rect 680997 531392 681002 531448
rect 681058 531392 681106 531448
rect 680997 531387 681106 531392
rect 681046 531216 681106 531387
rect 62113 531178 62179 531181
rect 62113 531176 64706 531178
rect 62113 531120 62118 531176
rect 62174 531120 64706 531176
rect 62113 531118 64706 531120
rect 62113 531115 62179 531118
rect 676029 530838 676095 530841
rect 676029 530836 676292 530838
rect 676029 530780 676034 530836
rect 676090 530780 676292 530836
rect 676029 530778 676292 530780
rect 676029 530775 676095 530778
rect 41454 530708 41460 530772
rect 41524 530770 41530 530772
rect 42609 530770 42675 530773
rect 41524 530768 42675 530770
rect 41524 530712 42614 530768
rect 42670 530712 42675 530768
rect 41524 530710 42675 530712
rect 41524 530708 41530 530710
rect 42609 530707 42675 530710
rect 62297 530634 62363 530637
rect 682377 530634 682443 530637
rect 62297 530632 64706 530634
rect 62297 530576 62302 530632
rect 62358 530576 64706 530632
rect 62297 530574 64706 530576
rect 62297 530571 62363 530574
rect 64646 529990 64706 530574
rect 682334 530632 682443 530634
rect 682334 530576 682382 530632
rect 682438 530576 682443 530632
rect 682334 530571 682443 530576
rect 682334 530400 682394 530571
rect 676029 530022 676095 530025
rect 676029 530020 676292 530022
rect 676029 529964 676034 530020
rect 676090 529964 676292 530020
rect 676029 529962 676292 529964
rect 676029 529959 676095 529962
rect 42793 529818 42859 529821
rect 45277 529818 45343 529821
rect 42793 529816 45343 529818
rect 42793 529760 42798 529816
rect 42854 529760 45282 529816
rect 45338 529760 45343 529816
rect 42793 529758 45343 529760
rect 42793 529755 42859 529758
rect 45277 529755 45343 529758
rect 676262 529413 676322 529584
rect 676213 529408 676322 529413
rect 676213 529352 676218 529408
rect 676274 529352 676322 529408
rect 676213 529350 676322 529352
rect 676213 529347 676279 529350
rect 676029 529206 676095 529209
rect 676029 529204 676292 529206
rect 676029 529148 676034 529204
rect 676090 529148 676292 529204
rect 676029 529146 676292 529148
rect 676029 529143 676095 529146
rect 41822 528940 41828 529004
rect 41892 529002 41898 529004
rect 42425 529002 42491 529005
rect 41892 529000 42491 529002
rect 41892 528944 42430 529000
rect 42486 528944 42491 529000
rect 41892 528942 42491 528944
rect 41892 528940 41898 528942
rect 42425 528939 42491 528942
rect 62113 528594 62179 528597
rect 64646 528594 64706 528808
rect 676029 528798 676095 528801
rect 676029 528796 676292 528798
rect 676029 528740 676034 528796
rect 676090 528740 676292 528796
rect 676029 528738 676292 528740
rect 676029 528735 676095 528738
rect 62113 528592 64706 528594
rect 62113 528536 62118 528592
rect 62174 528536 64706 528592
rect 62113 528534 64706 528536
rect 683205 528594 683271 528597
rect 683205 528592 683314 528594
rect 683205 528536 683210 528592
rect 683266 528536 683314 528592
rect 62113 528531 62179 528534
rect 683205 528531 683314 528536
rect 683254 528360 683314 528531
rect 63217 528050 63283 528053
rect 63217 528048 64706 528050
rect 63217 527992 63222 528048
rect 63278 527992 64706 528048
rect 63217 527990 64706 527992
rect 63217 527987 63283 527990
rect 64646 527626 64706 527990
rect 676029 527982 676095 527985
rect 676029 527980 676292 527982
rect 676029 527924 676034 527980
rect 676090 527924 676292 527980
rect 676029 527922 676292 527924
rect 676029 527919 676095 527922
rect 683573 527778 683639 527781
rect 683573 527776 683682 527778
rect 683573 527720 683578 527776
rect 683634 527720 683682 527776
rect 683573 527715 683682 527720
rect 683622 527544 683682 527715
rect 45185 527234 45251 527237
rect 42566 527232 45251 527234
rect 42566 527176 45190 527232
rect 45246 527176 45251 527232
rect 42566 527174 45251 527176
rect 42566 526829 42626 527174
rect 45185 527171 45251 527174
rect 62113 527098 62179 527101
rect 62113 527096 64706 527098
rect 62113 527040 62118 527096
rect 62174 527040 64706 527096
rect 62113 527038 64706 527040
rect 62113 527035 62179 527038
rect 42566 526824 42675 526829
rect 42566 526768 42614 526824
rect 42670 526768 42675 526824
rect 42566 526766 42675 526768
rect 42609 526763 42675 526766
rect 64646 526444 64706 527038
rect 674414 527036 674420 527100
rect 674484 527098 674490 527100
rect 676262 527098 676322 527136
rect 674484 527038 676322 527098
rect 674484 527036 674490 527038
rect 683389 526962 683455 526965
rect 683389 526960 683498 526962
rect 683389 526904 683394 526960
rect 683450 526904 683498 526960
rect 683389 526899 683498 526904
rect 683438 526728 683498 526899
rect 673637 526418 673703 526421
rect 673637 526416 676322 526418
rect 673637 526360 673642 526416
rect 673698 526360 676322 526416
rect 673637 526358 676322 526360
rect 673637 526355 673703 526358
rect 676262 526320 676322 526358
rect 677918 525741 677978 525912
rect 62481 525738 62547 525741
rect 62481 525736 64706 525738
rect 62481 525680 62486 525736
rect 62542 525680 64706 525736
rect 62481 525678 64706 525680
rect 62481 525675 62547 525678
rect 64646 525262 64706 525678
rect 677869 525736 677978 525741
rect 677869 525680 677874 525736
rect 677930 525680 677978 525736
rect 677869 525678 677978 525680
rect 677869 525675 677935 525678
rect 683070 524925 683130 525504
rect 683070 524920 683179 524925
rect 683070 524864 683118 524920
rect 683174 524864 683179 524920
rect 683070 524862 683179 524864
rect 683113 524859 683179 524862
rect 680310 524517 680370 524688
rect 680310 524512 680419 524517
rect 680310 524456 680358 524512
rect 680414 524456 680419 524512
rect 680310 524454 680419 524456
rect 680353 524451 680419 524454
rect 676990 503644 676996 503708
rect 677060 503706 677066 503708
rect 683205 503706 683271 503709
rect 677060 503704 683271 503706
rect 677060 503648 683210 503704
rect 683266 503648 683271 503704
rect 677060 503646 683271 503648
rect 677060 503644 677066 503646
rect 683205 503643 683271 503646
rect 676806 500924 676812 500988
rect 676876 500986 676882 500988
rect 683389 500986 683455 500989
rect 676876 500984 683455 500986
rect 676876 500928 683394 500984
rect 683450 500928 683455 500984
rect 676876 500926 683455 500928
rect 676876 500924 676882 500926
rect 683389 500923 683455 500926
rect 673821 492146 673887 492149
rect 673821 492144 676292 492146
rect 673821 492088 673826 492144
rect 673882 492088 676292 492144
rect 673821 492086 676292 492088
rect 673821 492083 673887 492086
rect 676029 491738 676095 491741
rect 676029 491736 676292 491738
rect 676029 491680 676034 491736
rect 676090 491680 676292 491736
rect 676029 491678 676292 491680
rect 676029 491675 676095 491678
rect 674005 491330 674071 491333
rect 674005 491328 676292 491330
rect 674005 491272 674010 491328
rect 674066 491272 676292 491328
rect 674005 491270 676292 491272
rect 674005 491267 674071 491270
rect 674005 490922 674071 490925
rect 674005 490920 676292 490922
rect 674005 490864 674010 490920
rect 674066 490864 676292 490920
rect 674005 490862 676292 490864
rect 674005 490859 674071 490862
rect 672901 490514 672967 490517
rect 672901 490512 676292 490514
rect 672901 490456 672906 490512
rect 672962 490456 676292 490512
rect 672901 490454 676292 490456
rect 672901 490451 672967 490454
rect 672717 490106 672783 490109
rect 672717 490104 676292 490106
rect 672717 490048 672722 490104
rect 672778 490048 676292 490104
rect 672717 490046 676292 490048
rect 672717 490043 672783 490046
rect 674005 489698 674071 489701
rect 674005 489696 676292 489698
rect 674005 489640 674010 489696
rect 674066 489640 676292 489696
rect 674005 489638 676292 489640
rect 674005 489635 674071 489638
rect 674005 489290 674071 489293
rect 674005 489288 676292 489290
rect 674005 489232 674010 489288
rect 674066 489232 676292 489288
rect 674005 489230 676292 489232
rect 674005 489227 674071 489230
rect 676024 488820 676030 488884
rect 676094 488882 676100 488884
rect 676094 488822 676292 488882
rect 676094 488820 676100 488822
rect 674005 488474 674071 488477
rect 674005 488472 676292 488474
rect 674005 488416 674010 488472
rect 674066 488416 676292 488472
rect 674005 488414 676292 488416
rect 674005 488411 674071 488414
rect 676170 488006 676292 488066
rect 675886 487868 675892 487932
rect 675956 487930 675962 487932
rect 676170 487930 676230 488006
rect 675956 487870 676230 487930
rect 675956 487868 675962 487870
rect 681181 487658 681247 487661
rect 681181 487656 681260 487658
rect 681181 487600 681186 487656
rect 681242 487600 681260 487656
rect 681181 487598 681260 487600
rect 681181 487595 681247 487598
rect 679617 487250 679683 487253
rect 679604 487248 679683 487250
rect 679604 487192 679622 487248
rect 679678 487192 679683 487248
rect 679604 487190 679683 487192
rect 679617 487187 679683 487190
rect 676029 486842 676095 486845
rect 676029 486840 676292 486842
rect 676029 486784 676034 486840
rect 676090 486784 676292 486840
rect 676029 486782 676292 486784
rect 676029 486779 676095 486782
rect 680997 486434 681063 486437
rect 680997 486432 681076 486434
rect 680997 486376 681002 486432
rect 681058 486376 681076 486432
rect 680997 486374 681076 486376
rect 680997 486371 681063 486374
rect 674005 486026 674071 486029
rect 674005 486024 676292 486026
rect 674005 485968 674010 486024
rect 674066 485968 676292 486024
rect 674005 485966 676292 485968
rect 674005 485963 674071 485966
rect 683205 485618 683271 485621
rect 683205 485616 683284 485618
rect 683205 485560 683210 485616
rect 683266 485560 683284 485616
rect 683205 485558 683284 485560
rect 683205 485555 683271 485558
rect 676029 485210 676095 485213
rect 676029 485208 676292 485210
rect 676029 485152 676034 485208
rect 676090 485152 676292 485208
rect 676029 485150 676292 485152
rect 676029 485147 676095 485150
rect 673085 484802 673151 484805
rect 673085 484800 676292 484802
rect 673085 484744 673090 484800
rect 673146 484744 676292 484800
rect 673085 484742 676292 484744
rect 673085 484739 673151 484742
rect 673637 484394 673703 484397
rect 673637 484392 676292 484394
rect 673637 484336 673642 484392
rect 673698 484336 676292 484392
rect 673637 484334 676292 484336
rect 673637 484331 673703 484334
rect 676029 483986 676095 483989
rect 676029 483984 676292 483986
rect 676029 483928 676034 483984
rect 676090 483928 676292 483984
rect 676029 483926 676292 483928
rect 676029 483923 676095 483926
rect 683389 483578 683455 483581
rect 683389 483576 683468 483578
rect 683389 483520 683394 483576
rect 683450 483520 683468 483576
rect 683389 483518 683468 483520
rect 683389 483515 683455 483518
rect 674005 483170 674071 483173
rect 674005 483168 676292 483170
rect 674005 483112 674010 483168
rect 674066 483112 676292 483168
rect 674005 483110 676292 483112
rect 674005 483107 674071 483110
rect 676029 482762 676095 482765
rect 676029 482760 676292 482762
rect 676029 482704 676034 482760
rect 676090 482704 676292 482760
rect 676029 482702 676292 482704
rect 676029 482699 676095 482702
rect 676029 482354 676095 482357
rect 676029 482352 676292 482354
rect 676029 482296 676034 482352
rect 676090 482296 676292 482352
rect 676029 482294 676292 482296
rect 676029 482291 676095 482294
rect 680353 481946 680419 481949
rect 680340 481944 680419 481946
rect 680340 481888 680358 481944
rect 680414 481888 680419 481944
rect 680340 481886 680419 481888
rect 680353 481883 680419 481886
rect 677182 481130 677242 481508
rect 683113 481130 683179 481133
rect 677182 481128 683179 481130
rect 677182 481100 683118 481128
rect 677212 481072 683118 481100
rect 683174 481072 683179 481128
rect 677212 481070 683179 481072
rect 683113 481067 683179 481070
rect 675845 480722 675911 480725
rect 675845 480720 676292 480722
rect 675845 480664 675850 480720
rect 675906 480664 676292 480720
rect 675845 480662 676292 480664
rect 675845 480659 675911 480662
rect 669773 455426 669839 455429
rect 673269 455426 673335 455429
rect 669773 455424 673335 455426
rect 669773 455368 669778 455424
rect 669834 455368 673274 455424
rect 673330 455368 673335 455424
rect 669773 455366 673335 455368
rect 669773 455363 669839 455366
rect 673269 455363 673335 455366
rect 673381 455290 673447 455293
rect 673862 455290 673868 455292
rect 673381 455288 673868 455290
rect 673381 455232 673386 455288
rect 673442 455232 673868 455288
rect 673381 455230 673868 455232
rect 673381 455227 673447 455230
rect 673862 455228 673868 455230
rect 673932 455228 673938 455292
rect 670601 455154 670667 455157
rect 673269 455154 673335 455157
rect 670601 455152 673335 455154
rect 670601 455096 670606 455152
rect 670662 455096 673274 455152
rect 673330 455096 673335 455152
rect 670601 455094 673335 455096
rect 670601 455091 670667 455094
rect 673269 455091 673335 455094
rect 672809 454882 672875 454885
rect 674281 454882 674347 454885
rect 672809 454880 674347 454882
rect 672809 454824 672814 454880
rect 672870 454824 674286 454880
rect 674342 454824 674347 454880
rect 672809 454822 674347 454824
rect 672809 454819 672875 454822
rect 674281 454819 674347 454822
rect 673039 454610 673105 454613
rect 674281 454610 674347 454613
rect 673039 454608 674347 454610
rect 673039 454552 673044 454608
rect 673100 454552 674286 454608
rect 674342 454552 674347 454608
rect 673039 454550 674347 454552
rect 673039 454547 673105 454550
rect 674281 454547 674347 454550
rect 672947 454338 673013 454341
rect 674281 454338 674347 454341
rect 672947 454336 674347 454338
rect 672947 454280 672952 454336
rect 673008 454280 674286 454336
rect 674342 454280 674347 454336
rect 672947 454278 674347 454280
rect 672947 454275 673013 454278
rect 674281 454275 674347 454278
rect 672257 453930 672323 453933
rect 674281 453930 674347 453933
rect 672257 453928 674347 453930
rect 672257 453872 672262 453928
rect 672318 453872 674286 453928
rect 674342 453872 674347 453928
rect 672257 453870 674347 453872
rect 672257 453867 672323 453870
rect 674281 453867 674347 453870
rect 45277 430946 45343 430949
rect 41492 430944 45343 430946
rect 41492 430888 45282 430944
rect 45338 430888 45343 430944
rect 41492 430886 45343 430888
rect 45277 430883 45343 430886
rect 47761 430538 47827 430541
rect 41492 430536 47827 430538
rect 41492 430480 47766 430536
rect 47822 430480 47827 430536
rect 41492 430478 47827 430480
rect 47761 430475 47827 430478
rect 35801 430130 35867 430133
rect 35788 430128 35867 430130
rect 35788 430072 35806 430128
rect 35862 430072 35867 430128
rect 35788 430070 35867 430072
rect 35801 430067 35867 430070
rect 45001 429722 45067 429725
rect 41492 429720 45067 429722
rect 41492 429664 45006 429720
rect 45062 429664 45067 429720
rect 41492 429662 45067 429664
rect 45001 429659 45067 429662
rect 45093 429314 45159 429317
rect 41492 429312 45159 429314
rect 41492 429256 45098 429312
rect 45154 429256 45159 429312
rect 41492 429254 45159 429256
rect 45093 429251 45159 429254
rect 44633 428906 44699 428909
rect 41492 428904 44699 428906
rect 41492 428848 44638 428904
rect 44694 428848 44699 428904
rect 41492 428846 44699 428848
rect 44633 428843 44699 428846
rect 35801 428498 35867 428501
rect 35788 428496 35867 428498
rect 35788 428440 35806 428496
rect 35862 428440 35867 428496
rect 35788 428438 35867 428440
rect 35801 428435 35867 428438
rect 44357 428090 44423 428093
rect 41492 428088 44423 428090
rect 41492 428032 44362 428088
rect 44418 428032 44423 428088
rect 41492 428030 44423 428032
rect 44357 428027 44423 428030
rect 44357 427682 44423 427685
rect 41492 427680 44423 427682
rect 41492 427624 44362 427680
rect 44418 427624 44423 427680
rect 41492 427622 44423 427624
rect 44357 427619 44423 427622
rect 43161 427410 43227 427413
rect 41784 427408 43227 427410
rect 41784 427352 43166 427408
rect 43222 427352 43227 427408
rect 41784 427350 43227 427352
rect 41784 427274 41844 427350
rect 43161 427347 43227 427350
rect 41492 427214 41844 427274
rect 42149 427138 42215 427141
rect 63309 427138 63375 427141
rect 42149 427136 63375 427138
rect 42149 427080 42154 427136
rect 42210 427080 63314 427136
rect 63370 427080 63375 427136
rect 42149 427078 63375 427080
rect 42149 427075 42215 427078
rect 63309 427075 63375 427078
rect 44173 426866 44239 426869
rect 41492 426864 44239 426866
rect 41492 426808 44178 426864
rect 44234 426808 44239 426864
rect 41492 426806 44239 426808
rect 44173 426803 44239 426806
rect 41137 426458 41203 426461
rect 41124 426456 41203 426458
rect 41124 426400 41142 426456
rect 41198 426400 41203 426456
rect 41124 426398 41203 426400
rect 41137 426395 41203 426398
rect 41965 426458 42031 426461
rect 42793 426458 42859 426461
rect 41965 426456 42859 426458
rect 41965 426400 41970 426456
rect 42026 426400 42798 426456
rect 42854 426400 42859 426456
rect 41965 426398 42859 426400
rect 41965 426395 42031 426398
rect 42793 426395 42859 426398
rect 40953 426050 41019 426053
rect 40940 426048 41019 426050
rect 40940 425992 40958 426048
rect 41014 425992 41019 426048
rect 40940 425990 41019 425992
rect 40953 425987 41019 425990
rect 39297 425642 39363 425645
rect 39284 425640 39363 425642
rect 39284 425584 39302 425640
rect 39358 425584 39363 425640
rect 39284 425582 39363 425584
rect 39297 425579 39363 425582
rect 42977 425234 43043 425237
rect 41492 425232 43043 425234
rect 41492 425176 42982 425232
rect 43038 425176 43043 425232
rect 41492 425174 43043 425176
rect 42977 425171 43043 425174
rect 32029 424826 32095 424829
rect 32029 424824 32108 424826
rect 32029 424768 32034 424824
rect 32090 424768 32108 424824
rect 32029 424766 32108 424768
rect 32029 424763 32095 424766
rect 34513 424418 34579 424421
rect 34500 424416 34579 424418
rect 34500 424360 34518 424416
rect 34574 424360 34579 424416
rect 34500 424358 34579 424360
rect 34513 424355 34579 424358
rect 33777 424010 33843 424013
rect 33764 424008 33843 424010
rect 33764 423952 33782 424008
rect 33838 423952 33843 424008
rect 33764 423950 33843 423952
rect 33777 423947 33843 423950
rect 41137 423602 41203 423605
rect 41124 423600 41203 423602
rect 41124 423544 41142 423600
rect 41198 423544 41203 423600
rect 41124 423542 41203 423544
rect 41137 423539 41203 423542
rect 41781 423604 41847 423605
rect 41781 423600 41828 423604
rect 41892 423602 41898 423604
rect 41781 423544 41786 423600
rect 41781 423540 41828 423544
rect 41892 423542 41938 423602
rect 41892 423540 41898 423542
rect 41781 423539 41847 423540
rect 44541 423194 44607 423197
rect 41492 423192 44607 423194
rect 41492 423136 44546 423192
rect 44602 423136 44607 423192
rect 41492 423134 44607 423136
rect 44541 423131 44607 423134
rect 43161 422786 43227 422789
rect 41492 422784 43227 422786
rect 41492 422728 43166 422784
rect 43222 422728 43227 422784
rect 41492 422726 43227 422728
rect 43161 422723 43227 422726
rect 41781 422378 41847 422381
rect 43805 422378 43871 422381
rect 41781 422376 43871 422378
rect 40910 422312 40970 422348
rect 41781 422320 41786 422376
rect 41842 422320 43810 422376
rect 43866 422320 43871 422376
rect 41781 422318 43871 422320
rect 41781 422315 41847 422318
rect 43805 422315 43871 422318
rect 40902 422248 40908 422312
rect 40972 422248 40978 422312
rect 41781 421970 41847 421973
rect 41492 421968 41847 421970
rect 41492 421912 41786 421968
rect 41842 421912 41847 421968
rect 41492 421910 41847 421912
rect 41781 421907 41847 421910
rect 41781 421562 41847 421565
rect 41492 421560 41847 421562
rect 41492 421504 41786 421560
rect 41842 421504 41847 421560
rect 41492 421502 41847 421504
rect 41781 421499 41847 421502
rect 43989 421154 44055 421157
rect 41492 421152 44055 421154
rect 41492 421096 43994 421152
rect 44050 421096 44055 421152
rect 41492 421094 44055 421096
rect 43989 421091 44055 421094
rect 45461 420746 45527 420749
rect 41492 420744 45527 420746
rect 41492 420688 45466 420744
rect 45522 420688 45527 420744
rect 41492 420686 45527 420688
rect 45461 420683 45527 420686
rect 41462 419930 41522 420308
rect 47577 419930 47643 419933
rect 41462 419928 47643 419930
rect 41462 419900 47582 419928
rect 41492 419872 47582 419900
rect 47638 419872 47643 419928
rect 41492 419870 47643 419872
rect 47577 419867 47643 419870
rect 40718 418644 40724 418708
rect 40788 418706 40794 418708
rect 41597 418706 41663 418709
rect 40788 418704 41663 418706
rect 40788 418648 41602 418704
rect 41658 418648 41663 418704
rect 40788 418646 41663 418648
rect 40788 418644 40794 418646
rect 41597 418643 41663 418646
rect 40534 418372 40540 418436
rect 40604 418434 40610 418436
rect 41781 418434 41847 418437
rect 40604 418432 41847 418434
rect 40604 418376 41786 418432
rect 41842 418376 41847 418432
rect 40604 418374 41847 418376
rect 40604 418372 40610 418374
rect 41781 418371 41847 418374
rect 39297 415306 39363 415309
rect 42006 415306 42012 415308
rect 39297 415304 42012 415306
rect 39297 415248 39302 415304
rect 39358 415248 42012 415304
rect 39297 415246 42012 415248
rect 39297 415243 39363 415246
rect 42006 415244 42012 415246
rect 42076 415244 42082 415308
rect 33777 414626 33843 414629
rect 41822 414626 41828 414628
rect 33777 414624 41828 414626
rect 33777 414568 33782 414624
rect 33838 414568 41828 414624
rect 33777 414566 41828 414568
rect 33777 414563 33843 414566
rect 41822 414564 41828 414566
rect 41892 414564 41898 414628
rect 42057 408098 42123 408101
rect 43989 408098 44055 408101
rect 42057 408096 44055 408098
rect 42057 408040 42062 408096
rect 42118 408040 43994 408096
rect 44050 408040 44055 408096
rect 42057 408038 44055 408040
rect 42057 408035 42123 408038
rect 43989 408035 44055 408038
rect 42425 407282 42491 407285
rect 44725 407282 44791 407285
rect 42425 407280 44791 407282
rect 42425 407224 42430 407280
rect 42486 407224 44730 407280
rect 44786 407224 44791 407280
rect 42425 407222 44791 407224
rect 42425 407219 42491 407222
rect 44725 407219 44791 407222
rect 40902 406948 40908 407012
rect 40972 407010 40978 407012
rect 41781 407010 41847 407013
rect 40972 407008 41847 407010
rect 40972 406952 41786 407008
rect 41842 406952 41847 407008
rect 40972 406950 41847 406952
rect 40972 406948 40978 406950
rect 41781 406947 41847 406950
rect 40534 406676 40540 406740
rect 40604 406738 40610 406740
rect 41781 406738 41847 406741
rect 40604 406736 41847 406738
rect 40604 406680 41786 406736
rect 41842 406680 41847 406736
rect 40604 406678 41847 406680
rect 40604 406676 40610 406678
rect 41781 406675 41847 406678
rect 42425 404970 42491 404973
rect 51441 404970 51507 404973
rect 42425 404968 51507 404970
rect 42425 404912 42430 404968
rect 42486 404912 51446 404968
rect 51502 404912 51507 404968
rect 42425 404910 51507 404912
rect 42425 404907 42491 404910
rect 51441 404907 51507 404910
rect 40718 404500 40724 404564
rect 40788 404562 40794 404564
rect 42241 404562 42307 404565
rect 40788 404560 42307 404562
rect 40788 404504 42246 404560
rect 42302 404504 42307 404560
rect 40788 404502 42307 404504
rect 40788 404500 40794 404502
rect 42241 404499 42307 404502
rect 62113 404154 62179 404157
rect 62113 404152 64706 404154
rect 62113 404096 62118 404152
rect 62174 404096 64706 404152
rect 62113 404094 64706 404096
rect 62113 404091 62179 404094
rect 64646 403550 64706 404094
rect 676262 403746 676322 403852
rect 663750 403686 676322 403746
rect 657537 403338 657603 403341
rect 663750 403338 663810 403686
rect 676262 403341 676322 403444
rect 657537 403336 663810 403338
rect 657537 403280 657542 403336
rect 657598 403280 663810 403336
rect 657537 403278 663810 403280
rect 676213 403336 676322 403341
rect 676213 403280 676218 403336
rect 676274 403280 676322 403336
rect 676213 403278 676322 403280
rect 657537 403275 657603 403278
rect 676213 403275 676279 403278
rect 676630 402933 676690 403036
rect 42333 402930 42399 402933
rect 44541 402930 44607 402933
rect 42333 402928 44607 402930
rect 42333 402872 42338 402928
rect 42394 402872 44546 402928
rect 44602 402872 44607 402928
rect 42333 402870 44607 402872
rect 42333 402867 42399 402870
rect 44541 402867 44607 402870
rect 676581 402928 676690 402933
rect 676581 402872 676586 402928
rect 676642 402872 676690 402928
rect 676581 402870 676690 402872
rect 676581 402867 676647 402870
rect 62113 402658 62179 402661
rect 62113 402656 64706 402658
rect 62113 402600 62118 402656
rect 62174 402600 64706 402656
rect 62113 402598 64706 402600
rect 62113 402595 62179 402598
rect 42241 402522 42307 402525
rect 43805 402522 43871 402525
rect 42241 402520 43871 402522
rect 42241 402464 42246 402520
rect 42302 402464 43810 402520
rect 43866 402464 43871 402520
rect 42241 402462 43871 402464
rect 42241 402459 42307 402462
rect 43805 402459 43871 402462
rect 64646 402368 64706 402598
rect 672625 402522 672691 402525
rect 676262 402522 676322 402628
rect 672625 402520 676322 402522
rect 672625 402464 672630 402520
rect 672686 402464 676322 402520
rect 672625 402462 676322 402464
rect 672625 402459 672691 402462
rect 674833 402250 674899 402253
rect 674833 402248 676292 402250
rect 674833 402192 674838 402248
rect 674894 402192 676292 402248
rect 674833 402190 676292 402192
rect 674833 402187 674899 402190
rect 672441 401978 672507 401981
rect 672441 401976 676322 401978
rect 672441 401920 672446 401976
rect 672502 401920 676322 401976
rect 672441 401918 676322 401920
rect 672441 401915 672507 401918
rect 676262 401812 676322 401918
rect 673177 401706 673243 401709
rect 674833 401706 674899 401709
rect 673177 401704 674899 401706
rect 673177 401648 673182 401704
rect 673238 401648 674838 401704
rect 674894 401648 674899 401704
rect 673177 401646 674899 401648
rect 673177 401643 673243 401646
rect 674833 401643 674899 401646
rect 673913 401434 673979 401437
rect 673913 401432 676292 401434
rect 673913 401376 673918 401432
rect 673974 401376 676292 401432
rect 673913 401374 676292 401376
rect 673913 401371 673979 401374
rect 677174 401236 677180 401300
rect 677244 401236 677250 401300
rect 62113 400754 62179 400757
rect 64646 400754 64706 401186
rect 677182 400996 677242 401236
rect 652017 400890 652083 400893
rect 676581 400890 676647 400893
rect 652017 400888 676647 400890
rect 652017 400832 652022 400888
rect 652078 400832 676586 400888
rect 676642 400832 676647 400888
rect 652017 400830 676647 400832
rect 652017 400827 652083 400830
rect 676581 400827 676647 400830
rect 62113 400752 64706 400754
rect 62113 400696 62118 400752
rect 62174 400696 64706 400752
rect 62113 400694 64706 400696
rect 62113 400691 62179 400694
rect 673361 400482 673427 400485
rect 676262 400482 676322 400588
rect 673361 400480 676322 400482
rect 673361 400424 673366 400480
rect 673422 400424 676322 400480
rect 673361 400422 676322 400424
rect 673361 400419 673427 400422
rect 676806 400420 676812 400484
rect 676876 400420 676882 400484
rect 63309 400210 63375 400213
rect 63309 400208 64706 400210
rect 63309 400152 63314 400208
rect 63370 400152 64706 400208
rect 676814 400180 676874 400420
rect 63309 400150 64706 400152
rect 63309 400147 63375 400150
rect 41454 400012 41460 400076
rect 41524 400074 41530 400076
rect 41781 400074 41847 400077
rect 41524 400072 41847 400074
rect 41524 400016 41786 400072
rect 41842 400016 41847 400072
rect 41524 400014 41847 400016
rect 41524 400012 41530 400014
rect 41781 400011 41847 400014
rect 64646 400004 64706 400150
rect 672809 399666 672875 399669
rect 676262 399666 676322 399772
rect 672809 399664 676322 399666
rect 672809 399608 672814 399664
rect 672870 399608 676322 399664
rect 672809 399606 676322 399608
rect 672809 399603 672875 399606
rect 41781 399396 41847 399397
rect 41781 399392 41828 399396
rect 41892 399394 41898 399396
rect 62113 399394 62179 399397
rect 676029 399394 676095 399397
rect 41781 399336 41786 399392
rect 41781 399332 41828 399336
rect 41892 399334 41938 399394
rect 62113 399392 64706 399394
rect 62113 399336 62118 399392
rect 62174 399336 64706 399392
rect 62113 399334 64706 399336
rect 41892 399332 41898 399334
rect 41781 399331 41847 399332
rect 62113 399331 62179 399334
rect 41965 398852 42031 398853
rect 41965 398848 42012 398852
rect 42076 398850 42082 398852
rect 41965 398792 41970 398848
rect 41965 398788 42012 398792
rect 42076 398790 42122 398850
rect 64646 398822 64706 399334
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 42076 398788 42082 398790
rect 676070 398788 676076 398852
rect 676140 398850 676146 398852
rect 676262 398850 676322 398956
rect 676140 398790 676322 398850
rect 676140 398788 676146 398790
rect 41965 398787 42031 398788
rect 679574 398445 679634 398548
rect 679574 398440 679683 398445
rect 679574 398384 679622 398440
rect 679678 398384 679683 398440
rect 679574 398382 679683 398384
rect 679617 398379 679683 398382
rect 62113 398306 62179 398309
rect 62113 398304 64706 398306
rect 62113 398248 62118 398304
rect 62174 398248 64706 398304
rect 62113 398246 64706 398248
rect 62113 398243 62179 398246
rect 64646 397640 64706 398246
rect 676262 398037 676322 398140
rect 676213 398032 676322 398037
rect 676213 397976 676218 398032
rect 676274 397976 676322 398032
rect 676213 397974 676322 397976
rect 676213 397971 676279 397974
rect 678286 397629 678346 397732
rect 678237 397624 678346 397629
rect 678237 397568 678242 397624
rect 678298 397568 678346 397624
rect 678237 397566 678346 397568
rect 678237 397563 678303 397566
rect 674741 397354 674807 397357
rect 674741 397352 676292 397354
rect 674741 397296 674746 397352
rect 674802 397296 676292 397352
rect 674741 397294 676292 397296
rect 674741 397291 674807 397294
rect 676262 396812 676322 396916
rect 676254 396748 676260 396812
rect 676324 396748 676330 396812
rect 652201 396674 652267 396677
rect 674557 396674 674623 396677
rect 652201 396672 674623 396674
rect 652201 396616 652206 396672
rect 652262 396616 674562 396672
rect 674618 396616 674623 396672
rect 652201 396614 674623 396616
rect 652201 396611 652267 396614
rect 674557 396611 674623 396614
rect 676446 396404 676506 396508
rect 676438 396340 676444 396404
rect 676508 396340 676514 396404
rect 676029 396130 676095 396133
rect 676029 396128 676292 396130
rect 676029 396072 676034 396128
rect 676090 396072 676292 396128
rect 676029 396070 676292 396072
rect 676029 396067 676095 396070
rect 42149 395722 42215 395725
rect 51073 395722 51139 395725
rect 42149 395720 51139 395722
rect 42149 395664 42154 395720
rect 42210 395664 51078 395720
rect 51134 395664 51139 395720
rect 42149 395662 51139 395664
rect 42149 395659 42215 395662
rect 51073 395659 51139 395662
rect 673729 395722 673795 395725
rect 673729 395720 676292 395722
rect 673729 395664 673734 395720
rect 673790 395664 676292 395720
rect 673729 395662 676292 395664
rect 673729 395659 673795 395662
rect 676630 395180 676690 395284
rect 676622 395116 676628 395180
rect 676692 395116 676698 395180
rect 672993 395042 673059 395045
rect 672993 395040 676322 395042
rect 672993 394984 672998 395040
rect 673054 394984 676322 395040
rect 672993 394982 676322 394984
rect 672993 394979 673059 394982
rect 676262 394876 676322 394982
rect 676262 394365 676322 394468
rect 676213 394360 676322 394365
rect 676213 394304 676218 394360
rect 676274 394304 676322 394360
rect 676213 394302 676322 394304
rect 676213 394299 676279 394302
rect 672625 393954 672691 393957
rect 676262 393954 676322 394060
rect 672625 393952 676322 393954
rect 672625 393896 672630 393952
rect 672686 393896 676322 393952
rect 672625 393894 676322 393896
rect 672625 393891 672691 393894
rect 671889 393682 671955 393685
rect 671889 393680 676292 393682
rect 671889 393624 671894 393680
rect 671950 393624 676292 393680
rect 671889 393622 676292 393624
rect 671889 393619 671955 393622
rect 675334 392804 675340 392868
rect 675404 392866 675410 392868
rect 676262 392866 676322 393244
rect 675404 392836 676322 392866
rect 675404 392806 676292 392836
rect 675404 392804 675410 392806
rect 670509 392594 670575 392597
rect 670509 392592 676322 392594
rect 670509 392536 670514 392592
rect 670570 392536 676322 392592
rect 670509 392534 676322 392536
rect 670509 392531 670575 392534
rect 676262 392428 676322 392534
rect 47761 387698 47827 387701
rect 41492 387696 47827 387698
rect 41492 387640 47766 387696
rect 47822 387640 47827 387696
rect 41492 387638 47827 387640
rect 47761 387635 47827 387638
rect 675886 387636 675892 387700
rect 675956 387698 675962 387700
rect 678237 387698 678303 387701
rect 675956 387696 678303 387698
rect 675956 387640 678242 387696
rect 678298 387640 678303 387696
rect 675956 387638 678303 387640
rect 675956 387636 675962 387638
rect 678237 387635 678303 387638
rect 41278 387157 41338 387260
rect 41278 387152 41387 387157
rect 41278 387096 41326 387152
rect 41382 387096 41387 387152
rect 41278 387094 41387 387096
rect 41321 387091 41387 387094
rect 41094 386749 41154 386852
rect 41094 386744 41203 386749
rect 41094 386688 41142 386744
rect 41198 386688 41203 386744
rect 41094 386686 41203 386688
rect 41137 386683 41203 386686
rect 45093 386474 45159 386477
rect 41492 386472 45159 386474
rect 41492 386416 45098 386472
rect 45154 386416 45159 386472
rect 41492 386414 45159 386416
rect 45093 386411 45159 386414
rect 40910 385933 40970 386036
rect 40910 385928 41019 385933
rect 40910 385872 40958 385928
rect 41014 385872 41019 385928
rect 40910 385870 41019 385872
rect 40953 385867 41019 385870
rect 41137 385930 41203 385933
rect 63217 385930 63283 385933
rect 41137 385928 63283 385930
rect 41137 385872 41142 385928
rect 41198 385872 63222 385928
rect 63278 385872 63283 385928
rect 41137 385870 63283 385872
rect 41137 385867 41203 385870
rect 63217 385867 63283 385870
rect 42793 385658 42859 385661
rect 41492 385656 42859 385658
rect 41492 385600 42798 385656
rect 42854 385600 42859 385656
rect 41492 385598 42859 385600
rect 42793 385595 42859 385598
rect 43253 385250 43319 385253
rect 41492 385248 43319 385250
rect 41492 385192 43258 385248
rect 43314 385192 43319 385248
rect 41492 385190 43319 385192
rect 43253 385187 43319 385190
rect 675753 384978 675819 384981
rect 676254 384978 676260 384980
rect 675753 384976 676260 384978
rect 675753 384920 675758 384976
rect 675814 384920 676260 384976
rect 675753 384918 676260 384920
rect 675753 384915 675819 384918
rect 676254 384916 676260 384918
rect 676324 384916 676330 384980
rect 44357 384842 44423 384845
rect 41492 384840 44423 384842
rect 41492 384784 44362 384840
rect 44418 384784 44423 384840
rect 41492 384782 44423 384784
rect 44357 384779 44423 384782
rect 45185 384434 45251 384437
rect 41492 384432 45251 384434
rect 41492 384376 45190 384432
rect 45246 384376 45251 384432
rect 41492 384374 45251 384376
rect 45185 384371 45251 384374
rect 44173 384026 44239 384029
rect 41492 384024 44239 384026
rect 41492 383968 44178 384024
rect 44234 383968 44239 384024
rect 41492 383966 44239 383968
rect 44173 383963 44239 383966
rect 45093 383618 45159 383621
rect 41492 383616 45159 383618
rect 41492 383560 45098 383616
rect 45154 383560 45159 383616
rect 41492 383558 45159 383560
rect 45093 383555 45159 383558
rect 41094 383077 41154 383180
rect 41094 383072 41203 383077
rect 41094 383016 41142 383072
rect 41198 383016 41203 383072
rect 41094 383014 41203 383016
rect 41137 383011 41203 383014
rect 654777 382938 654843 382941
rect 675109 382938 675175 382941
rect 654777 382936 675175 382938
rect 654777 382880 654782 382936
rect 654838 382880 675114 382936
rect 675170 382880 675175 382936
rect 654777 382878 675175 382880
rect 654777 382875 654843 382878
rect 675109 382875 675175 382878
rect 41278 382669 41338 382772
rect 41278 382664 41387 382669
rect 41278 382608 41326 382664
rect 41382 382608 41387 382664
rect 41278 382606 41387 382608
rect 41321 382603 41387 382606
rect 39990 382261 40050 382364
rect 39990 382256 40099 382261
rect 39990 382200 40038 382256
rect 40094 382200 40099 382256
rect 39990 382198 40099 382200
rect 40033 382195 40099 382198
rect 40953 382258 41019 382261
rect 44909 382258 44975 382261
rect 40953 382256 44975 382258
rect 40953 382200 40958 382256
rect 41014 382200 44914 382256
rect 44970 382200 44975 382256
rect 40953 382198 44975 382200
rect 40953 382195 41019 382198
rect 44909 382195 44975 382198
rect 675753 382258 675819 382261
rect 676438 382258 676444 382260
rect 675753 382256 676444 382258
rect 675753 382200 675758 382256
rect 675814 382200 676444 382256
rect 675753 382198 676444 382200
rect 675753 382195 675819 382198
rect 676438 382196 676444 382198
rect 676508 382196 676514 382260
rect 35390 381853 35450 381956
rect 35390 381848 35499 381853
rect 35390 381792 35438 381848
rect 35494 381792 35499 381848
rect 35390 381790 35499 381792
rect 35433 381787 35499 381790
rect 41137 381850 41203 381853
rect 41454 381850 41460 381852
rect 41137 381848 41460 381850
rect 41137 381792 41142 381848
rect 41198 381792 41460 381848
rect 41137 381790 41460 381792
rect 41137 381787 41203 381790
rect 41454 381788 41460 381790
rect 41524 381788 41530 381852
rect 41873 381578 41939 381581
rect 62481 381578 62547 381581
rect 41873 381576 62547 381578
rect 39254 381445 39314 381548
rect 41873 381520 41878 381576
rect 41934 381520 62486 381576
rect 62542 381520 62547 381576
rect 41873 381518 62547 381520
rect 41873 381515 41939 381518
rect 62481 381515 62547 381518
rect 39254 381440 39363 381445
rect 39254 381384 39302 381440
rect 39358 381384 39363 381440
rect 39254 381382 39363 381384
rect 39297 381379 39363 381382
rect 33918 381037 33978 381140
rect 33918 381032 34027 381037
rect 33918 380976 33966 381032
rect 34022 380976 34027 381032
rect 33918 380974 34027 380976
rect 33961 380971 34027 380974
rect 672993 381034 673059 381037
rect 675385 381034 675451 381037
rect 672993 381032 675451 381034
rect 672993 380976 672998 381032
rect 673054 380976 675390 381032
rect 675446 380976 675451 381032
rect 672993 380974 675451 380976
rect 672993 380971 673059 380974
rect 675385 380971 675451 380974
rect 42885 380762 42951 380765
rect 41492 380760 42951 380762
rect 41492 380704 42890 380760
rect 42946 380704 42951 380760
rect 41492 380702 42951 380704
rect 42885 380699 42951 380702
rect 44633 380354 44699 380357
rect 41492 380352 44699 380354
rect 41492 380296 44638 380352
rect 44694 380296 44699 380352
rect 41492 380294 44699 380296
rect 44633 380291 44699 380294
rect 41278 379813 41338 379916
rect 41278 379808 41387 379813
rect 41278 379752 41326 379808
rect 41382 379752 41387 379808
rect 41278 379750 41387 379752
rect 41321 379747 41387 379750
rect 41505 379810 41571 379813
rect 43805 379810 43871 379813
rect 41505 379808 43871 379810
rect 41505 379752 41510 379808
rect 41566 379752 43810 379808
rect 43866 379752 43871 379808
rect 41505 379750 43871 379752
rect 41505 379747 41571 379750
rect 43805 379747 43871 379750
rect 35758 379405 35818 379530
rect 35758 379400 35867 379405
rect 35758 379344 35806 379400
rect 35862 379344 35867 379400
rect 35758 379342 35867 379344
rect 35801 379339 35867 379342
rect 40033 379402 40099 379405
rect 41638 379402 41644 379404
rect 40033 379400 41644 379402
rect 40033 379344 40038 379400
rect 40094 379344 41644 379400
rect 40033 379342 41644 379344
rect 40033 379339 40099 379342
rect 41638 379340 41644 379342
rect 41708 379340 41714 379404
rect 40726 378996 40786 379100
rect 40718 378932 40724 378996
rect 40788 378932 40794 378996
rect 40542 378588 40602 378692
rect 40534 378524 40540 378588
rect 40604 378524 40610 378588
rect 675661 378586 675727 378589
rect 675886 378586 675892 378588
rect 675661 378584 675892 378586
rect 675661 378528 675666 378584
rect 675722 378528 675892 378584
rect 675661 378526 675892 378528
rect 675661 378523 675727 378526
rect 675886 378524 675892 378526
rect 675956 378524 675962 378588
rect 35758 378181 35818 378284
rect 35758 378176 35867 378181
rect 35758 378120 35806 378176
rect 35862 378120 35867 378176
rect 35758 378118 35867 378120
rect 35801 378115 35867 378118
rect 41689 378178 41755 378181
rect 43989 378178 44055 378181
rect 41689 378176 44055 378178
rect 41689 378120 41694 378176
rect 41750 378120 43994 378176
rect 44050 378120 44055 378176
rect 41689 378118 44055 378120
rect 41689 378115 41755 378118
rect 43989 378115 44055 378118
rect 40910 377772 40970 377876
rect 40902 377708 40908 377772
rect 40972 377708 40978 377772
rect 44265 377498 44331 377501
rect 41492 377496 44331 377498
rect 41492 377440 44270 377496
rect 44326 377440 44331 377496
rect 41492 377438 44331 377440
rect 44265 377435 44331 377438
rect 675753 377498 675819 377501
rect 676622 377498 676628 377500
rect 675753 377496 676628 377498
rect 675753 377440 675758 377496
rect 675814 377440 676628 377496
rect 675753 377438 676628 377440
rect 675753 377435 675819 377438
rect 676622 377436 676628 377438
rect 676692 377436 676698 377500
rect 35758 376549 35818 377060
rect 40401 376954 40467 376957
rect 43069 376954 43135 376957
rect 40401 376952 43135 376954
rect 40401 376896 40406 376952
rect 40462 376896 43074 376952
rect 43130 376896 43135 376952
rect 40401 376894 43135 376896
rect 40401 376891 40467 376894
rect 43069 376891 43135 376894
rect 35758 376544 35867 376549
rect 35758 376488 35806 376544
rect 35862 376488 35867 376544
rect 35758 376486 35867 376488
rect 41462 376546 41522 376652
rect 41462 376486 41890 376546
rect 35801 376483 35867 376486
rect 35801 376138 35867 376141
rect 41830 376138 41890 376486
rect 672625 376274 672691 376277
rect 675385 376274 675451 376277
rect 672625 376272 675451 376274
rect 672625 376216 672630 376272
rect 672686 376216 675390 376272
rect 675446 376216 675451 376272
rect 672625 376214 675451 376216
rect 672625 376211 672691 376214
rect 675385 376211 675451 376214
rect 46381 376138 46447 376141
rect 35801 376136 46447 376138
rect 35801 376080 35806 376136
rect 35862 376080 46386 376136
rect 46442 376080 46447 376136
rect 35801 376078 46447 376080
rect 35801 376075 35867 376078
rect 46381 376075 46447 376078
rect 673729 375458 673795 375461
rect 675109 375458 675175 375461
rect 673729 375456 675175 375458
rect 673729 375400 673734 375456
rect 673790 375400 675114 375456
rect 675170 375400 675175 375456
rect 673729 375398 675175 375400
rect 673729 375395 673795 375398
rect 675109 375395 675175 375398
rect 35433 374642 35499 374645
rect 41822 374642 41828 374644
rect 35433 374640 41828 374642
rect 35433 374584 35438 374640
rect 35494 374584 41828 374640
rect 35433 374582 41828 374584
rect 35433 374579 35499 374582
rect 41822 374580 41828 374582
rect 41892 374580 41898 374644
rect 652201 373962 652267 373965
rect 649950 373960 652267 373962
rect 649950 373904 652206 373960
rect 652262 373904 652267 373960
rect 649950 373902 652267 373904
rect 649950 373892 650010 373902
rect 652201 373899 652267 373902
rect 675753 373690 675819 373693
rect 676070 373690 676076 373692
rect 675753 373688 676076 373690
rect 675753 373632 675758 373688
rect 675814 373632 676076 373688
rect 675753 373630 676076 373632
rect 675753 373627 675819 373630
rect 676070 373628 676076 373630
rect 676140 373628 676146 373692
rect 651465 373282 651531 373285
rect 649950 373280 651531 373282
rect 649950 373224 651470 373280
rect 651526 373224 651531 373280
rect 649950 373222 651531 373224
rect 649950 372710 650010 373222
rect 651465 373219 651531 373222
rect 675109 372874 675175 372877
rect 675334 372874 675340 372876
rect 675109 372872 675340 372874
rect 675109 372816 675114 372872
rect 675170 372816 675340 372872
rect 675109 372814 675340 372816
rect 675109 372811 675175 372814
rect 675334 372812 675340 372814
rect 675404 372812 675410 372876
rect 652017 372194 652083 372197
rect 649950 372192 652083 372194
rect 649950 372136 652022 372192
rect 652078 372136 652083 372192
rect 649950 372134 652083 372136
rect 649950 371528 650010 372134
rect 652017 372131 652083 372134
rect 668577 371242 668643 371245
rect 675017 371242 675083 371245
rect 668577 371240 675083 371242
rect 668577 371184 668582 371240
rect 668638 371184 675022 371240
rect 675078 371184 675083 371240
rect 668577 371182 675083 371184
rect 668577 371179 668643 371182
rect 675017 371179 675083 371182
rect 651465 370698 651531 370701
rect 649950 370696 651531 370698
rect 649950 370640 651470 370696
rect 651526 370640 651531 370696
rect 649950 370638 651531 370640
rect 649950 370346 650010 370638
rect 651465 370635 651531 370638
rect 40902 364788 40908 364852
rect 40972 364850 40978 364852
rect 41781 364850 41847 364853
rect 40972 364848 41847 364850
rect 40972 364792 41786 364848
rect 41842 364792 41847 364848
rect 40972 364790 41847 364792
rect 40972 364788 40978 364790
rect 41781 364787 41847 364790
rect 40718 364108 40724 364172
rect 40788 364170 40794 364172
rect 41781 364170 41847 364173
rect 40788 364168 41847 364170
rect 40788 364112 41786 364168
rect 41842 364112 41847 364168
rect 40788 364110 41847 364112
rect 40788 364108 40794 364110
rect 41781 364107 41847 364110
rect 42149 363626 42215 363629
rect 43989 363626 44055 363629
rect 42149 363624 44055 363626
rect 42149 363568 42154 363624
rect 42210 363568 43994 363624
rect 44050 363568 44055 363624
rect 42149 363566 44055 363568
rect 42149 363563 42215 363566
rect 43989 363563 44055 363566
rect 42701 363082 42767 363085
rect 44633 363082 44699 363085
rect 42701 363080 44699 363082
rect 42701 363024 42706 363080
rect 42762 363024 44638 363080
rect 44694 363024 44699 363080
rect 42701 363022 44699 363024
rect 42701 363019 42767 363022
rect 44633 363019 44699 363022
rect 42701 362266 42767 362269
rect 51073 362266 51139 362269
rect 42701 362264 51139 362266
rect 42701 362208 42706 362264
rect 42762 362208 51078 362264
rect 51134 362208 51139 362264
rect 42701 362206 51139 362208
rect 42701 362203 42767 362206
rect 51073 362203 51139 362206
rect 62113 360906 62179 360909
rect 62113 360904 64706 360906
rect 62113 360848 62118 360904
rect 62174 360848 64706 360904
rect 62113 360846 64706 360848
rect 62113 360843 62179 360846
rect 64646 360328 64706 360846
rect 40534 360028 40540 360092
rect 40604 360090 40610 360092
rect 41781 360090 41847 360093
rect 40604 360088 41847 360090
rect 40604 360032 41786 360088
rect 41842 360032 41847 360088
rect 40604 360030 41847 360032
rect 40604 360028 40610 360030
rect 41781 360027 41847 360030
rect 42149 359954 42215 359957
rect 43805 359954 43871 359957
rect 42149 359952 43871 359954
rect 42149 359896 42154 359952
rect 42210 359896 43810 359952
rect 43866 359896 43871 359952
rect 42149 359894 43871 359896
rect 42149 359891 42215 359894
rect 43805 359891 43871 359894
rect 62113 359818 62179 359821
rect 62113 359816 64706 359818
rect 62113 359760 62118 359816
rect 62174 359760 64706 359816
rect 62113 359758 64706 359760
rect 62113 359755 62179 359758
rect 64646 359146 64706 359758
rect 42425 359002 42491 359005
rect 44449 359002 44515 359005
rect 42425 359000 44515 359002
rect 42425 358944 42430 359000
rect 42486 358944 44454 359000
rect 44510 358944 44515 359000
rect 42425 358942 44515 358944
rect 42425 358939 42491 358942
rect 44449 358939 44515 358942
rect 41873 358732 41939 358733
rect 41822 358730 41828 358732
rect 41782 358670 41828 358730
rect 41892 358728 41939 358732
rect 41934 358672 41939 358728
rect 41822 358668 41828 358670
rect 41892 358668 41939 358672
rect 41873 358667 41939 358668
rect 663750 358670 676292 358730
rect 654777 358594 654843 358597
rect 663750 358594 663810 358670
rect 654777 358592 663810 358594
rect 654777 358536 654782 358592
rect 654838 358536 663810 358592
rect 654777 358534 663810 358536
rect 654777 358531 654843 358534
rect 674097 358322 674163 358325
rect 674097 358320 676292 358322
rect 674097 358264 674102 358320
rect 674158 358264 676292 358320
rect 674097 358262 676292 358264
rect 674097 358259 674163 358262
rect 62113 357778 62179 357781
rect 64646 357778 64706 357964
rect 675937 357914 676003 357917
rect 675937 357912 676292 357914
rect 675937 357856 675942 357912
rect 675998 357856 676292 357912
rect 675937 357854 676292 357856
rect 675937 357851 676003 357854
rect 62113 357776 64706 357778
rect 62113 357720 62118 357776
rect 62174 357720 64706 357776
rect 62113 357718 64706 357720
rect 62113 357715 62179 357718
rect 673177 357506 673243 357509
rect 673177 357504 676292 357506
rect 673177 357448 673182 357504
rect 673238 357448 676292 357504
rect 673177 357446 676292 357448
rect 673177 357443 673243 357446
rect 63217 357370 63283 357373
rect 63217 357368 64706 357370
rect 63217 357312 63222 357368
rect 63278 357312 64706 357368
rect 63217 357310 64706 357312
rect 63217 357307 63283 357310
rect 41454 356900 41460 356964
rect 41524 356962 41530 356964
rect 41781 356962 41847 356965
rect 41524 356960 41847 356962
rect 41524 356904 41786 356960
rect 41842 356904 41847 356960
rect 41524 356902 41847 356904
rect 41524 356900 41530 356902
rect 41781 356899 41847 356902
rect 64646 356782 64706 357310
rect 673177 357098 673243 357101
rect 673177 357096 676292 357098
rect 673177 357040 673182 357096
rect 673238 357040 676292 357096
rect 673177 357038 676292 357040
rect 673177 357035 673243 357038
rect 675937 356826 676003 356829
rect 669270 356824 676003 356826
rect 669270 356768 675942 356824
rect 675998 356768 676003 356824
rect 669270 356766 676003 356768
rect 652017 356690 652083 356693
rect 669270 356690 669330 356766
rect 675937 356763 676003 356766
rect 652017 356688 669330 356690
rect 652017 356632 652022 356688
rect 652078 356632 669330 356688
rect 652017 356630 669330 356632
rect 676170 356630 676292 356690
rect 652017 356627 652083 356630
rect 673913 356554 673979 356557
rect 676170 356554 676230 356630
rect 673913 356552 676230 356554
rect 673913 356496 673918 356552
rect 673974 356496 676230 356552
rect 673913 356494 676230 356496
rect 673913 356491 673979 356494
rect 672533 356282 672599 356285
rect 672533 356280 676292 356282
rect 672533 356224 672538 356280
rect 672594 356224 676292 356280
rect 672533 356222 676292 356224
rect 672533 356219 672599 356222
rect 42425 356010 42491 356013
rect 44633 356010 44699 356013
rect 42425 356008 44699 356010
rect 42425 355952 42430 356008
rect 42486 355952 44638 356008
rect 44694 355952 44699 356008
rect 42425 355950 44699 355952
rect 42425 355947 42491 355950
rect 44633 355947 44699 355950
rect 62113 356010 62179 356013
rect 62113 356008 64706 356010
rect 62113 355952 62118 356008
rect 62174 355952 64706 356008
rect 62113 355950 64706 355952
rect 62113 355947 62179 355950
rect 41873 355740 41939 355741
rect 41822 355738 41828 355740
rect 41782 355678 41828 355738
rect 41892 355736 41939 355740
rect 41934 355680 41939 355736
rect 41822 355676 41828 355678
rect 41892 355676 41939 355680
rect 41873 355675 41939 355676
rect 64646 355600 64706 355950
rect 673361 355874 673427 355877
rect 673361 355872 676292 355874
rect 673361 355816 673366 355872
rect 673422 355816 676292 355872
rect 673361 355814 676292 355816
rect 673361 355811 673427 355814
rect 672349 355466 672415 355469
rect 672349 355464 676292 355466
rect 672349 355408 672354 355464
rect 672410 355408 676292 355464
rect 672349 355406 676292 355408
rect 672349 355403 672415 355406
rect 672809 355058 672875 355061
rect 672809 355056 676292 355058
rect 672809 355000 672814 355056
rect 672870 355000 676292 355056
rect 672809 354998 676292 355000
rect 672809 354995 672875 354998
rect 43437 354786 43503 354789
rect 44449 354786 44515 354789
rect 43437 354784 44515 354786
rect 43437 354728 43442 354784
rect 43498 354728 44454 354784
rect 44510 354728 44515 354784
rect 43437 354726 44515 354728
rect 43437 354723 43503 354726
rect 44449 354723 44515 354726
rect 673913 354650 673979 354653
rect 673913 354648 676292 354650
rect 673913 354592 673918 354648
rect 673974 354592 676292 354648
rect 673913 354590 676292 354592
rect 673913 354587 673979 354590
rect 43294 354452 43300 354516
rect 43364 354514 43370 354516
rect 44633 354514 44699 354517
rect 43364 354512 44699 354514
rect 43364 354456 44638 354512
rect 44694 354456 44699 354512
rect 43364 354454 44699 354456
rect 43364 354452 43370 354454
rect 44633 354451 44699 354454
rect 62481 354514 62547 354517
rect 62481 354512 64706 354514
rect 62481 354456 62486 354512
rect 62542 354456 64706 354512
rect 62481 354454 64706 354456
rect 62481 354451 62547 354454
rect 64646 354418 64706 354454
rect 45461 354378 45527 354381
rect 51717 354378 51783 354381
rect 45461 354376 51783 354378
rect 45461 354320 45466 354376
rect 45522 354320 51722 354376
rect 51778 354320 51783 354376
rect 45461 354318 51783 354320
rect 45461 354315 45527 354318
rect 51717 354315 51783 354318
rect 675518 354180 675524 354244
rect 675588 354242 675594 354244
rect 675588 354182 676292 354242
rect 675588 354180 675594 354182
rect 43621 354106 43687 354109
rect 45461 354106 45527 354109
rect 43621 354104 45527 354106
rect 43621 354048 43626 354104
rect 43682 354048 45466 354104
rect 45522 354048 45527 354104
rect 43621 354046 45527 354048
rect 43621 354043 43687 354046
rect 45461 354043 45527 354046
rect 675886 353772 675892 353836
rect 675956 353834 675962 353836
rect 675956 353774 676292 353834
rect 675956 353772 675962 353774
rect 45461 353426 45527 353429
rect 64321 353426 64387 353429
rect 45461 353424 64387 353426
rect 45461 353368 45466 353424
rect 45522 353368 64326 353424
rect 64382 353368 64387 353424
rect 45461 353366 64387 353368
rect 45461 353363 45527 353366
rect 64321 353363 64387 353366
rect 672165 353426 672231 353429
rect 672165 353424 676292 353426
rect 672165 353368 672170 353424
rect 672226 353368 676292 353424
rect 672165 353366 676292 353368
rect 672165 353363 672231 353366
rect 44173 353154 44239 353157
rect 45415 353154 45481 353157
rect 44173 353152 45481 353154
rect 44173 353096 44178 353152
rect 44234 353096 45420 353152
rect 45476 353096 45481 353152
rect 44173 353094 45481 353096
rect 44173 353091 44239 353094
rect 45415 353091 45481 353094
rect 675702 352956 675708 353020
rect 675772 353018 675778 353020
rect 675772 352958 676292 353018
rect 675772 352956 675778 352958
rect 674465 352610 674531 352613
rect 674465 352608 676292 352610
rect 674465 352552 674470 352608
rect 674526 352552 676292 352608
rect 674465 352550 676292 352552
rect 674465 352547 674531 352550
rect 674649 352202 674715 352205
rect 674649 352200 676292 352202
rect 674649 352144 674654 352200
rect 674710 352144 676292 352200
rect 674649 352142 676292 352144
rect 674649 352139 674715 352142
rect 675886 351732 675892 351796
rect 675956 351794 675962 351796
rect 675956 351734 676292 351794
rect 675956 351732 675962 351734
rect 674281 351386 674347 351389
rect 674281 351384 676292 351386
rect 674281 351328 674286 351384
rect 674342 351328 676292 351384
rect 674281 351326 676292 351328
rect 674281 351323 674347 351326
rect 652385 351114 652451 351117
rect 674097 351114 674163 351117
rect 652385 351112 674163 351114
rect 652385 351056 652390 351112
rect 652446 351056 674102 351112
rect 674158 351056 674163 351112
rect 652385 351054 674163 351056
rect 652385 351051 652451 351054
rect 674097 351051 674163 351054
rect 676029 350978 676095 350981
rect 676029 350976 676292 350978
rect 676029 350920 676034 350976
rect 676090 350920 676292 350976
rect 676029 350918 676292 350920
rect 676029 350915 676095 350918
rect 673545 350570 673611 350573
rect 673545 350568 676292 350570
rect 673545 350512 673550 350568
rect 673606 350512 676292 350568
rect 673545 350510 676292 350512
rect 673545 350507 673611 350510
rect 673361 350162 673427 350165
rect 673361 350160 676292 350162
rect 673361 350104 673366 350160
rect 673422 350104 676292 350160
rect 673361 350102 676292 350104
rect 673361 350099 673427 350102
rect 672993 349754 673059 349757
rect 672993 349752 676292 349754
rect 672993 349696 672998 349752
rect 673054 349696 676292 349752
rect 672993 349694 676292 349696
rect 672993 349691 673059 349694
rect 673729 349346 673795 349349
rect 673729 349344 676292 349346
rect 673729 349288 673734 349344
rect 673790 349288 676292 349344
rect 673729 349286 676292 349288
rect 673729 349283 673795 349286
rect 671705 348938 671771 348941
rect 671705 348936 676292 348938
rect 671705 348880 671710 348936
rect 671766 348880 676292 348936
rect 671705 348878 676292 348880
rect 671705 348875 671771 348878
rect 672717 348530 672783 348533
rect 672717 348528 676292 348530
rect 672717 348472 672722 348528
rect 672778 348472 676292 348528
rect 672717 348470 676292 348472
rect 672717 348467 672783 348470
rect 675334 347652 675340 347716
rect 675404 347714 675410 347716
rect 683070 347714 683130 348092
rect 675404 347684 683130 347714
rect 675404 347654 683100 347684
rect 675404 347652 675410 347654
rect 669405 347306 669471 347309
rect 669405 347304 676292 347306
rect 669405 347248 669410 347304
rect 669466 347248 676292 347304
rect 669405 347246 676292 347248
rect 669405 347243 669471 347246
rect 676029 346626 676095 346629
rect 676438 346626 676444 346628
rect 676029 346624 676444 346626
rect 676029 346568 676034 346624
rect 676090 346568 676444 346624
rect 676029 346566 676444 346568
rect 676029 346563 676095 346566
rect 676438 346564 676444 346566
rect 676508 346564 676514 346628
rect 40217 345538 40283 345541
rect 43253 345538 43319 345541
rect 40217 345536 43319 345538
rect 40217 345480 40222 345536
rect 40278 345480 43258 345536
rect 43314 345480 43319 345536
rect 40217 345478 43319 345480
rect 40217 345475 40283 345478
rect 43253 345475 43319 345478
rect 35758 344317 35818 344556
rect 35525 344314 35591 344317
rect 35525 344312 35634 344314
rect 35525 344256 35530 344312
rect 35586 344256 35634 344312
rect 35525 344251 35634 344256
rect 35758 344312 35867 344317
rect 35758 344256 35806 344312
rect 35862 344256 35867 344312
rect 35758 344254 35867 344256
rect 35801 344251 35867 344254
rect 40033 344314 40099 344317
rect 42190 344314 42196 344316
rect 40033 344312 42196 344314
rect 40033 344256 40038 344312
rect 40094 344256 42196 344312
rect 40033 344254 42196 344256
rect 40033 344251 40099 344254
rect 42190 344252 42196 344254
rect 42260 344252 42266 344316
rect 35574 344148 35634 344251
rect 32998 343501 33058 343740
rect 32998 343496 33107 343501
rect 32998 343440 33046 343496
rect 33102 343440 33107 343496
rect 32998 343438 33107 343440
rect 33041 343435 33107 343438
rect 44909 343362 44975 343365
rect 41492 343360 44975 343362
rect 41492 343304 44914 343360
rect 44970 343304 44975 343360
rect 41492 343302 44975 343304
rect 44909 343299 44975 343302
rect 44214 342954 44220 342956
rect 41492 342894 44220 342954
rect 44214 342892 44220 342894
rect 44284 342892 44290 342956
rect 35758 342277 35818 342516
rect 44582 342410 44588 342412
rect 42014 342350 44588 342410
rect 35758 342272 35867 342277
rect 35758 342216 35806 342272
rect 35862 342216 35867 342272
rect 35758 342214 35867 342216
rect 35801 342211 35867 342214
rect 42014 342138 42074 342350
rect 44582 342348 44588 342350
rect 44652 342348 44658 342412
rect 41492 342078 42074 342138
rect 42190 342076 42196 342140
rect 42260 342138 42266 342140
rect 42260 342078 55230 342138
rect 42260 342076 42266 342078
rect 40033 341866 40099 341869
rect 40033 341864 50354 341866
rect 40033 341808 40038 341864
rect 40094 341808 50354 341864
rect 40033 341806 50354 341808
rect 40033 341803 40099 341806
rect 35574 341461 35634 341700
rect 35574 341456 35683 341461
rect 35574 341400 35622 341456
rect 35678 341400 35683 341456
rect 35574 341398 35683 341400
rect 35617 341395 35683 341398
rect 40217 341458 40283 341461
rect 45461 341458 45527 341461
rect 40217 341456 45527 341458
rect 40217 341400 40222 341456
rect 40278 341400 45466 341456
rect 45522 341400 45527 341456
rect 40217 341398 45527 341400
rect 50294 341458 50354 341806
rect 55170 341730 55230 342078
rect 62389 341730 62455 341733
rect 55170 341728 62455 341730
rect 55170 341672 62394 341728
rect 62450 341672 62455 341728
rect 55170 341670 62455 341672
rect 62389 341667 62455 341670
rect 63309 341458 63375 341461
rect 50294 341456 63375 341458
rect 50294 341400 63314 341456
rect 63370 341400 63375 341456
rect 50294 341398 63375 341400
rect 40217 341395 40283 341398
rect 45461 341395 45527 341398
rect 63309 341395 63375 341398
rect 39806 341053 39866 341292
rect 35801 341050 35867 341053
rect 35758 341048 35867 341050
rect 35758 340992 35806 341048
rect 35862 340992 35867 341048
rect 35758 340987 35867 340992
rect 39806 341048 39915 341053
rect 39806 340992 39854 341048
rect 39910 340992 39915 341048
rect 39806 340990 39915 340992
rect 39849 340987 39915 340990
rect 40217 341050 40283 341053
rect 45093 341050 45159 341053
rect 40217 341048 45159 341050
rect 40217 340992 40222 341048
rect 40278 340992 45098 341048
rect 45154 340992 45159 341048
rect 40217 340990 45159 340992
rect 40217 340987 40283 340990
rect 45093 340987 45159 340990
rect 35758 340884 35818 340987
rect 40033 340642 40099 340645
rect 45277 340642 45343 340645
rect 40033 340640 45343 340642
rect 40033 340584 40038 340640
rect 40094 340584 45282 340640
rect 45338 340584 45343 340640
rect 40033 340582 45343 340584
rect 40033 340579 40099 340582
rect 45277 340579 45343 340582
rect 41462 340234 41522 340476
rect 42742 340234 42748 340236
rect 41462 340174 42748 340234
rect 42742 340172 42748 340174
rect 42812 340172 42818 340236
rect 675753 340234 675819 340237
rect 676254 340234 676260 340236
rect 675753 340232 676260 340234
rect 675753 340176 675758 340232
rect 675814 340176 676260 340232
rect 675753 340174 676260 340176
rect 675753 340171 675819 340174
rect 676254 340172 676260 340174
rect 676324 340172 676330 340236
rect 35574 339829 35634 340068
rect 35525 339824 35634 339829
rect 35801 339826 35867 339829
rect 35525 339768 35530 339824
rect 35586 339768 35634 339824
rect 35525 339766 35634 339768
rect 35758 339824 35867 339826
rect 35758 339768 35806 339824
rect 35862 339768 35867 339824
rect 35525 339763 35591 339766
rect 35758 339763 35867 339768
rect 39849 339826 39915 339829
rect 44398 339826 44404 339828
rect 39849 339824 44404 339826
rect 39849 339768 39854 339824
rect 39910 339768 44404 339824
rect 39849 339766 44404 339768
rect 39849 339763 39915 339766
rect 44398 339764 44404 339766
rect 44468 339764 44474 339828
rect 35758 339660 35818 339763
rect 675477 339420 675543 339421
rect 675477 339416 675524 339420
rect 675588 339418 675594 339420
rect 675477 339360 675482 339416
rect 675477 339356 675524 339360
rect 675588 339358 675634 339418
rect 675588 339356 675594 339358
rect 675477 339355 675543 339356
rect 46933 339282 46999 339285
rect 41492 339280 46999 339282
rect 41492 339224 46938 339280
rect 46994 339224 46999 339280
rect 41492 339222 46999 339224
rect 46933 339219 46999 339222
rect 35206 338605 35266 338844
rect 653397 338738 653463 338741
rect 674925 338738 674991 338741
rect 653397 338736 674991 338738
rect 653397 338680 653402 338736
rect 653458 338680 674930 338736
rect 674986 338680 674991 338736
rect 653397 338678 674991 338680
rect 653397 338675 653463 338678
rect 674925 338675 674991 338678
rect 35157 338600 35266 338605
rect 35157 338544 35162 338600
rect 35218 338544 35266 338600
rect 35157 338542 35266 338544
rect 35157 338539 35223 338542
rect 45645 338466 45711 338469
rect 41492 338464 45711 338466
rect 41492 338408 45650 338464
rect 45706 338408 45711 338464
rect 41492 338406 45711 338408
rect 45645 338403 45711 338406
rect 47117 338058 47183 338061
rect 41492 338056 47183 338058
rect 41492 338000 47122 338056
rect 47178 338000 47183 338056
rect 41492 337998 47183 338000
rect 47117 337995 47183 337998
rect 672165 338058 672231 338061
rect 675109 338058 675175 338061
rect 672165 338056 675175 338058
rect 672165 338000 672170 338056
rect 672226 338000 675114 338056
rect 675170 338000 675175 338056
rect 672165 337998 675175 338000
rect 672165 337995 672231 337998
rect 675109 337995 675175 337998
rect 675753 337922 675819 337925
rect 676070 337922 676076 337924
rect 675753 337920 676076 337922
rect 675753 337864 675758 337920
rect 675814 337864 676076 337920
rect 675753 337862 676076 337864
rect 675753 337859 675819 337862
rect 676070 337860 676076 337862
rect 676140 337860 676146 337924
rect 674281 337786 674347 337789
rect 675109 337786 675175 337789
rect 674281 337784 675175 337786
rect 674281 337728 674286 337784
rect 674342 337728 675114 337784
rect 675170 337728 675175 337784
rect 674281 337726 675175 337728
rect 674281 337723 674347 337726
rect 675109 337723 675175 337726
rect 42926 337650 42932 337652
rect 41492 337590 42932 337650
rect 42926 337588 42932 337590
rect 42996 337588 43002 337652
rect 40542 336972 40602 337212
rect 40534 336908 40540 336972
rect 40604 336908 40610 336972
rect 45461 336834 45527 336837
rect 41492 336832 45527 336834
rect 41492 336776 45466 336832
rect 45522 336776 45527 336832
rect 41492 336774 45527 336776
rect 45461 336771 45527 336774
rect 38837 336562 38903 336565
rect 41822 336562 41828 336564
rect 38837 336560 41828 336562
rect 38837 336504 38842 336560
rect 38898 336504 41828 336560
rect 38837 336502 41828 336504
rect 38837 336499 38903 336502
rect 41822 336500 41828 336502
rect 41892 336500 41898 336564
rect 675753 336562 675819 336565
rect 676438 336562 676444 336564
rect 675753 336560 676444 336562
rect 675753 336504 675758 336560
rect 675814 336504 676444 336560
rect 675753 336502 676444 336504
rect 675753 336499 675819 336502
rect 676438 336500 676444 336502
rect 676508 336500 676514 336564
rect 35758 336157 35818 336396
rect 35758 336152 35867 336157
rect 35758 336096 35806 336152
rect 35862 336096 35867 336152
rect 35758 336094 35867 336096
rect 35801 336091 35867 336094
rect 40910 335748 40970 335988
rect 673361 335882 673427 335885
rect 674925 335882 674991 335885
rect 673361 335880 674991 335882
rect 673361 335824 673366 335880
rect 673422 335824 674930 335880
rect 674986 335824 674991 335880
rect 673361 335822 674991 335824
rect 673361 335819 673427 335822
rect 674925 335819 674991 335822
rect 40902 335684 40908 335748
rect 40972 335684 40978 335748
rect 672993 335610 673059 335613
rect 675109 335610 675175 335613
rect 672993 335608 675175 335610
rect 40726 335340 40786 335580
rect 672993 335552 672998 335608
rect 673054 335552 675114 335608
rect 675170 335552 675175 335608
rect 672993 335550 675175 335552
rect 672993 335547 673059 335550
rect 675109 335547 675175 335550
rect 40718 335276 40724 335340
rect 40788 335276 40794 335340
rect 35574 334933 35634 335172
rect 35574 334928 35683 334933
rect 35574 334872 35622 334928
rect 35678 334872 35683 334928
rect 35574 334870 35683 334872
rect 35617 334867 35683 334870
rect 35758 334525 35818 334764
rect 43294 334596 43300 334660
rect 43364 334658 43370 334660
rect 43989 334658 44055 334661
rect 43364 334656 44055 334658
rect 43364 334600 43994 334656
rect 44050 334600 44055 334656
rect 43364 334598 44055 334600
rect 43364 334596 43370 334598
rect 43989 334595 44055 334598
rect 35758 334520 35867 334525
rect 35758 334464 35806 334520
rect 35862 334464 35867 334520
rect 35758 334462 35867 334464
rect 35801 334459 35867 334462
rect 40217 334522 40283 334525
rect 43161 334522 43227 334525
rect 40217 334520 43227 334522
rect 40217 334464 40222 334520
rect 40278 334464 43166 334520
rect 43222 334464 43227 334520
rect 40217 334462 43227 334464
rect 40217 334459 40283 334462
rect 43161 334459 43227 334462
rect 41462 334114 41522 334356
rect 44817 334114 44883 334117
rect 41462 334112 44883 334114
rect 41462 334056 44822 334112
rect 44878 334056 44883 334112
rect 41462 334054 44883 334056
rect 44817 334051 44883 334054
rect 41462 333298 41522 333948
rect 41462 333238 51090 333298
rect 36537 332890 36603 332893
rect 41454 332890 41460 332892
rect 36537 332888 41460 332890
rect 36537 332832 36542 332888
rect 36598 332832 41460 332888
rect 36537 332830 41460 332832
rect 36537 332827 36603 332830
rect 41454 332828 41460 332830
rect 41524 332828 41530 332892
rect 51030 332618 51090 333238
rect 673729 332754 673795 332757
rect 675109 332754 675175 332757
rect 673729 332752 675175 332754
rect 673729 332696 673734 332752
rect 673790 332696 675114 332752
rect 675170 332696 675175 332752
rect 673729 332694 675175 332696
rect 673729 332691 673795 332694
rect 675109 332691 675175 332694
rect 62481 332618 62547 332621
rect 51030 332616 62547 332618
rect 51030 332560 62486 332616
rect 62542 332560 62547 332616
rect 51030 332558 62547 332560
rect 62481 332555 62547 332558
rect 39389 332482 39455 332485
rect 42793 332482 42859 332485
rect 39389 332480 42859 332482
rect 39389 332424 39394 332480
rect 39450 332424 42798 332480
rect 42854 332424 42859 332480
rect 39389 332422 42859 332424
rect 39389 332419 39455 332422
rect 42793 332419 42859 332422
rect 35157 331802 35223 331805
rect 41638 331802 41644 331804
rect 35157 331800 41644 331802
rect 35157 331744 35162 331800
rect 35218 331744 41644 331800
rect 35157 331742 41644 331744
rect 35157 331739 35223 331742
rect 41638 331740 41644 331742
rect 41708 331740 41714 331804
rect 673545 331122 673611 331125
rect 675293 331122 675359 331125
rect 673545 331120 675359 331122
rect 673545 331064 673550 331120
rect 673606 331064 675298 331120
rect 675354 331064 675359 331120
rect 673545 331062 675359 331064
rect 673545 331059 673611 331062
rect 675293 331059 675359 331062
rect 652385 329762 652451 329765
rect 649950 329760 652451 329762
rect 649950 329704 652390 329760
rect 652446 329704 652451 329760
rect 649950 329702 652451 329704
rect 649950 329234 650010 329702
rect 652385 329699 652451 329702
rect 671705 329762 671771 329765
rect 675109 329762 675175 329765
rect 671705 329760 675175 329762
rect 671705 329704 671710 329760
rect 671766 329704 675114 329760
rect 675170 329704 675175 329760
rect 671705 329702 675175 329704
rect 671705 329699 671771 329702
rect 675109 329699 675175 329702
rect 651373 328130 651439 328133
rect 649950 328128 651439 328130
rect 649950 328072 651378 328128
rect 651434 328072 651439 328128
rect 649950 328070 651439 328072
rect 649950 328052 650010 328070
rect 651373 328067 651439 328070
rect 675017 327994 675083 327997
rect 675385 327996 675451 327997
rect 675334 327994 675340 327996
rect 675017 327992 675340 327994
rect 675404 327994 675451 327996
rect 675404 327992 675496 327994
rect 675017 327936 675022 327992
rect 675078 327936 675340 327992
rect 675446 327936 675496 327992
rect 675017 327934 675340 327936
rect 675017 327931 675083 327934
rect 675334 327932 675340 327934
rect 675404 327934 675496 327936
rect 675404 327932 675451 327934
rect 675385 327931 675451 327932
rect 652017 326906 652083 326909
rect 650502 326904 652083 326906
rect 650502 326900 652022 326904
rect 649980 326848 652022 326900
rect 652078 326848 652083 326904
rect 649980 326846 652083 326848
rect 649980 326840 650562 326846
rect 652017 326843 652083 326846
rect 674649 326906 674715 326909
rect 675385 326906 675451 326909
rect 674649 326904 675451 326906
rect 674649 326848 674654 326904
rect 674710 326848 675390 326904
rect 675446 326848 675451 326904
rect 674649 326846 675451 326848
rect 674649 326843 674715 326846
rect 675385 326843 675451 326846
rect 649950 325682 650010 325710
rect 651373 325682 651439 325685
rect 649950 325680 651439 325682
rect 649950 325624 651378 325680
rect 651434 325624 651439 325680
rect 649950 325622 651439 325624
rect 651373 325619 651439 325622
rect 675201 325682 675267 325685
rect 676622 325682 676628 325684
rect 675201 325680 676628 325682
rect 675201 325624 675206 325680
rect 675262 325624 676628 325680
rect 675201 325622 676628 325624
rect 675201 325619 675267 325622
rect 676622 325620 676628 325622
rect 676692 325620 676698 325684
rect 672901 325002 672967 325005
rect 675017 325002 675083 325005
rect 672901 325000 675083 325002
rect 672901 324944 672906 325000
rect 672962 324944 675022 325000
rect 675078 324944 675083 325000
rect 672901 324942 675083 324944
rect 672901 324939 672967 324942
rect 675017 324939 675083 324942
rect 41781 324868 41847 324869
rect 41781 324864 41828 324868
rect 41892 324866 41898 324868
rect 41781 324808 41786 324864
rect 41781 324804 41828 324808
rect 41892 324806 41938 324866
rect 41892 324804 41898 324806
rect 41781 324803 41847 324804
rect 42241 324322 42307 324325
rect 47117 324322 47183 324325
rect 42241 324320 47183 324322
rect 42241 324264 42246 324320
rect 42302 324264 47122 324320
rect 47178 324264 47183 324320
rect 42241 324262 47183 324264
rect 42241 324259 42307 324262
rect 47117 324259 47183 324262
rect 40902 321132 40908 321196
rect 40972 321194 40978 321196
rect 41781 321194 41847 321197
rect 40972 321192 41847 321194
rect 40972 321136 41786 321192
rect 41842 321136 41847 321192
rect 40972 321134 41847 321136
rect 40972 321132 40978 321134
rect 41781 321131 41847 321134
rect 42057 321194 42123 321197
rect 42977 321194 43043 321197
rect 42057 321192 43043 321194
rect 42057 321136 42062 321192
rect 42118 321136 42982 321192
rect 43038 321136 43043 321192
rect 42057 321134 43043 321136
rect 42057 321131 42123 321134
rect 42977 321131 43043 321134
rect 42425 320786 42491 320789
rect 62021 320786 62087 320789
rect 42425 320784 62087 320786
rect 42425 320728 42430 320784
rect 42486 320728 62026 320784
rect 62082 320728 62087 320784
rect 42425 320726 62087 320728
rect 42425 320723 42491 320726
rect 62021 320723 62087 320726
rect 42609 319426 42675 319429
rect 60365 319426 60431 319429
rect 42609 319424 60431 319426
rect 42609 319368 42614 319424
rect 42670 319368 60370 319424
rect 60426 319368 60431 319424
rect 42609 319366 60431 319368
rect 42609 319363 42675 319366
rect 60365 319363 60431 319366
rect 42425 319154 42491 319157
rect 45645 319154 45711 319157
rect 42425 319152 45711 319154
rect 42425 319096 42430 319152
rect 42486 319096 45650 319152
rect 45706 319096 45711 319152
rect 42425 319094 45711 319096
rect 42425 319091 42491 319094
rect 45645 319091 45711 319094
rect 40718 317324 40724 317388
rect 40788 317386 40794 317388
rect 41781 317386 41847 317389
rect 40788 317384 41847 317386
rect 40788 317328 41786 317384
rect 41842 317328 41847 317384
rect 40788 317326 41847 317328
rect 40788 317324 40794 317326
rect 41781 317323 41847 317326
rect 62021 317386 62087 317389
rect 62021 317384 64706 317386
rect 62021 317328 62026 317384
rect 62082 317328 64706 317384
rect 62021 317326 64706 317328
rect 62021 317323 62087 317326
rect 64646 317106 64706 317326
rect 40534 315964 40540 316028
rect 40604 316026 40610 316028
rect 41781 316026 41847 316029
rect 40604 316024 41847 316026
rect 40604 315968 41786 316024
rect 41842 315968 41847 316024
rect 40604 315966 41847 315968
rect 40604 315964 40610 315966
rect 41781 315963 41847 315966
rect 62113 316026 62179 316029
rect 62113 316024 64706 316026
rect 62113 315968 62118 316024
rect 62174 315968 64706 316024
rect 62113 315966 64706 315968
rect 62113 315963 62179 315966
rect 64646 315924 64706 315966
rect 41781 315620 41847 315621
rect 41781 315616 41828 315620
rect 41892 315618 41898 315620
rect 41781 315560 41786 315616
rect 41781 315556 41828 315560
rect 41892 315558 41938 315618
rect 41892 315556 41898 315558
rect 41781 315555 41847 315556
rect 62113 314802 62179 314805
rect 62113 314800 64706 314802
rect 62113 314744 62118 314800
rect 62174 314744 64706 314800
rect 62113 314742 64706 314744
rect 62113 314739 62179 314742
rect 42425 314666 42491 314669
rect 45461 314666 45527 314669
rect 42425 314664 45527 314666
rect 42425 314608 42430 314664
rect 42486 314608 45466 314664
rect 45522 314608 45527 314664
rect 42425 314606 45527 314608
rect 42425 314603 42491 314606
rect 45461 314603 45527 314606
rect 62297 314122 62363 314125
rect 62297 314120 64706 314122
rect 62297 314064 62302 314120
rect 62358 314064 64706 314120
rect 62297 314062 64706 314064
rect 62297 314059 62363 314062
rect 41454 313652 41460 313716
rect 41524 313714 41530 313716
rect 41781 313714 41847 313717
rect 41524 313712 41847 313714
rect 41524 313656 41786 313712
rect 41842 313656 41847 313712
rect 41524 313654 41847 313656
rect 41524 313652 41530 313654
rect 41781 313651 41847 313654
rect 64646 313560 64706 314062
rect 676213 313986 676279 313989
rect 676213 313984 676322 313986
rect 676213 313928 676218 313984
rect 676274 313928 676322 313984
rect 676213 313923 676322 313928
rect 676262 313684 676322 313923
rect 653397 313306 653463 313309
rect 653397 313304 676292 313306
rect 653397 313248 653402 313304
rect 653458 313248 676292 313304
rect 653397 313246 676292 313248
rect 653397 313243 653463 313246
rect 62389 313034 62455 313037
rect 674649 313034 674715 313037
rect 62389 313032 64706 313034
rect 62389 312976 62394 313032
rect 62450 312976 64706 313032
rect 62389 312974 64706 312976
rect 62389 312971 62455 312974
rect 42425 312762 42491 312765
rect 42926 312762 42932 312764
rect 42425 312760 42932 312762
rect 42425 312704 42430 312760
rect 42486 312704 42932 312760
rect 42425 312702 42932 312704
rect 42425 312699 42491 312702
rect 42926 312700 42932 312702
rect 42996 312700 43002 312764
rect 64646 312378 64706 312974
rect 674649 313032 675034 313034
rect 674649 312976 674654 313032
rect 674710 312976 675034 313032
rect 674649 312974 675034 312976
rect 674649 312971 674715 312974
rect 674974 312898 675034 312974
rect 674974 312838 676292 312898
rect 673361 312762 673427 312765
rect 674833 312762 674899 312765
rect 673361 312760 674899 312762
rect 673361 312704 673366 312760
rect 673422 312704 674838 312760
rect 674894 312704 674899 312760
rect 673361 312702 674899 312704
rect 673361 312699 673427 312702
rect 674833 312699 674899 312702
rect 673177 312490 673243 312493
rect 673177 312488 676292 312490
rect 673177 312432 673182 312488
rect 673238 312432 676292 312488
rect 673177 312430 676292 312432
rect 673177 312427 673243 312430
rect 674833 312082 674899 312085
rect 674833 312080 676292 312082
rect 674833 312024 674838 312080
rect 674894 312024 676292 312080
rect 674833 312022 676292 312024
rect 674833 312019 674899 312022
rect 660297 311946 660363 311949
rect 674649 311946 674715 311949
rect 660297 311944 674715 311946
rect 660297 311888 660302 311944
rect 660358 311888 674654 311944
rect 674710 311888 674715 311944
rect 660297 311886 674715 311888
rect 660297 311883 660363 311886
rect 674649 311883 674715 311886
rect 63309 311810 63375 311813
rect 63309 311808 64706 311810
rect 63309 311752 63314 311808
rect 63370 311752 64706 311808
rect 63309 311750 64706 311752
rect 63309 311747 63375 311750
rect 64646 311196 64706 311750
rect 672533 311674 672599 311677
rect 672533 311672 676292 311674
rect 672533 311616 672538 311672
rect 672594 311616 676292 311672
rect 672533 311614 676292 311616
rect 672533 311611 672599 311614
rect 673177 311266 673243 311269
rect 673177 311264 676292 311266
rect 673177 311208 673182 311264
rect 673238 311208 676292 311264
rect 673177 311206 676292 311208
rect 673177 311203 673243 311206
rect 672349 310858 672415 310861
rect 672349 310856 676292 310858
rect 672349 310800 672354 310856
rect 672410 310800 676292 310856
rect 672349 310798 676292 310800
rect 672349 310795 672415 310798
rect 42057 310450 42123 310453
rect 51073 310450 51139 310453
rect 42057 310448 51139 310450
rect 42057 310392 42062 310448
rect 42118 310392 51078 310448
rect 51134 310392 51139 310448
rect 42057 310390 51139 310392
rect 42057 310387 42123 310390
rect 51073 310387 51139 310390
rect 674189 310450 674255 310453
rect 674189 310448 676292 310450
rect 674189 310392 674194 310448
rect 674250 310392 676292 310448
rect 674189 310390 676292 310392
rect 674189 310387 674255 310390
rect 42425 310178 42491 310181
rect 46933 310178 46999 310181
rect 42425 310176 46999 310178
rect 42425 310120 42430 310176
rect 42486 310120 46938 310176
rect 46994 310120 46999 310176
rect 42425 310118 46999 310120
rect 42425 310115 42491 310118
rect 46933 310115 46999 310118
rect 674373 310042 674439 310045
rect 674373 310040 676292 310042
rect 674373 309984 674378 310040
rect 674434 309984 676292 310040
rect 674373 309982 676292 309984
rect 674373 309979 674439 309982
rect 652293 309906 652359 309909
rect 652293 309904 663810 309906
rect 652293 309848 652298 309904
rect 652354 309848 663810 309904
rect 652293 309846 663810 309848
rect 652293 309843 652359 309846
rect 663750 309362 663810 309846
rect 674649 309634 674715 309637
rect 674649 309632 676292 309634
rect 674649 309576 674654 309632
rect 674710 309576 676292 309632
rect 674649 309574 676292 309576
rect 674649 309571 674715 309574
rect 675845 309362 675911 309365
rect 663750 309360 675911 309362
rect 663750 309304 675850 309360
rect 675906 309304 675911 309360
rect 663750 309302 675911 309304
rect 675845 309299 675911 309302
rect 676032 309166 676292 309226
rect 675845 309090 675911 309093
rect 676032 309090 676092 309166
rect 675845 309088 676092 309090
rect 675845 309032 675850 309088
rect 675906 309032 676092 309088
rect 675845 309030 676092 309032
rect 675845 309027 675911 309030
rect 675886 308756 675892 308820
rect 675956 308818 675962 308820
rect 675956 308758 676292 308818
rect 675956 308756 675962 308758
rect 676029 308410 676095 308413
rect 676029 308408 676292 308410
rect 676029 308352 676034 308408
rect 676090 308352 676292 308408
rect 676029 308350 676292 308352
rect 676029 308347 676095 308350
rect 675017 308002 675083 308005
rect 675017 308000 676292 308002
rect 675017 307944 675022 308000
rect 675078 307944 676292 308000
rect 675017 307942 676292 307944
rect 675017 307939 675083 307942
rect 675385 307594 675451 307597
rect 675385 307592 676292 307594
rect 675385 307536 675390 307592
rect 675446 307536 676292 307592
rect 675385 307534 676292 307536
rect 675385 307531 675451 307534
rect 676029 307186 676095 307189
rect 676029 307184 676292 307186
rect 676029 307128 676034 307184
rect 676090 307128 676292 307184
rect 676029 307126 676292 307128
rect 676029 307123 676095 307126
rect 679617 306778 679683 306781
rect 679604 306776 679683 306778
rect 679604 306720 679622 306776
rect 679678 306720 679683 306776
rect 679604 306718 679683 306720
rect 679617 306715 679683 306718
rect 675845 306642 675911 306645
rect 676070 306642 676076 306644
rect 675845 306640 676076 306642
rect 675845 306584 675850 306640
rect 675906 306584 676076 306640
rect 675845 306582 676076 306584
rect 675845 306579 675911 306582
rect 676070 306580 676076 306582
rect 676140 306580 676146 306644
rect 674833 306370 674899 306373
rect 674833 306368 676292 306370
rect 674833 306312 674838 306368
rect 674894 306312 676292 306368
rect 674833 306310 676292 306312
rect 674833 306307 674899 306310
rect 676029 305962 676095 305965
rect 676029 305960 676292 305962
rect 676029 305904 676034 305960
rect 676090 305904 676292 305960
rect 676029 305902 676292 305904
rect 676029 305899 676095 305902
rect 674465 305554 674531 305557
rect 674465 305552 676292 305554
rect 674465 305496 674470 305552
rect 674526 305496 676292 305552
rect 674465 305494 676292 305496
rect 674465 305491 674531 305494
rect 673913 305146 673979 305149
rect 673913 305144 676292 305146
rect 673913 305088 673918 305144
rect 673974 305088 676292 305144
rect 673913 305086 676292 305088
rect 673913 305083 673979 305086
rect 676254 304914 676260 304978
rect 676324 304976 676330 304978
rect 676324 304916 676506 304976
rect 676324 304914 676330 304916
rect 676446 304708 676506 304916
rect 673085 304330 673151 304333
rect 673085 304328 676292 304330
rect 673085 304272 673090 304328
rect 673146 304272 676292 304328
rect 673085 304270 676292 304272
rect 673085 304267 673151 304270
rect 673729 303922 673795 303925
rect 673729 303920 676292 303922
rect 673729 303864 673734 303920
rect 673790 303864 676292 303920
rect 673729 303862 676292 303864
rect 673729 303859 673795 303862
rect 676029 303514 676095 303517
rect 676029 303512 676292 303514
rect 676029 303456 676034 303512
rect 676090 303456 676292 303512
rect 676029 303454 676292 303456
rect 676029 303451 676095 303454
rect 651373 303378 651439 303381
rect 649950 303376 651439 303378
rect 649950 303320 651378 303376
rect 651434 303320 651439 303376
rect 649950 303318 651439 303320
rect 649950 302776 650010 303318
rect 651373 303315 651439 303318
rect 675201 302970 675267 302973
rect 675845 302970 675911 302973
rect 675201 302968 675911 302970
rect 675201 302912 675206 302968
rect 675262 302912 675850 302968
rect 675906 302912 675911 302968
rect 675201 302910 675911 302912
rect 675201 302907 675267 302910
rect 675845 302907 675911 302910
rect 675886 302636 675892 302700
rect 675956 302698 675962 302700
rect 676262 302698 676322 303076
rect 675956 302668 676322 302698
rect 675956 302638 676292 302668
rect 675956 302636 675962 302638
rect 671521 302290 671587 302293
rect 671521 302288 676292 302290
rect 671521 302232 671526 302288
rect 671582 302232 676292 302288
rect 671521 302230 676292 302232
rect 671521 302227 671587 302230
rect 652293 302154 652359 302157
rect 649950 302152 652359 302154
rect 649950 302096 652298 302152
rect 652354 302096 652359 302152
rect 649950 302094 652359 302096
rect 649950 301594 650010 302094
rect 652293 302091 652359 302094
rect 669957 302018 670023 302021
rect 676029 302018 676095 302021
rect 669957 302016 676095 302018
rect 669957 301960 669962 302016
rect 670018 301960 676034 302016
rect 676090 301960 676095 302016
rect 669957 301958 676095 301960
rect 669957 301955 670023 301958
rect 676029 301955 676095 301958
rect 676213 301610 676279 301613
rect 676438 301610 676444 301612
rect 676213 301608 676444 301610
rect 676213 301552 676218 301608
rect 676274 301552 676444 301608
rect 676213 301550 676444 301552
rect 676213 301547 676279 301550
rect 676438 301548 676444 301550
rect 676508 301548 676514 301612
rect 53281 301338 53347 301341
rect 41492 301336 53347 301338
rect 41492 301280 53286 301336
rect 53342 301280 53347 301336
rect 41492 301278 53347 301280
rect 53281 301275 53347 301278
rect 41492 300870 41844 300930
rect 41784 300794 41844 300870
rect 41784 300734 51090 300794
rect 41137 300522 41203 300525
rect 41124 300520 41203 300522
rect 41124 300464 41142 300520
rect 41198 300464 41203 300520
rect 41124 300462 41203 300464
rect 41137 300459 41203 300462
rect 44214 300114 44220 300116
rect 41492 300054 44220 300114
rect 44214 300052 44220 300054
rect 44284 300052 44290 300116
rect 42885 299706 42951 299709
rect 41492 299704 42951 299706
rect 41492 299648 42890 299704
rect 42946 299648 42951 299704
rect 41492 299646 42951 299648
rect 42885 299643 42951 299646
rect 51030 299570 51090 300734
rect 651465 300658 651531 300661
rect 649950 300656 651531 300658
rect 649950 300600 651470 300656
rect 651526 300600 651531 300656
rect 649950 300598 651531 300600
rect 649950 300412 650010 300598
rect 651465 300595 651531 300598
rect 63309 299570 63375 299573
rect 51030 299568 63375 299570
rect 51030 299512 63314 299568
rect 63370 299512 63375 299568
rect 51030 299510 63375 299512
rect 63309 299507 63375 299510
rect 44582 299298 44588 299300
rect 41492 299238 44588 299298
rect 44582 299236 44588 299238
rect 44652 299236 44658 299300
rect 45001 298890 45067 298893
rect 41492 298888 45067 298890
rect 41492 298832 45006 298888
rect 45062 298832 45067 298888
rect 41492 298830 45067 298832
rect 45001 298827 45067 298830
rect 649950 298618 650010 299230
rect 652569 298618 652635 298621
rect 649950 298616 652635 298618
rect 649950 298560 652574 298616
rect 652630 298560 652635 298616
rect 649950 298558 652635 298560
rect 652569 298555 652635 298558
rect 44398 298482 44404 298484
rect 41492 298422 44404 298482
rect 44398 298420 44404 298422
rect 44468 298420 44474 298484
rect 44265 298074 44331 298077
rect 41492 298072 44331 298074
rect 41492 298016 44270 298072
rect 44326 298016 44331 298072
rect 41492 298014 44331 298016
rect 44265 298011 44331 298014
rect 42742 297666 42748 297668
rect 41492 297606 42748 297666
rect 42742 297604 42748 297606
rect 42812 297604 42818 297668
rect 649950 297530 650010 298048
rect 652109 297530 652175 297533
rect 649950 297528 652175 297530
rect 649950 297472 652114 297528
rect 652170 297472 652175 297528
rect 649950 297470 652175 297472
rect 652109 297467 652175 297470
rect 41965 297394 42031 297397
rect 62389 297394 62455 297397
rect 41965 297392 62455 297394
rect 41965 297336 41970 297392
rect 42026 297336 62394 297392
rect 62450 297336 62455 297392
rect 41965 297334 62455 297336
rect 41965 297331 42031 297334
rect 62389 297331 62455 297334
rect 675702 297332 675708 297396
rect 675772 297394 675778 297396
rect 676857 297394 676923 297397
rect 675772 297392 676923 297394
rect 675772 297336 676862 297392
rect 676918 297336 676923 297392
rect 675772 297334 676923 297336
rect 675772 297332 675778 297334
rect 676857 297331 676923 297334
rect 41492 297198 41844 297258
rect 41784 297122 41844 297198
rect 44541 297122 44607 297125
rect 41784 297120 44607 297122
rect 41784 297064 44546 297120
rect 44602 297064 44607 297120
rect 41784 297062 44607 297064
rect 44541 297059 44607 297062
rect 42190 296850 42196 296852
rect 41492 296790 42196 296850
rect 42190 296788 42196 296790
rect 42260 296788 42266 296852
rect 649950 296850 650010 296866
rect 651925 296850 651991 296853
rect 649950 296848 651991 296850
rect 649950 296792 651930 296848
rect 651986 296792 651991 296848
rect 649950 296790 651991 296792
rect 651925 296787 651991 296790
rect 675150 296652 675156 296716
rect 675220 296714 675226 296716
rect 675477 296714 675543 296717
rect 675220 296712 675543 296714
rect 675220 296656 675482 296712
rect 675538 296656 675543 296712
rect 675220 296654 675543 296656
rect 675220 296652 675226 296654
rect 675477 296651 675543 296654
rect 41321 296442 41387 296445
rect 41308 296440 41387 296442
rect 41308 296384 41326 296440
rect 41382 296384 41387 296440
rect 41308 296382 41387 296384
rect 41321 296379 41387 296382
rect 670969 296306 671035 296309
rect 675661 296306 675727 296309
rect 670969 296304 675727 296306
rect 670969 296248 670974 296304
rect 671030 296248 675666 296304
rect 675722 296248 675727 296304
rect 670969 296246 675727 296248
rect 670969 296243 671035 296246
rect 675661 296243 675727 296246
rect 40953 296034 41019 296037
rect 40940 296032 41019 296034
rect 40940 295976 40958 296032
rect 41014 295976 41019 296032
rect 40940 295974 41019 295976
rect 40953 295971 41019 295974
rect 675293 295898 675359 295901
rect 675661 295898 675727 295901
rect 675293 295896 675727 295898
rect 675293 295840 675298 295896
rect 675354 295840 675666 295896
rect 675722 295840 675727 295896
rect 675293 295838 675727 295840
rect 675293 295835 675359 295838
rect 675661 295835 675727 295838
rect 62113 295762 62179 295765
rect 62113 295760 64706 295762
rect 62113 295704 62118 295760
rect 62174 295704 64706 295760
rect 62113 295702 64706 295704
rect 62113 295699 62179 295702
rect 64646 295684 64706 295702
rect 39297 295626 39363 295629
rect 39284 295624 39363 295626
rect 39284 295568 39302 295624
rect 39358 295568 39363 295624
rect 39284 295566 39363 295568
rect 39297 295563 39363 295566
rect 649950 295354 650010 295684
rect 651649 295354 651715 295357
rect 649950 295352 651715 295354
rect 649950 295296 651654 295352
rect 651710 295296 651715 295352
rect 649950 295294 651715 295296
rect 651649 295291 651715 295294
rect 41137 295218 41203 295221
rect 41124 295216 41203 295218
rect 41124 295160 41142 295216
rect 41198 295160 41203 295216
rect 41124 295158 41203 295160
rect 41137 295155 41203 295158
rect 33777 294810 33843 294813
rect 33764 294808 33843 294810
rect 33764 294752 33782 294808
rect 33838 294752 33843 294808
rect 33764 294750 33843 294752
rect 33777 294747 33843 294750
rect 674833 294538 674899 294541
rect 675150 294538 675156 294540
rect 674833 294536 675156 294538
rect 37917 294402 37983 294405
rect 37917 294400 37996 294402
rect 37917 294344 37922 294400
rect 37978 294344 37996 294400
rect 37917 294342 37996 294344
rect 37917 294339 37983 294342
rect 62113 294130 62179 294133
rect 64646 294130 64706 294502
rect 649950 294266 650010 294502
rect 674833 294480 674838 294536
rect 674894 294480 675156 294536
rect 674833 294478 675156 294480
rect 674833 294475 674899 294478
rect 675150 294476 675156 294478
rect 675220 294476 675226 294540
rect 675753 294538 675819 294541
rect 676622 294538 676628 294540
rect 675753 294536 676628 294538
rect 675753 294480 675758 294536
rect 675814 294480 676628 294536
rect 675753 294478 676628 294480
rect 675753 294475 675819 294478
rect 676622 294476 676628 294478
rect 676692 294476 676698 294540
rect 651465 294266 651531 294269
rect 649950 294264 651531 294266
rect 649950 294208 651470 294264
rect 651526 294208 651531 294264
rect 649950 294206 651531 294208
rect 651465 294203 651531 294206
rect 62113 294128 64706 294130
rect 62113 294072 62118 294128
rect 62174 294072 64706 294128
rect 62113 294070 64706 294072
rect 62113 294067 62179 294070
rect 43161 293994 43227 293997
rect 41492 293992 43227 293994
rect 41492 293936 43166 293992
rect 43222 293936 43227 293992
rect 41492 293934 43227 293936
rect 43161 293931 43227 293934
rect 652845 293858 652911 293861
rect 670969 293858 671035 293861
rect 652845 293856 671035 293858
rect 652845 293800 652850 293856
rect 652906 293800 670974 293856
rect 671030 293800 671035 293856
rect 652845 293798 671035 293800
rect 652845 293795 652911 293798
rect 670969 293795 671035 293798
rect 45185 293586 45251 293589
rect 41492 293584 45251 293586
rect 41492 293528 45190 293584
rect 45246 293528 45251 293584
rect 41492 293526 45251 293528
rect 45185 293523 45251 293526
rect 43437 293178 43503 293181
rect 41492 293176 43503 293178
rect 41492 293120 43442 293176
rect 43498 293120 43503 293176
rect 41492 293118 43503 293120
rect 43437 293115 43503 293118
rect 42701 292770 42767 292773
rect 41492 292768 42767 292770
rect 41492 292712 42706 292768
rect 42762 292712 42767 292768
rect 41492 292710 42767 292712
rect 42701 292707 42767 292710
rect 62113 292770 62179 292773
rect 64646 292770 64706 293320
rect 62113 292768 64706 292770
rect 62113 292712 62118 292768
rect 62174 292712 64706 292768
rect 62113 292710 64706 292712
rect 649950 292770 650010 293320
rect 652385 292770 652451 292773
rect 649950 292768 652451 292770
rect 649950 292712 652390 292768
rect 652446 292712 652451 292768
rect 649950 292710 652451 292712
rect 62113 292707 62179 292710
rect 652385 292707 652451 292710
rect 40534 292528 40540 292592
rect 40604 292528 40610 292592
rect 40542 292332 40602 292528
rect 62389 292498 62455 292501
rect 62389 292496 64706 292498
rect 62389 292440 62394 292496
rect 62450 292440 64706 292496
rect 62389 292438 64706 292440
rect 62389 292435 62455 292438
rect 41781 292226 41847 292229
rect 42006 292226 42012 292228
rect 41781 292224 42012 292226
rect 41781 292168 41786 292224
rect 41842 292168 42012 292224
rect 41781 292166 42012 292168
rect 41781 292163 41847 292166
rect 42006 292164 42012 292166
rect 42076 292164 42082 292228
rect 64646 292138 64706 292438
rect 41822 291954 41828 291956
rect 41492 291894 41828 291954
rect 41822 291892 41828 291894
rect 41892 291892 41898 291956
rect 649950 291682 650010 292138
rect 651465 291682 651531 291685
rect 649950 291680 651531 291682
rect 649950 291624 651470 291680
rect 651526 291624 651531 291680
rect 649950 291622 651531 291624
rect 651465 291619 651531 291622
rect 41229 291546 41295 291549
rect 675753 291546 675819 291549
rect 676438 291546 676444 291548
rect 41229 291544 41308 291546
rect 41229 291488 41234 291544
rect 41290 291488 41308 291544
rect 41229 291486 41308 291488
rect 675753 291544 676444 291546
rect 675753 291488 675758 291544
rect 675814 291488 676444 291544
rect 675753 291486 676444 291488
rect 41229 291483 41295 291486
rect 675753 291483 675819 291486
rect 676438 291484 676444 291486
rect 676508 291484 676514 291548
rect 41965 291274 42031 291277
rect 43621 291274 43687 291277
rect 41965 291272 43687 291274
rect 41965 291216 41970 291272
rect 42026 291216 43626 291272
rect 43682 291216 43687 291272
rect 41965 291214 43687 291216
rect 41965 291211 42031 291214
rect 43621 291211 43687 291214
rect 41492 291078 41890 291138
rect 41830 291002 41890 291078
rect 49141 291002 49207 291005
rect 41830 291000 49207 291002
rect 41830 290944 49146 291000
rect 49202 290944 49207 291000
rect 41830 290942 49207 290944
rect 49141 290939 49207 290942
rect 62113 291002 62179 291005
rect 675753 291002 675819 291005
rect 676254 291002 676260 291004
rect 62113 291000 64154 291002
rect 62113 290944 62118 291000
rect 62174 290986 64154 291000
rect 675753 291000 676260 291002
rect 62174 290944 64676 290986
rect 62113 290942 64676 290944
rect 62113 290939 62179 290942
rect 64094 290926 64676 290942
rect 47577 290730 47643 290733
rect 41492 290728 47643 290730
rect 41492 290672 47582 290728
rect 47638 290672 47643 290728
rect 41492 290670 47643 290672
rect 47577 290667 47643 290670
rect 649950 290458 650010 290956
rect 675753 290944 675758 291000
rect 675814 290944 676260 291000
rect 675753 290942 676260 290944
rect 675753 290939 675819 290942
rect 676254 290940 676260 290942
rect 676324 290940 676330 291004
rect 651373 290458 651439 290461
rect 649950 290456 651439 290458
rect 649950 290400 651378 290456
rect 651434 290400 651439 290456
rect 649950 290398 651439 290400
rect 651373 290395 651439 290398
rect 651649 290458 651715 290461
rect 673729 290458 673795 290461
rect 651649 290456 673795 290458
rect 651649 290400 651654 290456
rect 651710 290400 673734 290456
rect 673790 290400 673795 290456
rect 651649 290398 673795 290400
rect 651649 290395 651715 290398
rect 673729 290395 673795 290398
rect 41781 290322 41847 290325
rect 41492 290320 41847 290322
rect 41492 290264 41786 290320
rect 41842 290264 41847 290320
rect 41492 290262 41847 290264
rect 41781 290259 41847 290262
rect 41822 289988 41828 290052
rect 41892 290050 41898 290052
rect 42190 290050 42196 290052
rect 41892 289990 42196 290050
rect 41892 289988 41898 289990
rect 42190 289988 42196 289990
rect 42260 289988 42266 290052
rect 63309 289778 63375 289781
rect 63309 289776 64706 289778
rect 63309 289720 63314 289776
rect 63370 289720 64706 289776
rect 63309 289718 64706 289720
rect 63309 289715 63375 289718
rect 40902 289172 40908 289236
rect 40972 289234 40978 289236
rect 41781 289234 41847 289237
rect 40972 289232 41847 289234
rect 40972 289176 41786 289232
rect 41842 289176 41847 289232
rect 40972 289174 41847 289176
rect 649950 289234 650010 289774
rect 652201 289234 652267 289237
rect 649950 289232 652267 289234
rect 649950 289176 652206 289232
rect 652262 289176 652267 289232
rect 649950 289174 652267 289176
rect 40972 289172 40978 289174
rect 41781 289171 41847 289174
rect 652201 289171 652267 289174
rect 651465 288690 651531 288693
rect 649950 288688 651531 288690
rect 649950 288632 651470 288688
rect 651526 288632 651531 288688
rect 649950 288630 651531 288632
rect 649950 288592 650010 288630
rect 651465 288627 651531 288630
rect 62389 288554 62455 288557
rect 64646 288554 64706 288592
rect 62389 288552 64706 288554
rect 62389 288496 62394 288552
rect 62450 288496 64706 288552
rect 62389 288494 64706 288496
rect 62389 288491 62455 288494
rect 673085 287874 673151 287877
rect 675109 287874 675175 287877
rect 673085 287872 675175 287874
rect 673085 287816 673090 287872
rect 673146 287816 675114 287872
rect 675170 287816 675175 287872
rect 673085 287814 675175 287816
rect 673085 287811 673151 287814
rect 675109 287811 675175 287814
rect 651465 287466 651531 287469
rect 649766 287464 651531 287466
rect 62297 287194 62363 287197
rect 64646 287194 64706 287410
rect 649766 287408 651470 287464
rect 651526 287408 651531 287464
rect 649766 287406 651531 287408
rect 651465 287403 651531 287406
rect 62297 287192 64706 287194
rect 62297 287136 62302 287192
rect 62358 287136 64706 287192
rect 62297 287134 64706 287136
rect 62297 287131 62363 287134
rect 673913 286922 673979 286925
rect 675109 286922 675175 286925
rect 673913 286920 675175 286922
rect 673913 286864 673918 286920
rect 673974 286864 675114 286920
rect 675170 286864 675175 286920
rect 673913 286862 675175 286864
rect 673913 286859 673979 286862
rect 675109 286859 675175 286862
rect 673545 286514 673611 286517
rect 675385 286514 675451 286517
rect 673545 286512 675451 286514
rect 673545 286456 673550 286512
rect 673606 286456 675390 286512
rect 675446 286456 675451 286512
rect 673545 286454 675451 286456
rect 673545 286451 673611 286454
rect 675385 286451 675451 286454
rect 63033 285970 63099 285973
rect 64646 285970 64706 286228
rect 63033 285968 64706 285970
rect 63033 285912 63038 285968
rect 63094 285912 64706 285968
rect 63033 285910 64706 285912
rect 649950 285970 650010 286228
rect 651465 285970 651531 285973
rect 649950 285968 651531 285970
rect 649950 285912 651470 285968
rect 651526 285912 651531 285968
rect 649950 285910 651531 285912
rect 63033 285907 63099 285910
rect 651465 285907 651531 285910
rect 42190 284820 42196 284884
rect 42260 284882 42266 284884
rect 42517 284882 42583 284885
rect 42260 284880 42583 284882
rect 42260 284824 42522 284880
rect 42578 284824 42583 284880
rect 42260 284822 42583 284824
rect 42260 284820 42266 284822
rect 42517 284819 42583 284822
rect 62113 284474 62179 284477
rect 64646 284474 64706 285046
rect 649950 284746 650010 285046
rect 651465 284746 651531 284749
rect 649950 284744 651531 284746
rect 649950 284688 651470 284744
rect 651526 284688 651531 284744
rect 649950 284686 651531 284688
rect 651465 284683 651531 284686
rect 62113 284472 64706 284474
rect 62113 284416 62118 284472
rect 62174 284416 64706 284472
rect 62113 284414 64706 284416
rect 62113 284411 62179 284414
rect 37917 284338 37983 284341
rect 41822 284338 41828 284340
rect 37917 284336 41828 284338
rect 37917 284280 37922 284336
rect 37978 284280 41828 284336
rect 37917 284278 41828 284280
rect 37917 284275 37983 284278
rect 41822 284276 41828 284278
rect 41892 284276 41898 284340
rect 62113 283250 62179 283253
rect 64646 283250 64706 283864
rect 62113 283248 64706 283250
rect 62113 283192 62118 283248
rect 62174 283192 64706 283248
rect 62113 283190 64706 283192
rect 649950 283250 650010 283864
rect 675753 283658 675819 283661
rect 676070 283658 676076 283660
rect 675753 283656 676076 283658
rect 675753 283600 675758 283656
rect 675814 283600 676076 283656
rect 675753 283598 676076 283600
rect 675753 283595 675819 283598
rect 676070 283596 676076 283598
rect 676140 283596 676146 283660
rect 652017 283522 652083 283525
rect 673913 283522 673979 283525
rect 652017 283520 673979 283522
rect 652017 283464 652022 283520
rect 652078 283464 673918 283520
rect 673974 283464 673979 283520
rect 652017 283462 673979 283464
rect 652017 283459 652083 283462
rect 673913 283459 673979 283462
rect 651465 283250 651531 283253
rect 649950 283248 651531 283250
rect 649950 283192 651470 283248
rect 651526 283192 651531 283248
rect 649950 283190 651531 283192
rect 62113 283187 62179 283190
rect 651465 283187 651531 283190
rect 675661 282706 675727 282709
rect 675886 282706 675892 282708
rect 675661 282704 675892 282706
rect 40902 282236 40908 282300
rect 40972 282298 40978 282300
rect 41781 282298 41847 282301
rect 40972 282296 41847 282298
rect 40972 282240 41786 282296
rect 41842 282240 41847 282296
rect 40972 282238 41847 282240
rect 40972 282236 40978 282238
rect 41781 282235 41847 282238
rect 62113 282162 62179 282165
rect 64646 282162 64706 282682
rect 62113 282160 64706 282162
rect 62113 282104 62118 282160
rect 62174 282104 64706 282160
rect 62113 282102 64706 282104
rect 649950 282162 650010 282682
rect 675661 282648 675666 282704
rect 675722 282648 675892 282704
rect 675661 282646 675892 282648
rect 675661 282643 675727 282646
rect 675886 282644 675892 282646
rect 675956 282644 675962 282708
rect 652017 282162 652083 282165
rect 649950 282160 652083 282162
rect 649950 282104 652022 282160
rect 652078 282104 652083 282160
rect 649950 282102 652083 282104
rect 62113 282099 62179 282102
rect 652017 282099 652083 282102
rect 42149 281756 42215 281757
rect 42149 281754 42196 281756
rect 42104 281752 42196 281754
rect 42104 281696 42154 281752
rect 42104 281694 42196 281696
rect 42149 281692 42196 281694
rect 42260 281692 42266 281756
rect 42149 281691 42215 281692
rect 675661 281620 675727 281621
rect 675661 281616 675708 281620
rect 675772 281618 675778 281620
rect 675661 281560 675666 281616
rect 675661 281556 675708 281560
rect 675772 281558 675818 281618
rect 675772 281556 675778 281558
rect 675661 281555 675727 281556
rect 63217 280938 63283 280941
rect 64646 280938 64706 281500
rect 63217 280936 64706 280938
rect 63217 280880 63222 280936
rect 63278 280880 64706 280936
rect 63217 280878 64706 280880
rect 649950 280938 650010 281500
rect 651465 280938 651531 280941
rect 649950 280936 651531 280938
rect 649950 280880 651470 280936
rect 651526 280880 651531 280936
rect 649950 280878 651531 280880
rect 63217 280875 63283 280878
rect 651465 280875 651531 280878
rect 62113 280394 62179 280397
rect 652569 280394 652635 280397
rect 62113 280392 64706 280394
rect 62113 280336 62118 280392
rect 62174 280336 64706 280392
rect 62113 280334 64706 280336
rect 62113 280331 62179 280334
rect 64646 280318 64706 280334
rect 649950 280392 652635 280394
rect 649950 280336 652574 280392
rect 652630 280336 652635 280392
rect 649950 280334 652635 280336
rect 649950 280318 650010 280334
rect 652569 280331 652635 280334
rect 42149 280260 42215 280261
rect 42149 280258 42196 280260
rect 42104 280256 42196 280258
rect 42104 280200 42154 280256
rect 42104 280198 42196 280200
rect 42149 280196 42196 280198
rect 42260 280196 42266 280260
rect 42149 280195 42215 280196
rect 42149 279714 42215 279717
rect 43437 279714 43503 279717
rect 42149 279712 43503 279714
rect 42149 279656 42154 279712
rect 42210 279656 43442 279712
rect 43498 279656 43503 279712
rect 42149 279654 43503 279656
rect 42149 279651 42215 279654
rect 43437 279651 43503 279654
rect 42190 278700 42196 278764
rect 42260 278762 42266 278764
rect 50521 278762 50587 278765
rect 42260 278760 50587 278762
rect 42260 278704 50526 278760
rect 50582 278704 50587 278760
rect 42260 278702 50587 278704
rect 42260 278700 42266 278702
rect 50521 278699 50587 278702
rect 60181 278762 60247 278765
rect 60181 278760 663810 278762
rect 60181 278704 60186 278760
rect 60242 278704 663810 278760
rect 60181 278702 663810 278704
rect 60181 278699 60247 278702
rect 42057 278490 42123 278493
rect 43621 278490 43687 278493
rect 42057 278488 43687 278490
rect 42057 278432 42062 278488
rect 42118 278432 43626 278488
rect 43682 278432 43687 278488
rect 42057 278430 43687 278432
rect 42057 278427 42123 278430
rect 43621 278427 43687 278430
rect 663750 278354 663810 278702
rect 671705 278626 671771 278629
rect 672901 278626 672967 278629
rect 671705 278624 672967 278626
rect 671705 278568 671710 278624
rect 671766 278568 672906 278624
rect 672962 278568 672967 278624
rect 671705 278566 672967 278568
rect 671705 278563 671771 278566
rect 672901 278563 672967 278566
rect 675109 278354 675175 278357
rect 663750 278352 675175 278354
rect 663750 278296 675114 278352
rect 675170 278296 675175 278352
rect 663750 278294 675175 278296
rect 675109 278291 675175 278294
rect 59997 278082 60063 278085
rect 675477 278082 675543 278085
rect 59997 278080 675543 278082
rect 59997 278024 60002 278080
rect 60058 278024 675482 278080
rect 675538 278024 675543 278080
rect 59997 278022 675543 278024
rect 59997 278019 60063 278022
rect 675477 278019 675543 278022
rect 42149 277946 42215 277949
rect 42793 277946 42859 277949
rect 42149 277944 42859 277946
rect 42149 277888 42154 277944
rect 42210 277888 42798 277944
rect 42854 277888 42859 277944
rect 42149 277886 42859 277888
rect 42149 277883 42215 277886
rect 42793 277883 42859 277886
rect 40718 277068 40724 277132
rect 40788 277130 40794 277132
rect 41781 277130 41847 277133
rect 40788 277128 41847 277130
rect 40788 277072 41786 277128
rect 41842 277072 41847 277128
rect 40788 277070 41847 277072
rect 40788 277068 40794 277070
rect 41781 277067 41847 277070
rect 53097 276722 53163 276725
rect 674925 276722 674991 276725
rect 53097 276720 674991 276722
rect 53097 276664 53102 276720
rect 53158 276664 674930 276720
rect 674986 276664 674991 276720
rect 53097 276662 674991 276664
rect 53097 276659 53163 276662
rect 674925 276659 674991 276662
rect 42793 275906 42859 275909
rect 57237 275906 57303 275909
rect 42793 275904 57303 275906
rect 42793 275848 42798 275904
rect 42854 275848 57242 275904
rect 57298 275848 57303 275904
rect 42793 275846 57303 275848
rect 42793 275843 42859 275846
rect 57237 275843 57303 275846
rect 40534 274212 40540 274276
rect 40604 274274 40610 274276
rect 41781 274274 41847 274277
rect 40604 274272 41847 274274
rect 40604 274216 41786 274272
rect 41842 274216 41847 274272
rect 40604 274214 41847 274216
rect 40604 274212 40610 274214
rect 41781 274211 41847 274214
rect 539317 274002 539383 274005
rect 545941 274002 546007 274005
rect 539317 274000 546007 274002
rect 539317 273944 539322 274000
rect 539378 273944 545946 274000
rect 546002 273944 546007 274000
rect 539317 273942 546007 273944
rect 539317 273939 539383 273942
rect 545941 273939 546007 273942
rect 43437 273866 43503 273869
rect 62205 273866 62271 273869
rect 43437 273864 62271 273866
rect 43437 273808 43442 273864
rect 43498 273808 62210 273864
rect 62266 273808 62271 273864
rect 43437 273806 62271 273808
rect 43437 273803 43503 273806
rect 62205 273803 62271 273806
rect 674925 273866 674991 273869
rect 675334 273866 675340 273868
rect 674925 273864 675340 273866
rect 674925 273808 674930 273864
rect 674986 273808 675340 273864
rect 674925 273806 675340 273808
rect 674925 273803 674991 273806
rect 675334 273804 675340 273806
rect 675404 273804 675410 273868
rect 42149 273050 42215 273053
rect 45185 273050 45251 273053
rect 42149 273048 45251 273050
rect 42149 272992 42154 273048
rect 42210 272992 45190 273048
rect 45246 272992 45251 273048
rect 42149 272990 45251 272992
rect 42149 272987 42215 272990
rect 45185 272987 45251 272990
rect 461025 272914 461091 272917
rect 466269 272914 466335 272917
rect 461025 272912 466335 272914
rect 461025 272856 461030 272912
rect 461086 272856 466274 272912
rect 466330 272856 466335 272912
rect 461025 272854 466335 272856
rect 461025 272851 461091 272854
rect 466269 272851 466335 272854
rect 460841 272642 460907 272645
rect 461853 272642 461919 272645
rect 460841 272640 461919 272642
rect 460841 272584 460846 272640
rect 460902 272584 461858 272640
rect 461914 272584 461919 272640
rect 460841 272582 461919 272584
rect 460841 272579 460907 272582
rect 461853 272579 461919 272582
rect 464705 272506 464771 272509
rect 470685 272506 470751 272509
rect 464705 272504 470751 272506
rect 464705 272448 464710 272504
rect 464766 272448 470690 272504
rect 470746 272448 470751 272504
rect 464705 272446 470751 272448
rect 464705 272443 464771 272446
rect 470685 272443 470751 272446
rect 536557 272506 536623 272509
rect 547689 272506 547755 272509
rect 536557 272504 547755 272506
rect 536557 272448 536562 272504
rect 536618 272448 547694 272504
rect 547750 272448 547755 272504
rect 536557 272446 547755 272448
rect 536557 272443 536623 272446
rect 547689 272443 547755 272446
rect 479517 272098 479583 272101
rect 480529 272098 480595 272101
rect 479517 272096 480595 272098
rect 479517 272040 479522 272096
rect 479578 272040 480534 272096
rect 480590 272040 480595 272096
rect 479517 272038 480595 272040
rect 479517 272035 479583 272038
rect 480529 272035 480595 272038
rect 547505 272098 547571 272101
rect 547873 272098 547939 272101
rect 547505 272096 547939 272098
rect 547505 272040 547510 272096
rect 547566 272040 547878 272096
rect 547934 272040 547939 272096
rect 547505 272038 547939 272040
rect 547505 272035 547571 272038
rect 547873 272035 547939 272038
rect 470593 271962 470659 271965
rect 478045 271962 478111 271965
rect 470593 271960 478111 271962
rect 470593 271904 470598 271960
rect 470654 271904 478050 271960
rect 478106 271904 478111 271960
rect 470593 271902 478111 271904
rect 470593 271899 470659 271902
rect 478045 271899 478111 271902
rect 501597 271962 501663 271965
rect 504541 271962 504607 271965
rect 501597 271960 504607 271962
rect 501597 271904 501602 271960
rect 501658 271904 504546 271960
rect 504602 271904 504607 271960
rect 501597 271902 504607 271904
rect 501597 271899 501663 271902
rect 504541 271899 504607 271902
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 530393 270194 530459 270197
rect 534073 270194 534139 270197
rect 530393 270192 534139 270194
rect 530393 270136 530398 270192
rect 530454 270136 534078 270192
rect 534134 270136 534139 270192
rect 530393 270134 534139 270136
rect 530393 270131 530459 270134
rect 534073 270131 534139 270134
rect 509233 269922 509299 269925
rect 516593 269922 516659 269925
rect 509233 269920 516659 269922
rect 509233 269864 509238 269920
rect 509294 269864 516598 269920
rect 516654 269864 516659 269920
rect 509233 269862 516659 269864
rect 509233 269859 509299 269862
rect 516593 269859 516659 269862
rect 41781 269788 41847 269789
rect 41781 269784 41828 269788
rect 41892 269786 41898 269788
rect 538029 269786 538095 269789
rect 541341 269786 541407 269789
rect 41781 269728 41786 269784
rect 41781 269724 41828 269728
rect 41892 269726 41938 269786
rect 538029 269784 541407 269786
rect 538029 269728 538034 269784
rect 538090 269728 541346 269784
rect 541402 269728 541407 269784
rect 538029 269726 541407 269728
rect 41892 269724 41898 269726
rect 41781 269723 41847 269724
rect 538029 269723 538095 269726
rect 541341 269723 541407 269726
rect 509141 269514 509207 269517
rect 509877 269514 509943 269517
rect 509141 269512 509943 269514
rect 509141 269456 509146 269512
rect 509202 269456 509882 269512
rect 509938 269456 509943 269512
rect 509141 269454 509943 269456
rect 509141 269451 509207 269454
rect 509877 269451 509943 269454
rect 41965 269108 42031 269109
rect 41965 269104 42012 269108
rect 42076 269106 42082 269108
rect 41965 269048 41970 269104
rect 41965 269044 42012 269048
rect 42076 269046 42122 269106
rect 42076 269044 42082 269046
rect 41965 269043 42031 269044
rect 665817 268562 665883 268565
rect 676262 268562 676322 268668
rect 665817 268560 676322 268562
rect 665817 268504 665822 268560
rect 665878 268504 676322 268560
rect 665817 268502 676322 268504
rect 665817 268499 665883 268502
rect 673913 268290 673979 268293
rect 673913 268288 676292 268290
rect 673913 268232 673918 268288
rect 673974 268232 676292 268288
rect 673913 268230 676292 268232
rect 673913 268227 673979 268230
rect 673729 267882 673795 267885
rect 673729 267880 676292 267882
rect 673729 267824 673734 267880
rect 673790 267824 676292 267880
rect 673729 267822 676292 267824
rect 673729 267819 673795 267822
rect 673361 267474 673427 267477
rect 673361 267472 676292 267474
rect 673361 267416 673366 267472
rect 673422 267416 676292 267472
rect 673361 267414 676292 267416
rect 673361 267411 673427 267414
rect 673913 267066 673979 267069
rect 673913 267064 676292 267066
rect 673913 267008 673918 267064
rect 673974 267008 676292 267064
rect 673913 267006 676292 267008
rect 673913 267003 673979 267006
rect 673177 266658 673243 266661
rect 673177 266656 676292 266658
rect 673177 266600 673182 266656
rect 673238 266600 676292 266656
rect 673177 266598 676292 266600
rect 673177 266595 673243 266598
rect 42149 266250 42215 266253
rect 51901 266250 51967 266253
rect 42149 266248 51967 266250
rect 42149 266192 42154 266248
rect 42210 266192 51906 266248
rect 51962 266192 51967 266248
rect 42149 266190 51967 266192
rect 42149 266187 42215 266190
rect 51901 266187 51967 266190
rect 674373 266250 674439 266253
rect 674373 266248 676292 266250
rect 674373 266192 674378 266248
rect 674434 266192 676292 266248
rect 674373 266190 676292 266192
rect 674373 266187 674439 266190
rect 674557 265842 674623 265845
rect 674557 265840 676292 265842
rect 674557 265784 674562 265840
rect 674618 265784 676292 265840
rect 674557 265782 676292 265784
rect 674557 265779 674623 265782
rect 672349 265434 672415 265437
rect 672349 265432 676292 265434
rect 672349 265376 672354 265432
rect 672410 265376 676292 265432
rect 672349 265374 676292 265376
rect 672349 265371 672415 265374
rect 674741 265026 674807 265029
rect 674741 265024 676292 265026
rect 674741 264968 674746 265024
rect 674802 264968 676292 265024
rect 674741 264966 676292 264968
rect 674741 264963 674807 264966
rect 673545 264618 673611 264621
rect 673545 264616 676292 264618
rect 673545 264560 673550 264616
rect 673606 264560 676292 264616
rect 673545 264558 676292 264560
rect 673545 264555 673611 264558
rect 55857 264210 55923 264213
rect 675109 264210 675175 264213
rect 55857 264208 675175 264210
rect 55857 264152 55862 264208
rect 55918 264152 675114 264208
rect 675170 264152 675175 264208
rect 55857 264150 675175 264152
rect 55857 264147 55923 264150
rect 675109 264147 675175 264150
rect 676446 264077 676506 264180
rect 676397 264072 676506 264077
rect 676397 264016 676402 264072
rect 676458 264016 676506 264072
rect 676397 264014 676506 264016
rect 676397 264011 676463 264014
rect 670325 263802 670391 263805
rect 670325 263800 676292 263802
rect 670325 263744 670330 263800
rect 670386 263744 676292 263800
rect 670325 263742 676292 263744
rect 670325 263739 670391 263742
rect 673177 263394 673243 263397
rect 673177 263392 676292 263394
rect 673177 263336 673182 263392
rect 673238 263336 676292 263392
rect 673177 263334 676292 263336
rect 673177 263331 673243 263334
rect 676262 262853 676322 262956
rect 676213 262848 676322 262853
rect 676213 262792 676218 262848
rect 676274 262792 676322 262848
rect 676213 262790 676322 262792
rect 676213 262787 676279 262790
rect 674465 262578 674531 262581
rect 674465 262576 676292 262578
rect 674465 262520 674470 262576
rect 674526 262520 676292 262576
rect 674465 262518 676292 262520
rect 674465 262515 674531 262518
rect 554405 262170 554471 262173
rect 552460 262168 554471 262170
rect 552460 262112 554410 262168
rect 554466 262112 554471 262168
rect 552460 262110 554471 262112
rect 554405 262107 554471 262110
rect 670969 262170 671035 262173
rect 670969 262168 676292 262170
rect 670969 262112 670974 262168
rect 671030 262112 676292 262168
rect 670969 262110 676292 262112
rect 670969 262107 671035 262110
rect 676998 261628 677058 261732
rect 676990 261564 676996 261628
rect 677060 261564 677066 261628
rect 676814 261220 676874 261324
rect 676806 261156 676812 261220
rect 676876 261156 676882 261220
rect 673729 260946 673795 260949
rect 673729 260944 676292 260946
rect 673729 260888 673734 260944
rect 673790 260888 676292 260944
rect 673729 260886 676292 260888
rect 673729 260883 673795 260886
rect 671705 260538 671771 260541
rect 671705 260536 676292 260538
rect 671705 260480 671710 260536
rect 671766 260480 676292 260536
rect 671705 260478 676292 260480
rect 671705 260475 671771 260478
rect 674373 260130 674439 260133
rect 674373 260128 676292 260130
rect 674373 260072 674378 260128
rect 674434 260072 676292 260128
rect 674373 260070 676292 260072
rect 674373 260067 674439 260070
rect 554313 259994 554379 259997
rect 552460 259992 554379 259994
rect 552460 259936 554318 259992
rect 554374 259936 554379 259992
rect 552460 259934 554379 259936
rect 554313 259931 554379 259934
rect 672993 259722 673059 259725
rect 672993 259720 676292 259722
rect 672993 259664 672998 259720
rect 673054 259664 676292 259720
rect 672993 259662 676292 259664
rect 672993 259659 673059 259662
rect 674097 259314 674163 259317
rect 674097 259312 676292 259314
rect 674097 259256 674102 259312
rect 674158 259256 676292 259312
rect 674097 259254 676292 259256
rect 674097 259251 674163 259254
rect 673269 258906 673335 258909
rect 673269 258904 676292 258906
rect 673269 258848 673274 258904
rect 673330 258848 676292 258904
rect 673269 258846 676292 258848
rect 673269 258843 673335 258846
rect 670141 258498 670207 258501
rect 670141 258496 676292 258498
rect 670141 258440 670146 258496
rect 670202 258440 676292 258496
rect 670141 258438 676292 258440
rect 670141 258435 670207 258438
rect 46381 258090 46447 258093
rect 675477 258092 675543 258093
rect 675477 258090 675524 258092
rect 41492 258088 46447 258090
rect 41492 258032 46386 258088
rect 46442 258032 46447 258088
rect 41492 258030 46447 258032
rect 675396 258088 675524 258090
rect 675588 258090 675594 258092
rect 675396 258032 675482 258088
rect 675588 258060 676292 258090
rect 675396 258030 675524 258032
rect 46381 258027 46447 258030
rect 675477 258028 675524 258030
rect 675588 258030 676322 258060
rect 675588 258028 675594 258030
rect 675477 258027 675543 258028
rect 553945 257818 554011 257821
rect 552460 257816 554011 257818
rect 552460 257760 553950 257816
rect 554006 257760 554011 257816
rect 552460 257758 554011 257760
rect 553945 257755 554011 257758
rect 676262 257652 676322 258030
rect 41462 257546 41522 257652
rect 41462 257486 51090 257546
rect 35574 257141 35634 257244
rect 35574 257136 35683 257141
rect 35574 257080 35622 257136
rect 35678 257080 35683 257136
rect 35574 257078 35683 257080
rect 35617 257075 35683 257078
rect 39481 257138 39547 257141
rect 42793 257138 42859 257141
rect 39481 257136 42859 257138
rect 39481 257080 39486 257136
rect 39542 257080 42798 257136
rect 42854 257080 42859 257136
rect 39481 257078 42859 257080
rect 39481 257075 39547 257078
rect 42793 257075 42859 257078
rect 35758 256733 35818 256836
rect 35758 256728 35867 256733
rect 35758 256672 35806 256728
rect 35862 256672 35867 256728
rect 35758 256670 35867 256672
rect 51030 256730 51090 257486
rect 670693 257274 670759 257277
rect 670693 257272 676292 257274
rect 670693 257216 670698 257272
rect 670754 257216 676292 257272
rect 670693 257214 676292 257216
rect 670693 257211 670759 257214
rect 60365 256730 60431 256733
rect 51030 256728 60431 256730
rect 51030 256672 60370 256728
rect 60426 256672 60431 256728
rect 51030 256670 60431 256672
rect 35801 256667 35867 256670
rect 60365 256667 60431 256670
rect 35758 256325 35818 256428
rect 35758 256320 35867 256325
rect 35758 256264 35806 256320
rect 35862 256264 35867 256320
rect 35758 256262 35867 256264
rect 35801 256259 35867 256262
rect 45001 256050 45067 256053
rect 41492 256048 45067 256050
rect 41492 255992 45006 256048
rect 45062 255992 45067 256048
rect 41492 255990 45067 255992
rect 45001 255987 45067 255990
rect 45645 255642 45711 255645
rect 554497 255642 554563 255645
rect 41492 255640 45711 255642
rect 41492 255584 45650 255640
rect 45706 255584 45711 255640
rect 41492 255582 45711 255584
rect 552460 255640 554563 255642
rect 552460 255584 554502 255640
rect 554558 255584 554563 255640
rect 552460 255582 554563 255584
rect 45645 255579 45711 255582
rect 554497 255579 554563 255582
rect 44265 255234 44331 255237
rect 41492 255232 44331 255234
rect 41492 255176 44270 255232
rect 44326 255176 44331 255232
rect 41492 255174 44331 255176
rect 44265 255171 44331 255174
rect 674925 254962 674991 254965
rect 675845 254962 675911 254965
rect 674925 254960 675911 254962
rect 674925 254904 674930 254960
rect 674986 254904 675850 254960
rect 675906 254904 675911 254960
rect 674925 254902 675911 254904
rect 674925 254899 674991 254902
rect 675845 254899 675911 254902
rect 44173 254826 44239 254829
rect 41492 254824 44239 254826
rect 41492 254768 44178 254824
rect 44234 254768 44239 254824
rect 41492 254766 44239 254768
rect 44173 254763 44239 254766
rect 44541 254418 44607 254421
rect 41492 254416 44607 254418
rect 41492 254360 44546 254416
rect 44602 254360 44607 254416
rect 41492 254358 44607 254360
rect 44541 254355 44607 254358
rect 46197 254010 46263 254013
rect 41492 254008 46263 254010
rect 41492 253952 46202 254008
rect 46258 253952 46263 254008
rect 41492 253950 46263 253952
rect 46197 253947 46263 253950
rect 35574 253469 35634 253572
rect 35574 253464 35683 253469
rect 35574 253408 35622 253464
rect 35678 253408 35683 253464
rect 35574 253406 35683 253408
rect 35617 253403 35683 253406
rect 40217 253466 40283 253469
rect 42793 253466 42859 253469
rect 554405 253466 554471 253469
rect 40217 253464 42859 253466
rect 40217 253408 40222 253464
rect 40278 253408 42798 253464
rect 42854 253408 42859 253464
rect 40217 253406 42859 253408
rect 552460 253464 554471 253466
rect 552460 253408 554410 253464
rect 554466 253408 554471 253464
rect 552460 253406 554471 253408
rect 40217 253403 40283 253406
rect 42793 253403 42859 253406
rect 554405 253403 554471 253406
rect 35758 253061 35818 253164
rect 35758 253056 35867 253061
rect 35758 253000 35806 253056
rect 35862 253000 35867 253056
rect 35758 252998 35867 253000
rect 35801 252995 35867 252998
rect 45921 252786 45987 252789
rect 41492 252784 45987 252786
rect 41492 252728 45926 252784
rect 45982 252728 45987 252784
rect 41492 252726 45987 252728
rect 45921 252723 45987 252726
rect 35758 252245 35818 252348
rect 35758 252240 35867 252245
rect 35758 252184 35806 252240
rect 35862 252184 35867 252240
rect 35758 252182 35867 252184
rect 35801 252179 35867 252182
rect 46933 251970 46999 251973
rect 41492 251968 46999 251970
rect 41492 251912 46938 251968
rect 46994 251912 46999 251968
rect 41492 251910 46999 251912
rect 46933 251907 46999 251910
rect 47117 251562 47183 251565
rect 41492 251560 47183 251562
rect 41492 251504 47122 251560
rect 47178 251504 47183 251560
rect 41492 251502 47183 251504
rect 47117 251499 47183 251502
rect 554129 251290 554195 251293
rect 552460 251288 554195 251290
rect 552460 251232 554134 251288
rect 554190 251232 554195 251288
rect 552460 251230 554195 251232
rect 554129 251227 554195 251230
rect 44541 251154 44607 251157
rect 41492 251152 44607 251154
rect 41492 251096 44546 251152
rect 44602 251096 44607 251152
rect 41492 251094 44607 251096
rect 44541 251091 44607 251094
rect 673085 250746 673151 250749
rect 675477 250746 675543 250749
rect 673085 250744 675543 250746
rect 35574 250613 35634 250716
rect 673085 250688 673090 250744
rect 673146 250688 675482 250744
rect 675538 250688 675543 250744
rect 673085 250686 675543 250688
rect 673085 250683 673151 250686
rect 675477 250683 675543 250686
rect 35574 250608 35683 250613
rect 35574 250552 35622 250608
rect 35678 250552 35683 250608
rect 35574 250550 35683 250552
rect 35617 250547 35683 250550
rect 675753 250338 675819 250341
rect 676990 250338 676996 250340
rect 675753 250336 676996 250338
rect 35758 250205 35818 250308
rect 675753 250280 675758 250336
rect 675814 250280 676996 250336
rect 675753 250278 676996 250280
rect 675753 250275 675819 250278
rect 676990 250276 676996 250278
rect 677060 250276 677066 250340
rect 35758 250200 35867 250205
rect 35758 250144 35806 250200
rect 35862 250144 35867 250200
rect 35758 250142 35867 250144
rect 35801 250139 35867 250142
rect 673085 250066 673151 250069
rect 675518 250066 675524 250068
rect 673085 250064 675524 250066
rect 673085 250008 673090 250064
rect 673146 250008 675524 250064
rect 673085 250006 675524 250008
rect 673085 250003 673151 250006
rect 675518 250004 675524 250006
rect 675588 250004 675594 250068
rect 40542 249796 40602 249900
rect 40534 249732 40540 249796
rect 40604 249732 40610 249796
rect 675334 249732 675340 249796
rect 675404 249732 675410 249796
rect 674925 249522 674991 249525
rect 675342 249522 675402 249732
rect 674925 249520 675402 249522
rect 40726 249388 40786 249492
rect 674925 249464 674930 249520
rect 674986 249464 675402 249520
rect 674925 249462 675402 249464
rect 674925 249459 674991 249462
rect 40718 249324 40724 249388
rect 40788 249324 40794 249388
rect 44357 249114 44423 249117
rect 554037 249114 554103 249117
rect 41492 249112 44423 249114
rect 41492 249056 44362 249112
rect 44418 249056 44423 249112
rect 41492 249054 44423 249056
rect 552460 249112 554103 249114
rect 552460 249056 554042 249112
rect 554098 249056 554103 249112
rect 552460 249054 554103 249056
rect 44357 249051 44423 249054
rect 554037 249051 554103 249054
rect 45001 248706 45067 248709
rect 41492 248704 45067 248706
rect 41492 248648 45006 248704
rect 45062 248648 45067 248704
rect 41492 248646 45067 248648
rect 45001 248643 45067 248646
rect 46381 248298 46447 248301
rect 41492 248296 46447 248298
rect 41492 248240 46386 248296
rect 46442 248240 46447 248296
rect 41492 248238 46447 248240
rect 46381 248235 46447 248238
rect 675293 248162 675359 248165
rect 666510 248160 675359 248162
rect 666510 248104 675298 248160
rect 675354 248104 675359 248160
rect 666510 248102 675359 248104
rect 664437 248026 664503 248029
rect 666510 248026 666570 248102
rect 675293 248099 675359 248102
rect 664437 248024 666570 248026
rect 664437 247968 664442 248024
rect 664498 247968 666570 248024
rect 664437 247966 666570 247968
rect 664437 247963 664503 247966
rect 35758 247757 35818 247860
rect 35758 247752 35867 247757
rect 35758 247696 35806 247752
rect 35862 247696 35867 247752
rect 35758 247694 35867 247696
rect 35801 247691 35867 247694
rect 50521 247482 50587 247485
rect 41492 247480 50587 247482
rect 41492 247424 50526 247480
rect 50582 247424 50587 247480
rect 41492 247422 50587 247424
rect 50521 247419 50587 247422
rect 34470 246941 34530 247044
rect 34421 246936 34530 246941
rect 553853 246938 553919 246941
rect 34421 246880 34426 246936
rect 34482 246880 34530 246936
rect 34421 246878 34530 246880
rect 552460 246936 553919 246938
rect 552460 246880 553858 246936
rect 553914 246880 553919 246936
rect 552460 246878 553919 246880
rect 34421 246875 34487 246878
rect 553853 246875 553919 246878
rect 673729 246666 673795 246669
rect 675293 246666 675359 246669
rect 673729 246664 675359 246666
rect 673729 246608 673734 246664
rect 673790 246608 675298 246664
rect 675354 246608 675359 246664
rect 673729 246606 675359 246608
rect 673729 246603 673795 246606
rect 675293 246603 675359 246606
rect 675753 246666 675819 246669
rect 676806 246666 676812 246668
rect 675753 246664 676812 246666
rect 675753 246608 675758 246664
rect 675814 246608 676812 246664
rect 675753 246606 676812 246608
rect 675753 246603 675819 246606
rect 676806 246604 676812 246606
rect 676876 246604 676882 246668
rect 672165 246258 672231 246261
rect 673310 246258 673316 246260
rect 672165 246256 673316 246258
rect 672165 246200 672170 246256
rect 672226 246200 673316 246256
rect 672165 246198 673316 246200
rect 672165 246195 672231 246198
rect 673310 246196 673316 246198
rect 673380 246196 673386 246260
rect 675109 246258 675175 246261
rect 675518 246258 675524 246260
rect 675109 246256 675524 246258
rect 675109 246200 675114 246256
rect 675170 246200 675524 246256
rect 675109 246198 675524 246200
rect 675109 246195 675175 246198
rect 675518 246196 675524 246198
rect 675588 246196 675594 246260
rect 40125 245714 40191 245717
rect 43621 245714 43687 245717
rect 40125 245712 43687 245714
rect 40125 245656 40130 245712
rect 40186 245656 43626 245712
rect 43682 245656 43687 245712
rect 40125 245654 43687 245656
rect 40125 245651 40191 245654
rect 43621 245651 43687 245654
rect 666553 245714 666619 245717
rect 667790 245714 667796 245716
rect 666553 245712 667796 245714
rect 666553 245656 666558 245712
rect 666614 245656 667796 245712
rect 666553 245654 667796 245656
rect 666553 245651 666619 245654
rect 667790 245652 667796 245654
rect 667860 245652 667866 245716
rect 672993 245714 673059 245717
rect 675293 245714 675359 245717
rect 672993 245712 675359 245714
rect 672993 245656 672998 245712
rect 673054 245656 675298 245712
rect 675354 245656 675359 245712
rect 672993 245654 675359 245656
rect 672993 245651 673059 245654
rect 675293 245651 675359 245654
rect 672993 245442 673059 245445
rect 675017 245442 675083 245445
rect 672993 245440 675083 245442
rect 672993 245384 672998 245440
rect 673054 245384 675022 245440
rect 675078 245384 675083 245440
rect 672993 245382 675083 245384
rect 672993 245379 673059 245382
rect 675017 245379 675083 245382
rect 553485 244762 553551 244765
rect 552460 244760 553551 244762
rect 552460 244704 553490 244760
rect 553546 244704 553551 244760
rect 552460 244702 553551 244704
rect 553485 244699 553551 244702
rect 39849 244082 39915 244085
rect 43437 244082 43503 244085
rect 39849 244080 43503 244082
rect 39849 244024 39854 244080
rect 39910 244024 43442 244080
rect 43498 244024 43503 244080
rect 39849 244022 43503 244024
rect 39849 244019 39915 244022
rect 43437 244019 43503 244022
rect 675385 243266 675451 243269
rect 674606 243264 675451 243266
rect 674606 243208 675390 243264
rect 675446 243208 675451 243264
rect 674606 243206 675451 243208
rect 674606 242997 674666 243206
rect 675385 243203 675451 243206
rect 674557 242992 674666 242997
rect 674557 242936 674562 242992
rect 674618 242936 674666 242992
rect 674557 242934 674666 242936
rect 674557 242931 674623 242934
rect 674097 242722 674163 242725
rect 675477 242722 675543 242725
rect 674097 242720 675543 242722
rect 674097 242664 674102 242720
rect 674158 242664 675482 242720
rect 675538 242664 675543 242720
rect 674097 242662 675543 242664
rect 674097 242659 674163 242662
rect 675477 242659 675543 242662
rect 553669 242586 553735 242589
rect 552460 242584 553735 242586
rect 552460 242528 553674 242584
rect 553730 242528 553735 242584
rect 552460 242526 553735 242528
rect 553669 242523 553735 242526
rect 674373 242178 674439 242181
rect 675477 242178 675543 242181
rect 674373 242176 675543 242178
rect 674373 242120 674378 242176
rect 674434 242120 675482 242176
rect 675538 242120 675543 242176
rect 674373 242118 675543 242120
rect 674373 242115 674439 242118
rect 675477 242115 675543 242118
rect 673545 241770 673611 241773
rect 676806 241770 676812 241772
rect 673545 241768 676812 241770
rect 673545 241712 673550 241768
rect 673606 241712 676812 241768
rect 673545 241710 676812 241712
rect 673545 241707 673611 241710
rect 676806 241708 676812 241710
rect 676876 241708 676882 241772
rect 673269 241498 673335 241501
rect 675477 241498 675543 241501
rect 673269 241496 675543 241498
rect 673269 241440 673274 241496
rect 673330 241440 675482 241496
rect 675538 241440 675543 241496
rect 673269 241438 675543 241440
rect 673269 241435 673335 241438
rect 675477 241435 675543 241438
rect 40677 240954 40743 240957
rect 43069 240954 43135 240957
rect 40677 240952 43135 240954
rect 40677 240896 40682 240952
rect 40738 240896 43074 240952
rect 43130 240896 43135 240952
rect 40677 240894 43135 240896
rect 40677 240891 40743 240894
rect 43069 240891 43135 240894
rect 554497 240410 554563 240413
rect 552460 240408 554563 240410
rect 552460 240352 554502 240408
rect 554558 240352 554563 240408
rect 552460 240350 554563 240352
rect 554497 240347 554563 240350
rect 671705 240274 671771 240277
rect 675477 240274 675543 240277
rect 671705 240272 675543 240274
rect 671705 240216 671710 240272
rect 671766 240216 675482 240272
rect 675538 240216 675543 240272
rect 671705 240214 675543 240216
rect 671705 240211 671771 240214
rect 675477 240211 675543 240214
rect 42057 240138 42123 240141
rect 47117 240138 47183 240141
rect 42057 240136 47183 240138
rect 42057 240080 42062 240136
rect 42118 240080 47122 240136
rect 47178 240080 47183 240136
rect 42057 240078 47183 240080
rect 42057 240075 42123 240078
rect 47117 240075 47183 240078
rect 670325 238642 670391 238645
rect 675477 238642 675543 238645
rect 670325 238640 675543 238642
rect 670325 238584 670330 238640
rect 670386 238584 675482 238640
rect 675538 238584 675543 238640
rect 670325 238582 675543 238584
rect 670325 238579 670391 238582
rect 675477 238579 675543 238582
rect 554313 238234 554379 238237
rect 552460 238232 554379 238234
rect 552460 238176 554318 238232
rect 554374 238176 554379 238232
rect 552460 238174 554379 238176
rect 554313 238171 554379 238174
rect 42006 238036 42012 238100
rect 42076 238098 42082 238100
rect 42517 238098 42583 238101
rect 42076 238096 42583 238098
rect 42076 238040 42522 238096
rect 42578 238040 42583 238096
rect 42076 238038 42583 238040
rect 42076 238036 42082 238038
rect 42517 238035 42583 238038
rect 675017 237282 675083 237285
rect 675477 237282 675543 237285
rect 675017 237280 675543 237282
rect 675017 237224 675022 237280
rect 675078 237224 675482 237280
rect 675538 237224 675543 237280
rect 675017 237222 675543 237224
rect 675017 237219 675083 237222
rect 675477 237219 675543 237222
rect 672257 237010 672323 237013
rect 673729 237010 673795 237013
rect 672257 237008 673795 237010
rect 672257 236952 672262 237008
rect 672318 236952 673734 237008
rect 673790 236952 673795 237008
rect 672257 236950 673795 236952
rect 672257 236947 672323 236950
rect 673729 236947 673795 236950
rect 40534 236540 40540 236604
rect 40604 236602 40610 236604
rect 41781 236602 41847 236605
rect 40604 236600 41847 236602
rect 40604 236544 41786 236600
rect 41842 236544 41847 236600
rect 40604 236542 41847 236544
rect 40604 236540 40610 236542
rect 41781 236539 41847 236542
rect 672947 236466 673013 236469
rect 674649 236466 674715 236469
rect 672947 236464 674715 236466
rect 672947 236408 672952 236464
rect 673008 236408 674654 236464
rect 674710 236408 674715 236464
rect 672947 236406 674715 236408
rect 672947 236403 673013 236406
rect 674649 236403 674715 236406
rect 670969 236194 671035 236197
rect 675477 236194 675543 236197
rect 670969 236192 675543 236194
rect 670969 236136 670974 236192
rect 671030 236136 675482 236192
rect 675538 236136 675543 236192
rect 670969 236134 675543 236136
rect 670969 236131 671035 236134
rect 675477 236131 675543 236134
rect 553761 236058 553827 236061
rect 552460 236056 553827 236058
rect 552460 236000 553766 236056
rect 553822 236000 553827 236056
rect 552460 235998 553827 236000
rect 553761 235995 553827 235998
rect 42425 235922 42491 235925
rect 46381 235922 46447 235925
rect 42425 235920 46447 235922
rect 42425 235864 42430 235920
rect 42486 235864 46386 235920
rect 46442 235864 46447 235920
rect 42425 235862 46447 235864
rect 42425 235859 42491 235862
rect 46381 235859 46447 235862
rect 675477 235516 675543 235517
rect 675477 235514 675524 235516
rect 675432 235512 675524 235514
rect 675432 235456 675482 235512
rect 675432 235454 675524 235456
rect 675477 235452 675524 235454
rect 675588 235452 675594 235516
rect 675477 235451 675543 235452
rect 40718 234636 40724 234700
rect 40788 234698 40794 234700
rect 41781 234698 41847 234701
rect 40788 234696 41847 234698
rect 40788 234640 41786 234696
rect 41842 234640 41847 234696
rect 40788 234638 41847 234640
rect 40788 234636 40794 234638
rect 41781 234635 41847 234638
rect 42425 234562 42491 234565
rect 45001 234562 45067 234565
rect 42425 234560 45067 234562
rect 42425 234504 42430 234560
rect 42486 234504 45006 234560
rect 45062 234504 45067 234560
rect 42425 234502 45067 234504
rect 42425 234499 42491 234502
rect 45001 234499 45067 234502
rect 670877 234018 670943 234021
rect 675845 234018 675911 234021
rect 670877 234016 675911 234018
rect 670877 233960 670882 234016
rect 670938 233960 675850 234016
rect 675906 233960 675911 234016
rect 670877 233958 675911 233960
rect 670877 233955 670943 233958
rect 675845 233955 675911 233958
rect 554405 233882 554471 233885
rect 552460 233880 554471 233882
rect 552460 233824 554410 233880
rect 554466 233824 554471 233880
rect 552460 233822 554471 233824
rect 554405 233819 554471 233822
rect 674097 232658 674163 232661
rect 675845 232658 675911 232661
rect 674097 232656 675911 232658
rect 674097 232600 674102 232656
rect 674158 232600 675850 232656
rect 675906 232600 675911 232656
rect 674097 232598 675911 232600
rect 674097 232595 674163 232598
rect 675845 232595 675911 232598
rect 668669 232522 668735 232525
rect 673545 232522 673611 232525
rect 668669 232520 673611 232522
rect 668669 232464 668674 232520
rect 668730 232464 673550 232520
rect 673606 232464 673611 232520
rect 668669 232462 673611 232464
rect 668669 232459 668735 232462
rect 673545 232459 673611 232462
rect 674097 232386 674163 232389
rect 676029 232386 676095 232389
rect 674097 232384 676095 232386
rect 674097 232328 674102 232384
rect 674158 232328 676034 232384
rect 676090 232328 676095 232384
rect 674097 232326 676095 232328
rect 674097 232323 674163 232326
rect 676029 232323 676095 232326
rect 42425 232250 42491 232253
rect 46933 232250 46999 232253
rect 42425 232248 46999 232250
rect 42425 232192 42430 232248
rect 42486 232192 46938 232248
rect 46994 232192 46999 232248
rect 42425 232190 46999 232192
rect 42425 232187 42491 232190
rect 46933 232187 46999 232190
rect 670734 231916 670740 231980
rect 670804 231978 670810 231980
rect 671889 231978 671955 231981
rect 670804 231976 671955 231978
rect 670804 231920 671894 231976
rect 671950 231920 671955 231976
rect 670804 231918 671955 231920
rect 670804 231916 670810 231918
rect 671889 231915 671955 231918
rect 42425 231842 42491 231845
rect 44357 231842 44423 231845
rect 42425 231840 44423 231842
rect 42425 231784 42430 231840
rect 42486 231784 44362 231840
rect 44418 231784 44423 231840
rect 42425 231782 44423 231784
rect 42425 231779 42491 231782
rect 44357 231779 44423 231782
rect 668301 231162 668367 231165
rect 45510 231160 668367 231162
rect 45510 231104 668306 231160
rect 668362 231104 668367 231160
rect 45510 231102 668367 231104
rect 43989 231026 44055 231029
rect 45510 231026 45570 231102
rect 668301 231099 668367 231102
rect 43989 231024 45570 231026
rect 43989 230968 43994 231024
rect 44050 230968 45570 231024
rect 43989 230966 45570 230968
rect 43989 230963 44055 230966
rect 144637 230482 144703 230485
rect 151077 230482 151143 230485
rect 144637 230480 151143 230482
rect 144637 230424 144642 230480
rect 144698 230424 151082 230480
rect 151138 230424 151143 230480
rect 144637 230422 151143 230424
rect 144637 230419 144703 230422
rect 151077 230419 151143 230422
rect 665817 230482 665883 230485
rect 674097 230482 674163 230485
rect 665817 230480 674163 230482
rect 665817 230424 665822 230480
rect 665878 230424 674102 230480
rect 674158 230424 674163 230480
rect 665817 230422 674163 230424
rect 665817 230419 665883 230422
rect 674097 230419 674163 230422
rect 150341 230210 150407 230213
rect 151905 230210 151971 230213
rect 150341 230208 151971 230210
rect 150341 230152 150346 230208
rect 150402 230152 151910 230208
rect 151966 230152 151971 230208
rect 150341 230150 151971 230152
rect 150341 230147 150407 230150
rect 151905 230147 151971 230150
rect 666001 230210 666067 230213
rect 673269 230210 673335 230213
rect 676581 230210 676647 230213
rect 666001 230208 673335 230210
rect 666001 230152 666006 230208
rect 666062 230152 673274 230208
rect 673330 230152 673335 230208
rect 666001 230150 673335 230152
rect 666001 230147 666067 230150
rect 673269 230147 673335 230150
rect 674974 230208 676647 230210
rect 674974 230152 676586 230208
rect 676642 230152 676647 230208
rect 674974 230150 676647 230152
rect 185393 229938 185459 229941
rect 186037 229938 186103 229941
rect 185393 229936 186103 229938
rect 185393 229880 185398 229936
rect 185454 229880 186042 229936
rect 186098 229880 186103 229936
rect 185393 229878 186103 229880
rect 185393 229875 185459 229878
rect 186037 229875 186103 229878
rect 144453 229802 144519 229805
rect 150525 229802 150591 229805
rect 144453 229800 150591 229802
rect 144453 229744 144458 229800
rect 144514 229744 150530 229800
rect 150586 229744 150591 229800
rect 144453 229742 150591 229744
rect 144453 229739 144519 229742
rect 150525 229739 150591 229742
rect 154021 229802 154087 229805
rect 160829 229802 160895 229805
rect 154021 229800 160895 229802
rect 154021 229744 154026 229800
rect 154082 229744 160834 229800
rect 160890 229744 160895 229800
rect 154021 229742 160895 229744
rect 154021 229739 154087 229742
rect 160829 229739 160895 229742
rect 663885 229802 663951 229805
rect 673453 229802 673519 229805
rect 663885 229800 673519 229802
rect 663885 229744 663890 229800
rect 663946 229744 673458 229800
rect 673514 229744 673519 229800
rect 663885 229742 673519 229744
rect 663885 229739 663951 229742
rect 673453 229739 673519 229742
rect 674097 229802 674163 229805
rect 674974 229802 675034 230150
rect 676581 230147 676647 230150
rect 674097 229800 675034 229802
rect 674097 229744 674102 229800
rect 674158 229744 675034 229800
rect 674097 229742 675034 229744
rect 674097 229739 674163 229742
rect 42425 229394 42491 229397
rect 43621 229394 43687 229397
rect 42425 229392 43687 229394
rect 42425 229336 42430 229392
rect 42486 229336 43626 229392
rect 43682 229336 43687 229392
rect 42425 229334 43687 229336
rect 42425 229331 42491 229334
rect 43621 229331 43687 229334
rect 145833 229394 145899 229397
rect 147949 229394 148015 229397
rect 145833 229392 148015 229394
rect 145833 229336 145838 229392
rect 145894 229336 147954 229392
rect 148010 229336 148015 229392
rect 145833 229334 148015 229336
rect 145833 229331 145899 229334
rect 147949 229331 148015 229334
rect 161289 229394 161355 229397
rect 161749 229394 161815 229397
rect 161289 229392 161815 229394
rect 161289 229336 161294 229392
rect 161350 229336 161754 229392
rect 161810 229336 161815 229392
rect 161289 229334 161815 229336
rect 161289 229331 161355 229334
rect 161749 229331 161815 229334
rect 151629 229258 151695 229261
rect 153653 229258 153719 229261
rect 151629 229256 153719 229258
rect 151629 229200 151634 229256
rect 151690 229200 153658 229256
rect 153714 229200 153719 229256
rect 151629 229198 153719 229200
rect 151629 229195 151695 229198
rect 153653 229195 153719 229198
rect 140037 229122 140103 229125
rect 143533 229122 143599 229125
rect 140037 229120 143599 229122
rect 140037 229064 140042 229120
rect 140098 229064 143538 229120
rect 143594 229064 143599 229120
rect 140037 229062 143599 229064
rect 140037 229059 140103 229062
rect 143533 229059 143599 229062
rect 41965 228988 42031 228989
rect 41965 228984 42012 228988
rect 42076 228986 42082 228988
rect 193029 228986 193095 228989
rect 195421 228986 195487 228989
rect 41965 228928 41970 228984
rect 41965 228924 42012 228928
rect 42076 228926 42122 228986
rect 193029 228984 195487 228986
rect 193029 228928 193034 228984
rect 193090 228928 195426 228984
rect 195482 228928 195487 228984
rect 193029 228926 195487 228928
rect 42076 228924 42082 228926
rect 41965 228923 42031 228924
rect 193029 228923 193095 228926
rect 195421 228923 195487 228926
rect 161427 228850 161493 228853
rect 164233 228850 164299 228853
rect 161427 228848 164299 228850
rect 161427 228792 161432 228848
rect 161488 228792 164238 228848
rect 164294 228792 164299 228848
rect 161427 228790 164299 228792
rect 161427 228787 161493 228790
rect 164233 228787 164299 228790
rect 173157 228850 173223 228853
rect 176101 228850 176167 228853
rect 173157 228848 176167 228850
rect 173157 228792 173162 228848
rect 173218 228792 176106 228848
rect 176162 228792 176167 228848
rect 173157 228790 176167 228792
rect 173157 228787 173223 228790
rect 176101 228787 176167 228790
rect 652201 228578 652267 228581
rect 675477 228580 675543 228581
rect 674230 228578 674236 228580
rect 652201 228576 674236 228578
rect 652201 228520 652206 228576
rect 652262 228520 674236 228576
rect 652201 228518 674236 228520
rect 652201 228515 652267 228518
rect 674230 228516 674236 228518
rect 674300 228516 674306 228580
rect 675477 228578 675524 228580
rect 675432 228576 675524 228578
rect 675432 228520 675482 228576
rect 675432 228518 675524 228520
rect 675477 228516 675524 228518
rect 675588 228516 675594 228580
rect 675477 228515 675543 228516
rect 153101 228442 153167 228445
rect 154389 228442 154455 228445
rect 153101 228440 154455 228442
rect 153101 228384 153106 228440
rect 153162 228384 154394 228440
rect 154450 228384 154455 228440
rect 153101 228382 154455 228384
rect 153101 228379 153167 228382
rect 154389 228379 154455 228382
rect 160001 228442 160067 228445
rect 161565 228442 161631 228445
rect 160001 228440 161631 228442
rect 160001 228384 160006 228440
rect 160062 228384 161570 228440
rect 161626 228384 161631 228440
rect 160001 228382 161631 228384
rect 160001 228379 160067 228382
rect 161565 228379 161631 228382
rect 146201 228034 146267 228037
rect 147121 228034 147187 228037
rect 146201 228032 147187 228034
rect 146201 227976 146206 228032
rect 146262 227976 147126 228032
rect 147182 227976 147187 228032
rect 146201 227974 147187 227976
rect 146201 227971 146267 227974
rect 147121 227971 147187 227974
rect 136633 227898 136699 227901
rect 141509 227898 141575 227901
rect 136633 227896 141575 227898
rect 136633 227840 136638 227896
rect 136694 227840 141514 227896
rect 141570 227840 141575 227896
rect 136633 227838 141575 227840
rect 136633 227835 136699 227838
rect 141509 227835 141575 227838
rect 175365 227626 175431 227629
rect 177205 227626 177271 227629
rect 175365 227624 177271 227626
rect 175365 227568 175370 227624
rect 175426 227568 177210 227624
rect 177266 227568 177271 227624
rect 175365 227566 177271 227568
rect 175365 227563 175431 227566
rect 177205 227563 177271 227566
rect 170765 227490 170831 227493
rect 171685 227490 171751 227493
rect 170765 227488 171751 227490
rect 170765 227432 170770 227488
rect 170826 227432 171690 227488
rect 171746 227432 171751 227488
rect 170765 227430 171751 227432
rect 170765 227427 170831 227430
rect 171685 227427 171751 227430
rect 161427 227354 161493 227357
rect 166901 227354 166967 227357
rect 161427 227352 166967 227354
rect 161427 227296 161432 227352
rect 161488 227296 166906 227352
rect 166962 227296 166967 227352
rect 161427 227294 166967 227296
rect 161427 227291 161493 227294
rect 166901 227291 166967 227294
rect 175917 227354 175983 227357
rect 176745 227354 176811 227357
rect 175917 227352 176811 227354
rect 175917 227296 175922 227352
rect 175978 227296 176750 227352
rect 176806 227296 176811 227352
rect 175917 227294 176811 227296
rect 175917 227291 175983 227294
rect 176745 227291 176811 227294
rect 169569 227218 169635 227221
rect 171087 227218 171153 227221
rect 169569 227216 171153 227218
rect 169569 227160 169574 227216
rect 169630 227160 171092 227216
rect 171148 227160 171153 227216
rect 169569 227158 171153 227160
rect 169569 227155 169635 227158
rect 171087 227155 171153 227158
rect 155861 227082 155927 227085
rect 161565 227082 161631 227085
rect 672625 227084 672691 227085
rect 672574 227082 672580 227084
rect 155861 227080 161631 227082
rect 155861 227024 155866 227080
rect 155922 227024 161570 227080
rect 161626 227024 161631 227080
rect 155861 227022 161631 227024
rect 672534 227022 672580 227082
rect 672644 227080 672691 227084
rect 672686 227024 672691 227080
rect 155861 227019 155927 227022
rect 161565 227019 161631 227022
rect 672574 227020 672580 227022
rect 672644 227020 672691 227024
rect 672625 227019 672691 227020
rect 674097 227082 674163 227085
rect 676397 227082 676463 227085
rect 674097 227080 676463 227082
rect 674097 227024 674102 227080
rect 674158 227024 676402 227080
rect 676458 227024 676463 227080
rect 674097 227022 676463 227024
rect 674097 227019 674163 227022
rect 676397 227019 676463 227022
rect 683205 227082 683271 227085
rect 683798 227082 683804 227084
rect 683205 227080 683804 227082
rect 683205 227024 683210 227080
rect 683266 227024 683804 227080
rect 683205 227022 683804 227024
rect 683205 227019 683271 227022
rect 683798 227020 683804 227022
rect 683868 227020 683874 227084
rect 652569 226946 652635 226949
rect 652569 226944 663810 226946
rect 652569 226888 652574 226944
rect 652630 226888 663810 226944
rect 652569 226886 663810 226888
rect 652569 226883 652635 226886
rect 663750 226810 663810 226886
rect 673545 226810 673611 226813
rect 676949 226810 677015 226813
rect 663750 226750 673010 226810
rect 42149 226674 42215 226677
rect 44541 226674 44607 226677
rect 42149 226672 44607 226674
rect 42149 226616 42154 226672
rect 42210 226616 44546 226672
rect 44602 226616 44607 226672
rect 42149 226614 44607 226616
rect 42149 226611 42215 226614
rect 44541 226611 44607 226614
rect 141601 226538 141667 226541
rect 142245 226538 142311 226541
rect 141601 226536 142311 226538
rect 141601 226480 141606 226536
rect 141662 226480 142250 226536
rect 142306 226480 142311 226536
rect 141601 226478 142311 226480
rect 672950 226538 673010 226750
rect 673545 226808 677015 226810
rect 673545 226752 673550 226808
rect 673606 226752 676954 226808
rect 677010 226752 677015 226808
rect 673545 226750 677015 226752
rect 673545 226747 673611 226750
rect 676949 226747 677015 226750
rect 674046 226538 674052 226540
rect 672950 226478 674052 226538
rect 141601 226475 141667 226478
rect 142245 226475 142311 226478
rect 674046 226476 674052 226478
rect 674116 226476 674122 226540
rect 653581 226402 653647 226405
rect 672717 226402 672783 226405
rect 653581 226400 672783 226402
rect 653581 226344 653586 226400
rect 653642 226344 672722 226400
rect 672778 226344 672783 226400
rect 653581 226342 672783 226344
rect 653581 226339 653647 226342
rect 672717 226339 672783 226342
rect 672597 226130 672663 226133
rect 674833 226130 674899 226133
rect 672597 226128 674899 226130
rect 672597 226072 672602 226128
rect 672658 226072 674838 226128
rect 674894 226072 674899 226128
rect 672597 226070 674899 226072
rect 672597 226067 672663 226070
rect 674833 226067 674899 226070
rect 148869 225994 148935 225997
rect 151905 225994 151971 225997
rect 148869 225992 151971 225994
rect 148869 225936 148874 225992
rect 148930 225936 151910 225992
rect 151966 225936 151971 225992
rect 148869 225934 151971 225936
rect 148869 225931 148935 225934
rect 151905 225931 151971 225934
rect 664437 225858 664503 225861
rect 672257 225858 672323 225861
rect 664437 225856 672323 225858
rect 664437 225800 664442 225856
rect 664498 225800 672262 225856
rect 672318 225800 672323 225856
rect 664437 225798 672323 225800
rect 664437 225795 664503 225798
rect 672257 225795 672323 225798
rect 42425 225722 42491 225725
rect 45921 225722 45987 225725
rect 42425 225720 45987 225722
rect 42425 225664 42430 225720
rect 42486 225664 45926 225720
rect 45982 225664 45987 225720
rect 42425 225662 45987 225664
rect 42425 225659 42491 225662
rect 45921 225659 45987 225662
rect 151721 225722 151787 225725
rect 157517 225722 157583 225725
rect 151721 225720 157583 225722
rect 151721 225664 151726 225720
rect 151782 225664 157522 225720
rect 157578 225664 157583 225720
rect 151721 225662 157583 225664
rect 151721 225659 151787 225662
rect 157517 225659 157583 225662
rect 672373 225722 672439 225725
rect 675477 225722 675543 225725
rect 672373 225720 675543 225722
rect 672373 225664 672378 225720
rect 672434 225664 675482 225720
rect 675538 225664 675543 225720
rect 672373 225662 675543 225664
rect 672373 225659 672439 225662
rect 675477 225659 675543 225662
rect 142107 225586 142173 225589
rect 147765 225586 147831 225589
rect 142107 225584 147831 225586
rect 142107 225528 142112 225584
rect 142168 225528 147770 225584
rect 147826 225528 147831 225584
rect 142107 225526 147831 225528
rect 142107 225523 142173 225526
rect 147765 225523 147831 225526
rect 659101 225586 659167 225589
rect 659101 225584 669330 225586
rect 659101 225528 659106 225584
rect 659162 225528 669330 225584
rect 659101 225526 669330 225528
rect 659101 225523 659167 225526
rect 669270 225314 669330 225526
rect 672149 225450 672215 225453
rect 675845 225450 675911 225453
rect 672149 225448 675911 225450
rect 672149 225392 672154 225448
rect 672210 225392 675850 225448
rect 675906 225392 675911 225448
rect 672149 225390 675911 225392
rect 672149 225387 672215 225390
rect 675845 225387 675911 225390
rect 672027 225314 672093 225317
rect 669270 225312 672093 225314
rect 669270 225256 672032 225312
rect 672088 225256 672093 225312
rect 669270 225254 672093 225256
rect 672027 225251 672093 225254
rect 654777 225042 654843 225045
rect 672441 225042 672507 225045
rect 654777 225040 672507 225042
rect 654777 224984 654782 225040
rect 654838 224984 672446 225040
rect 672502 224984 672507 225040
rect 654777 224982 672507 224984
rect 654777 224979 654843 224982
rect 672441 224979 672507 224982
rect 179321 224906 179387 224909
rect 181989 224906 182055 224909
rect 179321 224904 182055 224906
rect 179321 224848 179326 224904
rect 179382 224848 181994 224904
rect 182050 224848 182055 224904
rect 179321 224846 182055 224848
rect 179321 224843 179387 224846
rect 181989 224843 182055 224846
rect 557625 224770 557691 224773
rect 561949 224770 562015 224773
rect 557625 224768 562015 224770
rect 557625 224712 557630 224768
rect 557686 224712 561954 224768
rect 562010 224712 562015 224768
rect 557625 224710 562015 224712
rect 557625 224707 557691 224710
rect 561949 224707 562015 224710
rect 562133 224770 562199 224773
rect 563697 224770 563763 224773
rect 562133 224768 563763 224770
rect 562133 224712 562138 224768
rect 562194 224712 563702 224768
rect 563758 224712 563763 224768
rect 562133 224710 563763 224712
rect 562133 224707 562199 224710
rect 563697 224707 563763 224710
rect 671813 224770 671879 224773
rect 673545 224770 673611 224773
rect 671813 224768 673611 224770
rect 671813 224712 671818 224768
rect 671874 224712 673550 224768
rect 673606 224712 673611 224768
rect 671813 224710 673611 224712
rect 671813 224707 671879 224710
rect 673545 224707 673611 224710
rect 669998 224572 670004 224636
rect 670068 224634 670074 224636
rect 670325 224634 670391 224637
rect 670068 224632 670391 224634
rect 670068 224576 670330 224632
rect 670386 224576 670391 224632
rect 670068 224574 670391 224576
rect 670068 224572 670074 224574
rect 670325 224571 670391 224574
rect 41689 224498 41755 224501
rect 63217 224498 63283 224501
rect 41689 224496 63283 224498
rect 41689 224440 41694 224496
rect 41750 224440 63222 224496
rect 63278 224440 63283 224496
rect 41689 224438 63283 224440
rect 41689 224435 41755 224438
rect 63217 224435 63283 224438
rect 151629 224498 151695 224501
rect 152365 224498 152431 224501
rect 151629 224496 152431 224498
rect 151629 224440 151634 224496
rect 151690 224440 152370 224496
rect 152426 224440 152431 224496
rect 151629 224438 152431 224440
rect 151629 224435 151695 224438
rect 152365 224435 152431 224438
rect 543733 224498 543799 224501
rect 544285 224498 544351 224501
rect 543733 224496 544351 224498
rect 543733 224440 543738 224496
rect 543794 224440 544290 224496
rect 544346 224440 544351 224496
rect 543733 224438 544351 224440
rect 543733 224435 543799 224438
rect 544285 224435 544351 224438
rect 554865 224498 554931 224501
rect 556061 224498 556127 224501
rect 557625 224498 557691 224501
rect 554865 224496 557691 224498
rect 554865 224440 554870 224496
rect 554926 224440 556066 224496
rect 556122 224440 557630 224496
rect 557686 224440 557691 224496
rect 554865 224438 557691 224440
rect 554865 224435 554931 224438
rect 556061 224435 556127 224438
rect 557625 224435 557691 224438
rect 671521 224364 671587 224365
rect 671470 224362 671476 224364
rect 671430 224302 671476 224362
rect 671540 224360 671587 224364
rect 671582 224304 671587 224360
rect 671470 224300 671476 224302
rect 671540 224300 671587 224304
rect 671521 224299 671587 224300
rect 62665 224226 62731 224229
rect 591481 224226 591547 224229
rect 667749 224226 667815 224229
rect 62665 224224 591547 224226
rect 62665 224168 62670 224224
rect 62726 224168 591486 224224
rect 591542 224168 591547 224224
rect 62665 224166 591547 224168
rect 62665 224163 62731 224166
rect 591481 224163 591547 224166
rect 663750 224224 667815 224226
rect 663750 224168 667754 224224
rect 667810 224168 667815 224224
rect 663750 224166 667815 224168
rect 137277 223954 137343 223957
rect 142245 223954 142311 223957
rect 137277 223952 142311 223954
rect 137277 223896 137282 223952
rect 137338 223896 142250 223952
rect 142306 223896 142311 223952
rect 137277 223894 142311 223896
rect 137277 223891 137343 223894
rect 142245 223891 142311 223894
rect 142429 223954 142495 223957
rect 151629 223954 151695 223957
rect 142429 223952 151695 223954
rect 142429 223896 142434 223952
rect 142490 223896 151634 223952
rect 151690 223896 151695 223952
rect 142429 223894 151695 223896
rect 142429 223891 142495 223894
rect 151629 223891 151695 223894
rect 656157 223954 656223 223957
rect 663750 223954 663810 224166
rect 667749 224163 667815 224166
rect 656157 223952 663810 223954
rect 656157 223896 656162 223952
rect 656218 223896 663810 223952
rect 656157 223894 663810 223896
rect 670509 223956 670575 223957
rect 670509 223952 670556 223956
rect 670620 223954 670626 223956
rect 671475 223954 671541 223957
rect 672073 223954 672139 223957
rect 670509 223896 670514 223952
rect 656157 223891 656223 223894
rect 670509 223892 670556 223896
rect 670620 223894 670666 223954
rect 671475 223952 672139 223954
rect 671475 223896 671480 223952
rect 671536 223896 672078 223952
rect 672134 223896 672139 223952
rect 671475 223894 672139 223896
rect 670620 223892 670626 223894
rect 670509 223891 670575 223892
rect 671475 223891 671541 223894
rect 672073 223891 672139 223894
rect 683798 223756 683804 223820
rect 683868 223756 683874 223820
rect 657537 223682 657603 223685
rect 667013 223682 667079 223685
rect 670417 223684 670483 223685
rect 671521 223684 671587 223685
rect 670366 223682 670372 223684
rect 657537 223680 667079 223682
rect 657537 223624 657542 223680
rect 657598 223624 667018 223680
rect 667074 223624 667079 223680
rect 657537 223622 667079 223624
rect 670326 223622 670372 223682
rect 670436 223680 670483 223684
rect 670478 223624 670483 223680
rect 657537 223619 657603 223622
rect 667013 223619 667079 223622
rect 670366 223620 670372 223622
rect 670436 223620 670483 223624
rect 671470 223620 671476 223684
rect 671540 223682 671587 223684
rect 672625 223682 672691 223685
rect 673361 223682 673427 223685
rect 671540 223680 671632 223682
rect 671582 223624 671632 223680
rect 671540 223622 671632 223624
rect 672625 223680 673427 223682
rect 672625 223624 672630 223680
rect 672686 223624 673366 223680
rect 673422 223624 673427 223680
rect 672625 223622 673427 223624
rect 671540 223620 671587 223622
rect 670417 223619 670483 223620
rect 671521 223619 671587 223620
rect 672625 223619 672691 223622
rect 673361 223619 673427 223622
rect 42149 223546 42215 223549
rect 51717 223546 51783 223549
rect 42149 223544 51783 223546
rect 42149 223488 42154 223544
rect 42210 223488 51722 223544
rect 51778 223488 51783 223544
rect 42149 223486 51783 223488
rect 42149 223483 42215 223486
rect 51717 223483 51783 223486
rect 62849 223546 62915 223549
rect 62849 223544 582390 223546
rect 62849 223488 62854 223544
rect 62910 223488 582390 223544
rect 683806 223516 683866 223756
rect 62849 223486 582390 223488
rect 62849 223483 62915 223486
rect 582330 223410 582390 223486
rect 591982 223410 591988 223412
rect 582330 223350 591988 223410
rect 591982 223348 591988 223350
rect 592052 223348 592058 223412
rect 676029 223138 676095 223141
rect 676029 223136 676292 223138
rect 676029 223080 676034 223136
rect 676090 223080 676292 223136
rect 676029 223078 676292 223080
rect 676029 223075 676095 223078
rect 141969 222866 142035 222869
rect 142153 222866 142219 222869
rect 141969 222864 142219 222866
rect 141969 222808 141974 222864
rect 142030 222808 142158 222864
rect 142214 222808 142219 222864
rect 141969 222806 142219 222808
rect 141969 222803 142035 222806
rect 142153 222803 142219 222806
rect 653397 222866 653463 222869
rect 673085 222866 673151 222869
rect 653397 222864 673151 222866
rect 653397 222808 653402 222864
rect 653458 222808 673090 222864
rect 673146 222808 673151 222864
rect 653397 222806 673151 222808
rect 653397 222803 653463 222806
rect 673085 222803 673151 222806
rect 683389 222730 683455 222733
rect 683389 222728 683468 222730
rect 683389 222672 683394 222728
rect 683450 222672 683468 222728
rect 683389 222670 683468 222672
rect 683389 222667 683455 222670
rect 649574 222396 649580 222460
rect 649644 222458 649650 222460
rect 651966 222458 651972 222460
rect 649644 222398 651972 222458
rect 649644 222396 649650 222398
rect 651966 222396 651972 222398
rect 652036 222396 652042 222460
rect 658917 222322 658983 222325
rect 667013 222322 667079 222325
rect 658917 222320 667079 222322
rect 658917 222264 658922 222320
rect 658978 222264 667018 222320
rect 667074 222264 667079 222320
rect 658917 222262 667079 222264
rect 658917 222259 658983 222262
rect 667013 222259 667079 222262
rect 674005 222322 674071 222325
rect 674005 222320 676292 222322
rect 674005 222264 674010 222320
rect 674066 222264 676292 222320
rect 674005 222262 676292 222264
rect 674005 222259 674071 222262
rect 140773 222050 140839 222053
rect 141969 222050 142035 222053
rect 140773 222048 142035 222050
rect 140773 221992 140778 222048
rect 140834 221992 141974 222048
rect 142030 221992 142035 222048
rect 140773 221990 142035 221992
rect 140773 221987 140839 221990
rect 141969 221987 142035 221990
rect 533245 222050 533311 222053
rect 538489 222050 538555 222053
rect 533245 222048 538555 222050
rect 533245 221992 533250 222048
rect 533306 221992 538494 222048
rect 538550 221992 538555 222048
rect 533245 221990 538555 221992
rect 533245 221987 533311 221990
rect 538489 221987 538555 221990
rect 556797 222050 556863 222053
rect 557533 222050 557599 222053
rect 556797 222048 557599 222050
rect 556797 221992 556802 222048
rect 556858 221992 557538 222048
rect 557594 221992 557599 222048
rect 556797 221990 557599 221992
rect 556797 221987 556863 221990
rect 557533 221987 557599 221990
rect 559373 222050 559439 222053
rect 561489 222050 561555 222053
rect 559373 222048 561555 222050
rect 559373 221992 559378 222048
rect 559434 221992 561494 222048
rect 561550 221992 561555 222048
rect 559373 221990 561555 221992
rect 559373 221987 559439 221990
rect 561489 221987 561555 221990
rect 176285 221914 176351 221917
rect 177389 221914 177455 221917
rect 176285 221912 177455 221914
rect 176285 221856 176290 221912
rect 176346 221856 177394 221912
rect 177450 221856 177455 221912
rect 176285 221854 177455 221856
rect 176285 221851 176351 221854
rect 177389 221851 177455 221854
rect 676029 221914 676095 221917
rect 676029 221912 676292 221914
rect 676029 221856 676034 221912
rect 676090 221856 676292 221912
rect 676029 221854 676292 221856
rect 676029 221851 676095 221854
rect 161427 221778 161493 221781
rect 166993 221778 167059 221781
rect 161427 221776 167059 221778
rect 161427 221720 161432 221776
rect 161488 221720 166998 221776
rect 167054 221720 167059 221776
rect 161427 221718 167059 221720
rect 161427 221715 161493 221718
rect 166993 221715 167059 221718
rect 535729 221778 535795 221781
rect 538673 221778 538739 221781
rect 535729 221776 538739 221778
rect 535729 221720 535734 221776
rect 535790 221720 538678 221776
rect 538734 221720 538739 221776
rect 535729 221718 538739 221720
rect 535729 221715 535795 221718
rect 538673 221715 538739 221718
rect 545757 221778 545823 221781
rect 549253 221778 549319 221781
rect 545757 221776 549319 221778
rect 545757 221720 545762 221776
rect 545818 221720 549258 221776
rect 549314 221720 549319 221776
rect 545757 221718 549319 221720
rect 545757 221715 545823 221718
rect 549253 221715 549319 221718
rect 553301 221778 553367 221781
rect 557165 221778 557231 221781
rect 553301 221776 557231 221778
rect 553301 221720 553306 221776
rect 553362 221720 557170 221776
rect 557226 221720 557231 221776
rect 553301 221718 557231 221720
rect 553301 221715 553367 221718
rect 557165 221715 557231 221718
rect 563697 221778 563763 221781
rect 572621 221778 572687 221781
rect 563697 221776 572687 221778
rect 563697 221720 563702 221776
rect 563758 221720 572626 221776
rect 572682 221720 572687 221776
rect 563697 221718 572687 221720
rect 563697 221715 563763 221718
rect 572621 221715 572687 221718
rect 651465 221778 651531 221781
rect 668485 221778 668551 221781
rect 651465 221776 668551 221778
rect 651465 221720 651470 221776
rect 651526 221720 668490 221776
rect 668546 221720 668551 221776
rect 651465 221718 668551 221720
rect 651465 221715 651531 221718
rect 668485 221715 668551 221718
rect 671889 221778 671955 221781
rect 675661 221778 675727 221781
rect 671889 221776 675727 221778
rect 671889 221720 671894 221776
rect 671950 221720 675666 221776
rect 675722 221720 675727 221776
rect 671889 221718 675727 221720
rect 671889 221715 671955 221718
rect 675661 221715 675727 221718
rect 138289 221642 138355 221645
rect 141325 221642 141391 221645
rect 138289 221640 141391 221642
rect 138289 221584 138294 221640
rect 138350 221584 141330 221640
rect 141386 221584 141391 221640
rect 138289 221582 141391 221584
rect 138289 221579 138355 221582
rect 141325 221579 141391 221582
rect 171409 221506 171475 221509
rect 171961 221506 172027 221509
rect 171409 221504 172027 221506
rect 171409 221448 171414 221504
rect 171470 221448 171966 221504
rect 172022 221448 172027 221504
rect 171409 221446 172027 221448
rect 171409 221443 171475 221446
rect 171961 221443 172027 221446
rect 513557 221506 513623 221509
rect 599485 221506 599551 221509
rect 513557 221504 599551 221506
rect 513557 221448 513562 221504
rect 513618 221448 599490 221504
rect 599546 221448 599551 221504
rect 513557 221446 599551 221448
rect 513557 221443 513623 221446
rect 599485 221443 599551 221446
rect 649809 221506 649875 221509
rect 674833 221506 674899 221509
rect 649809 221504 674899 221506
rect 649809 221448 649814 221504
rect 649870 221448 674838 221504
rect 674894 221448 674899 221504
rect 649809 221446 674899 221448
rect 649809 221443 649875 221446
rect 674833 221443 674899 221446
rect 675017 221506 675083 221509
rect 675017 221504 676292 221506
rect 675017 221448 675022 221504
rect 675078 221448 676292 221504
rect 675017 221446 676292 221448
rect 675017 221443 675083 221446
rect 145557 221234 145623 221237
rect 146385 221234 146451 221237
rect 145557 221232 146451 221234
rect 145557 221176 145562 221232
rect 145618 221176 146390 221232
rect 146446 221176 146451 221232
rect 145557 221174 146451 221176
rect 145557 221171 145623 221174
rect 146385 221171 146451 221174
rect 515765 221234 515831 221237
rect 600865 221234 600931 221237
rect 515765 221232 600931 221234
rect 515765 221176 515770 221232
rect 515826 221176 600870 221232
rect 600926 221176 600931 221232
rect 515765 221174 600931 221176
rect 515765 221171 515831 221174
rect 600865 221171 600931 221174
rect 673177 221098 673243 221101
rect 673177 221096 676292 221098
rect 673177 221040 673182 221096
rect 673238 221040 676292 221096
rect 673177 221038 676292 221040
rect 673177 221035 673243 221038
rect 142107 220962 142173 220965
rect 151169 220962 151235 220965
rect 142107 220960 151235 220962
rect 142107 220904 142112 220960
rect 142168 220904 151174 220960
rect 151230 220904 151235 220960
rect 142107 220902 151235 220904
rect 142107 220899 142173 220902
rect 151169 220899 151235 220902
rect 158345 220962 158411 220965
rect 161565 220962 161631 220965
rect 158345 220960 161631 220962
rect 158345 220904 158350 220960
rect 158406 220904 161570 220960
rect 161626 220904 161631 220960
rect 158345 220902 161631 220904
rect 158345 220899 158411 220902
rect 161565 220899 161631 220902
rect 522665 220962 522731 220965
rect 618253 220962 618319 220965
rect 522665 220960 618319 220962
rect 522665 220904 522670 220960
rect 522726 220904 618258 220960
rect 618314 220904 618319 220960
rect 522665 220902 618319 220904
rect 522665 220899 522731 220902
rect 618253 220899 618319 220902
rect 177205 220826 177271 220829
rect 185117 220826 185183 220829
rect 177205 220824 185183 220826
rect 177205 220768 177210 220824
rect 177266 220768 185122 220824
rect 185178 220768 185183 220824
rect 177205 220766 185183 220768
rect 177205 220763 177271 220766
rect 185117 220763 185183 220766
rect 185945 220826 186011 220829
rect 190545 220826 190611 220829
rect 185945 220824 190611 220826
rect 185945 220768 185950 220824
rect 186006 220768 190550 220824
rect 190606 220768 190611 220824
rect 185945 220766 190611 220768
rect 185945 220763 186011 220766
rect 190545 220763 190611 220766
rect 654133 220826 654199 220829
rect 667749 220826 667815 220829
rect 670049 220828 670115 220829
rect 654133 220824 667815 220826
rect 654133 220768 654138 220824
rect 654194 220768 667754 220824
rect 667810 220768 667815 220824
rect 654133 220766 667815 220768
rect 654133 220763 654199 220766
rect 667749 220763 667815 220766
rect 669998 220764 670004 220828
rect 670068 220826 670115 220828
rect 670068 220824 670160 220826
rect 670110 220768 670160 220824
rect 670068 220766 670160 220768
rect 670068 220764 670115 220766
rect 670049 220763 670115 220764
rect 563053 220690 563119 220693
rect 563010 220688 563119 220690
rect 563010 220632 563058 220688
rect 563114 220632 563119 220688
rect 563010 220627 563119 220632
rect 582373 220690 582439 220693
rect 587525 220690 587591 220693
rect 582373 220688 587591 220690
rect 582373 220632 582378 220688
rect 582434 220632 587530 220688
rect 587586 220632 587591 220688
rect 582373 220630 587591 220632
rect 582373 220627 582439 220630
rect 587525 220627 587591 220630
rect 672901 220690 672967 220693
rect 672901 220688 676292 220690
rect 672901 220632 672906 220688
rect 672962 220632 676292 220688
rect 672901 220630 676292 220632
rect 672901 220627 672967 220630
rect 561765 220554 561831 220557
rect 563010 220554 563070 220627
rect 561765 220552 563070 220554
rect 561765 220496 561770 220552
rect 561826 220496 563070 220552
rect 561765 220494 563070 220496
rect 565629 220554 565695 220557
rect 574737 220554 574803 220557
rect 565629 220552 574803 220554
rect 565629 220496 565634 220552
rect 565690 220496 574742 220552
rect 574798 220496 574803 220552
rect 565629 220494 574803 220496
rect 561765 220491 561831 220494
rect 565629 220491 565695 220494
rect 574737 220491 574803 220494
rect 145649 220418 145715 220421
rect 148317 220418 148383 220421
rect 145649 220416 148383 220418
rect 145649 220360 145654 220416
rect 145710 220360 148322 220416
rect 148378 220360 148383 220416
rect 145649 220358 148383 220360
rect 145649 220355 145715 220358
rect 148317 220355 148383 220358
rect 670325 220418 670391 220421
rect 670550 220418 670556 220420
rect 670325 220416 670556 220418
rect 670325 220360 670330 220416
rect 670386 220360 670556 220416
rect 670325 220358 670556 220360
rect 670325 220355 670391 220358
rect 670550 220356 670556 220358
rect 670620 220356 670626 220420
rect 486969 220282 487035 220285
rect 611629 220282 611695 220285
rect 486969 220280 611695 220282
rect 486969 220224 486974 220280
rect 487030 220224 611634 220280
rect 611690 220224 611695 220280
rect 486969 220222 611695 220224
rect 486969 220219 487035 220222
rect 611629 220219 611695 220222
rect 673361 220282 673427 220285
rect 673361 220280 676292 220282
rect 673361 220224 673366 220280
rect 673422 220224 676292 220280
rect 673361 220222 676292 220224
rect 673361 220219 673427 220222
rect 515121 220010 515187 220013
rect 617149 220010 617215 220013
rect 515121 220008 617215 220010
rect 515121 219952 515126 220008
rect 515182 219952 617154 220008
rect 617210 219952 617215 220008
rect 515121 219950 617215 219952
rect 515121 219947 515187 219950
rect 617149 219947 617215 219950
rect 646037 219874 646103 219877
rect 675477 219874 675543 219877
rect 646037 219872 675543 219874
rect 646037 219816 646042 219872
rect 646098 219816 675482 219872
rect 675538 219816 675543 219872
rect 646037 219814 675543 219816
rect 646037 219811 646103 219814
rect 675477 219811 675543 219814
rect 676024 219812 676030 219876
rect 676094 219874 676100 219876
rect 676094 219814 676292 219874
rect 676094 219812 676100 219814
rect 492949 219738 493015 219741
rect 493685 219738 493751 219741
rect 612733 219738 612799 219741
rect 492949 219736 612799 219738
rect 492949 219680 492954 219736
rect 493010 219680 493690 219736
rect 493746 219680 612738 219736
rect 612794 219680 612799 219736
rect 492949 219678 612799 219680
rect 492949 219675 493015 219678
rect 493685 219675 493751 219678
rect 612733 219675 612799 219678
rect 168925 219466 168991 219469
rect 169753 219466 169819 219469
rect 168925 219464 169819 219466
rect 168925 219408 168930 219464
rect 168986 219408 169758 219464
rect 169814 219408 169819 219464
rect 168925 219406 169819 219408
rect 168925 219403 168991 219406
rect 169753 219403 169819 219406
rect 520181 219466 520247 219469
rect 618437 219466 618503 219469
rect 520181 219464 618503 219466
rect 520181 219408 520186 219464
rect 520242 219408 618442 219464
rect 618498 219408 618503 219464
rect 520181 219406 618503 219408
rect 520181 219403 520247 219406
rect 618437 219403 618503 219406
rect 667749 219466 667815 219469
rect 667749 219464 676292 219466
rect 667749 219408 667754 219464
rect 667810 219408 676292 219464
rect 667749 219406 676292 219408
rect 667749 219403 667815 219406
rect 194869 219330 194935 219333
rect 197813 219330 197879 219333
rect 194869 219328 197879 219330
rect 194869 219272 194874 219328
rect 194930 219272 197818 219328
rect 197874 219272 197879 219328
rect 194869 219270 197879 219272
rect 194869 219267 194935 219270
rect 197813 219267 197879 219270
rect 562041 219194 562107 219197
rect 562593 219194 562659 219197
rect 562041 219192 562659 219194
rect 562041 219136 562046 219192
rect 562102 219136 562598 219192
rect 562654 219136 562659 219192
rect 562041 219134 562659 219136
rect 562041 219131 562107 219134
rect 562593 219131 562659 219134
rect 564801 219058 564867 219061
rect 572667 219058 572733 219061
rect 564801 219056 572733 219058
rect 564801 219000 564806 219056
rect 564862 219000 572672 219056
rect 572728 219000 572733 219056
rect 564801 218998 572733 219000
rect 564801 218995 564867 218998
rect 572667 218995 572733 218998
rect 674833 219058 674899 219061
rect 674833 219056 676292 219058
rect 674833 219000 674838 219056
rect 674894 219000 676292 219056
rect 674833 218998 676292 219000
rect 674833 218995 674899 218998
rect 656709 218922 656775 218925
rect 666645 218922 666711 218925
rect 562918 218862 564634 218922
rect 180517 218786 180583 218789
rect 182265 218786 182331 218789
rect 180517 218784 182331 218786
rect 180517 218728 180522 218784
rect 180578 218728 182270 218784
rect 182326 218728 182331 218784
rect 180517 218726 182331 218728
rect 180517 218723 180583 218726
rect 182265 218723 182331 218726
rect 561765 218786 561831 218789
rect 562918 218786 562978 218862
rect 561765 218784 562978 218786
rect 561765 218728 561770 218784
rect 561826 218728 562978 218784
rect 561765 218726 562978 218728
rect 564574 218786 564634 218862
rect 656709 218920 666711 218922
rect 656709 218864 656714 218920
rect 656770 218864 666650 218920
rect 666706 218864 666711 218920
rect 656709 218862 666711 218864
rect 656709 218859 656775 218862
rect 666645 218859 666711 218862
rect 566457 218786 566523 218789
rect 564574 218784 566523 218786
rect 564574 218728 566462 218784
rect 566518 218728 566523 218784
rect 564574 218726 566523 218728
rect 561765 218723 561831 218726
rect 566457 218723 566523 218726
rect 563053 218650 563119 218653
rect 564157 218650 564223 218653
rect 563053 218648 564223 218650
rect 563053 218592 563058 218648
rect 563114 218592 564162 218648
rect 564218 218592 564223 218648
rect 563053 218590 564223 218592
rect 563053 218587 563119 218590
rect 564157 218587 564223 218590
rect 572345 218650 572411 218653
rect 574369 218650 574435 218653
rect 572345 218648 574435 218650
rect 572345 218592 572350 218648
rect 572406 218592 574374 218648
rect 574430 218592 574435 218648
rect 572345 218590 574435 218592
rect 572345 218587 572411 218590
rect 574369 218587 574435 218590
rect 648521 218650 648587 218653
rect 671889 218650 671955 218653
rect 648521 218648 671955 218650
rect 648521 218592 648526 218648
rect 648582 218592 671894 218648
rect 671950 218592 671955 218648
rect 648521 218590 671955 218592
rect 648521 218587 648587 218590
rect 671889 218587 671955 218590
rect 675518 218588 675524 218652
rect 675588 218650 675594 218652
rect 675588 218590 676292 218650
rect 675588 218588 675594 218590
rect 171409 218378 171475 218381
rect 171961 218378 172027 218381
rect 171409 218376 172027 218378
rect 171409 218320 171414 218376
rect 171470 218320 171966 218376
rect 172022 218320 172027 218376
rect 171409 218318 172027 218320
rect 171409 218315 171475 218318
rect 171961 218315 172027 218318
rect 494697 218378 494763 218381
rect 630673 218378 630739 218381
rect 494697 218376 630739 218378
rect 494697 218320 494702 218376
rect 494758 218320 630678 218376
rect 630734 218320 630739 218376
rect 494697 218318 630739 218320
rect 494697 218315 494763 218318
rect 630673 218315 630739 218318
rect 675017 218242 675083 218245
rect 675017 218240 676292 218242
rect 675017 218184 675022 218240
rect 675078 218184 676292 218240
rect 675017 218182 676292 218184
rect 675017 218179 675083 218182
rect 487797 218106 487863 218109
rect 623957 218106 624023 218109
rect 487797 218104 624023 218106
rect 487797 218048 487802 218104
rect 487858 218048 623962 218104
rect 624018 218048 624023 218104
rect 487797 218046 624023 218048
rect 487797 218043 487863 218046
rect 623957 218043 624023 218046
rect 669630 218044 669636 218108
rect 669700 218106 669706 218108
rect 670325 218106 670391 218109
rect 669700 218104 670391 218106
rect 669700 218048 670330 218104
rect 670386 218048 670391 218104
rect 669700 218046 670391 218048
rect 669700 218044 669706 218046
rect 670325 218043 670391 218046
rect 35525 217970 35591 217973
rect 58801 217970 58867 217973
rect 35525 217968 58867 217970
rect 35525 217912 35530 217968
rect 35586 217912 58806 217968
rect 58862 217912 58867 217968
rect 35525 217910 58867 217912
rect 35525 217907 35591 217910
rect 58801 217907 58867 217910
rect 674005 217970 674071 217973
rect 676029 217970 676095 217973
rect 674005 217968 676095 217970
rect 674005 217912 674010 217968
rect 674066 217912 676034 217968
rect 676090 217912 676095 217968
rect 674005 217910 676095 217912
rect 674005 217907 674071 217910
rect 676029 217907 676095 217910
rect 561305 217834 561371 217837
rect 574737 217834 574803 217837
rect 561305 217832 574803 217834
rect 561305 217776 561310 217832
rect 561366 217776 574742 217832
rect 574798 217776 574803 217832
rect 561305 217774 574803 217776
rect 561305 217771 561371 217774
rect 574737 217771 574803 217774
rect 666645 217834 666711 217837
rect 666645 217832 672826 217834
rect 666645 217776 666650 217832
rect 666706 217776 672826 217832
rect 666645 217774 672826 217776
rect 666645 217771 666711 217774
rect 510981 217564 511047 217565
rect 519997 217564 520063 217565
rect 510981 217562 511028 217564
rect 510936 217560 511028 217562
rect 510936 217504 510986 217560
rect 510936 217502 511028 217504
rect 510981 217500 511028 217502
rect 511092 217500 511098 217564
rect 519997 217562 520044 217564
rect 519952 217560 520044 217562
rect 519952 217504 520002 217560
rect 519952 217502 520044 217504
rect 519997 217500 520044 217502
rect 520108 217500 520114 217564
rect 531497 217562 531563 217565
rect 532509 217564 532575 217565
rect 532509 217562 532556 217564
rect 531497 217560 532556 217562
rect 531497 217504 531502 217560
rect 531558 217504 532514 217560
rect 531497 217502 532556 217504
rect 510981 217499 511047 217500
rect 519997 217499 520063 217500
rect 531497 217499 531563 217502
rect 532509 217500 532556 217502
rect 532620 217500 532626 217564
rect 560753 217562 560819 217565
rect 560937 217562 561003 217565
rect 563329 217562 563395 217565
rect 560753 217560 563395 217562
rect 560753 217504 560758 217560
rect 560814 217504 560942 217560
rect 560998 217504 563334 217560
rect 563390 217504 563395 217560
rect 560753 217502 563395 217504
rect 532509 217499 532575 217500
rect 560753 217499 560819 217502
rect 560937 217499 561003 217502
rect 563329 217499 563395 217502
rect 571977 217562 572043 217565
rect 574185 217562 574251 217565
rect 571977 217560 574251 217562
rect 571977 217504 571982 217560
rect 572038 217504 574190 217560
rect 574246 217504 574251 217560
rect 571977 217502 574251 217504
rect 571977 217499 572043 217502
rect 574185 217499 574251 217502
rect 653765 217562 653831 217565
rect 672073 217562 672139 217565
rect 653765 217560 672139 217562
rect 653765 217504 653770 217560
rect 653826 217504 672078 217560
rect 672134 217504 672139 217560
rect 653765 217502 672139 217504
rect 653765 217499 653831 217502
rect 672073 217499 672139 217502
rect 502241 217290 502307 217293
rect 595161 217290 595227 217293
rect 502241 217288 595227 217290
rect 502241 217232 502246 217288
rect 502302 217232 595166 217288
rect 595222 217232 595227 217288
rect 502241 217230 595227 217232
rect 502241 217227 502307 217230
rect 595161 217227 595227 217230
rect 651097 217290 651163 217293
rect 651097 217288 663810 217290
rect 651097 217232 651102 217288
rect 651158 217232 663810 217288
rect 651097 217230 663810 217232
rect 651097 217227 651163 217230
rect 488809 217154 488875 217157
rect 495157 217154 495223 217157
rect 488809 217152 491034 217154
rect 488809 217096 488814 217152
rect 488870 217096 491034 217152
rect 488809 217094 491034 217096
rect 488809 217091 488875 217094
rect 490974 216746 491034 217094
rect 495157 217152 499590 217154
rect 495157 217096 495162 217152
rect 495218 217096 499590 217152
rect 495157 217094 499590 217096
rect 495157 217091 495223 217094
rect 499530 217018 499590 217094
rect 595713 217018 595779 217021
rect 499530 217016 595779 217018
rect 499530 216960 595718 217016
rect 595774 216960 595779 217016
rect 499530 216958 595779 216960
rect 663750 217018 663810 217230
rect 669078 217228 669084 217292
rect 669148 217290 669154 217292
rect 669405 217290 669471 217293
rect 669148 217288 669471 217290
rect 669148 217232 669410 217288
rect 669466 217232 669471 217288
rect 669148 217230 669471 217232
rect 669148 217228 669154 217230
rect 669405 217227 669471 217230
rect 672766 217154 672826 217774
rect 676170 217774 676292 217834
rect 675702 217636 675708 217700
rect 675772 217698 675778 217700
rect 676170 217698 676230 217774
rect 675772 217638 676230 217698
rect 675772 217636 675778 217638
rect 672993 217426 673059 217429
rect 672993 217424 676292 217426
rect 672993 217368 672998 217424
rect 673054 217368 676292 217424
rect 672993 217366 676292 217368
rect 672993 217363 673059 217366
rect 672766 217094 676230 217154
rect 676170 217018 676230 217094
rect 663750 216958 669330 217018
rect 676170 216958 676292 217018
rect 595713 216955 595779 216958
rect 669270 216882 669330 216958
rect 673545 216882 673611 216885
rect 669270 216880 673611 216882
rect 669270 216824 673550 216880
rect 673606 216824 673611 216880
rect 669270 216822 673611 216824
rect 673545 216819 673611 216822
rect 575473 216746 575539 216749
rect 490974 216744 575539 216746
rect 490974 216688 575478 216744
rect 575534 216688 575539 216744
rect 490974 216686 575539 216688
rect 575473 216683 575539 216686
rect 670509 216610 670575 216613
rect 672993 216610 673059 216613
rect 670509 216608 673059 216610
rect 670509 216552 670514 216608
rect 670570 216552 672998 216608
rect 673054 216552 673059 216608
rect 670509 216550 673059 216552
rect 670509 216547 670575 216550
rect 672993 216547 673059 216550
rect 673545 216610 673611 216613
rect 673545 216608 676292 216610
rect 673545 216552 673550 216608
rect 673606 216552 676292 216608
rect 673545 216550 676292 216552
rect 673545 216547 673611 216550
rect 670325 216476 670391 216477
rect 670325 216474 670372 216476
rect 670280 216472 670372 216474
rect 670280 216416 670330 216472
rect 670280 216414 670372 216416
rect 670325 216412 670372 216414
rect 670436 216412 670442 216476
rect 670325 216411 670391 216412
rect 671889 216202 671955 216205
rect 669270 216200 671955 216202
rect 669270 216144 671894 216200
rect 671950 216144 671955 216200
rect 669270 216142 671955 216144
rect 520038 215868 520044 215932
rect 520108 215930 520114 215932
rect 617793 215930 617859 215933
rect 669270 215930 669330 216142
rect 671889 216139 671955 216142
rect 672073 216202 672139 216205
rect 672073 216200 676292 216202
rect 672073 216144 672078 216200
rect 672134 216144 676292 216200
rect 672073 216142 676292 216144
rect 672073 216139 672139 216142
rect 520108 215928 617859 215930
rect 520108 215872 617798 215928
rect 617854 215872 617859 215928
rect 520108 215870 617859 215872
rect 520108 215868 520114 215870
rect 617793 215867 617859 215870
rect 663750 215870 669330 215930
rect 511022 215596 511028 215660
rect 511092 215658 511098 215660
rect 599025 215658 599091 215661
rect 511092 215656 599091 215658
rect 511092 215600 599030 215656
rect 599086 215600 599091 215656
rect 511092 215598 599091 215600
rect 511092 215596 511098 215598
rect 599025 215595 599091 215598
rect 662413 215658 662479 215661
rect 663750 215658 663810 215870
rect 669814 215868 669820 215932
rect 669884 215930 669890 215932
rect 673545 215930 673611 215933
rect 669884 215928 673611 215930
rect 669884 215872 673550 215928
rect 673606 215872 673611 215928
rect 669884 215870 673611 215872
rect 669884 215868 669890 215870
rect 673545 215867 673611 215870
rect 673862 215868 673868 215932
rect 673932 215930 673938 215932
rect 676029 215930 676095 215933
rect 673932 215928 676095 215930
rect 673932 215872 676034 215928
rect 676090 215872 676095 215928
rect 673932 215870 676095 215872
rect 673932 215868 673938 215870
rect 676029 215867 676095 215870
rect 676170 215734 676292 215794
rect 662413 215656 663810 215658
rect 662413 215600 662418 215656
rect 662474 215600 663810 215656
rect 662413 215598 663810 215600
rect 666829 215658 666895 215661
rect 676170 215658 676230 215734
rect 666829 215656 676230 215658
rect 666829 215600 666834 215656
rect 666890 215600 676230 215656
rect 666829 215598 676230 215600
rect 662413 215595 662479 215598
rect 666829 215595 666895 215598
rect 532550 215324 532556 215388
rect 532620 215386 532626 215388
rect 621105 215386 621171 215389
rect 532620 215384 621171 215386
rect 532620 215328 621110 215384
rect 621166 215328 621171 215384
rect 532620 215326 621171 215328
rect 532620 215324 532626 215326
rect 621105 215323 621171 215326
rect 657905 215386 657971 215389
rect 670550 215386 670556 215388
rect 657905 215384 670556 215386
rect 657905 215328 657910 215384
rect 657966 215328 670556 215384
rect 657905 215326 670556 215328
rect 657905 215323 657971 215326
rect 670550 215324 670556 215326
rect 670620 215324 670626 215388
rect 671889 215386 671955 215389
rect 675661 215386 675727 215389
rect 671889 215384 675727 215386
rect 671889 215328 671894 215384
rect 671950 215328 675666 215384
rect 675722 215328 675727 215384
rect 671889 215326 675727 215328
rect 671889 215323 671955 215326
rect 675661 215323 675727 215326
rect 676262 215310 676322 215356
rect 675886 215188 675892 215252
rect 675956 215250 675962 215252
rect 676078 215250 676322 215310
rect 675956 215190 676138 215250
rect 675956 215188 675962 215190
rect 52453 215114 52519 215117
rect 53281 215114 53347 215117
rect 52453 215112 53347 215114
rect 52453 215056 52458 215112
rect 52514 215056 53286 215112
rect 53342 215056 53347 215112
rect 52453 215054 53347 215056
rect 52453 215051 52519 215054
rect 53281 215051 53347 215054
rect 674465 214978 674531 214981
rect 674465 214976 676292 214978
rect 35758 214709 35818 214948
rect 674465 214920 674470 214976
rect 674526 214920 676292 214976
rect 674465 214918 676292 214920
rect 674465 214915 674531 214918
rect 669405 214842 669471 214845
rect 669814 214842 669820 214844
rect 669405 214840 669820 214842
rect 669405 214784 669410 214840
rect 669466 214784 669820 214840
rect 669405 214782 669820 214784
rect 669405 214779 669471 214782
rect 669814 214780 669820 214782
rect 669884 214780 669890 214844
rect 35525 214706 35591 214709
rect 35525 214704 35634 214706
rect 35525 214648 35530 214704
rect 35586 214648 35634 214704
rect 35525 214643 35634 214648
rect 35758 214704 35867 214709
rect 35758 214648 35806 214704
rect 35862 214648 35867 214704
rect 35758 214646 35867 214648
rect 35801 214643 35867 214646
rect 35574 214540 35634 214643
rect 660389 214570 660455 214573
rect 660389 214568 663810 214570
rect 660389 214512 660394 214568
rect 660450 214512 663810 214568
rect 660389 214510 663810 214512
rect 660389 214507 660455 214510
rect 52453 214298 52519 214301
rect 41462 214296 52519 214298
rect 41462 214240 52458 214296
rect 52514 214240 52519 214296
rect 41462 214238 52519 214240
rect 41462 214132 41522 214238
rect 52453 214235 52519 214238
rect 575982 214026 576042 214404
rect 663750 214298 663810 214510
rect 675886 214508 675892 214572
rect 675956 214570 675962 214572
rect 675956 214510 676292 214570
rect 675956 214508 675962 214510
rect 675753 214434 675819 214437
rect 669270 214432 675819 214434
rect 669270 214376 675758 214432
rect 675814 214376 675819 214432
rect 669270 214374 675819 214376
rect 669270 214298 669330 214374
rect 675753 214371 675819 214374
rect 663750 214238 669330 214298
rect 673085 214162 673151 214165
rect 673085 214160 676292 214162
rect 673085 214104 673090 214160
rect 673146 214104 676292 214160
rect 673085 214102 676292 214104
rect 673085 214099 673151 214102
rect 578877 214026 578943 214029
rect 575982 214024 578943 214026
rect 575982 213968 578882 214024
rect 578938 213968 578943 214024
rect 575982 213966 578943 213968
rect 578877 213963 578943 213966
rect 674649 213754 674715 213757
rect 674649 213752 676292 213754
rect 35758 213485 35818 213724
rect 674649 213696 674654 213752
rect 674710 213696 676292 213752
rect 674649 213694 676292 213696
rect 674649 213691 674715 213694
rect 673862 213618 673868 213620
rect 663750 213558 673868 213618
rect 35758 213480 35867 213485
rect 35758 213424 35806 213480
rect 35862 213424 35867 213480
rect 35758 213422 35867 213424
rect 35801 213419 35867 213422
rect 39573 213482 39639 213485
rect 42793 213482 42859 213485
rect 39573 213480 42859 213482
rect 39573 213424 39578 213480
rect 39634 213424 42798 213480
rect 42854 213424 42859 213480
rect 39573 213422 42859 213424
rect 39573 213419 39639 213422
rect 42793 213419 42859 213422
rect 658733 213482 658799 213485
rect 663750 213482 663810 213558
rect 673862 213556 673868 213558
rect 673932 213556 673938 213620
rect 658733 213480 663810 213482
rect 658733 213424 658738 213480
rect 658794 213424 663810 213480
rect 658733 213422 663810 213424
rect 658733 213419 658799 213422
rect 672625 213346 672691 213349
rect 672625 213344 676292 213346
rect 672625 213288 672630 213344
rect 672686 213288 676292 213344
rect 672625 213286 676292 213288
rect 672625 213283 672691 213286
rect 661493 213210 661559 213213
rect 672441 213210 672507 213213
rect 661493 213208 672507 213210
rect 661493 213152 661498 213208
rect 661554 213152 672446 213208
rect 672502 213152 672507 213208
rect 661493 213150 672507 213152
rect 661493 213147 661559 213150
rect 672441 213147 672507 213150
rect 45645 212938 45711 212941
rect 41492 212936 45711 212938
rect 41492 212880 45650 212936
rect 45706 212880 45711 212936
rect 41492 212878 45711 212880
rect 45645 212875 45711 212878
rect 675293 212530 675359 212533
rect 675702 212530 675708 212532
rect 675293 212528 675708 212530
rect 675293 212472 675298 212528
rect 675354 212472 675708 212528
rect 675293 212470 675708 212472
rect 675293 212467 675359 212470
rect 675702 212468 675708 212470
rect 675772 212530 675778 212532
rect 683070 212530 683130 212908
rect 675772 212500 683130 212530
rect 675772 212470 683100 212500
rect 675772 212468 675778 212470
rect 44173 212122 44239 212125
rect 41492 212120 44239 212122
rect 41492 212064 44178 212120
rect 44234 212064 44239 212120
rect 41492 212062 44239 212064
rect 44173 212059 44239 212062
rect 575982 211714 576042 212228
rect 672441 212122 672507 212125
rect 672441 212120 676292 212122
rect 672441 212064 672446 212120
rect 672502 212064 676292 212120
rect 672441 212062 676292 212064
rect 672441 212059 672507 212062
rect 578509 211714 578575 211717
rect 575982 211712 578575 211714
rect 575982 211656 578514 211712
rect 578570 211656 578575 211712
rect 575982 211654 578575 211656
rect 578509 211651 578575 211654
rect 46197 211306 46263 211309
rect 41492 211304 46263 211306
rect 41492 211248 46202 211304
rect 46258 211248 46263 211304
rect 41492 211246 46263 211248
rect 46197 211243 46263 211246
rect 670141 211170 670207 211173
rect 670366 211170 670372 211172
rect 670141 211168 670372 211170
rect 670141 211112 670146 211168
rect 670202 211112 670372 211168
rect 670141 211110 670372 211112
rect 670141 211107 670207 211110
rect 670366 211108 670372 211110
rect 670436 211108 670442 211172
rect 35758 210221 35818 210460
rect 35758 210216 35867 210221
rect 35758 210160 35806 210216
rect 35862 210160 35867 210216
rect 35758 210158 35867 210160
rect 35801 210155 35867 210158
rect 41822 210082 41828 210084
rect 41492 210022 41828 210082
rect 41822 210020 41828 210022
rect 41892 210020 41898 210084
rect 575982 209810 576042 210052
rect 579521 209810 579587 209813
rect 575982 209808 579587 209810
rect 575982 209752 579526 209808
rect 579582 209752 579587 209808
rect 575982 209750 579587 209752
rect 579521 209747 579587 209750
rect 35574 209405 35634 209644
rect 35574 209400 35683 209405
rect 35574 209344 35622 209400
rect 35678 209344 35683 209400
rect 35574 209342 35683 209344
rect 35617 209339 35683 209342
rect 40125 209402 40191 209405
rect 42977 209402 43043 209405
rect 40125 209400 43043 209402
rect 40125 209344 40130 209400
rect 40186 209344 42982 209400
rect 43038 209344 43043 209400
rect 40125 209342 43043 209344
rect 40125 209339 40191 209342
rect 42977 209339 43043 209342
rect 35758 208997 35818 209236
rect 35758 208992 35867 208997
rect 35758 208936 35806 208992
rect 35862 208936 35867 208992
rect 35758 208934 35867 208936
rect 35801 208931 35867 208934
rect 46933 208858 46999 208861
rect 41492 208856 46999 208858
rect 41492 208800 46938 208856
rect 46994 208800 46999 208856
rect 41492 208798 46999 208800
rect 46933 208795 46999 208798
rect 44357 208450 44423 208453
rect 41492 208448 44423 208450
rect 41492 208392 44362 208448
rect 44418 208392 44423 208448
rect 41492 208390 44423 208392
rect 44357 208387 44423 208390
rect 40033 208178 40099 208181
rect 41638 208178 41644 208180
rect 40033 208176 41644 208178
rect 40033 208120 40038 208176
rect 40094 208120 41644 208176
rect 40033 208118 41644 208120
rect 40033 208115 40099 208118
rect 41638 208116 41644 208118
rect 41708 208116 41714 208180
rect 589457 208042 589523 208045
rect 589457 208040 592572 208042
rect 35758 207773 35818 208012
rect 589457 207984 589462 208040
rect 589518 207984 592572 208040
rect 589457 207982 592572 207984
rect 589457 207979 589523 207982
rect 35758 207768 35867 207773
rect 35758 207712 35806 207768
rect 35862 207712 35867 207768
rect 35758 207710 35867 207712
rect 35801 207707 35867 207710
rect 39757 207770 39823 207773
rect 43805 207770 43871 207773
rect 39757 207768 43871 207770
rect 39757 207712 39762 207768
rect 39818 207712 43810 207768
rect 43866 207712 43871 207768
rect 39757 207710 43871 207712
rect 39757 207707 39823 207710
rect 43805 207707 43871 207710
rect 40542 207364 40602 207604
rect 575982 207498 576042 207876
rect 579521 207498 579587 207501
rect 575982 207496 579587 207498
rect 575982 207440 579526 207496
rect 579582 207440 579587 207496
rect 575982 207438 579587 207440
rect 579521 207435 579587 207438
rect 40534 207300 40540 207364
rect 40604 207300 40610 207364
rect 44173 207226 44239 207229
rect 41492 207224 44239 207226
rect 41492 207168 44178 207224
rect 44234 207168 44239 207224
rect 41492 207166 44239 207168
rect 44173 207163 44239 207166
rect 40125 206954 40191 206957
rect 42793 206954 42859 206957
rect 40125 206952 42859 206954
rect 40125 206896 40130 206952
rect 40186 206896 42798 206952
rect 42854 206896 42859 206952
rect 40125 206894 42859 206896
rect 40125 206891 40191 206894
rect 42793 206891 42859 206894
rect 674230 206892 674236 206956
rect 674300 206954 674306 206956
rect 675201 206954 675267 206957
rect 674300 206952 675267 206954
rect 674300 206896 675206 206952
rect 675262 206896 675267 206952
rect 674300 206894 675267 206896
rect 674300 206892 674306 206894
rect 675201 206891 675267 206894
rect 40726 206548 40786 206788
rect 40718 206484 40724 206548
rect 40788 206484 40794 206548
rect 589457 206410 589523 206413
rect 589457 206408 592572 206410
rect 35801 206138 35867 206141
rect 40910 206140 40970 206380
rect 589457 206352 589462 206408
rect 589518 206352 592572 206408
rect 589457 206350 592572 206352
rect 589457 206347 589523 206350
rect 35758 206136 35867 206138
rect 35758 206080 35806 206136
rect 35862 206080 35867 206136
rect 35758 206075 35867 206080
rect 40902 206076 40908 206140
rect 40972 206076 40978 206140
rect 35758 205972 35818 206075
rect 579521 205866 579587 205869
rect 575798 205864 579587 205866
rect 575798 205808 579526 205864
rect 579582 205808 579587 205864
rect 575798 205806 579587 205808
rect 575798 205700 575858 205806
rect 579521 205803 579587 205806
rect 669262 205668 669268 205732
rect 669332 205730 669338 205732
rect 669630 205730 669636 205732
rect 669332 205670 669636 205730
rect 669332 205668 669338 205670
rect 669630 205668 669636 205670
rect 669700 205668 669706 205732
rect 44541 205594 44607 205597
rect 41492 205592 44607 205594
rect 41492 205536 44546 205592
rect 44602 205536 44607 205592
rect 41492 205534 44607 205536
rect 44541 205531 44607 205534
rect 669262 205396 669268 205460
rect 669332 205458 669338 205460
rect 669630 205458 669636 205460
rect 669332 205398 669636 205458
rect 669332 205396 669338 205398
rect 669630 205396 669636 205398
rect 669700 205396 669706 205460
rect 35574 204917 35634 205156
rect 35574 204912 35683 204917
rect 35574 204856 35622 204912
rect 35678 204856 35683 204912
rect 35574 204854 35683 204856
rect 35617 204851 35683 204854
rect 40217 204914 40283 204917
rect 43253 204914 43319 204917
rect 40217 204912 43319 204914
rect 40217 204856 40222 204912
rect 40278 204856 43258 204912
rect 43314 204856 43319 204912
rect 40217 204854 43319 204856
rect 40217 204851 40283 204854
rect 43253 204851 43319 204854
rect 589457 204778 589523 204781
rect 589457 204776 592572 204778
rect 35758 204509 35818 204748
rect 589457 204720 589462 204776
rect 589518 204720 592572 204776
rect 589457 204718 592572 204720
rect 589457 204715 589523 204718
rect 35758 204504 35867 204509
rect 35758 204448 35806 204504
rect 35862 204448 35867 204504
rect 35758 204446 35867 204448
rect 35801 204443 35867 204446
rect 46197 204370 46263 204373
rect 41492 204368 46263 204370
rect 41492 204312 46202 204368
rect 46258 204312 46263 204368
rect 41492 204310 46263 204312
rect 46197 204307 46263 204310
rect 674925 204234 674991 204237
rect 675385 204234 675451 204237
rect 674925 204232 675451 204234
rect 674925 204176 674930 204232
rect 674986 204176 675390 204232
rect 675446 204176 675451 204232
rect 674925 204174 675451 204176
rect 674925 204171 674991 204174
rect 675385 204171 675451 204174
rect 41689 204098 41755 204101
rect 43989 204098 44055 204101
rect 668301 204098 668367 204101
rect 41689 204096 44055 204098
rect 41689 204040 41694 204096
rect 41750 204040 43994 204096
rect 44050 204040 44055 204096
rect 41689 204038 44055 204040
rect 41689 204035 41755 204038
rect 43989 204035 44055 204038
rect 666694 204096 668367 204098
rect 666694 204040 668306 204096
rect 668362 204040 668367 204096
rect 666694 204038 668367 204040
rect 666694 204030 666754 204038
rect 668301 204035 668367 204038
rect 666356 203970 666754 204030
rect 35758 203693 35818 203932
rect 35758 203688 35867 203693
rect 35758 203632 35806 203688
rect 35862 203632 35867 203688
rect 35758 203630 35867 203632
rect 35801 203627 35867 203630
rect 41505 203690 41571 203693
rect 43621 203690 43687 203693
rect 41505 203688 43687 203690
rect 41505 203632 41510 203688
rect 41566 203632 43626 203688
rect 43682 203632 43687 203688
rect 41505 203630 43687 203632
rect 41505 203627 41571 203630
rect 43621 203627 43687 203630
rect 575982 203282 576042 203524
rect 578325 203282 578391 203285
rect 575982 203280 578391 203282
rect 575982 203224 578330 203280
rect 578386 203224 578391 203280
rect 575982 203222 578391 203224
rect 578325 203219 578391 203222
rect 589457 203146 589523 203149
rect 589457 203144 592572 203146
rect 589457 203088 589462 203144
rect 589518 203088 592572 203144
rect 589457 203086 592572 203088
rect 589457 203083 589523 203086
rect 669405 202874 669471 202877
rect 674925 202874 674991 202877
rect 669405 202872 674991 202874
rect 669405 202816 669410 202872
rect 669466 202816 674930 202872
rect 674986 202816 674991 202872
rect 669405 202814 674991 202816
rect 669405 202811 669471 202814
rect 674925 202811 674991 202814
rect 675753 202738 675819 202741
rect 676254 202738 676260 202740
rect 675753 202736 676260 202738
rect 675753 202680 675758 202736
rect 675814 202680 676260 202736
rect 675753 202678 676260 202680
rect 675753 202675 675819 202678
rect 676254 202676 676260 202678
rect 676324 202676 676330 202740
rect 589457 201514 589523 201517
rect 589457 201512 592572 201514
rect 589457 201456 589462 201512
rect 589518 201456 592572 201512
rect 589457 201454 592572 201456
rect 589457 201451 589523 201454
rect 672073 201378 672139 201381
rect 675477 201378 675543 201381
rect 672073 201376 675543 201378
rect 575982 200834 576042 201348
rect 672073 201320 672078 201376
rect 672134 201320 675482 201376
rect 675538 201320 675543 201376
rect 672073 201318 675543 201320
rect 672073 201315 672139 201318
rect 675477 201315 675543 201318
rect 672441 201106 672507 201109
rect 672441 201104 673010 201106
rect 672441 201048 672446 201104
rect 672502 201048 673010 201104
rect 672441 201046 673010 201048
rect 672441 201043 672507 201046
rect 578785 200834 578851 200837
rect 672533 200836 672599 200837
rect 672533 200834 672580 200836
rect 575982 200832 578851 200834
rect 575982 200776 578790 200832
rect 578846 200776 578851 200832
rect 575982 200774 578851 200776
rect 672488 200832 672580 200834
rect 672488 200776 672538 200832
rect 672488 200774 672580 200776
rect 578785 200771 578851 200774
rect 672533 200772 672580 200774
rect 672644 200772 672650 200836
rect 672533 200771 672599 200772
rect 672950 200701 673010 201046
rect 672901 200696 673010 200701
rect 672901 200640 672906 200696
rect 672962 200640 673010 200696
rect 672901 200638 673010 200640
rect 672901 200635 672967 200638
rect 675753 200018 675819 200021
rect 676438 200018 676444 200020
rect 675753 200016 676444 200018
rect 675753 199960 675758 200016
rect 675814 199960 676444 200016
rect 675753 199958 676444 199960
rect 675753 199955 675819 199958
rect 676438 199956 676444 199958
rect 676508 199956 676514 200020
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 673085 199746 673151 199749
rect 674925 199746 674991 199749
rect 673085 199744 674991 199746
rect 673085 199688 673090 199744
rect 673146 199688 674930 199744
rect 674986 199688 674991 199744
rect 673085 199686 674991 199688
rect 673085 199683 673151 199686
rect 674925 199683 674991 199686
rect 668945 199202 669011 199205
rect 666694 199200 669011 199202
rect 575982 198930 576042 199172
rect 666694 199144 668950 199200
rect 669006 199144 669011 199200
rect 666694 199142 669011 199144
rect 666694 199134 666754 199142
rect 668945 199139 669011 199142
rect 666356 199074 666754 199134
rect 579521 198930 579587 198933
rect 575982 198928 579587 198930
rect 575982 198872 579526 198928
rect 579582 198872 579587 198928
rect 575982 198870 579587 198872
rect 579521 198867 579587 198870
rect 37917 198794 37983 198797
rect 42006 198794 42012 198796
rect 37917 198792 42012 198794
rect 37917 198736 37922 198792
rect 37978 198736 42012 198792
rect 37917 198734 42012 198736
rect 37917 198731 37983 198734
rect 42006 198732 42012 198734
rect 42076 198732 42082 198796
rect 668393 198794 668459 198797
rect 670734 198794 670740 198796
rect 668393 198792 670740 198794
rect 668393 198736 668398 198792
rect 668454 198736 670740 198792
rect 668393 198734 670740 198736
rect 668393 198731 668459 198734
rect 670734 198732 670740 198734
rect 670804 198732 670810 198796
rect 666829 198522 666895 198525
rect 675109 198522 675175 198525
rect 666829 198520 675175 198522
rect 666829 198464 666834 198520
rect 666890 198464 675114 198520
rect 675170 198464 675175 198520
rect 666829 198462 675175 198464
rect 666829 198459 666895 198462
rect 675109 198459 675175 198462
rect 590377 198250 590443 198253
rect 670509 198250 670575 198253
rect 675477 198250 675543 198253
rect 590377 198248 592572 198250
rect 590377 198192 590382 198248
rect 590438 198192 592572 198248
rect 590377 198190 592572 198192
rect 670509 198248 675543 198250
rect 670509 198192 670514 198248
rect 670570 198192 675482 198248
rect 675538 198192 675543 198248
rect 670509 198190 675543 198192
rect 590377 198187 590443 198190
rect 670509 198187 670575 198190
rect 675477 198187 675543 198190
rect 673177 197842 673243 197845
rect 676806 197842 676812 197844
rect 673177 197840 676812 197842
rect 673177 197784 673182 197840
rect 673238 197784 676812 197840
rect 673177 197782 676812 197784
rect 673177 197779 673243 197782
rect 676806 197780 676812 197782
rect 676876 197780 676882 197844
rect 42425 197298 42491 197301
rect 44357 197298 44423 197301
rect 42425 197296 44423 197298
rect 42425 197240 42430 197296
rect 42486 197240 44362 197296
rect 44418 197240 44423 197296
rect 42425 197238 44423 197240
rect 42425 197235 42491 197238
rect 44357 197235 44423 197238
rect 674465 197162 674531 197165
rect 675385 197162 675451 197165
rect 674465 197160 675451 197162
rect 674465 197104 674470 197160
rect 674526 197104 675390 197160
rect 675446 197104 675451 197160
rect 674465 197102 675451 197104
rect 674465 197099 674531 197102
rect 675385 197099 675451 197102
rect 575982 196482 576042 196996
rect 589457 196618 589523 196621
rect 589457 196616 592572 196618
rect 589457 196560 589462 196616
rect 589518 196560 592572 196616
rect 589457 196558 592572 196560
rect 589457 196555 589523 196558
rect 578509 196482 578575 196485
rect 575982 196480 578575 196482
rect 575982 196424 578514 196480
rect 578570 196424 578575 196480
rect 575982 196422 578575 196424
rect 578509 196419 578575 196422
rect 669262 196012 669268 196076
rect 669332 196074 669338 196076
rect 669630 196074 669636 196076
rect 669332 196014 669636 196074
rect 669332 196012 669338 196014
rect 669630 196012 669636 196014
rect 669700 196012 669706 196076
rect 41965 195804 42031 195805
rect 41965 195800 42012 195804
rect 42076 195802 42082 195804
rect 41965 195744 41970 195800
rect 41965 195740 42012 195744
rect 42076 195742 42122 195802
rect 42076 195740 42082 195742
rect 41965 195739 42031 195740
rect 41781 195260 41847 195261
rect 41781 195256 41828 195260
rect 41892 195258 41898 195260
rect 41781 195200 41786 195256
rect 41781 195196 41828 195200
rect 41892 195198 41938 195258
rect 41892 195196 41898 195198
rect 41781 195195 41847 195196
rect 40902 194924 40908 194988
rect 40972 194986 40978 194988
rect 42241 194986 42307 194989
rect 579521 194986 579587 194989
rect 40972 194984 42307 194986
rect 40972 194928 42246 194984
rect 42302 194928 42307 194984
rect 40972 194926 42307 194928
rect 40972 194924 40978 194926
rect 42241 194923 42307 194926
rect 575798 194984 579587 194986
rect 575798 194928 579526 194984
rect 579582 194928 579587 194984
rect 575798 194926 579587 194928
rect 575798 194820 575858 194926
rect 579521 194923 579587 194926
rect 589273 194986 589339 194989
rect 589273 194984 592572 194986
rect 589273 194928 589278 194984
rect 589334 194928 592572 194984
rect 589273 194926 592572 194928
rect 589273 194923 589339 194926
rect 675753 194578 675819 194581
rect 676622 194578 676628 194580
rect 675753 194576 676628 194578
rect 675753 194520 675758 194576
rect 675814 194520 676628 194576
rect 675753 194518 676628 194520
rect 675753 194515 675819 194518
rect 676622 194516 676628 194518
rect 676692 194516 676698 194580
rect 668117 194306 668183 194309
rect 666694 194304 668183 194306
rect 666694 194248 668122 194304
rect 668178 194248 668183 194304
rect 666694 194246 668183 194248
rect 666694 194238 666754 194246
rect 668117 194243 668183 194246
rect 666356 194178 666754 194238
rect 40718 193428 40724 193492
rect 40788 193490 40794 193492
rect 41781 193490 41847 193493
rect 40788 193488 41847 193490
rect 40788 193432 41786 193488
rect 41842 193432 41847 193488
rect 40788 193430 41847 193432
rect 40788 193428 40794 193430
rect 41781 193427 41847 193430
rect 589457 193354 589523 193357
rect 589457 193352 592572 193354
rect 589457 193296 589462 193352
rect 589518 193296 592572 193352
rect 589457 193294 592572 193296
rect 589457 193291 589523 193294
rect 675753 193218 675819 193221
rect 676070 193218 676076 193220
rect 675753 193216 676076 193218
rect 675753 193160 675758 193216
rect 675814 193160 676076 193216
rect 675753 193158 676076 193160
rect 675753 193155 675819 193158
rect 676070 193156 676076 193158
rect 676140 193156 676146 193220
rect 675661 192810 675727 192813
rect 675886 192810 675892 192812
rect 675661 192808 675892 192810
rect 675661 192752 675666 192808
rect 675722 192752 675892 192808
rect 675661 192750 675892 192752
rect 675661 192747 675727 192750
rect 675886 192748 675892 192750
rect 675956 192748 675962 192812
rect 575982 192266 576042 192644
rect 579521 192266 579587 192269
rect 575982 192264 579587 192266
rect 575982 192208 579526 192264
rect 579582 192208 579587 192264
rect 575982 192206 579587 192208
rect 579521 192203 579587 192206
rect 589457 191722 589523 191725
rect 669037 191722 669103 191725
rect 669446 191722 669452 191724
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 669037 191720 669452 191722
rect 669037 191664 669042 191720
rect 669098 191664 669452 191720
rect 669037 191662 669452 191664
rect 589457 191659 589523 191662
rect 669037 191659 669103 191662
rect 669446 191660 669452 191662
rect 669516 191660 669522 191724
rect 42057 191586 42123 191589
rect 43989 191586 44055 191589
rect 42057 191584 44055 191586
rect 42057 191528 42062 191584
rect 42118 191528 43994 191584
rect 44050 191528 44055 191584
rect 42057 191526 44055 191528
rect 42057 191523 42123 191526
rect 43989 191523 44055 191526
rect 579521 190770 579587 190773
rect 575798 190768 579587 190770
rect 575798 190712 579526 190768
rect 579582 190712 579587 190768
rect 575798 190710 579587 190712
rect 42425 190498 42491 190501
rect 44541 190498 44607 190501
rect 42425 190496 44607 190498
rect 42425 190440 42430 190496
rect 42486 190440 44546 190496
rect 44602 190440 44607 190496
rect 575798 190468 575858 190710
rect 579521 190707 579587 190710
rect 42425 190438 44607 190440
rect 42425 190435 42491 190438
rect 44541 190435 44607 190438
rect 590561 190090 590627 190093
rect 590561 190088 592572 190090
rect 590561 190032 590566 190088
rect 590622 190032 592572 190088
rect 590561 190030 592572 190032
rect 590561 190027 590627 190030
rect 669221 189410 669287 189413
rect 666694 189408 669287 189410
rect 666694 189352 669226 189408
rect 669282 189352 669287 189408
rect 666694 189350 669287 189352
rect 666694 189342 666754 189350
rect 669221 189347 669287 189350
rect 666356 189282 666754 189342
rect 675334 189076 675340 189140
rect 675404 189138 675410 189140
rect 676121 189138 676187 189141
rect 675404 189136 676187 189138
rect 675404 189080 676126 189136
rect 676182 189080 676187 189136
rect 675404 189078 676187 189080
rect 675404 189076 675410 189078
rect 676121 189075 676187 189078
rect 666645 188866 666711 188869
rect 675109 188866 675175 188869
rect 666645 188864 675175 188866
rect 666645 188808 666650 188864
rect 666706 188808 675114 188864
rect 675170 188808 675175 188864
rect 666645 188806 675175 188808
rect 666645 188803 666711 188806
rect 675109 188803 675175 188806
rect 589641 188458 589707 188461
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 589641 188395 589707 188398
rect 575982 188050 576042 188292
rect 579521 188050 579587 188053
rect 575982 188048 579587 188050
rect 575982 187992 579526 188048
rect 579582 187992 579587 188048
rect 575982 187990 579587 187992
rect 579521 187987 579587 187990
rect 42425 187642 42491 187645
rect 46933 187642 46999 187645
rect 42425 187640 46999 187642
rect 42425 187584 42430 187640
rect 42486 187584 46938 187640
rect 46994 187584 46999 187640
rect 42425 187582 46999 187584
rect 42425 187579 42491 187582
rect 46933 187579 46999 187582
rect 42425 186826 42491 186829
rect 44173 186826 44239 186829
rect 42425 186824 44239 186826
rect 42425 186768 42430 186824
rect 42486 186768 44178 186824
rect 44234 186768 44239 186824
rect 42425 186766 44239 186768
rect 42425 186763 42491 186766
rect 44173 186763 44239 186766
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 40534 186356 40540 186420
rect 40604 186418 40610 186420
rect 41781 186418 41847 186421
rect 40604 186416 41847 186418
rect 40604 186360 41786 186416
rect 41842 186360 41847 186416
rect 40604 186358 41847 186360
rect 40604 186356 40610 186358
rect 41781 186355 41847 186358
rect 579521 186282 579587 186285
rect 575798 186280 579587 186282
rect 575798 186224 579526 186280
rect 579582 186224 579587 186280
rect 575798 186222 579587 186224
rect 575798 186116 575858 186222
rect 579521 186219 579587 186222
rect 41454 185948 41460 186012
rect 41524 186010 41530 186012
rect 41781 186010 41847 186013
rect 41524 186008 41847 186010
rect 41524 185952 41786 186008
rect 41842 185952 41847 186008
rect 41524 185950 41847 185952
rect 41524 185948 41530 185950
rect 41781 185947 41847 185950
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 667933 184514 667999 184517
rect 666694 184512 667999 184514
rect 666694 184456 667938 184512
rect 667994 184456 667999 184512
rect 666694 184454 667999 184456
rect 666694 184446 666754 184454
rect 667933 184451 667999 184454
rect 666356 184386 666754 184446
rect 579521 184378 579587 184381
rect 575798 184376 579587 184378
rect 575798 184320 579526 184376
rect 579582 184320 579587 184376
rect 575798 184318 579587 184320
rect 575798 183940 575858 184318
rect 579521 184315 579587 184318
rect 589457 183562 589523 183565
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 589457 183499 589523 183502
rect 42425 183018 42491 183021
rect 43805 183018 43871 183021
rect 42425 183016 43871 183018
rect 42425 182960 42430 183016
rect 42486 182960 43810 183016
rect 43866 182960 43871 183016
rect 42425 182958 43871 182960
rect 42425 182955 42491 182958
rect 43805 182955 43871 182958
rect 579521 181930 579587 181933
rect 575798 181928 579587 181930
rect 575798 181872 579526 181928
rect 579582 181872 579587 181928
rect 575798 181870 579587 181872
rect 575798 181764 575858 181870
rect 579521 181867 579587 181870
rect 590561 181930 590627 181933
rect 590561 181928 592572 181930
rect 590561 181872 590566 181928
rect 590622 181872 592572 181928
rect 590561 181870 592572 181872
rect 590561 181867 590627 181870
rect 672533 181658 672599 181661
rect 673126 181658 673132 181660
rect 672533 181656 673132 181658
rect 672533 181600 672538 181656
rect 672594 181600 673132 181656
rect 672533 181598 673132 181600
rect 672533 181595 672599 181598
rect 673126 181596 673132 181598
rect 673196 181596 673202 181660
rect 667565 181386 667631 181389
rect 675293 181386 675359 181389
rect 667565 181384 675359 181386
rect 667565 181328 667570 181384
rect 667626 181328 675298 181384
rect 675354 181328 675359 181384
rect 667565 181326 675359 181328
rect 667565 181323 667631 181326
rect 675293 181323 675359 181326
rect 589641 180298 589707 180301
rect 589641 180296 592572 180298
rect 589641 180240 589646 180296
rect 589702 180240 592572 180296
rect 589641 180238 592572 180240
rect 589641 180235 589707 180238
rect 578785 180162 578851 180165
rect 575798 180160 578851 180162
rect 575798 180104 578790 180160
rect 578846 180104 578851 180160
rect 575798 180102 578851 180104
rect 575798 179588 575858 180102
rect 578785 180099 578851 180102
rect 668158 179618 668164 179620
rect 666694 179558 668164 179618
rect 666694 179550 666754 179558
rect 668158 179556 668164 179558
rect 668228 179556 668234 179620
rect 666356 179490 666754 179550
rect 673310 179420 673316 179484
rect 673380 179482 673386 179484
rect 675477 179482 675543 179485
rect 673380 179480 675543 179482
rect 673380 179424 675482 179480
rect 675538 179424 675543 179480
rect 673380 179422 675543 179424
rect 673380 179420 673386 179422
rect 675477 179419 675543 179422
rect 42057 179346 42123 179349
rect 47761 179346 47827 179349
rect 42057 179344 47827 179346
rect 42057 179288 42062 179344
rect 42118 179288 47766 179344
rect 47822 179288 47827 179344
rect 42057 179286 47827 179288
rect 42057 179283 42123 179286
rect 47761 179283 47827 179286
rect 675293 179074 675359 179077
rect 675293 179072 676322 179074
rect 675293 179016 675298 179072
rect 675354 179016 676322 179072
rect 675293 179014 676322 179016
rect 675293 179011 675359 179014
rect 667381 178802 667447 178805
rect 675661 178802 675727 178805
rect 667381 178800 675727 178802
rect 667381 178744 667386 178800
rect 667442 178744 675666 178800
rect 675722 178744 675727 178800
rect 667381 178742 675727 178744
rect 667381 178739 667447 178742
rect 675661 178739 675727 178742
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 676262 178500 676322 179014
rect 675477 178122 675543 178125
rect 675477 178120 676292 178122
rect 675477 178064 675482 178120
rect 675538 178064 676292 178120
rect 675477 178062 676292 178064
rect 675477 178059 675543 178062
rect 668209 177986 668275 177989
rect 666694 177984 668275 177986
rect 666694 177928 668214 177984
rect 668270 177928 668275 177984
rect 666694 177926 668275 177928
rect 666694 177918 666754 177926
rect 668209 177923 668275 177926
rect 670785 177986 670851 177989
rect 671337 177986 671403 177989
rect 670785 177984 671403 177986
rect 670785 177928 670790 177984
rect 670846 177928 671342 177984
rect 671398 177928 671403 177984
rect 670785 177926 671403 177928
rect 670785 177923 670851 177926
rect 671337 177923 671403 177926
rect 666356 177858 666754 177918
rect 579521 177714 579587 177717
rect 575798 177712 579587 177714
rect 575798 177656 579526 177712
rect 579582 177656 579587 177712
rect 575798 177654 579587 177656
rect 575798 177412 575858 177654
rect 579521 177651 579587 177654
rect 675661 177714 675727 177717
rect 675661 177712 676292 177714
rect 675661 177656 675666 177712
rect 675722 177656 676292 177712
rect 675661 177654 676292 177656
rect 675661 177651 675727 177654
rect 673913 177306 673979 177309
rect 673913 177304 676292 177306
rect 673913 177248 673918 177304
rect 673974 177248 676292 177304
rect 673913 177246 676292 177248
rect 673913 177243 673979 177246
rect 589641 177034 589707 177037
rect 589641 177032 592572 177034
rect 589641 176976 589646 177032
rect 589702 176976 592572 177032
rect 589641 176974 592572 176976
rect 589641 176971 589707 176974
rect 673913 176898 673979 176901
rect 673913 176896 676292 176898
rect 673913 176840 673918 176896
rect 673974 176840 676292 176896
rect 673913 176838 676292 176840
rect 673913 176835 673979 176838
rect 676806 176608 676812 176672
rect 676876 176608 676882 176672
rect 676814 176460 676874 176608
rect 674649 176082 674715 176085
rect 674649 176080 676292 176082
rect 674649 176024 674654 176080
rect 674710 176024 676292 176080
rect 674649 176022 676292 176024
rect 674649 176019 674715 176022
rect 673361 175674 673427 175677
rect 673361 175672 676292 175674
rect 673361 175616 673366 175672
rect 673422 175616 676292 175672
rect 673361 175614 676292 175616
rect 673361 175611 673427 175614
rect 589457 175402 589523 175405
rect 589457 175400 592572 175402
rect 589457 175344 589462 175400
rect 589518 175344 592572 175400
rect 589457 175342 592572 175344
rect 589457 175339 589523 175342
rect 674465 175266 674531 175269
rect 674465 175264 676292 175266
rect 575982 175130 576042 175236
rect 674465 175208 674470 175264
rect 674526 175208 676292 175264
rect 674465 175206 676292 175208
rect 674465 175203 674531 175206
rect 578785 175130 578851 175133
rect 575982 175128 578851 175130
rect 575982 175072 578790 175128
rect 578846 175072 578851 175128
rect 575982 175070 578851 175072
rect 578785 175067 578851 175070
rect 667749 174994 667815 174997
rect 667749 174992 669330 174994
rect 667749 174936 667754 174992
rect 667810 174936 669330 174992
rect 667749 174934 669330 174936
rect 667749 174931 667815 174934
rect 669270 174858 669330 174934
rect 669270 174798 676292 174858
rect 667933 174722 667999 174725
rect 666694 174720 667999 174722
rect 666694 174664 667938 174720
rect 667994 174664 667999 174720
rect 666694 174662 667999 174664
rect 666694 174654 666754 174662
rect 667933 174659 667999 174662
rect 666356 174594 666754 174654
rect 673269 174450 673335 174453
rect 673269 174448 676292 174450
rect 673269 174392 673274 174448
rect 673330 174392 676292 174448
rect 673269 174390 676292 174392
rect 673269 174387 673335 174390
rect 676029 174042 676095 174045
rect 676029 174040 676292 174042
rect 676029 173984 676034 174040
rect 676090 173984 676292 174040
rect 676029 173982 676292 173984
rect 676029 173979 676095 173982
rect 589457 173770 589523 173773
rect 589457 173768 592572 173770
rect 589457 173712 589462 173768
rect 589518 173712 592572 173768
rect 589457 173710 592572 173712
rect 589457 173707 589523 173710
rect 675702 173572 675708 173636
rect 675772 173634 675778 173636
rect 675772 173574 676292 173634
rect 675772 173572 675778 173574
rect 578417 173498 578483 173501
rect 575798 173496 578483 173498
rect 575798 173440 578422 173496
rect 578478 173440 578483 173496
rect 575798 173438 578483 173440
rect 575798 173060 575858 173438
rect 578417 173435 578483 173438
rect 679617 173226 679683 173229
rect 679604 173224 679683 173226
rect 679604 173168 679622 173224
rect 679678 173168 679683 173224
rect 679604 173166 679683 173168
rect 679617 173163 679683 173166
rect 666356 172962 666938 173022
rect 666878 172954 666938 172962
rect 674097 172954 674163 172957
rect 666878 172952 674163 172954
rect 666878 172896 674102 172952
rect 674158 172896 674163 172952
rect 666878 172894 674163 172896
rect 674097 172891 674163 172894
rect 680997 172818 681063 172821
rect 680997 172816 681076 172818
rect 680997 172760 681002 172816
rect 681058 172760 681076 172816
rect 680997 172758 681076 172760
rect 680997 172755 681063 172758
rect 675518 172348 675524 172412
rect 675588 172410 675594 172412
rect 675588 172350 676292 172410
rect 675588 172348 675594 172350
rect 673545 172274 673611 172277
rect 674097 172274 674163 172277
rect 673545 172272 674163 172274
rect 673545 172216 673550 172272
rect 673606 172216 674102 172272
rect 674158 172216 674163 172272
rect 673545 172214 674163 172216
rect 673545 172211 673611 172214
rect 674097 172211 674163 172214
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 671889 172002 671955 172005
rect 671889 172000 676292 172002
rect 671889 171944 671894 172000
rect 671950 171944 676292 172000
rect 671889 171942 676292 171944
rect 671889 171939 671955 171942
rect 673453 171594 673519 171597
rect 673453 171592 676292 171594
rect 673453 171536 673458 171592
rect 673514 171536 676292 171592
rect 673453 171534 676292 171536
rect 673453 171531 673519 171534
rect 669589 171186 669655 171189
rect 669589 171184 676292 171186
rect 669589 171128 669594 171184
rect 669650 171128 676292 171184
rect 669589 171126 676292 171128
rect 669589 171123 669655 171126
rect 578233 171050 578299 171053
rect 575798 171048 578299 171050
rect 575798 170992 578238 171048
rect 578294 170992 578299 171048
rect 575798 170990 578299 170992
rect 575798 170884 575858 170990
rect 578233 170987 578299 170990
rect 675886 170716 675892 170780
rect 675956 170778 675962 170780
rect 675956 170718 676292 170778
rect 675956 170716 675962 170718
rect 589641 170506 589707 170509
rect 589641 170504 592572 170506
rect 589641 170448 589646 170504
rect 589702 170448 592572 170504
rect 589641 170446 592572 170448
rect 589641 170443 589707 170446
rect 670601 170370 670667 170373
rect 670601 170368 676292 170370
rect 670601 170312 670606 170368
rect 670662 170312 676292 170368
rect 670601 170310 676292 170312
rect 670601 170307 670667 170310
rect 675894 169902 676292 169962
rect 666356 169698 666754 169758
rect 666694 169690 666754 169698
rect 667933 169690 667999 169693
rect 675894 169692 675954 169902
rect 666694 169688 667999 169690
rect 666694 169632 667938 169688
rect 667994 169632 667999 169688
rect 666694 169630 667999 169632
rect 667933 169627 667999 169630
rect 675886 169628 675892 169692
rect 675956 169628 675962 169692
rect 669773 169554 669839 169557
rect 675518 169554 675524 169556
rect 669773 169552 675524 169554
rect 669773 169496 669778 169552
rect 669834 169496 675524 169552
rect 669773 169494 675524 169496
rect 669773 169491 669839 169494
rect 675518 169492 675524 169494
rect 675588 169492 675594 169556
rect 676397 169554 676463 169557
rect 676397 169552 676476 169554
rect 676397 169496 676402 169552
rect 676458 169496 676476 169552
rect 676397 169494 676476 169496
rect 676397 169491 676463 169494
rect 578693 169282 578759 169285
rect 575798 169280 578759 169282
rect 575798 169224 578698 169280
rect 578754 169224 578759 169280
rect 575798 169222 578759 169224
rect 575798 168708 575858 169222
rect 578693 169219 578759 169222
rect 672073 169146 672139 169149
rect 672073 169144 676292 169146
rect 672073 169088 672078 169144
rect 672134 169088 676292 169144
rect 672073 169086 676292 169088
rect 672073 169083 672139 169086
rect 589457 168874 589523 168877
rect 589457 168872 592572 168874
rect 589457 168816 589462 168872
rect 589518 168816 592572 168872
rect 589457 168814 592572 168816
rect 589457 168811 589523 168814
rect 673177 168738 673243 168741
rect 673177 168736 676292 168738
rect 673177 168680 673182 168736
rect 673238 168680 676292 168736
rect 673177 168678 676292 168680
rect 673177 168675 673243 168678
rect 672533 168330 672599 168333
rect 672533 168328 676292 168330
rect 672533 168272 672538 168328
rect 672594 168272 676292 168328
rect 672533 168270 676292 168272
rect 672533 168267 672599 168270
rect 672257 168194 672323 168197
rect 666694 168192 672323 168194
rect 666694 168136 672262 168192
rect 672318 168136 672323 168192
rect 666694 168134 672323 168136
rect 666694 168126 666754 168134
rect 672257 168131 672323 168134
rect 666356 168066 666754 168126
rect 683113 167922 683179 167925
rect 683100 167920 683179 167922
rect 683100 167864 683118 167920
rect 683174 167864 683179 167920
rect 683100 167862 683179 167864
rect 683113 167859 683179 167862
rect 675334 167452 675340 167516
rect 675404 167514 675410 167516
rect 675845 167514 675911 167517
rect 675404 167512 676292 167514
rect 675404 167456 675850 167512
rect 675906 167456 676292 167512
rect 675404 167454 676292 167456
rect 675404 167452 675410 167454
rect 675845 167451 675911 167454
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 676170 167046 676292 167106
rect 578233 166970 578299 166973
rect 575798 166968 578299 166970
rect 575798 166912 578238 166968
rect 578294 166912 578299 166968
rect 575798 166910 578299 166912
rect 575798 166532 575858 166910
rect 578233 166907 578299 166910
rect 672165 166970 672231 166973
rect 676170 166970 676230 167046
rect 672165 166968 676230 166970
rect 672165 166912 672170 166968
rect 672226 166912 676230 166968
rect 672165 166910 676230 166912
rect 672165 166907 672231 166910
rect 676397 166428 676463 166429
rect 676397 166424 676444 166428
rect 676508 166426 676514 166428
rect 676397 166368 676402 166424
rect 676397 166364 676444 166368
rect 676508 166366 676554 166426
rect 676508 166364 676514 166366
rect 676397 166363 676463 166364
rect 589457 165610 589523 165613
rect 589457 165608 592572 165610
rect 589457 165552 589462 165608
rect 589518 165552 592572 165608
rect 589457 165550 592572 165552
rect 589457 165547 589523 165550
rect 668025 164930 668091 164933
rect 666694 164928 668091 164930
rect 666694 164872 668030 164928
rect 668086 164872 668091 164928
rect 666694 164870 668091 164872
rect 666694 164862 666754 164870
rect 668025 164867 668091 164870
rect 666356 164802 666754 164862
rect 579521 164522 579587 164525
rect 575798 164520 579587 164522
rect 575798 164464 579526 164520
rect 579582 164464 579587 164520
rect 575798 164462 579587 164464
rect 575798 164356 575858 164462
rect 579521 164459 579587 164462
rect 589457 163978 589523 163981
rect 589457 163976 592572 163978
rect 589457 163920 589462 163976
rect 589518 163920 592572 163976
rect 589457 163918 592572 163920
rect 589457 163915 589523 163918
rect 668761 163298 668827 163301
rect 666694 163296 668827 163298
rect 666694 163240 668766 163296
rect 668822 163240 668827 163296
rect 666694 163238 668827 163240
rect 666694 163230 666754 163238
rect 668761 163235 668827 163238
rect 666356 163170 666754 163230
rect 579337 162754 579403 162757
rect 575798 162752 579403 162754
rect 575798 162696 579342 162752
rect 579398 162696 579403 162752
rect 575798 162694 579403 162696
rect 575798 162180 575858 162694
rect 579337 162691 579403 162694
rect 589457 162346 589523 162349
rect 668853 162346 668919 162349
rect 674097 162346 674163 162349
rect 589457 162344 592572 162346
rect 589457 162288 589462 162344
rect 589518 162288 592572 162344
rect 589457 162286 592572 162288
rect 668853 162344 674163 162346
rect 668853 162288 668858 162344
rect 668914 162288 674102 162344
rect 674158 162288 674163 162344
rect 668853 162286 674163 162288
rect 589457 162283 589523 162286
rect 668853 162283 668919 162286
rect 674097 162283 674163 162286
rect 674097 162074 674163 162077
rect 683113 162074 683179 162077
rect 674097 162072 683179 162074
rect 674097 162016 674102 162072
rect 674158 162016 683118 162072
rect 683174 162016 683179 162072
rect 674097 162014 683179 162016
rect 674097 162011 674163 162014
rect 683113 162011 683179 162014
rect 675017 161394 675083 161397
rect 676029 161394 676095 161397
rect 675017 161392 676095 161394
rect 675017 161336 675022 161392
rect 675078 161336 676034 161392
rect 676090 161336 676095 161392
rect 675017 161334 676095 161336
rect 675017 161331 675083 161334
rect 676029 161331 676095 161334
rect 673126 161060 673132 161124
rect 673196 161122 673202 161124
rect 675477 161122 675543 161125
rect 673196 161120 675543 161122
rect 673196 161064 675482 161120
rect 675538 161064 675543 161120
rect 673196 161062 675543 161064
rect 673196 161060 673202 161062
rect 675477 161059 675543 161062
rect 589457 160714 589523 160717
rect 589457 160712 592572 160714
rect 589457 160656 589462 160712
rect 589518 160656 592572 160712
rect 589457 160654 592572 160656
rect 589457 160651 589523 160654
rect 668209 160034 668275 160037
rect 666694 160032 668275 160034
rect 575982 159898 576042 160004
rect 666694 159976 668214 160032
rect 668270 159976 668275 160032
rect 666694 159974 668275 159976
rect 666694 159966 666754 159974
rect 668209 159971 668275 159974
rect 673545 160034 673611 160037
rect 675385 160034 675451 160037
rect 673545 160032 675451 160034
rect 673545 159976 673550 160032
rect 673606 159976 675390 160032
rect 675446 159976 675451 160032
rect 673545 159974 675451 159976
rect 673545 159971 673611 159974
rect 675385 159971 675451 159974
rect 666356 159906 666754 159966
rect 578233 159898 578299 159901
rect 575982 159896 578299 159898
rect 575982 159840 578238 159896
rect 578294 159840 578299 159896
rect 575982 159838 578299 159840
rect 578233 159835 578299 159838
rect 589457 159082 589523 159085
rect 668761 159082 668827 159085
rect 673729 159082 673795 159085
rect 589457 159080 592572 159082
rect 589457 159024 589462 159080
rect 589518 159024 592572 159080
rect 589457 159022 592572 159024
rect 668761 159080 673795 159082
rect 668761 159024 668766 159080
rect 668822 159024 673734 159080
rect 673790 159024 673795 159080
rect 668761 159022 673795 159024
rect 589457 159019 589523 159022
rect 668761 159019 668827 159022
rect 673729 159019 673795 159022
rect 578417 158402 578483 158405
rect 668761 158402 668827 158405
rect 575798 158400 578483 158402
rect 575798 158344 578422 158400
rect 578478 158344 578483 158400
rect 575798 158342 578483 158344
rect 575798 157828 575858 158342
rect 578417 158339 578483 158342
rect 666694 158400 668827 158402
rect 666694 158344 668766 158400
rect 668822 158344 668827 158400
rect 666694 158342 668827 158344
rect 666694 158334 666754 158342
rect 668761 158339 668827 158342
rect 666356 158274 666754 158334
rect 589273 157450 589339 157453
rect 589273 157448 592572 157450
rect 589273 157392 589278 157448
rect 589334 157392 592572 157448
rect 589273 157390 592572 157392
rect 589273 157387 589339 157390
rect 578877 155954 578943 155957
rect 575798 155952 578943 155954
rect 575798 155896 578882 155952
rect 578938 155896 578943 155952
rect 575798 155894 578943 155896
rect 575798 155652 575858 155894
rect 578877 155891 578943 155894
rect 589457 155818 589523 155821
rect 675753 155818 675819 155821
rect 676438 155818 676444 155820
rect 589457 155816 592572 155818
rect 589457 155760 589462 155816
rect 589518 155760 592572 155816
rect 589457 155758 592572 155760
rect 675753 155816 676444 155818
rect 675753 155760 675758 155816
rect 675814 155760 676444 155816
rect 675753 155758 676444 155760
rect 589457 155755 589523 155758
rect 675753 155755 675819 155758
rect 676438 155756 676444 155758
rect 676508 155756 676514 155820
rect 675385 155546 675451 155549
rect 676622 155546 676628 155548
rect 675385 155544 676628 155546
rect 675385 155488 675390 155544
rect 675446 155488 676628 155544
rect 675385 155486 676628 155488
rect 675385 155483 675451 155486
rect 676622 155484 676628 155486
rect 676692 155484 676698 155548
rect 668209 155138 668275 155141
rect 666694 155136 668275 155138
rect 666694 155080 668214 155136
rect 668270 155080 668275 155136
rect 666694 155078 668275 155080
rect 666694 155070 666754 155078
rect 668209 155075 668275 155078
rect 666356 155010 666754 155070
rect 669589 154458 669655 154461
rect 675109 154458 675175 154461
rect 669589 154456 675175 154458
rect 669589 154400 669594 154456
rect 669650 154400 675114 154456
rect 675170 154400 675175 154456
rect 669589 154398 675175 154400
rect 669589 154395 669655 154398
rect 675109 154395 675175 154398
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 578325 153642 578391 153645
rect 575798 153640 578391 153642
rect 575798 153584 578330 153640
rect 578386 153584 578391 153640
rect 575798 153582 578391 153584
rect 575798 153476 575858 153582
rect 578325 153579 578391 153582
rect 666356 153378 666938 153438
rect 666878 153370 666938 153378
rect 666878 153310 673470 153370
rect 673410 153234 673470 153310
rect 674281 153234 674347 153237
rect 673410 153232 674347 153234
rect 673410 153176 674286 153232
rect 674342 153176 674347 153232
rect 673410 153174 674347 153176
rect 674281 153171 674347 153174
rect 672349 152690 672415 152693
rect 675109 152690 675175 152693
rect 672349 152688 675175 152690
rect 672349 152632 672354 152688
rect 672410 152632 675114 152688
rect 675170 152632 675175 152688
rect 672349 152630 675175 152632
rect 672349 152627 672415 152630
rect 675109 152627 675175 152630
rect 589457 152554 589523 152557
rect 589457 152552 592572 152554
rect 589457 152496 589462 152552
rect 589518 152496 592572 152552
rect 589457 152494 592572 152496
rect 589457 152491 589523 152494
rect 578233 151738 578299 151741
rect 575798 151736 578299 151738
rect 575798 151680 578238 151736
rect 578294 151680 578299 151736
rect 575798 151678 578299 151680
rect 575798 151300 575858 151678
rect 578233 151675 578299 151678
rect 675753 151466 675819 151469
rect 676254 151466 676260 151468
rect 675753 151464 676260 151466
rect 675753 151408 675758 151464
rect 675814 151408 676260 151464
rect 675753 151406 676260 151408
rect 675753 151403 675819 151406
rect 676254 151404 676260 151406
rect 676324 151404 676330 151468
rect 673177 151330 673243 151333
rect 675109 151330 675175 151333
rect 673177 151328 675175 151330
rect 673177 151272 673182 151328
rect 673238 151272 675114 151328
rect 675170 151272 675175 151328
rect 673177 151270 675175 151272
rect 673177 151267 673243 151270
rect 675109 151267 675175 151270
rect 590009 150922 590075 150925
rect 590009 150920 592572 150922
rect 590009 150864 590014 150920
rect 590070 150864 592572 150920
rect 590009 150862 592572 150864
rect 590009 150859 590075 150862
rect 669773 150378 669839 150381
rect 674925 150378 674991 150381
rect 669773 150376 674991 150378
rect 669773 150320 669778 150376
rect 669834 150320 674930 150376
rect 674986 150320 674991 150376
rect 669773 150318 674991 150320
rect 669773 150315 669839 150318
rect 674925 150315 674991 150318
rect 666356 150114 666754 150174
rect 666694 150106 666754 150114
rect 671705 150106 671771 150109
rect 666694 150104 671771 150106
rect 666694 150048 671710 150104
rect 671766 150048 671771 150104
rect 666694 150046 671771 150048
rect 671705 150043 671771 150046
rect 578877 149698 578943 149701
rect 575798 149696 578943 149698
rect 575798 149640 578882 149696
rect 578938 149640 578943 149696
rect 575798 149638 578943 149640
rect 575798 149124 575858 149638
rect 578877 149635 578943 149638
rect 589457 149290 589523 149293
rect 589457 149288 592572 149290
rect 589457 149232 589462 149288
rect 589518 149232 592572 149288
rect 589457 149230 592572 149232
rect 589457 149227 589523 149230
rect 668853 148610 668919 148613
rect 666694 148608 668919 148610
rect 666694 148552 668858 148608
rect 668914 148552 668919 148608
rect 666694 148550 668919 148552
rect 666694 148542 666754 148550
rect 668853 148547 668919 148550
rect 666356 148482 666754 148542
rect 675753 148474 675819 148477
rect 676070 148474 676076 148476
rect 675753 148472 676076 148474
rect 675753 148416 675758 148472
rect 675814 148416 676076 148472
rect 675753 148414 676076 148416
rect 675753 148411 675819 148414
rect 676070 148412 676076 148414
rect 676140 148412 676146 148476
rect 588537 147658 588603 147661
rect 670601 147658 670667 147661
rect 675109 147658 675175 147661
rect 675385 147660 675451 147661
rect 588537 147656 592572 147658
rect 588537 147600 588542 147656
rect 588598 147600 592572 147656
rect 588537 147598 592572 147600
rect 670601 147656 675175 147658
rect 670601 147600 670606 147656
rect 670662 147600 675114 147656
rect 675170 147600 675175 147656
rect 670601 147598 675175 147600
rect 588537 147595 588603 147598
rect 670601 147595 670667 147598
rect 675109 147595 675175 147598
rect 675334 147596 675340 147660
rect 675404 147658 675451 147660
rect 675404 147656 675496 147658
rect 675446 147600 675496 147656
rect 675404 147598 675496 147600
rect 675404 147596 675451 147598
rect 675385 147595 675451 147596
rect 579521 147522 579587 147525
rect 575798 147520 579587 147522
rect 575798 147464 579526 147520
rect 579582 147464 579587 147520
rect 575798 147462 579587 147464
rect 575798 146948 575858 147462
rect 579521 147459 579587 147462
rect 589457 146026 589523 146029
rect 589457 146024 592572 146026
rect 589457 145968 589462 146024
rect 589518 145968 592572 146024
rect 589457 145966 592572 145968
rect 589457 145963 589523 145966
rect 668761 145346 668827 145349
rect 666694 145344 668827 145346
rect 666694 145288 668766 145344
rect 668822 145288 668827 145344
rect 666694 145286 668827 145288
rect 666694 145278 666754 145286
rect 668761 145283 668827 145286
rect 666356 145218 666754 145278
rect 671981 144938 672047 144941
rect 675109 144938 675175 144941
rect 671981 144936 675175 144938
rect 671981 144880 671986 144936
rect 672042 144880 675114 144936
rect 675170 144880 675175 144936
rect 671981 144878 675175 144880
rect 671981 144875 672047 144878
rect 675109 144875 675175 144878
rect 575982 144666 576042 144772
rect 579245 144666 579311 144669
rect 575982 144664 579311 144666
rect 575982 144608 579250 144664
rect 579306 144608 579311 144664
rect 575982 144606 579311 144608
rect 579245 144603 579311 144606
rect 589457 144394 589523 144397
rect 589457 144392 592572 144394
rect 589457 144336 589462 144392
rect 589518 144336 592572 144392
rect 589457 144334 592572 144336
rect 589457 144331 589523 144334
rect 668393 143714 668459 143717
rect 666694 143712 668459 143714
rect 666694 143656 668398 143712
rect 668454 143656 668459 143712
rect 666694 143654 668459 143656
rect 666694 143646 666754 143654
rect 668393 143651 668459 143654
rect 666356 143586 666754 143646
rect 579521 143034 579587 143037
rect 575798 143032 579587 143034
rect 575798 142976 579526 143032
rect 579582 142976 579587 143032
rect 575798 142974 579587 142976
rect 575798 142596 575858 142974
rect 579521 142971 579587 142974
rect 589825 142762 589891 142765
rect 589825 142760 592572 142762
rect 589825 142704 589830 142760
rect 589886 142704 592572 142760
rect 589825 142702 592572 142704
rect 589825 142699 589891 142702
rect 589457 141130 589523 141133
rect 589457 141128 592572 141130
rect 589457 141072 589462 141128
rect 589518 141072 592572 141128
rect 589457 141070 592572 141072
rect 589457 141067 589523 141070
rect 578601 140586 578667 140589
rect 575798 140584 578667 140586
rect 575798 140528 578606 140584
rect 578662 140528 578667 140584
rect 575798 140526 578667 140528
rect 575798 140420 575858 140526
rect 578601 140523 578667 140526
rect 669262 140450 669268 140452
rect 666694 140390 669268 140450
rect 666694 140382 666754 140390
rect 669262 140388 669268 140390
rect 669332 140388 669338 140452
rect 666356 140322 666754 140382
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 578601 138818 578667 138821
rect 668577 138818 668643 138821
rect 575798 138816 578667 138818
rect 575798 138760 578606 138816
rect 578662 138760 578667 138816
rect 575798 138758 578667 138760
rect 575798 138244 575858 138758
rect 578601 138755 578667 138758
rect 666694 138816 668643 138818
rect 666694 138760 668582 138816
rect 668638 138760 668643 138816
rect 666694 138758 668643 138760
rect 666694 138750 666754 138758
rect 668577 138755 668643 138758
rect 666356 138690 666754 138750
rect 589457 137866 589523 137869
rect 589457 137864 592572 137866
rect 589457 137808 589462 137864
rect 589518 137808 592572 137864
rect 589457 137806 592572 137808
rect 589457 137803 589523 137806
rect 578877 136642 578943 136645
rect 575798 136640 578943 136642
rect 575798 136584 578882 136640
rect 578938 136584 578943 136640
rect 575798 136582 578943 136584
rect 575798 136068 575858 136582
rect 578877 136579 578943 136582
rect 589457 136234 589523 136237
rect 589457 136232 592572 136234
rect 589457 136176 589462 136232
rect 589518 136176 592572 136232
rect 589457 136174 592572 136176
rect 589457 136171 589523 136174
rect 669037 135554 669103 135557
rect 666694 135552 669103 135554
rect 666694 135496 669042 135552
rect 669098 135496 669103 135552
rect 666694 135494 669103 135496
rect 666694 135486 666754 135494
rect 669037 135491 669103 135494
rect 666356 135426 666754 135486
rect 590377 134602 590443 134605
rect 667197 134602 667263 134605
rect 676029 134602 676095 134605
rect 590377 134600 592572 134602
rect 590377 134544 590382 134600
rect 590438 134544 592572 134600
rect 590377 134542 592572 134544
rect 667197 134600 676095 134602
rect 667197 134544 667202 134600
rect 667258 134544 676034 134600
rect 676090 134544 676095 134600
rect 667197 134542 676095 134544
rect 590377 134539 590443 134542
rect 667197 134539 667263 134542
rect 676029 134539 676095 134542
rect 579521 134466 579587 134469
rect 575798 134464 579587 134466
rect 575798 134408 579526 134464
rect 579582 134408 579587 134464
rect 575798 134406 579587 134408
rect 575798 133892 575858 134406
rect 579521 134403 579587 134406
rect 666356 133794 666754 133854
rect 666694 133786 666754 133794
rect 667933 133786 667999 133789
rect 666694 133784 667999 133786
rect 666694 133728 667938 133784
rect 667994 133728 667999 133784
rect 666694 133726 667999 133728
rect 667933 133723 667999 133726
rect 672533 133378 672599 133381
rect 672533 133376 676292 133378
rect 672533 133320 672538 133376
rect 672594 133320 676292 133376
rect 672533 133318 676292 133320
rect 672533 133315 672599 133318
rect 589457 132970 589523 132973
rect 589457 132968 592572 132970
rect 589457 132912 589462 132968
rect 589518 132912 592572 132968
rect 589457 132910 592572 132912
rect 589457 132907 589523 132910
rect 667790 132908 667796 132972
rect 667860 132970 667866 132972
rect 667860 132910 676292 132970
rect 667860 132908 667866 132910
rect 667013 132698 667079 132701
rect 672533 132698 672599 132701
rect 667013 132696 672599 132698
rect 667013 132640 667018 132696
rect 667074 132640 672538 132696
rect 672594 132640 672599 132696
rect 667013 132638 672599 132640
rect 667013 132635 667079 132638
rect 672533 132635 672599 132638
rect 676029 132562 676095 132565
rect 676029 132560 676292 132562
rect 676029 132504 676034 132560
rect 676090 132504 676292 132560
rect 676029 132502 676292 132504
rect 676029 132499 676095 132502
rect 579061 132290 579127 132293
rect 575798 132288 579127 132290
rect 575798 132232 579066 132288
rect 579122 132232 579127 132288
rect 575798 132230 579127 132232
rect 575798 131716 575858 132230
rect 579061 132227 579127 132230
rect 673913 132154 673979 132157
rect 673913 132152 676292 132154
rect 673913 132096 673918 132152
rect 673974 132096 676292 132152
rect 673913 132094 676292 132096
rect 673913 132091 673979 132094
rect 672533 131746 672599 131749
rect 672533 131744 676292 131746
rect 672533 131688 672538 131744
rect 672594 131688 676292 131744
rect 672533 131686 676292 131688
rect 672533 131683 672599 131686
rect 589457 131338 589523 131341
rect 674649 131338 674715 131341
rect 589457 131336 592572 131338
rect 589457 131280 589462 131336
rect 589518 131280 592572 131336
rect 589457 131278 592572 131280
rect 674649 131336 676292 131338
rect 674649 131280 674654 131336
rect 674710 131280 676292 131336
rect 674649 131278 676292 131280
rect 589457 131275 589523 131278
rect 674649 131275 674715 131278
rect 668853 131202 668919 131205
rect 672349 131202 672415 131205
rect 668853 131200 672415 131202
rect 668853 131144 668858 131200
rect 668914 131144 672354 131200
rect 672410 131144 672415 131200
rect 668853 131142 672415 131144
rect 668853 131139 668919 131142
rect 672349 131139 672415 131142
rect 671337 130930 671403 130933
rect 671337 130928 676292 130930
rect 671337 130872 671342 130928
rect 671398 130872 676292 130928
rect 671337 130870 676292 130872
rect 671337 130867 671403 130870
rect 668669 130658 668735 130661
rect 666694 130656 668735 130658
rect 666694 130600 668674 130656
rect 668730 130600 668735 130656
rect 666694 130598 668735 130600
rect 666694 130590 666754 130598
rect 668669 130595 668735 130598
rect 666356 130530 666754 130590
rect 674465 130522 674531 130525
rect 674465 130520 676292 130522
rect 674465 130464 674470 130520
rect 674526 130464 676292 130520
rect 674465 130462 676292 130464
rect 674465 130459 674531 130462
rect 676213 130250 676279 130253
rect 676213 130248 676322 130250
rect 676213 130192 676218 130248
rect 676274 130192 676322 130248
rect 676213 130187 676322 130192
rect 676262 130084 676322 130187
rect 578877 129706 578943 129709
rect 575798 129704 578943 129706
rect 575798 129648 578882 129704
rect 578938 129648 578943 129704
rect 575798 129646 578943 129648
rect 575798 129540 575858 129646
rect 578877 129643 578943 129646
rect 588537 129706 588603 129709
rect 673361 129706 673427 129709
rect 588537 129704 592572 129706
rect 588537 129648 588542 129704
rect 588598 129648 592572 129704
rect 588537 129646 592572 129648
rect 673361 129704 676292 129706
rect 673361 129648 673366 129704
rect 673422 129648 676292 129704
rect 673361 129646 676292 129648
rect 588537 129643 588603 129646
rect 673361 129643 673427 129646
rect 669957 129298 670023 129301
rect 669957 129296 676292 129298
rect 669957 129240 669962 129296
rect 670018 129240 676292 129296
rect 669957 129238 676292 129240
rect 669957 129235 670023 129238
rect 667933 129026 667999 129029
rect 666694 129024 667999 129026
rect 666694 128968 667938 129024
rect 667994 128968 667999 129024
rect 666694 128966 667999 128968
rect 666694 128958 666754 128966
rect 667933 128963 667999 128966
rect 666356 128898 666754 128958
rect 675845 128890 675911 128893
rect 675845 128888 676292 128890
rect 675845 128832 675850 128888
rect 675906 128832 676292 128888
rect 675845 128830 676292 128832
rect 675845 128827 675911 128830
rect 673177 128482 673243 128485
rect 673177 128480 676292 128482
rect 673177 128424 673182 128480
rect 673238 128424 676292 128480
rect 673177 128422 676292 128424
rect 673177 128419 673243 128422
rect 589457 128074 589523 128077
rect 589457 128072 592572 128074
rect 589457 128016 589462 128072
rect 589518 128016 592572 128072
rect 589457 128014 592572 128016
rect 589457 128011 589523 128014
rect 579521 127938 579587 127941
rect 575798 127936 579587 127938
rect 575798 127880 579526 127936
rect 579582 127880 579587 127936
rect 575798 127878 579587 127880
rect 575798 127364 575858 127878
rect 579521 127875 579587 127878
rect 676446 127805 676506 128044
rect 668577 127802 668643 127805
rect 676213 127802 676279 127805
rect 668577 127800 676279 127802
rect 668577 127744 668582 127800
rect 668638 127744 676218 127800
rect 676274 127744 676279 127800
rect 668577 127742 676279 127744
rect 668577 127739 668643 127742
rect 676213 127739 676279 127742
rect 676397 127800 676506 127805
rect 676397 127744 676402 127800
rect 676458 127744 676506 127800
rect 676397 127742 676506 127744
rect 676397 127739 676463 127742
rect 676446 127396 676506 127636
rect 676438 127332 676444 127396
rect 676508 127332 676514 127396
rect 668393 126986 668459 126989
rect 672901 126986 672967 126989
rect 668393 126984 672967 126986
rect 668393 126928 668398 126984
rect 668454 126928 672906 126984
rect 672962 126928 672967 126984
rect 668393 126926 672967 126928
rect 668393 126923 668459 126926
rect 672901 126923 672967 126926
rect 676070 126924 676076 126988
rect 676140 126986 676146 126988
rect 676262 126986 676322 127228
rect 676140 126926 676322 126986
rect 676140 126924 676146 126926
rect 671981 126578 672047 126581
rect 676262 126578 676322 126820
rect 671981 126576 676322 126578
rect 671981 126520 671986 126576
rect 672042 126520 676322 126576
rect 671981 126518 676322 126520
rect 671981 126515 672047 126518
rect 589917 126442 589983 126445
rect 589917 126440 592572 126442
rect 589917 126384 589922 126440
rect 589978 126384 592572 126440
rect 589917 126382 592572 126384
rect 589917 126379 589983 126382
rect 682334 126173 682394 126412
rect 682334 126168 682443 126173
rect 682334 126112 682382 126168
rect 682438 126112 682443 126168
rect 682334 126110 682443 126112
rect 682377 126107 682443 126110
rect 683254 125765 683314 126004
rect 669221 125762 669287 125765
rect 666694 125760 669287 125762
rect 666694 125704 669226 125760
rect 669282 125704 669287 125760
rect 666694 125702 669287 125704
rect 683254 125760 683363 125765
rect 683254 125704 683302 125760
rect 683358 125704 683363 125760
rect 683254 125702 683363 125704
rect 666694 125694 666754 125702
rect 669221 125699 669287 125702
rect 683297 125699 683363 125702
rect 666356 125634 666754 125694
rect 681046 125357 681106 125596
rect 578325 125354 578391 125357
rect 575798 125352 578391 125354
rect 575798 125296 578330 125352
rect 578386 125296 578391 125352
rect 575798 125294 578391 125296
rect 575798 125188 575858 125294
rect 578325 125291 578391 125294
rect 680997 125352 681106 125357
rect 680997 125296 681002 125352
rect 681058 125296 681106 125352
rect 680997 125294 681106 125296
rect 680997 125291 681063 125294
rect 674373 125218 674439 125221
rect 674373 125216 676292 125218
rect 674373 125160 674378 125216
rect 674434 125160 676292 125216
rect 674373 125158 676292 125160
rect 674373 125155 674439 125158
rect 589457 124810 589523 124813
rect 673913 124810 673979 124813
rect 589457 124808 592572 124810
rect 589457 124752 589462 124808
rect 589518 124752 592572 124808
rect 589457 124750 592572 124752
rect 673913 124808 676292 124810
rect 673913 124752 673918 124808
rect 673974 124752 676292 124808
rect 673913 124750 676292 124752
rect 589457 124747 589523 124750
rect 673913 124747 673979 124750
rect 676254 124476 676260 124540
rect 676324 124476 676330 124540
rect 676262 124372 676322 124476
rect 672717 124130 672783 124133
rect 666694 124128 672783 124130
rect 666694 124072 672722 124128
rect 672778 124072 672783 124128
rect 666694 124070 672783 124072
rect 666694 124062 666754 124070
rect 672717 124067 672783 124070
rect 666356 124002 666754 124062
rect 672950 123934 676292 123994
rect 672717 123858 672783 123861
rect 672950 123858 673010 123934
rect 672717 123856 673010 123858
rect 672717 123800 672722 123856
rect 672778 123800 673010 123856
rect 672717 123798 673010 123800
rect 672717 123795 672783 123798
rect 578417 123586 578483 123589
rect 575798 123584 578483 123586
rect 575798 123528 578422 123584
rect 578478 123528 578483 123584
rect 575798 123526 578483 123528
rect 575798 123012 575858 123526
rect 578417 123523 578483 123526
rect 674649 123586 674715 123589
rect 674649 123584 676292 123586
rect 674649 123528 674654 123584
rect 674710 123528 676292 123584
rect 674649 123526 676292 123528
rect 674649 123523 674715 123526
rect 589457 123178 589523 123181
rect 672901 123178 672967 123181
rect 589457 123176 592572 123178
rect 589457 123120 589462 123176
rect 589518 123120 592572 123176
rect 589457 123118 592572 123120
rect 672901 123176 676292 123178
rect 672901 123120 672906 123176
rect 672962 123120 676292 123176
rect 672901 123118 676292 123120
rect 589457 123115 589523 123118
rect 672901 123115 672967 123118
rect 670141 122770 670207 122773
rect 670141 122768 676292 122770
rect 670141 122712 670146 122768
rect 670202 122712 676292 122768
rect 670141 122710 676292 122712
rect 670141 122707 670207 122710
rect 675334 122300 675340 122364
rect 675404 122362 675410 122364
rect 675404 122302 676292 122362
rect 675404 122300 675410 122302
rect 676262 121682 676322 121924
rect 675894 121622 676322 121682
rect 590009 121546 590075 121549
rect 590009 121544 592572 121546
rect 590009 121488 590014 121544
rect 590070 121488 592572 121544
rect 590009 121486 592572 121488
rect 590009 121483 590075 121486
rect 578877 121410 578943 121413
rect 575798 121408 578943 121410
rect 575798 121352 578882 121408
rect 578938 121352 578943 121408
rect 575798 121350 578943 121352
rect 575798 120836 575858 121350
rect 578877 121347 578943 121350
rect 668393 120866 668459 120869
rect 666694 120864 668459 120866
rect 666694 120808 668398 120864
rect 668454 120808 668459 120864
rect 666694 120806 668459 120808
rect 666694 120798 666754 120806
rect 668393 120803 668459 120806
rect 666356 120738 666754 120798
rect 668945 120730 669011 120733
rect 675894 120730 675954 121622
rect 668945 120728 675954 120730
rect 668945 120672 668950 120728
rect 669006 120672 675954 120728
rect 668945 120670 675954 120672
rect 668945 120667 669011 120670
rect 676806 119988 676812 120052
rect 676876 120050 676882 120052
rect 683297 120050 683363 120053
rect 676876 120048 683363 120050
rect 676876 119992 683302 120048
rect 683358 119992 683363 120048
rect 676876 119990 683363 119992
rect 676876 119988 676882 119990
rect 683297 119987 683363 119990
rect 589641 119914 589707 119917
rect 589641 119912 592572 119914
rect 589641 119856 589646 119912
rect 589702 119856 592572 119912
rect 589641 119854 592572 119856
rect 589641 119851 589707 119854
rect 668761 119234 668827 119237
rect 666694 119232 668827 119234
rect 666694 119176 668766 119232
rect 668822 119176 668827 119232
rect 666694 119174 668827 119176
rect 666694 119166 666754 119174
rect 668761 119171 668827 119174
rect 666356 119106 666754 119166
rect 575982 118418 576042 118660
rect 578509 118418 578575 118421
rect 575982 118416 578575 118418
rect 575982 118360 578514 118416
rect 578570 118360 578575 118416
rect 575982 118358 578575 118360
rect 578509 118355 578575 118358
rect 590101 118282 590167 118285
rect 590101 118280 592572 118282
rect 590101 118224 590106 118280
rect 590162 118224 592572 118280
rect 590101 118222 592572 118224
rect 590101 118219 590167 118222
rect 666356 117474 666938 117534
rect 666878 117466 666938 117474
rect 674097 117466 674163 117469
rect 666878 117464 674163 117466
rect 666878 117408 674102 117464
rect 674158 117408 674163 117464
rect 666878 117406 674163 117408
rect 674097 117403 674163 117406
rect 675702 117268 675708 117332
rect 675772 117330 675778 117332
rect 680997 117330 681063 117333
rect 675772 117328 681063 117330
rect 675772 117272 681002 117328
rect 681058 117272 681063 117328
rect 675772 117270 681063 117272
rect 675772 117268 675778 117270
rect 680997 117267 681063 117270
rect 579521 116922 579587 116925
rect 575798 116920 579587 116922
rect 575798 116864 579526 116920
rect 579582 116864 579587 116920
rect 575798 116862 579587 116864
rect 575798 116484 575858 116862
rect 579521 116859 579587 116862
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 682377 116106 682443 116109
rect 675342 116104 682443 116106
rect 675342 116048 682382 116104
rect 682438 116048 682443 116104
rect 675342 116046 682443 116048
rect 666356 115842 666754 115902
rect 666694 115834 666754 115842
rect 675342 115837 675402 116046
rect 682377 116043 682443 116046
rect 672165 115834 672231 115837
rect 666694 115832 672231 115834
rect 666694 115776 672170 115832
rect 672226 115776 672231 115832
rect 666694 115774 672231 115776
rect 672165 115771 672231 115774
rect 675293 115832 675402 115837
rect 675293 115776 675298 115832
rect 675354 115776 675402 115832
rect 675293 115774 675402 115776
rect 675293 115771 675359 115774
rect 675017 115290 675083 115293
rect 675385 115290 675451 115293
rect 675017 115288 675451 115290
rect 675017 115232 675022 115288
rect 675078 115232 675390 115288
rect 675446 115232 675451 115288
rect 675017 115230 675451 115232
rect 675017 115227 675083 115230
rect 675385 115227 675451 115230
rect 675753 115288 675819 115293
rect 675753 115232 675758 115288
rect 675814 115232 675819 115288
rect 675753 115227 675819 115232
rect 590285 115018 590351 115021
rect 590285 115016 592572 115018
rect 590285 114960 590290 115016
rect 590346 114960 592572 115016
rect 590285 114958 592572 114960
rect 590285 114955 590351 114958
rect 674046 114956 674052 115020
rect 674116 115018 674122 115020
rect 675756 115018 675816 115227
rect 674116 114958 675816 115018
rect 674116 114956 674122 114958
rect 579245 114474 579311 114477
rect 575798 114472 579311 114474
rect 575798 114416 579250 114472
rect 579306 114416 579311 114472
rect 575798 114414 579311 114416
rect 575798 114308 575858 114414
rect 579245 114411 579311 114414
rect 672901 114338 672967 114341
rect 666694 114336 672967 114338
rect 666694 114280 672906 114336
rect 672962 114280 672967 114336
rect 666694 114278 672967 114280
rect 666694 114270 666754 114278
rect 672901 114275 672967 114278
rect 666356 114210 666754 114270
rect 589457 113386 589523 113389
rect 589457 113384 592572 113386
rect 589457 113328 589462 113384
rect 589518 113328 592572 113384
rect 589457 113326 592572 113328
rect 589457 113323 589523 113326
rect 668117 112706 668183 112709
rect 666694 112704 668183 112706
rect 666694 112648 668122 112704
rect 668178 112648 668183 112704
rect 666694 112646 668183 112648
rect 666694 112638 666754 112646
rect 668117 112643 668183 112646
rect 666356 112578 666754 112638
rect 579521 112570 579587 112573
rect 575798 112568 579587 112570
rect 575798 112512 579526 112568
rect 579582 112512 579587 112568
rect 575798 112510 579587 112512
rect 575798 112132 575858 112510
rect 579521 112507 579587 112510
rect 675753 112434 675819 112437
rect 676438 112434 676444 112436
rect 675753 112432 676444 112434
rect 675753 112376 675758 112432
rect 675814 112376 676444 112432
rect 675753 112374 676444 112376
rect 675753 112371 675819 112374
rect 676438 112372 676444 112374
rect 676508 112372 676514 112436
rect 589457 111754 589523 111757
rect 675753 111754 675819 111757
rect 676806 111754 676812 111756
rect 589457 111752 592572 111754
rect 589457 111696 589462 111752
rect 589518 111696 592572 111752
rect 589457 111694 592572 111696
rect 675753 111752 676812 111754
rect 675753 111696 675758 111752
rect 675814 111696 676812 111752
rect 675753 111694 676812 111696
rect 589457 111691 589523 111694
rect 675753 111691 675819 111694
rect 676806 111692 676812 111694
rect 676876 111692 676882 111756
rect 675753 111348 675819 111349
rect 675702 111284 675708 111348
rect 675772 111346 675819 111348
rect 675772 111344 675864 111346
rect 675814 111288 675864 111344
rect 675772 111286 675864 111288
rect 675772 111284 675819 111286
rect 675753 111283 675819 111284
rect 668945 111074 669011 111077
rect 666694 111072 669011 111074
rect 666694 111016 668950 111072
rect 669006 111016 669011 111072
rect 666694 111014 669011 111016
rect 666694 111006 666754 111014
rect 668945 111011 669011 111014
rect 666356 110946 666754 111006
rect 675753 110394 675819 110397
rect 676254 110394 676260 110396
rect 675753 110392 676260 110394
rect 675753 110336 675758 110392
rect 675814 110336 676260 110392
rect 675753 110334 676260 110336
rect 675753 110331 675819 110334
rect 676254 110332 676260 110334
rect 676324 110332 676330 110396
rect 579337 110122 579403 110125
rect 575798 110120 579403 110122
rect 575798 110064 579342 110120
rect 579398 110064 579403 110120
rect 575798 110062 579403 110064
rect 575798 109956 575858 110062
rect 579337 110059 579403 110062
rect 589273 110122 589339 110125
rect 589273 110120 592572 110122
rect 589273 110064 589278 110120
rect 589334 110064 592572 110120
rect 589273 110062 592572 110064
rect 589273 110059 589339 110062
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 578325 108354 578391 108357
rect 575798 108352 578391 108354
rect 575798 108296 578330 108352
rect 578386 108296 578391 108352
rect 575798 108294 578391 108296
rect 575798 107780 575858 108294
rect 578325 108291 578391 108294
rect 675753 108218 675819 108221
rect 676070 108218 676076 108220
rect 675753 108216 676076 108218
rect 675753 108160 675758 108216
rect 675814 108160 676076 108216
rect 675753 108158 676076 108160
rect 675753 108155 675819 108158
rect 676070 108156 676076 108158
rect 676140 108156 676146 108220
rect 668393 107810 668459 107813
rect 666694 107808 668459 107810
rect 666694 107752 668398 107808
rect 668454 107752 668459 107808
rect 666694 107750 668459 107752
rect 666694 107742 666754 107750
rect 668393 107747 668459 107750
rect 666356 107682 666754 107742
rect 673913 106994 673979 106997
rect 675385 106994 675451 106997
rect 673913 106992 675451 106994
rect 673913 106936 673918 106992
rect 673974 106936 675390 106992
rect 675446 106936 675451 106992
rect 673913 106934 675451 106936
rect 673913 106931 673979 106934
rect 675385 106931 675451 106934
rect 589825 106858 589891 106861
rect 589825 106856 592572 106858
rect 589825 106800 589830 106856
rect 589886 106800 592572 106856
rect 589825 106798 592572 106800
rect 589825 106795 589891 106798
rect 672717 106314 672783 106317
rect 675109 106314 675175 106317
rect 672717 106312 675175 106314
rect 672717 106256 672722 106312
rect 672778 106256 675114 106312
rect 675170 106256 675175 106312
rect 672717 106254 675175 106256
rect 672717 106251 672783 106254
rect 675109 106251 675175 106254
rect 672349 106178 672415 106181
rect 666694 106176 672415 106178
rect 666694 106120 672354 106176
rect 672410 106120 672415 106176
rect 666694 106118 672415 106120
rect 666694 106110 666754 106118
rect 672349 106115 672415 106118
rect 666356 106050 666754 106110
rect 579061 105906 579127 105909
rect 575798 105904 579127 105906
rect 575798 105848 579066 105904
rect 579122 105848 579127 105904
rect 575798 105846 579127 105848
rect 575798 105604 575858 105846
rect 579061 105843 579127 105846
rect 589457 105226 589523 105229
rect 589457 105224 592572 105226
rect 589457 105168 589462 105224
rect 589518 105168 592572 105224
rect 589457 105166 592572 105168
rect 589457 105163 589523 105166
rect 667933 104546 667999 104549
rect 666694 104544 667999 104546
rect 666694 104488 667938 104544
rect 667994 104488 667999 104544
rect 666694 104486 667999 104488
rect 666694 104478 666754 104486
rect 667933 104483 667999 104486
rect 666356 104418 666754 104478
rect 588721 103594 588787 103597
rect 588721 103592 592572 103594
rect 588721 103536 588726 103592
rect 588782 103536 592572 103592
rect 588721 103534 592572 103536
rect 588721 103531 588787 103534
rect 673361 103458 673427 103461
rect 675109 103458 675175 103461
rect 673361 103456 675175 103458
rect 575982 103322 576042 103428
rect 673361 103400 673366 103456
rect 673422 103400 675114 103456
rect 675170 103400 675175 103456
rect 673361 103398 675175 103400
rect 673361 103395 673427 103398
rect 675109 103395 675175 103398
rect 579521 103322 579587 103325
rect 575982 103320 579587 103322
rect 575982 103264 579526 103320
rect 579582 103264 579587 103320
rect 575982 103262 579587 103264
rect 579521 103259 579587 103262
rect 668577 102914 668643 102917
rect 666694 102912 668643 102914
rect 666694 102856 668582 102912
rect 668638 102856 668643 102912
rect 666694 102854 668643 102856
rect 666694 102846 666754 102854
rect 668577 102851 668643 102854
rect 666356 102786 666754 102846
rect 589457 101962 589523 101965
rect 675385 101964 675451 101965
rect 675334 101962 675340 101964
rect 589457 101960 592572 101962
rect 589457 101904 589462 101960
rect 589518 101904 592572 101960
rect 589457 101902 592572 101904
rect 673410 101902 675340 101962
rect 675404 101962 675451 101964
rect 675404 101960 675496 101962
rect 675446 101904 675496 101960
rect 589457 101899 589523 101902
rect 673410 101826 673470 101902
rect 675334 101900 675340 101902
rect 675404 101902 675496 101904
rect 675404 101900 675451 101902
rect 675385 101899 675451 101900
rect 596130 101766 673470 101826
rect 579521 101690 579587 101693
rect 575798 101688 579587 101690
rect 575798 101632 579526 101688
rect 579582 101632 579587 101688
rect 575798 101630 579587 101632
rect 575798 101252 575858 101630
rect 579521 101627 579587 101630
rect 591481 101690 591547 101693
rect 596130 101690 596190 101766
rect 591481 101688 596190 101690
rect 591481 101632 591486 101688
rect 591542 101632 596190 101688
rect 591481 101630 596190 101632
rect 591481 101627 591547 101630
rect 671981 99378 672047 99381
rect 675293 99378 675359 99381
rect 671981 99376 675359 99378
rect 671981 99320 671986 99376
rect 672042 99320 675298 99376
rect 675354 99320 675359 99376
rect 671981 99318 675359 99320
rect 671981 99315 672047 99318
rect 675293 99315 675359 99318
rect 578601 99242 578667 99245
rect 575798 99240 578667 99242
rect 575798 99184 578606 99240
rect 578662 99184 578667 99240
rect 575798 99182 578667 99184
rect 575798 99076 575858 99182
rect 578601 99179 578667 99182
rect 578325 97474 578391 97477
rect 575798 97472 578391 97474
rect 575798 97416 578330 97472
rect 578386 97416 578391 97472
rect 575798 97414 578391 97416
rect 575798 96900 575858 97414
rect 578325 97411 578391 97414
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 641989 96522 642055 96525
rect 647182 96522 647188 96524
rect 641989 96520 647188 96522
rect 641989 96464 641994 96520
rect 642050 96464 647188 96520
rect 641989 96462 647188 96464
rect 641989 96459 642055 96462
rect 647182 96460 647188 96462
rect 647252 96460 647258 96524
rect 633934 95372 633940 95436
rect 634004 95434 634010 95436
rect 635733 95434 635799 95437
rect 634004 95432 635799 95434
rect 634004 95376 635738 95432
rect 635794 95376 635799 95432
rect 634004 95374 635799 95376
rect 634004 95372 634010 95374
rect 635733 95371 635799 95374
rect 579521 95026 579587 95029
rect 575798 95024 579587 95026
rect 575798 94968 579526 95024
rect 579582 94968 579587 95024
rect 575798 94966 579587 94968
rect 575798 94724 575858 94966
rect 579521 94963 579587 94966
rect 647141 95026 647207 95029
rect 647141 95024 647434 95026
rect 647141 94968 647146 95024
rect 647202 94968 647434 95024
rect 647141 94966 647434 94968
rect 647141 94963 647207 94966
rect 626441 94482 626507 94485
rect 626441 94480 628268 94482
rect 626441 94424 626446 94480
rect 626502 94424 628268 94480
rect 647374 94452 647434 94966
rect 626441 94422 628268 94424
rect 626441 94419 626507 94422
rect 654593 94210 654659 94213
rect 654593 94208 656788 94210
rect 654593 94152 654598 94208
rect 654654 94152 656788 94208
rect 654593 94150 656788 94152
rect 654593 94147 654659 94150
rect 626257 93666 626323 93669
rect 626257 93664 628268 93666
rect 626257 93608 626262 93664
rect 626318 93608 628268 93664
rect 626257 93606 628268 93608
rect 626257 93603 626323 93606
rect 655421 93394 655487 93397
rect 665173 93394 665239 93397
rect 655421 93392 656788 93394
rect 655421 93336 655426 93392
rect 655482 93336 656788 93392
rect 655421 93334 656788 93336
rect 663596 93392 665239 93394
rect 663596 93336 665178 93392
rect 665234 93336 665239 93392
rect 663596 93334 665239 93336
rect 655421 93331 655487 93334
rect 665173 93331 665239 93334
rect 578509 93122 578575 93125
rect 575798 93120 578575 93122
rect 575798 93064 578514 93120
rect 578570 93064 578575 93120
rect 575798 93062 578575 93064
rect 575798 92548 575858 93062
rect 578509 93059 578575 93062
rect 650310 93060 650316 93124
rect 650380 93122 650386 93124
rect 650380 93062 656818 93122
rect 650380 93060 650386 93062
rect 626441 92850 626507 92853
rect 626441 92848 628268 92850
rect 626441 92792 626446 92848
rect 626502 92792 628268 92848
rect 626441 92790 628268 92792
rect 626441 92787 626507 92790
rect 656758 92548 656818 93062
rect 663701 92850 663767 92853
rect 663382 92848 663767 92850
rect 663382 92792 663706 92848
rect 663762 92792 663767 92848
rect 663382 92790 663767 92792
rect 663382 92548 663442 92790
rect 663701 92787 663767 92790
rect 647509 92442 647575 92445
rect 647509 92440 647618 92442
rect 647509 92384 647514 92440
rect 647570 92384 647618 92440
rect 647509 92379 647618 92384
rect 625797 92034 625863 92037
rect 625797 92032 628268 92034
rect 625797 91976 625802 92032
rect 625858 91976 628268 92032
rect 647558 92004 647618 92379
rect 625797 91974 628268 91976
rect 625797 91971 625863 91974
rect 665357 91762 665423 91765
rect 663596 91760 665423 91762
rect 663596 91704 665362 91760
rect 665418 91704 665423 91760
rect 663596 91702 665423 91704
rect 665357 91699 665423 91702
rect 654317 91490 654383 91493
rect 654317 91488 656788 91490
rect 654317 91432 654322 91488
rect 654378 91432 656788 91488
rect 654317 91430 656788 91432
rect 654317 91427 654383 91430
rect 626441 91218 626507 91221
rect 626441 91216 628268 91218
rect 626441 91160 626446 91216
rect 626502 91160 628268 91216
rect 626441 91158 628268 91160
rect 626441 91155 626507 91158
rect 579061 90946 579127 90949
rect 575798 90944 579127 90946
rect 575798 90888 579066 90944
rect 579122 90888 579127 90944
rect 575798 90886 579127 90888
rect 575798 90372 575858 90886
rect 579061 90883 579127 90886
rect 655421 90674 655487 90677
rect 665541 90674 665607 90677
rect 655421 90672 656788 90674
rect 655421 90616 655426 90672
rect 655482 90616 656788 90672
rect 655421 90614 656788 90616
rect 663596 90672 665607 90674
rect 663596 90616 665546 90672
rect 665602 90616 665607 90672
rect 663596 90614 665607 90616
rect 655421 90611 655487 90614
rect 665541 90611 665607 90614
rect 626441 90402 626507 90405
rect 626441 90400 628268 90402
rect 626441 90344 626446 90400
rect 626502 90344 628268 90400
rect 626441 90342 628268 90344
rect 626441 90339 626507 90342
rect 655789 89858 655855 89861
rect 664161 89858 664227 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 655789 89798 656788 89800
rect 663596 89856 664227 89858
rect 663596 89800 664166 89856
rect 664222 89800 664227 89856
rect 663596 89798 664227 89800
rect 655789 89795 655855 89798
rect 664161 89795 664227 89798
rect 626441 89586 626507 89589
rect 648245 89586 648311 89589
rect 626441 89584 628268 89586
rect 626441 89528 626446 89584
rect 626502 89528 628268 89584
rect 626441 89526 628268 89528
rect 648140 89584 648311 89586
rect 648140 89528 648250 89584
rect 648306 89528 648311 89584
rect 648140 89526 648311 89528
rect 626441 89523 626507 89526
rect 648245 89523 648311 89526
rect 664345 89042 664411 89045
rect 663596 89040 664411 89042
rect 663596 88984 664350 89040
rect 664406 88984 664411 89040
rect 663596 88982 664411 88984
rect 664345 88979 664411 88982
rect 624969 88362 625035 88365
rect 628238 88362 628298 88740
rect 624969 88360 628298 88362
rect 624969 88304 624974 88360
rect 625030 88304 628298 88360
rect 624969 88302 628298 88304
rect 624969 88299 625035 88302
rect 575982 88090 576042 88196
rect 579521 88090 579587 88093
rect 575982 88088 579587 88090
rect 575982 88032 579526 88088
rect 579582 88032 579587 88088
rect 575982 88030 579587 88032
rect 579521 88027 579587 88030
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 626257 87138 626323 87141
rect 649993 87138 650059 87141
rect 626257 87136 628268 87138
rect 626257 87080 626262 87136
rect 626318 87080 628268 87136
rect 626257 87078 628268 87080
rect 648140 87136 650059 87138
rect 648140 87080 649998 87136
rect 650054 87080 650059 87136
rect 648140 87078 650059 87080
rect 626257 87075 626323 87078
rect 649993 87075 650059 87078
rect 579337 86458 579403 86461
rect 575798 86456 579403 86458
rect 575798 86400 579342 86456
rect 579398 86400 579403 86456
rect 575798 86398 579403 86400
rect 575798 86020 575858 86398
rect 579337 86395 579403 86398
rect 626441 86322 626507 86325
rect 626441 86320 628268 86322
rect 626441 86264 626446 86320
rect 626502 86264 628268 86320
rect 626441 86262 628268 86264
rect 626441 86259 626507 86262
rect 625337 85506 625403 85509
rect 625337 85504 628268 85506
rect 625337 85448 625342 85504
rect 625398 85448 628268 85504
rect 625337 85446 628268 85448
rect 625337 85443 625403 85446
rect 626441 84690 626507 84693
rect 650545 84690 650611 84693
rect 626441 84688 628268 84690
rect 626441 84632 626446 84688
rect 626502 84632 628268 84688
rect 626441 84630 628268 84632
rect 648140 84688 650611 84690
rect 648140 84632 650550 84688
rect 650606 84632 650611 84688
rect 648140 84630 650611 84632
rect 626441 84627 626507 84630
rect 650545 84627 650611 84630
rect 579153 84010 579219 84013
rect 575798 84008 579219 84010
rect 575798 83952 579158 84008
rect 579214 83952 579219 84008
rect 575798 83950 579219 83952
rect 575798 83844 575858 83950
rect 579153 83947 579219 83950
rect 625797 83874 625863 83877
rect 625797 83872 628268 83874
rect 625797 83816 625802 83872
rect 625858 83816 628268 83872
rect 625797 83814 628268 83816
rect 625797 83811 625863 83814
rect 628741 83330 628807 83333
rect 628741 83328 628850 83330
rect 628741 83272 628746 83328
rect 628802 83272 628850 83328
rect 628741 83267 628850 83272
rect 628790 83028 628850 83267
rect 579061 82242 579127 82245
rect 650361 82242 650427 82245
rect 575798 82240 579127 82242
rect 575798 82184 579066 82240
rect 579122 82184 579127 82240
rect 648140 82240 650427 82242
rect 575798 82182 579127 82184
rect 575798 81668 575858 82182
rect 579061 82179 579127 82182
rect 628790 81698 628850 82212
rect 648140 82184 650366 82240
rect 650422 82184 650427 82240
rect 648140 82182 650427 82184
rect 650361 82179 650427 82182
rect 629201 81698 629267 81701
rect 628790 81696 629267 81698
rect 628790 81640 629206 81696
rect 629262 81640 629267 81696
rect 628790 81638 629267 81640
rect 629201 81635 629267 81638
rect 578877 80066 578943 80069
rect 575798 80064 578943 80066
rect 575798 80008 578882 80064
rect 578938 80008 578943 80064
rect 575798 80006 578943 80008
rect 575798 79492 575858 80006
rect 578877 80003 578943 80006
rect 633893 78572 633959 78573
rect 633893 78570 633940 78572
rect 633848 78568 633940 78570
rect 633848 78512 633898 78568
rect 633848 78510 633940 78512
rect 633893 78508 633940 78510
rect 634004 78508 634010 78572
rect 633893 78507 633959 78508
rect 637062 78162 637068 78164
rect 625110 78102 637068 78162
rect 579521 77890 579587 77893
rect 575798 77888 579587 77890
rect 575798 77832 579526 77888
rect 579582 77832 579587 77888
rect 575798 77830 579587 77832
rect 575798 77316 575858 77830
rect 579521 77827 579587 77830
rect 581637 77890 581703 77893
rect 625110 77890 625170 78102
rect 637062 78100 637068 78102
rect 637132 78162 637138 78164
rect 639597 78162 639663 78165
rect 637132 78160 639663 78162
rect 637132 78104 639602 78160
rect 639658 78104 639663 78160
rect 637132 78102 639663 78104
rect 637132 78100 637138 78102
rect 639597 78099 639663 78102
rect 581637 77888 625170 77890
rect 581637 77832 581642 77888
rect 581698 77832 625170 77888
rect 581637 77830 625170 77832
rect 581637 77827 581703 77830
rect 624417 77346 624483 77349
rect 633893 77346 633959 77349
rect 624417 77344 633959 77346
rect 624417 77288 624422 77344
rect 624478 77288 633898 77344
rect 633954 77288 633959 77344
rect 624417 77286 633959 77288
rect 624417 77283 624483 77286
rect 633893 77283 633959 77286
rect 578233 75578 578299 75581
rect 575798 75576 578299 75578
rect 575798 75520 578238 75576
rect 578294 75520 578299 75576
rect 575798 75518 578299 75520
rect 575798 75140 575858 75518
rect 578233 75515 578299 75518
rect 646129 74218 646195 74221
rect 646086 74216 646195 74218
rect 646086 74160 646134 74216
rect 646190 74160 646195 74216
rect 646086 74155 646195 74160
rect 646086 73848 646146 74155
rect 579061 73130 579127 73133
rect 575798 73128 579127 73130
rect 575798 73072 579066 73128
rect 579122 73072 579127 73128
rect 575798 73070 579127 73072
rect 575798 72964 575858 73070
rect 579061 73067 579127 73070
rect 646313 71770 646379 71773
rect 646270 71768 646379 71770
rect 646270 71712 646318 71768
rect 646374 71712 646379 71768
rect 646270 71707 646379 71712
rect 646270 71400 646330 71707
rect 579061 71226 579127 71229
rect 575798 71224 579127 71226
rect 575798 71168 579066 71224
rect 579122 71168 579127 71224
rect 575798 71166 579127 71168
rect 575798 70788 575858 71166
rect 579061 71163 579127 71166
rect 646638 68914 646698 68952
rect 647233 68914 647299 68917
rect 646638 68912 647299 68914
rect 646638 68856 647238 68912
rect 647294 68856 647299 68912
rect 646638 68854 647299 68856
rect 647233 68851 647299 68854
rect 646497 67146 646563 67149
rect 646454 67144 646563 67146
rect 646454 67088 646502 67144
rect 646558 67088 646563 67144
rect 646454 67083 646563 67088
rect 646454 66504 646514 67083
rect 646129 64426 646195 64429
rect 646086 64424 646195 64426
rect 646086 64368 646134 64424
rect 646190 64368 646195 64424
rect 646086 64363 646195 64368
rect 646086 64056 646146 64363
rect 648613 62114 648679 62117
rect 646638 62112 648679 62114
rect 646638 62056 648618 62112
rect 648674 62056 648679 62112
rect 646638 62054 648679 62056
rect 646638 61608 646698 62054
rect 648613 62051 648679 62054
rect 647233 59258 647299 59261
rect 646638 59256 647299 59258
rect 646638 59200 647238 59256
rect 647294 59200 647299 59256
rect 646638 59198 647299 59200
rect 646638 59160 646698 59198
rect 647233 59195 647299 59198
rect 648797 57354 648863 57357
rect 646638 57352 648863 57354
rect 646638 57296 648802 57352
rect 648858 57296 648863 57352
rect 646638 57294 648863 57296
rect 646638 56712 646698 57294
rect 648797 57291 648863 57294
rect 460790 54980 460796 55044
rect 460860 55042 460866 55044
rect 576117 55042 576183 55045
rect 460860 55040 576183 55042
rect 460860 54984 576122 55040
rect 576178 54984 576183 55040
rect 460860 54982 576183 54984
rect 460860 54980 460866 54982
rect 576117 54979 576183 54982
rect 462630 54708 462636 54772
rect 462700 54770 462706 54772
rect 580257 54770 580323 54773
rect 462700 54768 580323 54770
rect 462700 54712 580262 54768
rect 580318 54712 580323 54768
rect 462700 54710 580323 54712
rect 462700 54708 462706 54710
rect 580257 54707 580323 54710
rect 578877 54498 578943 54501
rect 466410 54496 578943 54498
rect 466410 54440 578882 54496
rect 578938 54440 578943 54496
rect 466410 54438 578943 54440
rect 466410 54226 466470 54438
rect 578877 54435 578943 54438
rect 577497 54226 577563 54229
rect 459878 54166 466470 54226
rect 476070 54224 577563 54226
rect 476070 54168 577502 54224
rect 577558 54168 577563 54224
rect 476070 54166 577563 54168
rect 459878 53685 459938 54166
rect 460790 53892 460796 53956
rect 460860 53892 460866 53956
rect 476070 53954 476130 54166
rect 577497 54163 577563 54166
rect 461718 53894 476130 53954
rect 460798 53685 460858 53892
rect 461718 53685 461778 53894
rect 459829 53680 459938 53685
rect 459829 53624 459834 53680
rect 459890 53624 459938 53680
rect 459829 53622 459938 53624
rect 460749 53680 460858 53685
rect 460749 53624 460754 53680
rect 460810 53624 460858 53680
rect 460749 53622 460858 53624
rect 461669 53680 461778 53685
rect 462589 53684 462655 53685
rect 462589 53682 462636 53684
rect 461669 53624 461674 53680
rect 461730 53624 461778 53680
rect 461669 53622 461778 53624
rect 462544 53680 462636 53682
rect 462544 53624 462594 53680
rect 462544 53622 462636 53624
rect 459829 53619 459895 53622
rect 460749 53619 460815 53622
rect 461669 53619 461735 53622
rect 462589 53620 462636 53622
rect 462700 53620 462706 53684
rect 462589 53619 462655 53620
rect 460381 53410 460447 53413
rect 465441 53410 465507 53413
rect 460381 53408 465507 53410
rect 460381 53352 460386 53408
rect 460442 53352 465446 53408
rect 465502 53352 465507 53408
rect 460381 53350 465507 53352
rect 460381 53347 460447 53350
rect 465441 53347 465507 53350
rect 518750 48860 518756 48924
rect 518820 48922 518826 48924
rect 549989 48922 550055 48925
rect 518820 48920 550055 48922
rect 518820 48864 549994 48920
rect 550050 48864 550055 48920
rect 518820 48862 550055 48864
rect 518820 48860 518826 48862
rect 549989 48859 550055 48862
rect 661585 48512 661651 48515
rect 661480 48510 661651 48512
rect 661480 48454 661590 48510
rect 661646 48454 661651 48510
rect 661480 48452 661651 48454
rect 661585 48449 661651 48452
rect 529606 48044 529612 48108
rect 529676 48106 529682 48108
rect 553669 48106 553735 48109
rect 529676 48104 553735 48106
rect 529676 48048 553674 48104
rect 553730 48048 553735 48104
rect 529676 48046 553735 48048
rect 529676 48044 529682 48046
rect 553669 48043 553735 48046
rect 515438 47772 515444 47836
rect 515508 47834 515514 47836
rect 522941 47834 523007 47837
rect 515508 47832 523007 47834
rect 515508 47776 522946 47832
rect 523002 47776 523007 47832
rect 515508 47774 523007 47776
rect 515508 47772 515514 47774
rect 522941 47771 523007 47774
rect 526478 47772 526484 47836
rect 526548 47834 526554 47836
rect 552013 47834 552079 47837
rect 526548 47832 552079 47834
rect 526548 47776 552018 47832
rect 552074 47776 552079 47832
rect 526548 47774 552079 47776
rect 526548 47772 526554 47774
rect 552013 47771 552079 47774
rect 520958 47500 520964 47564
rect 521028 47562 521034 47564
rect 547873 47562 547939 47565
rect 521028 47560 547939 47562
rect 521028 47504 547878 47560
rect 547934 47504 547939 47560
rect 521028 47502 547939 47504
rect 521028 47500 521034 47502
rect 547873 47499 547939 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 522062 47228 522068 47292
rect 522132 47290 522138 47292
rect 545665 47290 545731 47293
rect 522132 47288 545731 47290
rect 522132 47232 545670 47288
rect 545726 47232 545731 47288
rect 522132 47230 545731 47232
rect 522132 47228 522138 47230
rect 545665 47227 545731 47230
rect 458173 47018 458239 47021
rect 465073 47018 465139 47021
rect 458173 47016 465139 47018
rect 458173 46960 458178 47016
rect 458234 46960 465078 47016
rect 465134 46960 465139 47016
rect 458173 46958 465139 46960
rect 458173 46955 458239 46958
rect 465073 46955 465139 46958
rect 458357 46746 458423 46749
rect 465257 46746 465323 46749
rect 458357 46744 465323 46746
rect 458357 46688 458362 46744
rect 458418 46688 465262 46744
rect 465318 46688 465323 46744
rect 458357 46686 465323 46688
rect 458357 46683 458423 46686
rect 465257 46683 465323 46686
rect 130377 44298 130443 44301
rect 132769 44298 132835 44301
rect 142613 44298 142679 44301
rect 130377 44296 132835 44298
rect 130377 44240 130382 44296
rect 130438 44240 132774 44296
rect 132830 44240 132835 44296
rect 130377 44238 132835 44240
rect 130377 44235 130443 44238
rect 132769 44235 132835 44238
rect 142110 44296 142679 44298
rect 142110 44240 142618 44296
rect 142674 44240 142679 44296
rect 142110 44238 142679 44240
rect 141734 43964 141740 44028
rect 141804 44026 141810 44028
rect 142110 44026 142170 44238
rect 142613 44235 142679 44238
rect 461342 44236 461348 44300
rect 461412 44298 461418 44300
rect 461945 44298 462011 44301
rect 461412 44296 462011 44298
rect 461412 44240 461950 44296
rect 462006 44240 462011 44296
rect 461412 44238 462011 44240
rect 461412 44236 461418 44238
rect 461945 44235 462011 44238
rect 463693 44300 463759 44301
rect 463693 44296 463740 44300
rect 463804 44298 463810 44300
rect 463693 44240 463698 44296
rect 463693 44236 463740 44240
rect 463804 44238 463850 44298
rect 463804 44236 463810 44238
rect 464102 44236 464108 44300
rect 464172 44298 464178 44300
rect 464705 44298 464771 44301
rect 464172 44296 464771 44298
rect 464172 44240 464710 44296
rect 464766 44240 464771 44296
rect 464172 44238 464771 44240
rect 464172 44236 464178 44238
rect 463693 44235 463759 44236
rect 464705 44235 464771 44238
rect 255865 44162 255931 44165
rect 460105 44162 460171 44165
rect 255865 44160 460171 44162
rect 255865 44104 255870 44160
rect 255926 44104 460110 44160
rect 460166 44104 460171 44160
rect 255865 44102 460171 44104
rect 255865 44099 255931 44102
rect 460105 44099 460171 44102
rect 462865 44026 462931 44029
rect 141804 43966 142170 44026
rect 460890 44024 462931 44026
rect 460890 43968 462870 44024
rect 462926 43968 462931 44024
rect 460890 43966 462931 43968
rect 141804 43964 141810 43966
rect 419717 43890 419783 43893
rect 440233 43890 440299 43893
rect 419717 43888 440299 43890
rect 419717 43832 419722 43888
rect 419778 43832 440238 43888
rect 440294 43832 440299 43888
rect 419717 43830 440299 43832
rect 419717 43827 419783 43830
rect 440233 43827 440299 43830
rect 441061 43890 441127 43893
rect 460890 43890 460950 43966
rect 462865 43963 462931 43966
rect 441061 43888 460950 43890
rect 441061 43832 441066 43888
rect 441122 43832 460950 43888
rect 441061 43830 460950 43832
rect 441061 43827 441127 43830
rect 460749 43482 460815 43485
rect 471053 43482 471119 43485
rect 460749 43480 471119 43482
rect 460749 43424 460754 43480
rect 460810 43424 471058 43480
rect 471114 43424 471119 43480
rect 460749 43422 471119 43424
rect 460749 43419 460815 43422
rect 471053 43419 471119 43422
rect 462681 43210 462747 43213
rect 465809 43210 465875 43213
rect 462681 43208 465875 43210
rect 462681 43152 462686 43208
rect 462742 43152 465814 43208
rect 465870 43152 465875 43208
rect 462681 43150 465875 43152
rect 462681 43147 462747 43150
rect 465809 43147 465875 43150
rect 461761 42938 461827 42941
rect 463969 42938 464035 42941
rect 461761 42936 464035 42938
rect 461761 42880 461766 42936
rect 461822 42880 463974 42936
rect 464030 42880 464035 42936
rect 461761 42878 464035 42880
rect 461761 42875 461827 42878
rect 463969 42875 464035 42878
rect 518801 42804 518867 42805
rect 518750 42802 518756 42804
rect 518710 42742 518756 42802
rect 518820 42800 518867 42804
rect 518862 42744 518867 42800
rect 518750 42740 518756 42742
rect 518820 42740 518867 42744
rect 518801 42739 518867 42740
rect 460933 42394 460999 42397
rect 447090 42392 460999 42394
rect 447090 42336 460938 42392
rect 460994 42336 460999 42392
rect 447090 42334 460999 42336
rect 416681 42258 416747 42261
rect 446213 42258 446279 42261
rect 447090 42258 447150 42334
rect 460933 42331 460999 42334
rect 416681 42256 427830 42258
rect 416681 42200 416686 42256
rect 416742 42200 427830 42256
rect 416681 42198 427830 42200
rect 416681 42195 416747 42198
rect 415577 42124 415643 42125
rect 415526 42122 415532 42124
rect 415486 42062 415532 42122
rect 415596 42120 415643 42124
rect 415638 42064 415643 42120
rect 415526 42060 415532 42062
rect 415596 42060 415643 42064
rect 415577 42059 415643 42060
rect 361941 41852 362007 41853
rect 361941 41848 361988 41852
rect 362052 41850 362058 41852
rect 365161 41850 365227 41853
rect 365662 41850 365668 41852
rect 361941 41792 361946 41848
rect 361941 41788 361988 41792
rect 362052 41790 362098 41850
rect 365161 41848 365668 41850
rect 365161 41792 365166 41848
rect 365222 41792 365668 41848
rect 365161 41790 365668 41792
rect 362052 41788 362058 41790
rect 361941 41787 362007 41788
rect 365161 41787 365227 41790
rect 365662 41788 365668 41790
rect 365732 41788 365738 41852
rect 403014 41788 403020 41852
rect 403084 41850 403090 41852
rect 421966 41850 421972 41852
rect 403084 41790 421972 41850
rect 403084 41788 403090 41790
rect 421966 41788 421972 41790
rect 422036 41788 422042 41852
rect 427770 41578 427830 42198
rect 446213 42256 447150 42258
rect 446213 42200 446218 42256
rect 446274 42200 447150 42256
rect 446213 42198 447150 42200
rect 446213 42195 446279 42198
rect 515397 42124 515463 42125
rect 520917 42124 520983 42125
rect 522021 42124 522087 42125
rect 526437 42124 526503 42125
rect 529565 42124 529631 42125
rect 515397 42122 515444 42124
rect 515352 42120 515444 42122
rect 515352 42064 515402 42120
rect 515352 42062 515444 42064
rect 515397 42060 515444 42062
rect 515508 42060 515514 42124
rect 520917 42122 520964 42124
rect 520872 42120 520964 42122
rect 520872 42064 520922 42120
rect 520872 42062 520964 42064
rect 520917 42060 520964 42062
rect 521028 42060 521034 42124
rect 522021 42122 522068 42124
rect 521976 42120 522068 42122
rect 521976 42064 522026 42120
rect 521976 42062 522068 42064
rect 522021 42060 522068 42062
rect 522132 42060 522138 42124
rect 526437 42122 526484 42124
rect 526392 42120 526484 42122
rect 526392 42064 526442 42120
rect 526392 42062 526484 42064
rect 526437 42060 526484 42062
rect 526548 42060 526554 42124
rect 529565 42122 529612 42124
rect 529520 42120 529612 42122
rect 529520 42064 529570 42120
rect 529520 42062 529612 42064
rect 529565 42060 529612 42062
rect 529676 42060 529682 42124
rect 515397 42059 515463 42060
rect 520917 42059 520983 42060
rect 522021 42059 522087 42060
rect 526437 42059 526503 42060
rect 529565 42059 529631 42060
rect 441838 41788 441844 41852
rect 441908 41850 441914 41852
rect 460790 41850 460796 41852
rect 441908 41790 460796 41850
rect 441908 41788 441914 41790
rect 460790 41788 460796 41790
rect 460860 41788 460866 41852
rect 460974 41788 460980 41852
rect 461044 41850 461050 41852
rect 464102 41850 464108 41852
rect 461044 41790 464108 41850
rect 461044 41788 461050 41790
rect 464102 41788 464108 41790
rect 464172 41788 464178 41852
rect 446213 41578 446279 41581
rect 427770 41576 446279 41578
rect 427770 41520 446218 41576
rect 446274 41520 446279 41576
rect 427770 41518 446279 41520
rect 446213 41515 446279 41518
rect 141693 40356 141759 40357
rect 141693 40352 141740 40356
rect 141804 40354 141810 40356
rect 141693 40296 141698 40352
rect 141693 40292 141740 40296
rect 141804 40294 141850 40354
rect 141804 40292 141810 40294
rect 141693 40291 141759 40292
<< via3 >>
rect 675892 892196 675956 892260
rect 675892 887708 675956 887772
rect 675708 885804 675772 885868
rect 675524 880636 675588 880700
rect 676444 880364 676508 880428
rect 675340 878460 675404 878524
rect 675340 874108 675404 874172
rect 676444 872748 676508 872812
rect 676260 869756 676324 869820
rect 675708 865676 675772 865740
rect 676076 865404 676140 865468
rect 675892 864860 675956 864924
rect 41828 813180 41892 813244
rect 42012 811956 42076 812020
rect 40540 805564 40604 805628
rect 40908 805216 40972 805220
rect 40908 805160 40958 805216
rect 40958 805160 40972 805216
rect 40908 805156 40972 805160
rect 40724 804884 40788 804948
rect 41644 804672 41708 804676
rect 41644 804616 41658 804672
rect 41658 804616 41708 804672
rect 41644 804612 41708 804616
rect 41092 800532 41156 800596
rect 41092 794412 41156 794476
rect 40908 793460 40972 793524
rect 40724 791964 40788 792028
rect 40540 789516 40604 789580
rect 41644 789244 41708 789308
rect 41460 788836 41524 788900
rect 41828 788624 41892 788628
rect 41828 788568 41878 788624
rect 41878 788568 41892 788624
rect 41828 788564 41892 788568
rect 676076 788020 676140 788084
rect 674420 786660 674484 786724
rect 675340 786720 675404 786724
rect 675340 786664 675390 786720
rect 675390 786664 675404 786720
rect 675340 786660 675404 786664
rect 41644 769796 41708 769860
rect 41460 767348 41524 767412
rect 40724 766532 40788 766596
rect 40540 765308 40604 765372
rect 40908 764900 40972 764964
rect 41828 757692 41892 757756
rect 40356 757284 40420 757348
rect 40908 755788 40972 755852
rect 40356 754972 40420 755036
rect 40540 749396 40604 749460
rect 40724 746812 40788 746876
rect 41828 745316 41892 745380
rect 41460 745044 41524 745108
rect 41644 744772 41708 744836
rect 674236 743276 674300 743340
rect 674604 738108 674668 738172
rect 675340 730824 675404 730828
rect 675340 730768 675354 730824
rect 675354 730768 675404 730824
rect 675340 730764 675404 730768
rect 676812 729812 676876 729876
rect 676076 726548 676140 726612
rect 674420 726276 674484 726340
rect 41828 725792 41892 725796
rect 41828 725736 41842 725792
rect 41842 725736 41892 725792
rect 41828 725732 41892 725736
rect 41828 723072 41892 723076
rect 41828 723016 41842 723072
rect 41842 723016 41892 723072
rect 41828 723012 41892 723016
rect 674052 721712 674116 721716
rect 674052 721656 674066 721712
rect 674066 721656 674116 721712
rect 674052 721652 674116 721656
rect 675340 721516 675404 721580
rect 674052 719808 674116 719812
rect 674052 719752 674066 719808
rect 674066 719752 674116 719808
rect 674052 719748 674116 719752
rect 40540 718524 40604 718588
rect 40724 718252 40788 718316
rect 41828 716892 41892 716956
rect 42748 714580 42812 714644
rect 42380 714444 42444 714508
rect 42196 713900 42260 713964
rect 42196 710424 42260 710428
rect 42196 710368 42246 710424
rect 42246 710368 42260 710424
rect 42196 710364 42260 710368
rect 42748 710016 42812 710020
rect 42748 709960 42762 710016
rect 42762 709960 42812 710016
rect 42748 709956 42812 709960
rect 40724 709412 40788 709476
rect 40540 707916 40604 707980
rect 42196 707916 42260 707980
rect 42380 706208 42444 706212
rect 42380 706152 42430 706208
rect 42430 706152 42444 706208
rect 42380 706148 42444 706152
rect 42196 704244 42260 704308
rect 41828 701796 41892 701860
rect 41644 701524 41708 701588
rect 41460 700436 41524 700500
rect 675524 696824 675588 696828
rect 675524 696768 675538 696824
rect 675538 696768 675588 696824
rect 675524 696764 675588 696768
rect 674420 694588 674484 694652
rect 675340 686216 675404 686220
rect 675340 686160 675354 686216
rect 675354 686160 675404 686216
rect 675340 686156 675404 686160
rect 675524 685884 675588 685948
rect 41092 683402 41156 683466
rect 674236 682620 674300 682684
rect 40540 678928 40604 678992
rect 41828 678872 41892 678876
rect 41828 678816 41842 678872
rect 41842 678816 41892 678872
rect 41828 678812 41892 678816
rect 40724 677750 40788 677754
rect 40724 677694 40774 677750
rect 40774 677694 40788 677750
rect 40724 677690 40788 677694
rect 676076 676364 676140 676428
rect 41828 672692 41892 672756
rect 42196 671468 42260 671532
rect 40908 670924 40972 670988
rect 40908 667388 40972 667452
rect 42196 666632 42260 666636
rect 42196 666576 42210 666632
rect 42210 666576 42260 666632
rect 42196 666572 42260 666576
rect 676812 665756 676876 665820
rect 40540 665348 40604 665412
rect 40724 665076 40788 665140
rect 674604 662356 674668 662420
rect 41644 658548 41708 658612
rect 41828 658336 41892 658340
rect 41828 658280 41842 658336
rect 41842 658280 41892 658336
rect 41828 658276 41892 658280
rect 41460 657188 41524 657252
rect 674236 652836 674300 652900
rect 674788 646036 674852 646100
rect 41460 640596 41524 640660
rect 674788 640248 674852 640252
rect 674788 640192 674838 640248
rect 674838 640192 674852 640248
rect 674788 640188 674852 640192
rect 676076 637468 676140 637532
rect 40540 635292 40604 635356
rect 40724 634884 40788 634948
rect 675156 631348 675220 631412
rect 676076 631348 676140 631412
rect 41644 629852 41708 629916
rect 41828 629172 41892 629236
rect 40724 621964 40788 622028
rect 40540 620740 40604 620804
rect 674420 618972 674484 619036
rect 676812 617068 676876 617132
rect 673868 616116 673932 616180
rect 41460 615980 41524 616044
rect 41828 615436 41892 615500
rect 41828 613456 41892 613460
rect 41828 613400 41878 613456
rect 41878 613400 41892 613456
rect 41828 613396 41892 613400
rect 40540 612308 40604 612372
rect 674420 602924 674484 602988
rect 40540 601972 40604 602036
rect 42748 598436 42812 598500
rect 42012 597212 42076 597276
rect 42748 597000 42812 597004
rect 42748 596944 42798 597000
rect 42798 596944 42812 597000
rect 42748 596940 42812 596944
rect 675340 595368 675404 595372
rect 675340 595312 675390 595368
rect 675390 595312 675404 595368
rect 675340 595308 675404 595312
rect 41828 593948 41892 594012
rect 675156 593132 675220 593196
rect 40724 592486 40788 592550
rect 41828 592316 41892 592380
rect 42196 592044 42260 592108
rect 675340 591500 675404 591564
rect 676076 591364 676140 591428
rect 674236 591092 674300 591156
rect 676076 586196 676140 586260
rect 41828 585108 41892 585172
rect 41092 584836 41156 584900
rect 40356 584564 40420 584628
rect 40356 580212 40420 580276
rect 41092 579940 41156 580004
rect 42196 579396 42260 579460
rect 673684 578580 673748 578644
rect 42012 578308 42076 578372
rect 673500 577900 673564 577964
rect 40908 577764 40972 577828
rect 676812 576812 676876 576876
rect 40724 574636 40788 574700
rect 41460 573956 41524 574020
rect 40540 573412 40604 573476
rect 42196 573472 42260 573476
rect 42196 573416 42210 573472
rect 42210 573416 42260 573472
rect 42196 573412 42260 573416
rect 42012 572656 42076 572660
rect 42012 572600 42062 572656
rect 42062 572600 42076 572656
rect 42012 572596 42076 572600
rect 41644 571508 41708 571572
rect 41828 570208 41892 570212
rect 41828 570152 41842 570208
rect 41842 570152 41892 570208
rect 41828 570148 41892 570152
rect 675340 561912 675404 561916
rect 675340 561856 675390 561912
rect 675390 561856 675404 561912
rect 675340 561852 675404 561856
rect 41092 558724 41156 558788
rect 41092 557488 41156 557552
rect 676260 554644 676324 554708
rect 674052 554160 674116 554164
rect 674052 554104 674102 554160
rect 674102 554104 674116 554160
rect 674052 554100 674116 554104
rect 41828 553964 41892 554028
rect 676812 553828 676876 553892
rect 674052 552876 674116 552940
rect 41828 552740 41892 552804
rect 674052 550428 674116 550492
rect 42196 549476 42260 549540
rect 675340 548388 675404 548452
rect 676996 548252 677060 548316
rect 674052 547844 674116 547908
rect 676260 547572 676324 547636
rect 676076 546756 676140 546820
rect 40724 545592 40788 545596
rect 40724 545536 40774 545592
rect 40774 545536 40788 545592
rect 40724 545532 40788 545536
rect 40540 545260 40604 545324
rect 42196 545260 42260 545324
rect 41828 542268 41892 542332
rect 40724 535196 40788 535260
rect 40540 533292 40604 533356
rect 41644 531660 41708 531724
rect 41460 530708 41524 530772
rect 41828 528940 41892 529004
rect 674420 527036 674484 527100
rect 676996 503644 677060 503708
rect 676812 500924 676876 500988
rect 676030 488820 676094 488884
rect 675892 487868 675956 487932
rect 673868 455228 673932 455292
rect 41828 423600 41892 423604
rect 41828 423544 41842 423600
rect 41842 423544 41892 423600
rect 41828 423540 41892 423544
rect 40908 422248 40972 422312
rect 40724 418644 40788 418708
rect 40540 418372 40604 418436
rect 42012 415244 42076 415308
rect 41828 414564 41892 414628
rect 40908 406948 40972 407012
rect 40540 406676 40604 406740
rect 40724 404500 40788 404564
rect 677180 401236 677244 401300
rect 676812 400420 676876 400484
rect 41460 400012 41524 400076
rect 41828 399392 41892 399396
rect 41828 399336 41842 399392
rect 41842 399336 41892 399392
rect 41828 399332 41892 399336
rect 42012 398848 42076 398852
rect 42012 398792 42026 398848
rect 42026 398792 42076 398848
rect 42012 398788 42076 398792
rect 676076 398788 676140 398852
rect 676260 396748 676324 396812
rect 676444 396340 676508 396404
rect 676628 395116 676692 395180
rect 675340 392804 675404 392868
rect 675892 387636 675956 387700
rect 676260 384916 676324 384980
rect 676444 382196 676508 382260
rect 41460 381788 41524 381852
rect 41644 379340 41708 379404
rect 40724 378932 40788 378996
rect 40540 378524 40604 378588
rect 675892 378524 675956 378588
rect 40908 377708 40972 377772
rect 676628 377436 676692 377500
rect 41828 374580 41892 374644
rect 676076 373628 676140 373692
rect 675340 372812 675404 372876
rect 40908 364788 40972 364852
rect 40724 364108 40788 364172
rect 40540 360028 40604 360092
rect 41828 358728 41892 358732
rect 41828 358672 41878 358728
rect 41878 358672 41892 358728
rect 41828 358668 41892 358672
rect 41460 356900 41524 356964
rect 41828 355736 41892 355740
rect 41828 355680 41878 355736
rect 41878 355680 41892 355736
rect 41828 355676 41892 355680
rect 43300 354452 43364 354516
rect 675524 354180 675588 354244
rect 675892 353772 675956 353836
rect 675708 352956 675772 353020
rect 675892 351732 675956 351796
rect 675340 347652 675404 347716
rect 676444 346564 676508 346628
rect 42196 344252 42260 344316
rect 44220 342892 44284 342956
rect 44588 342348 44652 342412
rect 42196 342076 42260 342140
rect 42748 340172 42812 340236
rect 676260 340172 676324 340236
rect 44404 339764 44468 339828
rect 675524 339416 675588 339420
rect 675524 339360 675538 339416
rect 675538 339360 675588 339416
rect 675524 339356 675588 339360
rect 676076 337860 676140 337924
rect 42932 337588 42996 337652
rect 40540 336908 40604 336972
rect 41828 336500 41892 336564
rect 676444 336500 676508 336564
rect 40908 335684 40972 335748
rect 40724 335276 40788 335340
rect 43300 334596 43364 334660
rect 41460 332828 41524 332892
rect 41644 331740 41708 331804
rect 675340 327992 675404 327996
rect 675340 327936 675390 327992
rect 675390 327936 675404 327992
rect 675340 327932 675404 327936
rect 676628 325620 676692 325684
rect 41828 324864 41892 324868
rect 41828 324808 41842 324864
rect 41842 324808 41892 324864
rect 41828 324804 41892 324808
rect 40908 321132 40972 321196
rect 40724 317324 40788 317388
rect 40540 315964 40604 316028
rect 41828 315616 41892 315620
rect 41828 315560 41842 315616
rect 41842 315560 41892 315616
rect 41828 315556 41892 315560
rect 41460 313652 41524 313716
rect 42932 312700 42996 312764
rect 675892 308756 675956 308820
rect 676076 306580 676140 306644
rect 676260 304914 676324 304978
rect 675892 302636 675956 302700
rect 676444 301548 676508 301612
rect 44220 300052 44284 300116
rect 44588 299236 44652 299300
rect 44404 298420 44468 298484
rect 42748 297604 42812 297668
rect 675708 297332 675772 297396
rect 42196 296788 42260 296852
rect 675156 296652 675220 296716
rect 675156 294476 675220 294540
rect 676628 294476 676692 294540
rect 40540 292528 40604 292592
rect 42012 292164 42076 292228
rect 41828 291892 41892 291956
rect 676444 291484 676508 291548
rect 676260 290940 676324 291004
rect 41828 289988 41892 290052
rect 42196 289988 42260 290052
rect 40908 289172 40972 289236
rect 42196 284820 42260 284884
rect 41828 284276 41892 284340
rect 676076 283596 676140 283660
rect 40908 282236 40972 282300
rect 675892 282644 675956 282708
rect 42196 281752 42260 281756
rect 42196 281696 42210 281752
rect 42210 281696 42260 281752
rect 42196 281692 42260 281696
rect 675708 281616 675772 281620
rect 675708 281560 675722 281616
rect 675722 281560 675772 281616
rect 675708 281556 675772 281560
rect 42196 280256 42260 280260
rect 42196 280200 42210 280256
rect 42210 280200 42260 280256
rect 42196 280196 42260 280200
rect 42196 278700 42260 278764
rect 40724 277068 40788 277132
rect 40540 274212 40604 274276
rect 675340 273804 675404 273868
rect 41460 270404 41524 270468
rect 41828 269784 41892 269788
rect 41828 269728 41842 269784
rect 41842 269728 41892 269784
rect 41828 269724 41892 269728
rect 42012 269104 42076 269108
rect 42012 269048 42026 269104
rect 42026 269048 42076 269104
rect 42012 269044 42076 269048
rect 676996 261564 677060 261628
rect 676812 261156 676876 261220
rect 675524 258088 675588 258092
rect 675524 258032 675538 258088
rect 675538 258032 675588 258088
rect 675524 258028 675588 258032
rect 676996 250276 677060 250340
rect 675524 250004 675588 250068
rect 40540 249732 40604 249796
rect 675340 249732 675404 249796
rect 40724 249324 40788 249388
rect 676812 246604 676876 246668
rect 673316 246196 673380 246260
rect 675524 246196 675588 246260
rect 667796 245652 667860 245716
rect 676812 241708 676876 241772
rect 42012 238036 42076 238100
rect 40540 236540 40604 236604
rect 675524 235512 675588 235516
rect 675524 235456 675538 235512
rect 675538 235456 675588 235512
rect 675524 235452 675588 235456
rect 40724 234636 40788 234700
rect 670740 231916 670804 231980
rect 42012 228984 42076 228988
rect 42012 228928 42026 228984
rect 42026 228928 42076 228984
rect 42012 228924 42076 228928
rect 674236 228516 674300 228580
rect 675524 228576 675588 228580
rect 675524 228520 675538 228576
rect 675538 228520 675588 228576
rect 675524 228516 675588 228520
rect 672580 227080 672644 227084
rect 672580 227024 672630 227080
rect 672630 227024 672644 227080
rect 672580 227020 672644 227024
rect 683804 227020 683868 227084
rect 674052 226476 674116 226540
rect 670004 224572 670068 224636
rect 671476 224360 671540 224364
rect 671476 224304 671526 224360
rect 671526 224304 671540 224360
rect 671476 224300 671540 224304
rect 670556 223952 670620 223956
rect 670556 223896 670570 223952
rect 670570 223896 670620 223952
rect 670556 223892 670620 223896
rect 683804 223756 683868 223820
rect 670372 223680 670436 223684
rect 670372 223624 670422 223680
rect 670422 223624 670436 223680
rect 670372 223620 670436 223624
rect 671476 223680 671540 223684
rect 671476 223624 671526 223680
rect 671526 223624 671540 223680
rect 671476 223620 671540 223624
rect 591988 223348 592052 223412
rect 649580 222396 649644 222460
rect 651972 222396 652036 222460
rect 670004 220824 670068 220828
rect 670004 220768 670054 220824
rect 670054 220768 670068 220824
rect 670004 220764 670068 220768
rect 670556 220356 670620 220420
rect 676030 219812 676094 219876
rect 675524 218588 675588 218652
rect 669636 218044 669700 218108
rect 511028 217560 511092 217564
rect 511028 217504 511042 217560
rect 511042 217504 511092 217560
rect 511028 217500 511092 217504
rect 520044 217560 520108 217564
rect 520044 217504 520058 217560
rect 520058 217504 520108 217560
rect 520044 217500 520108 217504
rect 532556 217560 532620 217564
rect 532556 217504 532570 217560
rect 532570 217504 532620 217560
rect 532556 217500 532620 217504
rect 669084 217228 669148 217292
rect 675708 217636 675772 217700
rect 670372 216472 670436 216476
rect 670372 216416 670386 216472
rect 670386 216416 670436 216472
rect 670372 216412 670436 216416
rect 520044 215868 520108 215932
rect 511028 215596 511092 215660
rect 669820 215868 669884 215932
rect 673868 215868 673932 215932
rect 532556 215324 532620 215388
rect 670556 215324 670620 215388
rect 675892 215188 675956 215252
rect 669820 214780 669884 214844
rect 675892 214508 675956 214572
rect 673868 213556 673932 213620
rect 675708 212468 675772 212532
rect 670372 211108 670436 211172
rect 41828 210020 41892 210084
rect 41644 208116 41708 208180
rect 40540 207300 40604 207364
rect 674236 206892 674300 206956
rect 40724 206484 40788 206548
rect 40908 206076 40972 206140
rect 669268 205668 669332 205732
rect 669636 205668 669700 205732
rect 669268 205396 669332 205460
rect 669636 205396 669700 205460
rect 676260 202676 676324 202740
rect 672580 200832 672644 200836
rect 672580 200776 672594 200832
rect 672594 200776 672644 200832
rect 672580 200772 672644 200776
rect 676444 199956 676508 200020
rect 42012 198732 42076 198796
rect 670740 198732 670804 198796
rect 676812 197780 676876 197844
rect 669268 196012 669332 196076
rect 669636 196012 669700 196076
rect 42012 195800 42076 195804
rect 42012 195744 42026 195800
rect 42026 195744 42076 195800
rect 42012 195740 42076 195744
rect 41828 195256 41892 195260
rect 41828 195200 41842 195256
rect 41842 195200 41892 195256
rect 41828 195196 41892 195200
rect 40908 194924 40972 194988
rect 676628 194516 676692 194580
rect 40724 193428 40788 193492
rect 676076 193156 676140 193220
rect 675892 192748 675956 192812
rect 669452 191660 669516 191724
rect 675340 189076 675404 189140
rect 40540 186356 40604 186420
rect 41460 185948 41524 186012
rect 673132 181596 673196 181660
rect 668164 179556 668228 179620
rect 673316 179420 673380 179484
rect 676812 176608 676876 176672
rect 675708 173572 675772 173636
rect 675524 172348 675588 172412
rect 675892 170716 675956 170780
rect 675892 169628 675956 169692
rect 675524 169492 675588 169556
rect 675340 167452 675404 167516
rect 676444 166424 676508 166428
rect 676444 166368 676458 166424
rect 676458 166368 676508 166424
rect 676444 166364 676508 166368
rect 673132 161060 673196 161124
rect 676444 155756 676508 155820
rect 676628 155484 676692 155548
rect 676260 151404 676324 151468
rect 676076 148412 676140 148476
rect 675340 147656 675404 147660
rect 675340 147600 675390 147656
rect 675390 147600 675404 147656
rect 675340 147596 675404 147600
rect 669268 140388 669332 140452
rect 667796 132908 667860 132972
rect 676444 127332 676508 127396
rect 676076 126924 676140 126988
rect 676260 124476 676324 124540
rect 675340 122300 675404 122364
rect 676812 119988 676876 120052
rect 675708 117268 675772 117332
rect 674052 114956 674116 115020
rect 676444 112372 676508 112436
rect 676812 111692 676876 111756
rect 675708 111344 675772 111348
rect 675708 111288 675758 111344
rect 675758 111288 675772 111344
rect 675708 111284 675772 111288
rect 676260 110332 676324 110396
rect 676076 108156 676140 108220
rect 675340 101960 675404 101964
rect 675340 101904 675390 101960
rect 675390 101904 675404 101960
rect 675340 101900 675404 101904
rect 637252 96868 637316 96932
rect 647188 96460 647252 96524
rect 633940 95372 634004 95436
rect 650316 93060 650380 93124
rect 633940 78568 634004 78572
rect 633940 78512 633954 78568
rect 633954 78512 634004 78568
rect 633940 78508 634004 78512
rect 637068 78100 637132 78164
rect 460796 54980 460860 55044
rect 462636 54708 462700 54772
rect 460796 53892 460860 53956
rect 462636 53680 462700 53684
rect 462636 53624 462650 53680
rect 462650 53624 462700 53680
rect 462636 53620 462700 53624
rect 518756 48860 518820 48924
rect 529612 48044 529676 48108
rect 515444 47772 515508 47836
rect 526484 47772 526548 47836
rect 520964 47500 521028 47564
rect 522068 47228 522132 47292
rect 141740 43964 141804 44028
rect 461348 44236 461412 44300
rect 463740 44296 463804 44300
rect 463740 44240 463754 44296
rect 463754 44240 463804 44296
rect 463740 44236 463804 44240
rect 464108 44236 464172 44300
rect 518756 42800 518820 42804
rect 518756 42744 518806 42800
rect 518806 42744 518820 42800
rect 518756 42740 518820 42744
rect 415532 42120 415596 42124
rect 415532 42064 415582 42120
rect 415582 42064 415596 42120
rect 415532 42060 415596 42064
rect 361988 41848 362052 41852
rect 361988 41792 362002 41848
rect 362002 41792 362052 41848
rect 361988 41788 362052 41792
rect 365668 41788 365732 41852
rect 403020 41788 403084 41852
rect 421972 41788 422036 41852
rect 515444 42120 515508 42124
rect 515444 42064 515458 42120
rect 515458 42064 515508 42120
rect 515444 42060 515508 42064
rect 520964 42120 521028 42124
rect 520964 42064 520978 42120
rect 520978 42064 521028 42120
rect 520964 42060 521028 42064
rect 522068 42120 522132 42124
rect 522068 42064 522082 42120
rect 522082 42064 522132 42120
rect 522068 42060 522132 42064
rect 526484 42120 526548 42124
rect 526484 42064 526498 42120
rect 526498 42064 526548 42120
rect 526484 42060 526548 42064
rect 529612 42120 529676 42124
rect 529612 42064 529626 42120
rect 529626 42064 529676 42120
rect 529612 42060 529676 42064
rect 441844 41788 441908 41852
rect 460796 41788 460860 41852
rect 460980 41788 461044 41852
rect 464108 41788 464172 41852
rect 141740 40352 141804 40356
rect 141740 40296 141754 40352
rect 141754 40296 141804 40352
rect 141740 40292 141804 40296
<< metal4 >>
rect 675891 892260 675957 892261
rect 675891 892196 675892 892260
rect 675956 892196 675957 892260
rect 675891 892195 675957 892196
rect 675894 891510 675954 892195
rect 675710 891450 675954 891510
rect 675710 887090 675770 891450
rect 675891 887772 675957 887773
rect 675891 887708 675892 887772
rect 675956 887770 675957 887772
rect 675956 887710 676322 887770
rect 675956 887708 675957 887710
rect 675891 887707 675957 887708
rect 675710 887030 675954 887090
rect 675707 885868 675773 885869
rect 675707 885804 675708 885868
rect 675772 885804 675773 885868
rect 675707 885803 675773 885804
rect 675523 880700 675589 880701
rect 675523 880636 675524 880700
rect 675588 880636 675589 880700
rect 675523 880635 675589 880636
rect 675339 878524 675405 878525
rect 675339 878460 675340 878524
rect 675404 878460 675405 878524
rect 675339 878459 675405 878460
rect 675342 874173 675402 878459
rect 675339 874172 675405 874173
rect 675339 874108 675340 874172
rect 675404 874108 675405 874172
rect 675339 874107 675405 874108
rect 675526 872190 675586 880635
rect 675710 876890 675770 885803
rect 675894 881850 675954 887030
rect 675894 881790 676138 881850
rect 675710 876830 675954 876890
rect 675526 872130 675770 872190
rect 675710 865741 675770 872130
rect 675707 865740 675773 865741
rect 675707 865676 675708 865740
rect 675772 865676 675773 865740
rect 675707 865675 675773 865676
rect 675894 864925 675954 876830
rect 676078 865469 676138 881790
rect 676262 869821 676322 887710
rect 676443 880428 676509 880429
rect 676443 880364 676444 880428
rect 676508 880364 676509 880428
rect 676443 880363 676509 880364
rect 676446 872813 676506 880363
rect 676443 872812 676509 872813
rect 676443 872748 676444 872812
rect 676508 872748 676509 872812
rect 676443 872747 676509 872748
rect 676259 869820 676325 869821
rect 676259 869756 676260 869820
rect 676324 869756 676325 869820
rect 676259 869755 676325 869756
rect 676075 865468 676141 865469
rect 676075 865404 676076 865468
rect 676140 865404 676141 865468
rect 676075 865403 676141 865404
rect 675891 864924 675957 864925
rect 675891 864860 675892 864924
rect 675956 864860 675957 864924
rect 675891 864859 675957 864860
rect 41827 813244 41893 813245
rect 41827 813180 41828 813244
rect 41892 813180 41893 813244
rect 41827 813179 41893 813180
rect 41830 812970 41890 813179
rect 41462 812910 41890 812970
rect 40539 805628 40605 805629
rect 40539 805564 40540 805628
rect 40604 805564 40605 805628
rect 40539 805563 40605 805564
rect 40542 789581 40602 805563
rect 40907 805220 40973 805221
rect 40907 805156 40908 805220
rect 40972 805156 40973 805220
rect 40907 805155 40973 805156
rect 40723 804948 40789 804949
rect 40723 804884 40724 804948
rect 40788 804884 40789 804948
rect 40723 804883 40789 804884
rect 40726 792029 40786 804883
rect 40910 793525 40970 805155
rect 41091 800596 41157 800597
rect 41091 800532 41092 800596
rect 41156 800532 41157 800596
rect 41091 800531 41157 800532
rect 41094 794477 41154 800531
rect 41091 794476 41157 794477
rect 41091 794412 41092 794476
rect 41156 794412 41157 794476
rect 41091 794411 41157 794412
rect 40907 793524 40973 793525
rect 40907 793460 40908 793524
rect 40972 793460 40973 793524
rect 40907 793459 40973 793460
rect 40723 792028 40789 792029
rect 40723 791964 40724 792028
rect 40788 791964 40789 792028
rect 40723 791963 40789 791964
rect 40539 789580 40605 789581
rect 40539 789516 40540 789580
rect 40604 789516 40605 789580
rect 40539 789515 40605 789516
rect 41462 788901 41522 812910
rect 42011 812020 42077 812021
rect 42011 811956 42012 812020
rect 42076 811956 42077 812020
rect 42011 811955 42077 811956
rect 41643 804676 41709 804677
rect 41643 804612 41644 804676
rect 41708 804612 41709 804676
rect 41643 804611 41709 804612
rect 41646 789309 41706 804611
rect 42014 794910 42074 811955
rect 41830 794850 42074 794910
rect 41643 789308 41709 789309
rect 41643 789244 41644 789308
rect 41708 789244 41709 789308
rect 41643 789243 41709 789244
rect 41459 788900 41525 788901
rect 41459 788836 41460 788900
rect 41524 788836 41525 788900
rect 41459 788835 41525 788836
rect 41830 788629 41890 794850
rect 41827 788628 41893 788629
rect 41827 788564 41828 788628
rect 41892 788564 41893 788628
rect 41827 788563 41893 788564
rect 676075 788084 676141 788085
rect 676075 788020 676076 788084
rect 676140 788020 676141 788084
rect 676075 788019 676141 788020
rect 674419 786724 674485 786725
rect 674419 786660 674420 786724
rect 674484 786660 674485 786724
rect 674419 786659 674485 786660
rect 675339 786724 675405 786725
rect 675339 786660 675340 786724
rect 675404 786660 675405 786724
rect 675339 786659 675405 786660
rect 41643 769860 41709 769861
rect 41643 769796 41644 769860
rect 41708 769796 41709 769860
rect 41643 769795 41709 769796
rect 41459 767412 41525 767413
rect 41459 767348 41460 767412
rect 41524 767348 41525 767412
rect 41459 767347 41525 767348
rect 40723 766596 40789 766597
rect 40723 766532 40724 766596
rect 40788 766532 40789 766596
rect 40723 766531 40789 766532
rect 40539 765372 40605 765373
rect 40539 765308 40540 765372
rect 40604 765308 40605 765372
rect 40539 765307 40605 765308
rect 40355 757348 40421 757349
rect 40355 757284 40356 757348
rect 40420 757284 40421 757348
rect 40355 757283 40421 757284
rect 40358 755037 40418 757283
rect 40355 755036 40421 755037
rect 40355 754972 40356 755036
rect 40420 754972 40421 755036
rect 40355 754971 40421 754972
rect 40542 749461 40602 765307
rect 40539 749460 40605 749461
rect 40539 749396 40540 749460
rect 40604 749396 40605 749460
rect 40539 749395 40605 749396
rect 40726 746877 40786 766531
rect 40907 764964 40973 764965
rect 40907 764900 40908 764964
rect 40972 764900 40973 764964
rect 40907 764899 40973 764900
rect 40910 755853 40970 764899
rect 40907 755852 40973 755853
rect 40907 755788 40908 755852
rect 40972 755788 40973 755852
rect 40907 755787 40973 755788
rect 40723 746876 40789 746877
rect 40723 746812 40724 746876
rect 40788 746812 40789 746876
rect 40723 746811 40789 746812
rect 41462 745109 41522 767347
rect 41459 745108 41525 745109
rect 41459 745044 41460 745108
rect 41524 745044 41525 745108
rect 41459 745043 41525 745044
rect 41646 744837 41706 769795
rect 41827 757756 41893 757757
rect 41827 757692 41828 757756
rect 41892 757692 41893 757756
rect 41827 757691 41893 757692
rect 41830 745381 41890 757691
rect 41827 745380 41893 745381
rect 41827 745316 41828 745380
rect 41892 745316 41893 745380
rect 41827 745315 41893 745316
rect 41643 744836 41709 744837
rect 41643 744772 41644 744836
rect 41708 744772 41709 744836
rect 41643 744771 41709 744772
rect 674235 743340 674301 743341
rect 674235 743276 674236 743340
rect 674300 743276 674301 743340
rect 674235 743275 674301 743276
rect 41827 725796 41893 725797
rect 41827 725732 41828 725796
rect 41892 725732 41893 725796
rect 41827 725731 41893 725732
rect 41830 725250 41890 725731
rect 41462 725190 41890 725250
rect 40539 718588 40605 718589
rect 40539 718524 40540 718588
rect 40604 718524 40605 718588
rect 40539 718523 40605 718524
rect 40542 707981 40602 718523
rect 40723 718316 40789 718317
rect 40723 718252 40724 718316
rect 40788 718252 40789 718316
rect 40723 718251 40789 718252
rect 40726 709477 40786 718251
rect 40723 709476 40789 709477
rect 40723 709412 40724 709476
rect 40788 709412 40789 709476
rect 40723 709411 40789 709412
rect 40539 707980 40605 707981
rect 40539 707916 40540 707980
rect 40604 707916 40605 707980
rect 40539 707915 40605 707916
rect 41462 700501 41522 725190
rect 41827 723076 41893 723077
rect 41827 723012 41828 723076
rect 41892 723012 41893 723076
rect 41827 723011 41893 723012
rect 41830 717630 41890 723011
rect 674051 721716 674117 721717
rect 674051 721652 674052 721716
rect 674116 721652 674117 721716
rect 674051 721651 674117 721652
rect 674054 719813 674114 721651
rect 674051 719812 674117 719813
rect 674051 719748 674052 719812
rect 674116 719748 674117 719812
rect 674051 719747 674117 719748
rect 41646 717570 41890 717630
rect 41646 701589 41706 717570
rect 41827 716956 41893 716957
rect 41827 716892 41828 716956
rect 41892 716892 41893 716956
rect 41827 716891 41893 716892
rect 41830 701861 41890 716891
rect 42747 714644 42813 714645
rect 42747 714580 42748 714644
rect 42812 714580 42813 714644
rect 42747 714579 42813 714580
rect 42379 714508 42445 714509
rect 42379 714444 42380 714508
rect 42444 714444 42445 714508
rect 42379 714443 42445 714444
rect 42195 713964 42261 713965
rect 42195 713900 42196 713964
rect 42260 713900 42261 713964
rect 42195 713899 42261 713900
rect 42198 710429 42258 713899
rect 42195 710428 42261 710429
rect 42195 710364 42196 710428
rect 42260 710364 42261 710428
rect 42195 710363 42261 710364
rect 42195 707980 42261 707981
rect 42195 707916 42196 707980
rect 42260 707916 42261 707980
rect 42195 707915 42261 707916
rect 42198 704309 42258 707915
rect 42382 706213 42442 714443
rect 42750 710021 42810 714579
rect 42747 710020 42813 710021
rect 42747 709956 42748 710020
rect 42812 709956 42813 710020
rect 42747 709955 42813 709956
rect 42379 706212 42445 706213
rect 42379 706148 42380 706212
rect 42444 706148 42445 706212
rect 42379 706147 42445 706148
rect 42195 704308 42261 704309
rect 42195 704244 42196 704308
rect 42260 704244 42261 704308
rect 42195 704243 42261 704244
rect 41827 701860 41893 701861
rect 41827 701796 41828 701860
rect 41892 701796 41893 701860
rect 41827 701795 41893 701796
rect 41643 701588 41709 701589
rect 41643 701524 41644 701588
rect 41708 701524 41709 701588
rect 41643 701523 41709 701524
rect 41459 700500 41525 700501
rect 41459 700436 41460 700500
rect 41524 700436 41525 700500
rect 41459 700435 41525 700436
rect 41091 683466 41157 683467
rect 41091 683402 41092 683466
rect 41156 683402 41157 683466
rect 41091 683401 41157 683402
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40542 665413 40602 678927
rect 40723 677754 40789 677755
rect 40723 677690 40724 677754
rect 40788 677690 40789 677754
rect 40723 677689 40789 677690
rect 40539 665412 40605 665413
rect 40539 665348 40540 665412
rect 40604 665348 40605 665412
rect 40539 665347 40605 665348
rect 40726 665141 40786 677689
rect 41094 676230 41154 683401
rect 674238 682685 674298 743275
rect 674422 726341 674482 786659
rect 674603 738172 674669 738173
rect 674603 738108 674604 738172
rect 674668 738108 674669 738172
rect 674603 738107 674669 738108
rect 674419 726340 674485 726341
rect 674419 726276 674420 726340
rect 674484 726276 674485 726340
rect 674419 726275 674485 726276
rect 674419 694652 674485 694653
rect 674419 694588 674420 694652
rect 674484 694588 674485 694652
rect 674419 694587 674485 694588
rect 674235 682684 674301 682685
rect 674235 682620 674236 682684
rect 674300 682620 674301 682684
rect 674235 682619 674301 682620
rect 41827 678876 41893 678877
rect 41827 678812 41828 678876
rect 41892 678812 41893 678876
rect 41827 678811 41893 678812
rect 41830 678330 41890 678811
rect 41646 678270 41890 678330
rect 41094 676170 41522 676230
rect 40907 670988 40973 670989
rect 40907 670924 40908 670988
rect 40972 670924 40973 670988
rect 40907 670923 40973 670924
rect 40910 667453 40970 670923
rect 40907 667452 40973 667453
rect 40907 667388 40908 667452
rect 40972 667388 40973 667452
rect 40907 667387 40973 667388
rect 40723 665140 40789 665141
rect 40723 665076 40724 665140
rect 40788 665076 40789 665140
rect 40723 665075 40789 665076
rect 41462 657253 41522 676170
rect 41646 658613 41706 678270
rect 41827 672756 41893 672757
rect 41827 672692 41828 672756
rect 41892 672692 41893 672756
rect 41827 672691 41893 672692
rect 41643 658612 41709 658613
rect 41643 658548 41644 658612
rect 41708 658548 41709 658612
rect 41643 658547 41709 658548
rect 41830 658341 41890 672691
rect 42195 671532 42261 671533
rect 42195 671468 42196 671532
rect 42260 671468 42261 671532
rect 42195 671467 42261 671468
rect 42198 666637 42258 671467
rect 42195 666636 42261 666637
rect 42195 666572 42196 666636
rect 42260 666572 42261 666636
rect 42195 666571 42261 666572
rect 41827 658340 41893 658341
rect 41827 658276 41828 658340
rect 41892 658276 41893 658340
rect 41827 658275 41893 658276
rect 41459 657252 41525 657253
rect 41459 657188 41460 657252
rect 41524 657188 41525 657252
rect 41459 657187 41525 657188
rect 674235 652900 674301 652901
rect 674235 652836 674236 652900
rect 674300 652836 674301 652900
rect 674235 652835 674301 652836
rect 41459 640660 41525 640661
rect 41459 640596 41460 640660
rect 41524 640596 41525 640660
rect 41459 640595 41525 640596
rect 40539 635356 40605 635357
rect 40539 635292 40540 635356
rect 40604 635292 40605 635356
rect 40539 635291 40605 635292
rect 40542 620805 40602 635291
rect 40723 634948 40789 634949
rect 40723 634884 40724 634948
rect 40788 634884 40789 634948
rect 40723 634883 40789 634884
rect 40726 622029 40786 634883
rect 40723 622028 40789 622029
rect 40723 621964 40724 622028
rect 40788 621964 40789 622028
rect 40723 621963 40789 621964
rect 40539 620804 40605 620805
rect 40539 620740 40540 620804
rect 40604 620740 40605 620804
rect 40539 620739 40605 620740
rect 41462 616045 41522 640595
rect 41643 629916 41709 629917
rect 41643 629852 41644 629916
rect 41708 629852 41709 629916
rect 41643 629851 41709 629852
rect 41459 616044 41525 616045
rect 41459 615980 41460 616044
rect 41524 615980 41525 616044
rect 41459 615979 41525 615980
rect 41646 615090 41706 629851
rect 41827 629236 41893 629237
rect 41827 629172 41828 629236
rect 41892 629172 41893 629236
rect 41827 629171 41893 629172
rect 41830 615501 41890 629171
rect 673867 616180 673933 616181
rect 673867 616116 673868 616180
rect 673932 616116 673933 616180
rect 673867 616115 673933 616116
rect 41827 615500 41893 615501
rect 41827 615436 41828 615500
rect 41892 615436 41893 615500
rect 41827 615435 41893 615436
rect 41646 615030 41890 615090
rect 41830 613461 41890 615030
rect 41827 613460 41893 613461
rect 41827 613396 41828 613460
rect 41892 613396 41893 613460
rect 41827 613395 41893 613396
rect 40539 612372 40605 612373
rect 40539 612308 40540 612372
rect 40604 612308 40605 612372
rect 40539 612307 40605 612308
rect 40542 602037 40602 612307
rect 40539 602036 40605 602037
rect 40539 601972 40540 602036
rect 40604 601972 40605 602036
rect 40539 601971 40605 601972
rect 42747 598500 42813 598501
rect 42747 598436 42748 598500
rect 42812 598436 42813 598500
rect 42747 598435 42813 598436
rect 42011 597276 42077 597277
rect 42011 597212 42012 597276
rect 42076 597212 42077 597276
rect 42011 597211 42077 597212
rect 41827 594012 41893 594013
rect 41827 594010 41828 594012
rect 40542 593950 41828 594010
rect 40355 584628 40421 584629
rect 40355 584564 40356 584628
rect 40420 584564 40421 584628
rect 40355 584563 40421 584564
rect 40358 580277 40418 584563
rect 40355 580276 40421 580277
rect 40355 580212 40356 580276
rect 40420 580212 40421 580276
rect 40355 580211 40421 580212
rect 40542 573477 40602 593950
rect 41827 593948 41828 593950
rect 41892 593948 41893 594012
rect 41827 593947 41893 593948
rect 40723 592550 40789 592551
rect 40723 592486 40724 592550
rect 40788 592486 40789 592550
rect 40723 592485 40789 592486
rect 40726 574701 40786 592485
rect 41827 592380 41893 592381
rect 41827 592316 41828 592380
rect 41892 592316 41893 592380
rect 41827 592315 41893 592316
rect 41830 592050 41890 592315
rect 41462 591990 41890 592050
rect 41462 591970 41522 591990
rect 40910 591910 41522 591970
rect 40910 577829 40970 591910
rect 42014 587890 42074 597211
rect 42750 597005 42810 598435
rect 42747 597004 42813 597005
rect 42747 596940 42748 597004
rect 42812 596940 42813 597004
rect 42747 596939 42813 596940
rect 42195 592108 42261 592109
rect 42195 592044 42196 592108
rect 42260 592044 42261 592108
rect 42195 592043 42261 592044
rect 41462 587830 42074 587890
rect 41091 584900 41157 584901
rect 41091 584836 41092 584900
rect 41156 584836 41157 584900
rect 41091 584835 41157 584836
rect 41094 580005 41154 584835
rect 41091 580004 41157 580005
rect 41091 579940 41092 580004
rect 41156 579940 41157 580004
rect 41091 579939 41157 579940
rect 40907 577828 40973 577829
rect 40907 577764 40908 577828
rect 40972 577764 40973 577828
rect 40907 577763 40973 577764
rect 40723 574700 40789 574701
rect 40723 574636 40724 574700
rect 40788 574636 40789 574700
rect 40723 574635 40789 574636
rect 41462 574021 41522 587830
rect 42198 587210 42258 592043
rect 41646 587150 42258 587210
rect 41459 574020 41525 574021
rect 41459 573956 41460 574020
rect 41524 573956 41525 574020
rect 41459 573955 41525 573956
rect 40539 573476 40605 573477
rect 40539 573412 40540 573476
rect 40604 573412 40605 573476
rect 40539 573411 40605 573412
rect 41646 571573 41706 587150
rect 41827 585172 41893 585173
rect 41827 585108 41828 585172
rect 41892 585108 41893 585172
rect 41827 585107 41893 585108
rect 41643 571572 41709 571573
rect 41643 571508 41644 571572
rect 41708 571508 41709 571572
rect 41643 571507 41709 571508
rect 41830 570213 41890 585107
rect 42195 579460 42261 579461
rect 42195 579396 42196 579460
rect 42260 579396 42261 579460
rect 42195 579395 42261 579396
rect 42011 578372 42077 578373
rect 42011 578308 42012 578372
rect 42076 578308 42077 578372
rect 42011 578307 42077 578308
rect 42014 572661 42074 578307
rect 42198 573477 42258 579395
rect 673683 578644 673749 578645
rect 673683 578580 673684 578644
rect 673748 578580 673749 578644
rect 673683 578579 673749 578580
rect 673686 578370 673746 578579
rect 673502 578310 673746 578370
rect 673502 577965 673562 578310
rect 673499 577964 673565 577965
rect 673499 577900 673500 577964
rect 673564 577900 673565 577964
rect 673499 577899 673565 577900
rect 42195 573476 42261 573477
rect 42195 573412 42196 573476
rect 42260 573412 42261 573476
rect 42195 573411 42261 573412
rect 42011 572660 42077 572661
rect 42011 572596 42012 572660
rect 42076 572596 42077 572660
rect 42011 572595 42077 572596
rect 41827 570212 41893 570213
rect 41827 570148 41828 570212
rect 41892 570148 41893 570212
rect 41827 570147 41893 570148
rect 41091 558788 41157 558789
rect 41091 558724 41092 558788
rect 41156 558724 41157 558788
rect 41091 558723 41157 558724
rect 41094 557553 41154 558723
rect 41091 557552 41157 557553
rect 41091 557488 41092 557552
rect 41156 557488 41157 557552
rect 41091 557487 41157 557488
rect 41827 554028 41893 554029
rect 41827 553964 41828 554028
rect 41892 553964 41893 554028
rect 41827 553963 41893 553964
rect 41830 553410 41890 553963
rect 41462 553350 41890 553410
rect 40723 545596 40789 545597
rect 40723 545532 40724 545596
rect 40788 545532 40789 545596
rect 40723 545531 40789 545532
rect 40539 545324 40605 545325
rect 40539 545260 40540 545324
rect 40604 545260 40605 545324
rect 40539 545259 40605 545260
rect 40542 533357 40602 545259
rect 40726 535261 40786 545531
rect 40723 535260 40789 535261
rect 40723 535196 40724 535260
rect 40788 535196 40789 535260
rect 40723 535195 40789 535196
rect 40539 533356 40605 533357
rect 40539 533292 40540 533356
rect 40604 533292 40605 533356
rect 40539 533291 40605 533292
rect 41462 530773 41522 553350
rect 41827 552804 41893 552805
rect 41827 552740 41828 552804
rect 41892 552740 41893 552804
rect 41827 552739 41893 552740
rect 41830 543750 41890 552739
rect 42195 549540 42261 549541
rect 42195 549476 42196 549540
rect 42260 549476 42261 549540
rect 42195 549475 42261 549476
rect 42198 545325 42258 549475
rect 42195 545324 42261 545325
rect 42195 545260 42196 545324
rect 42260 545260 42261 545324
rect 42195 545259 42261 545260
rect 41646 543690 41890 543750
rect 41646 531725 41706 543690
rect 41827 542332 41893 542333
rect 41827 542268 41828 542332
rect 41892 542268 41893 542332
rect 41827 542267 41893 542268
rect 41643 531724 41709 531725
rect 41643 531660 41644 531724
rect 41708 531660 41709 531724
rect 41643 531659 41709 531660
rect 41459 530772 41525 530773
rect 41459 530708 41460 530772
rect 41524 530708 41525 530772
rect 41459 530707 41525 530708
rect 41830 529005 41890 542267
rect 41827 529004 41893 529005
rect 41827 528940 41828 529004
rect 41892 528940 41893 529004
rect 41827 528939 41893 528940
rect 673870 455293 673930 616115
rect 674238 591157 674298 652835
rect 674422 619037 674482 694587
rect 674606 662421 674666 738107
rect 675342 730829 675402 786659
rect 675339 730828 675405 730829
rect 675339 730764 675340 730828
rect 675404 730764 675405 730828
rect 675339 730763 675405 730764
rect 676078 726613 676138 788019
rect 676811 729876 676877 729877
rect 676811 729812 676812 729876
rect 676876 729812 676877 729876
rect 676811 729811 676877 729812
rect 676075 726612 676141 726613
rect 676075 726548 676076 726612
rect 676140 726548 676141 726612
rect 676075 726547 676141 726548
rect 675339 721580 675405 721581
rect 675339 721516 675340 721580
rect 675404 721516 675405 721580
rect 675339 721515 675405 721516
rect 675342 686221 675402 721515
rect 675523 696828 675589 696829
rect 675523 696764 675524 696828
rect 675588 696764 675589 696828
rect 675523 696763 675589 696764
rect 675339 686220 675405 686221
rect 675339 686156 675340 686220
rect 675404 686156 675405 686220
rect 675339 686155 675405 686156
rect 675526 685949 675586 696763
rect 675523 685948 675589 685949
rect 675523 685884 675524 685948
rect 675588 685884 675589 685948
rect 675523 685883 675589 685884
rect 676075 676428 676141 676429
rect 676075 676364 676076 676428
rect 676140 676364 676141 676428
rect 676075 676363 676141 676364
rect 674603 662420 674669 662421
rect 674603 662356 674604 662420
rect 674668 662356 674669 662420
rect 674603 662355 674669 662356
rect 674787 646100 674853 646101
rect 674787 646036 674788 646100
rect 674852 646036 674853 646100
rect 674787 646035 674853 646036
rect 674790 640253 674850 646035
rect 674787 640252 674853 640253
rect 674787 640188 674788 640252
rect 674852 640188 674853 640252
rect 674787 640187 674853 640188
rect 676078 637533 676138 676363
rect 676814 665821 676874 729811
rect 676811 665820 676877 665821
rect 676811 665756 676812 665820
rect 676876 665756 676877 665820
rect 676811 665755 676877 665756
rect 676075 637532 676141 637533
rect 676075 637468 676076 637532
rect 676140 637468 676141 637532
rect 676075 637467 676141 637468
rect 675155 631412 675221 631413
rect 675155 631348 675156 631412
rect 675220 631348 675221 631412
rect 675155 631347 675221 631348
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 674419 619036 674485 619037
rect 674419 618972 674420 619036
rect 674484 618972 674485 619036
rect 674419 618971 674485 618972
rect 674419 602988 674485 602989
rect 674419 602924 674420 602988
rect 674484 602924 674485 602988
rect 674419 602923 674485 602924
rect 674235 591156 674301 591157
rect 674235 591092 674236 591156
rect 674300 591092 674301 591156
rect 674235 591091 674301 591092
rect 674051 554164 674117 554165
rect 674051 554100 674052 554164
rect 674116 554100 674117 554164
rect 674051 554099 674117 554100
rect 674054 552941 674114 554099
rect 674051 552940 674117 552941
rect 674051 552876 674052 552940
rect 674116 552876 674117 552940
rect 674051 552875 674117 552876
rect 674051 550492 674117 550493
rect 674051 550428 674052 550492
rect 674116 550428 674117 550492
rect 674051 550427 674117 550428
rect 674054 547909 674114 550427
rect 674051 547908 674117 547909
rect 674051 547844 674052 547908
rect 674116 547844 674117 547908
rect 674051 547843 674117 547844
rect 674422 527101 674482 602923
rect 675158 593197 675218 631347
rect 675339 595372 675405 595373
rect 675339 595308 675340 595372
rect 675404 595308 675405 595372
rect 675339 595307 675405 595308
rect 675155 593196 675221 593197
rect 675155 593132 675156 593196
rect 675220 593132 675221 593196
rect 675155 593131 675221 593132
rect 675342 591565 675402 595307
rect 675339 591564 675405 591565
rect 675339 591500 675340 591564
rect 675404 591500 675405 591564
rect 675339 591499 675405 591500
rect 676078 591429 676138 631347
rect 676811 617132 676877 617133
rect 676811 617068 676812 617132
rect 676876 617068 676877 617132
rect 676811 617067 676877 617068
rect 676075 591428 676141 591429
rect 676075 591364 676076 591428
rect 676140 591364 676141 591428
rect 676075 591363 676141 591364
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675339 561916 675405 561917
rect 675339 561852 675340 561916
rect 675404 561852 675405 561916
rect 675339 561851 675405 561852
rect 675342 548453 675402 561851
rect 675339 548452 675405 548453
rect 675339 548388 675340 548452
rect 675404 548388 675405 548452
rect 675339 548387 675405 548388
rect 676078 546821 676138 586195
rect 676814 576877 676874 617067
rect 676811 576876 676877 576877
rect 676811 576812 676812 576876
rect 676876 576812 676877 576876
rect 676811 576811 676877 576812
rect 676259 554708 676325 554709
rect 676259 554644 676260 554708
rect 676324 554644 676325 554708
rect 676259 554643 676325 554644
rect 676262 547637 676322 554643
rect 676811 553892 676877 553893
rect 676811 553828 676812 553892
rect 676876 553828 676877 553892
rect 676811 553827 676877 553828
rect 676259 547636 676325 547637
rect 676259 547572 676260 547636
rect 676324 547572 676325 547636
rect 676259 547571 676325 547572
rect 676075 546820 676141 546821
rect 676075 546756 676076 546820
rect 676140 546756 676141 546820
rect 676075 546755 676141 546756
rect 674419 527100 674485 527101
rect 674419 527036 674420 527100
rect 674484 527036 674485 527100
rect 674419 527035 674485 527036
rect 676814 500989 676874 553827
rect 676995 548316 677061 548317
rect 676995 548252 676996 548316
rect 677060 548252 677061 548316
rect 676995 548251 677061 548252
rect 676998 503709 677058 548251
rect 676995 503708 677061 503709
rect 676995 503644 676996 503708
rect 677060 503644 677061 503708
rect 676995 503643 677061 503644
rect 676811 500988 676877 500989
rect 676811 500924 676812 500988
rect 676876 500924 676877 500988
rect 676811 500923 676877 500924
rect 676029 488884 676095 488885
rect 676029 488820 676030 488884
rect 676094 488820 676095 488884
rect 676029 488819 676095 488820
rect 676032 488610 676092 488819
rect 676032 488550 677242 488610
rect 675891 487932 675957 487933
rect 675891 487868 675892 487932
rect 675956 487930 675957 487932
rect 675956 487870 676322 487930
rect 675956 487868 675957 487870
rect 675891 487867 675957 487868
rect 676262 483030 676322 487870
rect 676262 482970 676874 483030
rect 673867 455292 673933 455293
rect 673867 455228 673868 455292
rect 673932 455228 673933 455292
rect 673867 455227 673933 455228
rect 41827 423604 41893 423605
rect 41827 423540 41828 423604
rect 41892 423540 41893 423604
rect 41827 423539 41893 423540
rect 40907 422312 40973 422313
rect 40907 422248 40908 422312
rect 40972 422248 40973 422312
rect 40907 422247 40973 422248
rect 40723 418708 40789 418709
rect 40723 418644 40724 418708
rect 40788 418644 40789 418708
rect 40723 418643 40789 418644
rect 40539 418436 40605 418437
rect 40539 418372 40540 418436
rect 40604 418372 40605 418436
rect 40539 418371 40605 418372
rect 40542 406741 40602 418371
rect 40539 406740 40605 406741
rect 40539 406676 40540 406740
rect 40604 406676 40605 406740
rect 40539 406675 40605 406676
rect 40726 404565 40786 418643
rect 40910 407013 40970 422247
rect 41830 418170 41890 423539
rect 41462 418110 41890 418170
rect 40907 407012 40973 407013
rect 40907 406948 40908 407012
rect 40972 406948 40973 407012
rect 40907 406947 40973 406948
rect 40723 404564 40789 404565
rect 40723 404500 40724 404564
rect 40788 404500 40789 404564
rect 40723 404499 40789 404500
rect 41462 400077 41522 418110
rect 42011 415308 42077 415309
rect 42011 415244 42012 415308
rect 42076 415244 42077 415308
rect 42011 415243 42077 415244
rect 41827 414628 41893 414629
rect 41827 414564 41828 414628
rect 41892 414564 41893 414628
rect 41827 414563 41893 414564
rect 41459 400076 41525 400077
rect 41459 400012 41460 400076
rect 41524 400012 41525 400076
rect 41459 400011 41525 400012
rect 41830 399397 41890 414563
rect 41827 399396 41893 399397
rect 41827 399332 41828 399396
rect 41892 399332 41893 399396
rect 41827 399331 41893 399332
rect 42014 398853 42074 415243
rect 676814 400485 676874 482970
rect 677182 401301 677242 488550
rect 677179 401300 677245 401301
rect 677179 401236 677180 401300
rect 677244 401236 677245 401300
rect 677179 401235 677245 401236
rect 676811 400484 676877 400485
rect 676811 400420 676812 400484
rect 676876 400420 676877 400484
rect 676811 400419 676877 400420
rect 42011 398852 42077 398853
rect 42011 398788 42012 398852
rect 42076 398788 42077 398852
rect 42011 398787 42077 398788
rect 676075 398852 676141 398853
rect 676075 398788 676076 398852
rect 676140 398788 676141 398852
rect 676075 398787 676141 398788
rect 675339 392868 675405 392869
rect 675339 392804 675340 392868
rect 675404 392804 675405 392868
rect 675339 392803 675405 392804
rect 41459 381852 41525 381853
rect 41459 381788 41460 381852
rect 41524 381788 41525 381852
rect 41459 381787 41525 381788
rect 40723 378996 40789 378997
rect 40723 378932 40724 378996
rect 40788 378932 40789 378996
rect 40723 378931 40789 378932
rect 40539 378588 40605 378589
rect 40539 378524 40540 378588
rect 40604 378524 40605 378588
rect 40539 378523 40605 378524
rect 40542 360093 40602 378523
rect 40726 364173 40786 378931
rect 40907 377772 40973 377773
rect 40907 377708 40908 377772
rect 40972 377708 40973 377772
rect 40907 377707 40973 377708
rect 40910 364853 40970 377707
rect 40907 364852 40973 364853
rect 40907 364788 40908 364852
rect 40972 364788 40973 364852
rect 40907 364787 40973 364788
rect 40723 364172 40789 364173
rect 40723 364108 40724 364172
rect 40788 364108 40789 364172
rect 40723 364107 40789 364108
rect 40539 360092 40605 360093
rect 40539 360028 40540 360092
rect 40604 360028 40605 360092
rect 40539 360027 40605 360028
rect 41462 356965 41522 381787
rect 41643 379404 41709 379405
rect 41643 379340 41644 379404
rect 41708 379340 41709 379404
rect 41643 379339 41709 379340
rect 41646 358050 41706 379339
rect 41827 374644 41893 374645
rect 41827 374580 41828 374644
rect 41892 374580 41893 374644
rect 41827 374579 41893 374580
rect 41830 358733 41890 374579
rect 675342 372877 675402 392803
rect 675891 387700 675957 387701
rect 675891 387636 675892 387700
rect 675956 387636 675957 387700
rect 675891 387635 675957 387636
rect 675894 378589 675954 387635
rect 675891 378588 675957 378589
rect 675891 378524 675892 378588
rect 675956 378524 675957 378588
rect 675891 378523 675957 378524
rect 676078 373693 676138 398787
rect 676259 396812 676325 396813
rect 676259 396748 676260 396812
rect 676324 396748 676325 396812
rect 676259 396747 676325 396748
rect 676262 384981 676322 396747
rect 676443 396404 676509 396405
rect 676443 396340 676444 396404
rect 676508 396340 676509 396404
rect 676443 396339 676509 396340
rect 676259 384980 676325 384981
rect 676259 384916 676260 384980
rect 676324 384916 676325 384980
rect 676259 384915 676325 384916
rect 676446 382261 676506 396339
rect 676627 395180 676693 395181
rect 676627 395116 676628 395180
rect 676692 395116 676693 395180
rect 676627 395115 676693 395116
rect 676443 382260 676509 382261
rect 676443 382196 676444 382260
rect 676508 382196 676509 382260
rect 676443 382195 676509 382196
rect 676630 377501 676690 395115
rect 676627 377500 676693 377501
rect 676627 377436 676628 377500
rect 676692 377436 676693 377500
rect 676627 377435 676693 377436
rect 676075 373692 676141 373693
rect 676075 373628 676076 373692
rect 676140 373628 676141 373692
rect 676075 373627 676141 373628
rect 675339 372876 675405 372877
rect 675339 372812 675340 372876
rect 675404 372812 675405 372876
rect 675339 372811 675405 372812
rect 41827 358732 41893 358733
rect 41827 358668 41828 358732
rect 41892 358668 41893 358732
rect 41827 358667 41893 358668
rect 41646 357990 41890 358050
rect 41459 356964 41525 356965
rect 41459 356900 41460 356964
rect 41524 356900 41525 356964
rect 41459 356899 41525 356900
rect 41830 355741 41890 357990
rect 41827 355740 41893 355741
rect 41827 355676 41828 355740
rect 41892 355676 41893 355740
rect 41827 355675 41893 355676
rect 43299 354516 43365 354517
rect 43299 354452 43300 354516
rect 43364 354452 43365 354516
rect 43299 354451 43365 354452
rect 42195 344316 42261 344317
rect 42195 344252 42196 344316
rect 42260 344252 42261 344316
rect 42195 344251 42261 344252
rect 42198 342141 42258 344251
rect 42195 342140 42261 342141
rect 42195 342076 42196 342140
rect 42260 342076 42261 342140
rect 42195 342075 42261 342076
rect 42747 340236 42813 340237
rect 42747 340172 42748 340236
rect 42812 340172 42813 340236
rect 42747 340171 42813 340172
rect 40539 336972 40605 336973
rect 40539 336908 40540 336972
rect 40604 336908 40605 336972
rect 40539 336907 40605 336908
rect 40542 316029 40602 336907
rect 41827 336564 41893 336565
rect 41827 336500 41828 336564
rect 41892 336500 41893 336564
rect 41827 336499 41893 336500
rect 40907 335748 40973 335749
rect 40907 335684 40908 335748
rect 40972 335684 40973 335748
rect 40907 335683 40973 335684
rect 40723 335340 40789 335341
rect 40723 335276 40724 335340
rect 40788 335276 40789 335340
rect 40723 335275 40789 335276
rect 40726 317389 40786 335275
rect 40910 321197 40970 335683
rect 41459 332892 41525 332893
rect 41459 332828 41460 332892
rect 41524 332828 41525 332892
rect 41459 332827 41525 332828
rect 40907 321196 40973 321197
rect 40907 321132 40908 321196
rect 40972 321132 40973 321196
rect 40907 321131 40973 321132
rect 40723 317388 40789 317389
rect 40723 317324 40724 317388
rect 40788 317324 40789 317388
rect 40723 317323 40789 317324
rect 40539 316028 40605 316029
rect 40539 315964 40540 316028
rect 40604 315964 40605 316028
rect 40539 315963 40605 315964
rect 41462 313717 41522 332827
rect 41643 331804 41709 331805
rect 41643 331740 41644 331804
rect 41708 331740 41709 331804
rect 41643 331739 41709 331740
rect 41646 316050 41706 331739
rect 41830 324869 41890 336499
rect 41827 324868 41893 324869
rect 41827 324804 41828 324868
rect 41892 324804 41893 324868
rect 41827 324803 41893 324804
rect 41646 315990 41890 316050
rect 41830 315621 41890 315990
rect 41827 315620 41893 315621
rect 41827 315556 41828 315620
rect 41892 315556 41893 315620
rect 41827 315555 41893 315556
rect 41459 313716 41525 313717
rect 41459 313652 41460 313716
rect 41524 313652 41525 313716
rect 41459 313651 41525 313652
rect 42750 297669 42810 340171
rect 42931 337652 42997 337653
rect 42931 337588 42932 337652
rect 42996 337588 42997 337652
rect 42931 337587 42997 337588
rect 42934 312765 42994 337587
rect 43302 334661 43362 354451
rect 675523 354244 675589 354245
rect 675523 354180 675524 354244
rect 675588 354180 675589 354244
rect 675523 354179 675589 354180
rect 675339 347716 675405 347717
rect 675339 347652 675340 347716
rect 675404 347652 675405 347716
rect 675339 347651 675405 347652
rect 44219 342956 44285 342957
rect 44219 342892 44220 342956
rect 44284 342892 44285 342956
rect 44219 342891 44285 342892
rect 43299 334660 43365 334661
rect 43299 334596 43300 334660
rect 43364 334596 43365 334660
rect 43299 334595 43365 334596
rect 42931 312764 42997 312765
rect 42931 312700 42932 312764
rect 42996 312700 42997 312764
rect 42931 312699 42997 312700
rect 44222 300117 44282 342891
rect 44587 342412 44653 342413
rect 44587 342348 44588 342412
rect 44652 342348 44653 342412
rect 44587 342347 44653 342348
rect 44403 339828 44469 339829
rect 44403 339764 44404 339828
rect 44468 339764 44469 339828
rect 44403 339763 44469 339764
rect 44219 300116 44285 300117
rect 44219 300052 44220 300116
rect 44284 300052 44285 300116
rect 44219 300051 44285 300052
rect 44406 298485 44466 339763
rect 44590 299301 44650 342347
rect 675342 327997 675402 347651
rect 675526 339421 675586 354179
rect 675891 353836 675957 353837
rect 675891 353772 675892 353836
rect 675956 353772 675957 353836
rect 675891 353771 675957 353772
rect 675894 353290 675954 353771
rect 675894 353230 676690 353290
rect 675707 353020 675773 353021
rect 675707 352956 675708 353020
rect 675772 352956 675773 353020
rect 675707 352955 675773 352956
rect 675710 349210 675770 352955
rect 675891 351796 675957 351797
rect 675891 351732 675892 351796
rect 675956 351732 675957 351796
rect 675891 351731 675957 351732
rect 675894 349890 675954 351731
rect 675894 349830 676322 349890
rect 675710 349150 676138 349210
rect 675523 339420 675589 339421
rect 675523 339356 675524 339420
rect 675588 339356 675589 339420
rect 675523 339355 675589 339356
rect 676078 337925 676138 349150
rect 676262 340237 676322 349830
rect 676443 346628 676509 346629
rect 676443 346564 676444 346628
rect 676508 346564 676509 346628
rect 676443 346563 676509 346564
rect 676259 340236 676325 340237
rect 676259 340172 676260 340236
rect 676324 340172 676325 340236
rect 676259 340171 676325 340172
rect 676075 337924 676141 337925
rect 676075 337860 676076 337924
rect 676140 337860 676141 337924
rect 676075 337859 676141 337860
rect 676446 336565 676506 346563
rect 676443 336564 676509 336565
rect 676443 336500 676444 336564
rect 676508 336500 676509 336564
rect 676443 336499 676509 336500
rect 675339 327996 675405 327997
rect 675339 327932 675340 327996
rect 675404 327932 675405 327996
rect 675339 327931 675405 327932
rect 676630 325685 676690 353230
rect 676627 325684 676693 325685
rect 676627 325620 676628 325684
rect 676692 325620 676693 325684
rect 676627 325619 676693 325620
rect 675891 308820 675957 308821
rect 675891 308756 675892 308820
rect 675956 308756 675957 308820
rect 675891 308755 675957 308756
rect 675894 303650 675954 308755
rect 676075 306644 676141 306645
rect 676075 306580 676076 306644
rect 676140 306580 676141 306644
rect 676075 306579 676141 306580
rect 676078 306390 676138 306579
rect 676078 306330 676874 306390
rect 676259 304978 676325 304979
rect 676259 304914 676260 304978
rect 676324 304914 676325 304978
rect 676259 304913 676325 304914
rect 675894 303590 676138 303650
rect 675891 302700 675957 302701
rect 675891 302636 675892 302700
rect 675956 302636 675957 302700
rect 675891 302635 675957 302636
rect 44587 299300 44653 299301
rect 44587 299236 44588 299300
rect 44652 299236 44653 299300
rect 44587 299235 44653 299236
rect 44403 298484 44469 298485
rect 44403 298420 44404 298484
rect 44468 298420 44469 298484
rect 44403 298419 44469 298420
rect 42747 297668 42813 297669
rect 42747 297604 42748 297668
rect 42812 297604 42813 297668
rect 42747 297603 42813 297604
rect 675707 297396 675773 297397
rect 675707 297332 675708 297396
rect 675772 297332 675773 297396
rect 675707 297331 675773 297332
rect 42195 296852 42261 296853
rect 42195 296788 42196 296852
rect 42260 296788 42261 296852
rect 42195 296787 42261 296788
rect 40539 292592 40605 292593
rect 40539 292528 40540 292592
rect 40604 292528 40605 292592
rect 40539 292527 40605 292528
rect 40542 274277 40602 292527
rect 42011 292228 42077 292229
rect 42011 292164 42012 292228
rect 42076 292164 42077 292228
rect 42011 292163 42077 292164
rect 41827 291956 41893 291957
rect 41827 291892 41828 291956
rect 41892 291892 41893 291956
rect 41827 291891 41893 291892
rect 41830 291410 41890 291891
rect 40726 291350 41890 291410
rect 40726 277133 40786 291350
rect 41827 290052 41893 290053
rect 41827 289988 41828 290052
rect 41892 289988 41893 290052
rect 41827 289987 41893 289988
rect 41830 289830 41890 289987
rect 41462 289770 41890 289830
rect 40907 289236 40973 289237
rect 40907 289172 40908 289236
rect 40972 289172 40973 289236
rect 40907 289171 40973 289172
rect 40910 282301 40970 289171
rect 40907 282300 40973 282301
rect 40907 282236 40908 282300
rect 40972 282236 40973 282300
rect 40907 282235 40973 282236
rect 40723 277132 40789 277133
rect 40723 277068 40724 277132
rect 40788 277068 40789 277132
rect 40723 277067 40789 277068
rect 40539 274276 40605 274277
rect 40539 274212 40540 274276
rect 40604 274212 40605 274276
rect 40539 274211 40605 274212
rect 41462 270469 41522 289770
rect 41827 284340 41893 284341
rect 41827 284276 41828 284340
rect 41892 284276 41893 284340
rect 41827 284275 41893 284276
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 41830 269789 41890 284275
rect 41827 269788 41893 269789
rect 41827 269724 41828 269788
rect 41892 269724 41893 269788
rect 41827 269723 41893 269724
rect 42014 269109 42074 292163
rect 42198 290053 42258 296787
rect 675155 296716 675221 296717
rect 675155 296652 675156 296716
rect 675220 296652 675221 296716
rect 675155 296651 675221 296652
rect 675158 294541 675218 296651
rect 675155 294540 675221 294541
rect 675155 294476 675156 294540
rect 675220 294476 675221 294540
rect 675155 294475 675221 294476
rect 42195 290052 42261 290053
rect 42195 289988 42196 290052
rect 42260 289988 42261 290052
rect 42195 289987 42261 289988
rect 42195 284884 42261 284885
rect 42195 284820 42196 284884
rect 42260 284820 42261 284884
rect 42195 284819 42261 284820
rect 42198 281757 42258 284819
rect 42195 281756 42261 281757
rect 42195 281692 42196 281756
rect 42260 281692 42261 281756
rect 42195 281691 42261 281692
rect 675710 281621 675770 297331
rect 675894 282709 675954 302635
rect 676078 283661 676138 303590
rect 676262 291005 676322 304913
rect 676443 301612 676509 301613
rect 676443 301548 676444 301612
rect 676508 301548 676509 301612
rect 676443 301547 676509 301548
rect 676446 291549 676506 301547
rect 676814 298110 676874 306330
rect 676630 298050 676874 298110
rect 676630 294541 676690 298050
rect 676627 294540 676693 294541
rect 676627 294476 676628 294540
rect 676692 294476 676693 294540
rect 676627 294475 676693 294476
rect 676443 291548 676509 291549
rect 676443 291484 676444 291548
rect 676508 291484 676509 291548
rect 676443 291483 676509 291484
rect 676259 291004 676325 291005
rect 676259 290940 676260 291004
rect 676324 290940 676325 291004
rect 676259 290939 676325 290940
rect 676075 283660 676141 283661
rect 676075 283596 676076 283660
rect 676140 283596 676141 283660
rect 676075 283595 676141 283596
rect 675891 282708 675957 282709
rect 675891 282644 675892 282708
rect 675956 282644 675957 282708
rect 675891 282643 675957 282644
rect 675707 281620 675773 281621
rect 675707 281556 675708 281620
rect 675772 281556 675773 281620
rect 675707 281555 675773 281556
rect 42195 280260 42261 280261
rect 42195 280196 42196 280260
rect 42260 280196 42261 280260
rect 42195 280195 42261 280196
rect 42198 278765 42258 280195
rect 42195 278764 42261 278765
rect 42195 278700 42196 278764
rect 42260 278700 42261 278764
rect 42195 278699 42261 278700
rect 675339 273868 675405 273869
rect 675339 273804 675340 273868
rect 675404 273804 675405 273868
rect 675339 273803 675405 273804
rect 42011 269108 42077 269109
rect 42011 269044 42012 269108
rect 42076 269044 42077 269108
rect 42011 269043 42077 269044
rect 675342 249797 675402 273803
rect 676995 261628 677061 261629
rect 676995 261564 676996 261628
rect 677060 261564 677061 261628
rect 676995 261563 677061 261564
rect 676811 261220 676877 261221
rect 676811 261156 676812 261220
rect 676876 261156 676877 261220
rect 676811 261155 676877 261156
rect 675523 258092 675589 258093
rect 675523 258028 675524 258092
rect 675588 258028 675589 258092
rect 675523 258027 675589 258028
rect 675526 250069 675586 258027
rect 675523 250068 675589 250069
rect 675523 250004 675524 250068
rect 675588 250004 675589 250068
rect 675523 250003 675589 250004
rect 40539 249796 40605 249797
rect 40539 249732 40540 249796
rect 40604 249732 40605 249796
rect 40539 249731 40605 249732
rect 675339 249796 675405 249797
rect 675339 249732 675340 249796
rect 675404 249732 675405 249796
rect 675339 249731 675405 249732
rect 40542 236605 40602 249731
rect 40723 249388 40789 249389
rect 40723 249324 40724 249388
rect 40788 249324 40789 249388
rect 40723 249323 40789 249324
rect 40539 236604 40605 236605
rect 40539 236540 40540 236604
rect 40604 236540 40605 236604
rect 40539 236539 40605 236540
rect 40726 234701 40786 249323
rect 676814 246669 676874 261155
rect 676998 250341 677058 261563
rect 676995 250340 677061 250341
rect 676995 250276 676996 250340
rect 677060 250276 677061 250340
rect 676995 250275 677061 250276
rect 676811 246668 676877 246669
rect 676811 246604 676812 246668
rect 676876 246604 676877 246668
rect 676811 246603 676877 246604
rect 673315 246260 673381 246261
rect 673315 246196 673316 246260
rect 673380 246196 673381 246260
rect 673315 246195 673381 246196
rect 675523 246260 675589 246261
rect 675523 246196 675524 246260
rect 675588 246196 675589 246260
rect 675523 246195 675589 246196
rect 667795 245716 667861 245717
rect 667795 245652 667796 245716
rect 667860 245652 667861 245716
rect 667795 245651 667861 245652
rect 42011 238100 42077 238101
rect 42011 238036 42012 238100
rect 42076 238036 42077 238100
rect 42011 238035 42077 238036
rect 40723 234700 40789 234701
rect 40723 234636 40724 234700
rect 40788 234636 40789 234700
rect 40723 234635 40789 234636
rect 42014 228989 42074 238035
rect 42011 228988 42077 228989
rect 42011 228924 42012 228988
rect 42076 228924 42077 228988
rect 42011 228923 42077 228924
rect 649582 222461 649642 222582
rect 651974 222461 652034 222582
rect 649579 222460 649645 222461
rect 649579 222396 649580 222460
rect 649644 222396 649645 222460
rect 649579 222395 649645 222396
rect 651971 222460 652037 222461
rect 651971 222396 651972 222460
rect 652036 222396 652037 222460
rect 651971 222395 652037 222396
rect 511027 217564 511093 217565
rect 511027 217500 511028 217564
rect 511092 217500 511093 217564
rect 511027 217499 511093 217500
rect 520043 217564 520109 217565
rect 520043 217500 520044 217564
rect 520108 217500 520109 217564
rect 520043 217499 520109 217500
rect 532555 217564 532621 217565
rect 532555 217500 532556 217564
rect 532620 217500 532621 217564
rect 532555 217499 532621 217500
rect 511030 215661 511090 217499
rect 520046 215933 520106 217499
rect 520043 215932 520109 215933
rect 520043 215868 520044 215932
rect 520108 215868 520109 215932
rect 520043 215867 520109 215868
rect 511027 215660 511093 215661
rect 511027 215596 511028 215660
rect 511092 215596 511093 215660
rect 511027 215595 511093 215596
rect 532558 215389 532618 217499
rect 532555 215388 532621 215389
rect 532555 215324 532556 215388
rect 532620 215324 532621 215388
rect 532555 215323 532621 215324
rect 41827 210084 41893 210085
rect 41827 210020 41828 210084
rect 41892 210020 41893 210084
rect 41827 210019 41893 210020
rect 41643 208180 41709 208181
rect 41643 208116 41644 208180
rect 41708 208116 41709 208180
rect 41643 208115 41709 208116
rect 40539 207364 40605 207365
rect 40539 207300 40540 207364
rect 40604 207300 40605 207364
rect 40539 207299 40605 207300
rect 40542 186421 40602 207299
rect 40723 206548 40789 206549
rect 40723 206484 40724 206548
rect 40788 206484 40789 206548
rect 40723 206483 40789 206484
rect 40726 193493 40786 206483
rect 40907 206140 40973 206141
rect 40907 206076 40908 206140
rect 40972 206076 40973 206140
rect 40907 206075 40973 206076
rect 40910 194989 40970 206075
rect 41646 200130 41706 208115
rect 41462 200070 41706 200130
rect 40907 194988 40973 194989
rect 40907 194924 40908 194988
rect 40972 194924 40973 194988
rect 40907 194923 40973 194924
rect 40723 193492 40789 193493
rect 40723 193428 40724 193492
rect 40788 193428 40789 193492
rect 40723 193427 40789 193428
rect 40539 186420 40605 186421
rect 40539 186356 40540 186420
rect 40604 186356 40605 186420
rect 40539 186355 40605 186356
rect 41462 186013 41522 200070
rect 41830 195261 41890 210019
rect 42011 198796 42077 198797
rect 42011 198732 42012 198796
rect 42076 198732 42077 198796
rect 42011 198731 42077 198732
rect 42014 195805 42074 198731
rect 42011 195804 42077 195805
rect 42011 195740 42012 195804
rect 42076 195740 42077 195804
rect 42011 195739 42077 195740
rect 41827 195260 41893 195261
rect 41827 195196 41828 195260
rect 41892 195196 41893 195260
rect 41827 195195 41893 195196
rect 41459 186012 41525 186013
rect 41459 185948 41460 186012
rect 41524 185948 41525 186012
rect 41459 185947 41525 185948
rect 667798 132973 667858 245651
rect 670739 231980 670805 231981
rect 670739 231916 670740 231980
rect 670804 231916 670805 231980
rect 670739 231915 670805 231916
rect 670003 224636 670069 224637
rect 670003 224572 670004 224636
rect 670068 224572 670069 224636
rect 670003 224571 670069 224572
rect 668166 179621 668226 222582
rect 670006 220829 670066 224571
rect 670555 223956 670621 223957
rect 670555 223892 670556 223956
rect 670620 223892 670621 223956
rect 670555 223891 670621 223892
rect 670371 223684 670437 223685
rect 670371 223620 670372 223684
rect 670436 223620 670437 223684
rect 670371 223619 670437 223620
rect 670003 220828 670069 220829
rect 670003 220764 670004 220828
rect 670068 220764 670069 220828
rect 670003 220763 670069 220764
rect 670374 219450 670434 223619
rect 670558 220421 670618 223891
rect 670555 220420 670621 220421
rect 670555 220356 670556 220420
rect 670620 220356 670621 220420
rect 670555 220355 670621 220356
rect 670374 219390 670618 219450
rect 669635 218108 669701 218109
rect 669635 218044 669636 218108
rect 669700 218044 669701 218108
rect 669635 218043 669701 218044
rect 669083 217292 669149 217293
rect 669083 217228 669084 217292
rect 669148 217228 669149 217292
rect 669083 217227 669149 217228
rect 669086 212550 669146 217227
rect 669086 212490 669514 212550
rect 669267 205732 669333 205733
rect 669267 205668 669268 205732
rect 669332 205668 669333 205732
rect 669267 205667 669333 205668
rect 669270 205461 669330 205667
rect 669267 205460 669333 205461
rect 669267 205396 669268 205460
rect 669332 205396 669333 205460
rect 669267 205395 669333 205396
rect 669267 196076 669333 196077
rect 669267 196012 669268 196076
rect 669332 196012 669333 196076
rect 669267 196011 669333 196012
rect 669270 186330 669330 196011
rect 669454 191725 669514 212490
rect 669638 205733 669698 218043
rect 670371 216476 670437 216477
rect 670371 216412 670372 216476
rect 670436 216412 670437 216476
rect 670371 216411 670437 216412
rect 669819 215932 669885 215933
rect 669819 215868 669820 215932
rect 669884 215868 669885 215932
rect 669819 215867 669885 215868
rect 669822 214845 669882 215867
rect 669819 214844 669885 214845
rect 669819 214780 669820 214844
rect 669884 214780 669885 214844
rect 669819 214779 669885 214780
rect 670374 211173 670434 216411
rect 670558 215389 670618 219390
rect 670555 215388 670621 215389
rect 670555 215324 670556 215388
rect 670620 215324 670621 215388
rect 670555 215323 670621 215324
rect 670371 211172 670437 211173
rect 670371 211108 670372 211172
rect 670436 211108 670437 211172
rect 670371 211107 670437 211108
rect 669635 205732 669701 205733
rect 669635 205668 669636 205732
rect 669700 205668 669701 205732
rect 669635 205667 669701 205668
rect 669635 205460 669701 205461
rect 669635 205396 669636 205460
rect 669700 205396 669701 205460
rect 669635 205395 669701 205396
rect 669638 196077 669698 205395
rect 670742 198797 670802 231915
rect 672579 227084 672645 227085
rect 672579 227020 672580 227084
rect 672644 227020 672645 227084
rect 672579 227019 672645 227020
rect 671475 224364 671541 224365
rect 671475 224300 671476 224364
rect 671540 224300 671541 224364
rect 671475 224299 671541 224300
rect 671478 223685 671538 224299
rect 671475 223684 671541 223685
rect 671475 223620 671476 223684
rect 671540 223620 671541 223684
rect 671475 223619 671541 223620
rect 672582 200837 672642 227019
rect 672579 200836 672645 200837
rect 672579 200772 672580 200836
rect 672644 200772 672645 200836
rect 672579 200771 672645 200772
rect 670739 198796 670805 198797
rect 670739 198732 670740 198796
rect 670804 198732 670805 198796
rect 670739 198731 670805 198732
rect 669635 196076 669701 196077
rect 669635 196012 669636 196076
rect 669700 196012 669701 196076
rect 669635 196011 669701 196012
rect 669451 191724 669517 191725
rect 669451 191660 669452 191724
rect 669516 191660 669517 191724
rect 669451 191659 669517 191660
rect 669270 186270 669514 186330
rect 668163 179620 668229 179621
rect 668163 179556 668164 179620
rect 668228 179556 668229 179620
rect 668163 179555 668229 179556
rect 669454 157350 669514 186270
rect 673131 181660 673197 181661
rect 673131 181596 673132 181660
rect 673196 181596 673197 181660
rect 673131 181595 673197 181596
rect 673134 161125 673194 181595
rect 673318 179485 673378 246195
rect 675526 235517 675586 246195
rect 676811 241772 676877 241773
rect 676811 241708 676812 241772
rect 676876 241708 676877 241772
rect 676811 241707 676877 241708
rect 675523 235516 675589 235517
rect 675523 235452 675524 235516
rect 675588 235452 675589 235516
rect 675523 235451 675589 235452
rect 674235 228580 674301 228581
rect 674235 228516 674236 228580
rect 674300 228516 674301 228580
rect 674235 228515 674301 228516
rect 675523 228580 675589 228581
rect 675523 228516 675524 228580
rect 675588 228516 675589 228580
rect 675523 228515 675589 228516
rect 674051 226540 674117 226541
rect 674051 226476 674052 226540
rect 674116 226476 674117 226540
rect 674051 226475 674117 226476
rect 673867 215932 673933 215933
rect 673867 215868 673868 215932
rect 673932 215868 673933 215932
rect 673867 215867 673933 215868
rect 673870 213621 673930 215867
rect 673867 213620 673933 213621
rect 673867 213556 673868 213620
rect 673932 213556 673933 213620
rect 673867 213555 673933 213556
rect 673315 179484 673381 179485
rect 673315 179420 673316 179484
rect 673380 179420 673381 179484
rect 673315 179419 673381 179420
rect 673131 161124 673197 161125
rect 673131 161060 673132 161124
rect 673196 161060 673197 161124
rect 673131 161059 673197 161060
rect 669270 157290 669514 157350
rect 669270 140453 669330 157290
rect 669267 140452 669333 140453
rect 669267 140388 669268 140452
rect 669332 140388 669333 140452
rect 669267 140387 669333 140388
rect 667795 132972 667861 132973
rect 667795 132908 667796 132972
rect 667860 132908 667861 132972
rect 667795 132907 667861 132908
rect 674054 115021 674114 226475
rect 674238 206957 674298 228515
rect 675526 224970 675586 228515
rect 675342 224910 675586 224970
rect 674235 206956 674301 206957
rect 674235 206892 674236 206956
rect 674300 206892 674301 206956
rect 674235 206891 674301 206892
rect 675342 189141 675402 224910
rect 676814 220010 676874 241707
rect 683803 227084 683869 227085
rect 683803 227020 683804 227084
rect 683868 227020 683869 227084
rect 683803 227019 683869 227020
rect 683806 223821 683866 227019
rect 683803 223820 683869 223821
rect 683803 223756 683804 223820
rect 683868 223756 683869 223820
rect 683803 223755 683869 223756
rect 676078 219950 676874 220010
rect 676078 219877 676138 219950
rect 676029 219876 676138 219877
rect 676029 219812 676030 219876
rect 676094 219814 676138 219876
rect 676094 219812 676095 219814
rect 676029 219811 676095 219812
rect 675523 218652 675589 218653
rect 675523 218588 675524 218652
rect 675588 218588 675589 218652
rect 675523 218587 675589 218588
rect 675526 213210 675586 218587
rect 675707 217700 675773 217701
rect 675707 217636 675708 217700
rect 675772 217636 675773 217700
rect 675707 217635 675773 217636
rect 675710 213890 675770 217635
rect 675891 215252 675957 215253
rect 675891 215188 675892 215252
rect 675956 215250 675957 215252
rect 675956 215190 676690 215250
rect 675956 215188 675957 215190
rect 675891 215187 675957 215188
rect 675891 214572 675957 214573
rect 675891 214508 675892 214572
rect 675956 214570 675957 214572
rect 675956 214510 676506 214570
rect 675956 214508 675957 214510
rect 675891 214507 675957 214508
rect 675710 213830 676322 213890
rect 675526 213150 676138 213210
rect 675707 212532 675773 212533
rect 675707 212468 675708 212532
rect 675772 212468 675773 212532
rect 675707 212467 675773 212468
rect 675710 205650 675770 212467
rect 675710 205590 675954 205650
rect 675894 192813 675954 205590
rect 676078 193221 676138 213150
rect 676262 202741 676322 213830
rect 676259 202740 676325 202741
rect 676259 202676 676260 202740
rect 676324 202676 676325 202740
rect 676259 202675 676325 202676
rect 676446 200021 676506 214510
rect 676443 200020 676509 200021
rect 676443 199956 676444 200020
rect 676508 199956 676509 200020
rect 676443 199955 676509 199956
rect 676630 194581 676690 215190
rect 676811 197844 676877 197845
rect 676811 197780 676812 197844
rect 676876 197780 676877 197844
rect 676811 197779 676877 197780
rect 676627 194580 676693 194581
rect 676627 194516 676628 194580
rect 676692 194516 676693 194580
rect 676627 194515 676693 194516
rect 676075 193220 676141 193221
rect 676075 193156 676076 193220
rect 676140 193156 676141 193220
rect 676075 193155 676141 193156
rect 675891 192812 675957 192813
rect 675891 192748 675892 192812
rect 675956 192748 675957 192812
rect 675891 192747 675957 192748
rect 675339 189140 675405 189141
rect 675339 189076 675340 189140
rect 675404 189076 675405 189140
rect 675339 189075 675405 189076
rect 676814 176673 676874 197779
rect 676811 176672 676877 176673
rect 676811 176608 676812 176672
rect 676876 176608 676877 176672
rect 676811 176607 676877 176608
rect 675707 173636 675773 173637
rect 675707 173572 675708 173636
rect 675772 173572 675773 173636
rect 675707 173571 675773 173572
rect 675523 172412 675589 172413
rect 675523 172348 675524 172412
rect 675588 172348 675589 172412
rect 675523 172347 675589 172348
rect 675526 169557 675586 172347
rect 675523 169556 675589 169557
rect 675523 169492 675524 169556
rect 675588 169492 675589 169556
rect 675523 169491 675589 169492
rect 675339 167516 675405 167517
rect 675339 167452 675340 167516
rect 675404 167452 675405 167516
rect 675339 167451 675405 167452
rect 675342 147661 675402 167451
rect 675710 167010 675770 173571
rect 675891 170780 675957 170781
rect 675891 170716 675892 170780
rect 675956 170716 675957 170780
rect 675891 170715 675957 170716
rect 675894 170370 675954 170715
rect 675894 170310 676690 170370
rect 675891 169692 675957 169693
rect 675891 169628 675892 169692
rect 675956 169690 675957 169692
rect 675956 169630 676322 169690
rect 675956 169628 675957 169630
rect 675891 169627 675957 169628
rect 675710 166950 676138 167010
rect 676078 148477 676138 166950
rect 676262 151469 676322 169630
rect 676443 166428 676509 166429
rect 676443 166364 676444 166428
rect 676508 166364 676509 166428
rect 676443 166363 676509 166364
rect 676446 155821 676506 166363
rect 676443 155820 676509 155821
rect 676443 155756 676444 155820
rect 676508 155756 676509 155820
rect 676443 155755 676509 155756
rect 676630 155549 676690 170310
rect 676627 155548 676693 155549
rect 676627 155484 676628 155548
rect 676692 155484 676693 155548
rect 676627 155483 676693 155484
rect 676259 151468 676325 151469
rect 676259 151404 676260 151468
rect 676324 151404 676325 151468
rect 676259 151403 676325 151404
rect 676075 148476 676141 148477
rect 676075 148412 676076 148476
rect 676140 148412 676141 148476
rect 676075 148411 676141 148412
rect 675339 147660 675405 147661
rect 675339 147596 675340 147660
rect 675404 147596 675405 147660
rect 675339 147595 675405 147596
rect 676443 127396 676509 127397
rect 676443 127332 676444 127396
rect 676508 127332 676509 127396
rect 676443 127331 676509 127332
rect 676075 126988 676141 126989
rect 676075 126924 676076 126988
rect 676140 126924 676141 126988
rect 676075 126923 676141 126924
rect 675339 122364 675405 122365
rect 675339 122300 675340 122364
rect 675404 122300 675405 122364
rect 675339 122299 675405 122300
rect 674051 115020 674117 115021
rect 674051 114956 674052 115020
rect 674116 114956 674117 115020
rect 674051 114955 674117 114956
rect 675342 101965 675402 122299
rect 675707 117332 675773 117333
rect 675707 117268 675708 117332
rect 675772 117268 675773 117332
rect 675707 117267 675773 117268
rect 675710 111349 675770 117267
rect 675707 111348 675773 111349
rect 675707 111284 675708 111348
rect 675772 111284 675773 111348
rect 675707 111283 675773 111284
rect 676078 108221 676138 126923
rect 676259 124540 676325 124541
rect 676259 124476 676260 124540
rect 676324 124476 676325 124540
rect 676259 124475 676325 124476
rect 676262 110397 676322 124475
rect 676446 112437 676506 127331
rect 676811 120052 676877 120053
rect 676811 119988 676812 120052
rect 676876 119988 676877 120052
rect 676811 119987 676877 119988
rect 676443 112436 676509 112437
rect 676443 112372 676444 112436
rect 676508 112372 676509 112436
rect 676443 112371 676509 112372
rect 676814 111757 676874 119987
rect 676811 111756 676877 111757
rect 676811 111692 676812 111756
rect 676876 111692 676877 111756
rect 676811 111691 676877 111692
rect 676259 110396 676325 110397
rect 676259 110332 676260 110396
rect 676324 110332 676325 110396
rect 676259 110331 676325 110332
rect 676075 108220 676141 108221
rect 676075 108156 676076 108220
rect 676140 108156 676141 108220
rect 676075 108155 676141 108156
rect 675339 101964 675405 101965
rect 675339 101900 675340 101964
rect 675404 101900 675405 101964
rect 675339 101899 675405 101900
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 633939 95436 634005 95437
rect 633939 95372 633940 95436
rect 634004 95372 634005 95436
rect 633939 95371 634005 95372
rect 633942 78573 634002 95371
rect 637254 84210 637314 96867
rect 647187 96524 647253 96525
rect 647187 96460 647188 96524
rect 647252 96460 647253 96524
rect 647187 96459 647253 96460
rect 647190 94298 647250 96459
rect 650318 93125 650378 93382
rect 650315 93124 650381 93125
rect 650315 93060 650316 93124
rect 650380 93060 650381 93124
rect 650315 93059 650381 93060
rect 637070 84150 637314 84210
rect 633939 78572 634005 78573
rect 633939 78508 633940 78572
rect 634004 78508 634005 78572
rect 633939 78507 634005 78508
rect 637070 78165 637130 84150
rect 637067 78164 637133 78165
rect 637067 78100 637068 78164
rect 637132 78100 637133 78164
rect 637067 78099 637133 78100
rect 460795 55044 460861 55045
rect 460795 54980 460796 55044
rect 460860 54980 460861 55044
rect 460795 54979 460861 54980
rect 460798 53957 460858 54979
rect 462635 54772 462701 54773
rect 462635 54708 462636 54772
rect 462700 54708 462701 54772
rect 462635 54707 462701 54708
rect 460795 53956 460861 53957
rect 460795 53892 460796 53956
rect 460860 53892 460861 53956
rect 460795 53891 460861 53892
rect 462638 53685 462698 54707
rect 462635 53684 462701 53685
rect 462635 53620 462636 53684
rect 462700 53620 462701 53684
rect 462635 53619 462701 53620
rect 518755 48924 518821 48925
rect 518755 48860 518756 48924
rect 518820 48860 518821 48924
rect 518755 48859 518821 48860
rect 515443 47836 515509 47837
rect 515443 47772 515444 47836
rect 515508 47772 515509 47836
rect 515443 47771 515509 47772
rect 461347 44300 461413 44301
rect 461347 44236 461348 44300
rect 461412 44236 461413 44300
rect 461347 44235 461413 44236
rect 463739 44300 463805 44301
rect 463739 44236 463740 44300
rect 463804 44236 463805 44300
rect 463739 44235 463805 44236
rect 464107 44300 464173 44301
rect 464107 44236 464108 44300
rect 464172 44236 464173 44300
rect 464107 44235 464173 44236
rect 141739 44028 141805 44029
rect 141739 43964 141740 44028
rect 141804 43964 141805 44028
rect 141739 43963 141805 43964
rect 141742 40357 141802 43963
rect 415531 42124 415597 42125
rect 415531 42060 415532 42124
rect 415596 42060 415597 42124
rect 415531 42059 415597 42060
rect 365667 41852 365733 41853
rect 365667 41788 365668 41852
rect 365732 41788 365733 41852
rect 365667 41787 365733 41788
rect 365670 41258 365730 41787
rect 403019 41852 403085 41853
rect 403019 41850 403020 41852
rect 402802 41790 403020 41850
rect 403019 41788 403020 41790
rect 403084 41788 403085 41852
rect 403019 41787 403085 41788
rect 415534 40578 415594 42059
rect 421971 41852 422037 41853
rect 421971 41788 421972 41852
rect 422036 41850 422037 41852
rect 422036 41790 422162 41850
rect 422036 41788 422037 41790
rect 421971 41787 422037 41788
rect 441843 41852 441909 41853
rect 441843 41850 441844 41852
rect 441626 41790 441844 41850
rect 441843 41788 441844 41790
rect 441908 41788 441909 41852
rect 441843 41787 441909 41788
rect 460795 41852 460861 41853
rect 460795 41788 460796 41852
rect 460860 41850 460861 41852
rect 460979 41852 461045 41853
rect 460979 41850 460980 41852
rect 460860 41790 460980 41850
rect 460860 41788 460861 41790
rect 460795 41787 460861 41788
rect 460979 41788 460980 41790
rect 461044 41788 461045 41852
rect 460979 41787 461045 41788
rect 461350 40578 461410 44235
rect 463742 41938 463802 44235
rect 464110 41853 464170 44235
rect 515446 42125 515506 47771
rect 518758 42805 518818 48859
rect 529611 48108 529677 48109
rect 529611 48044 529612 48108
rect 529676 48044 529677 48108
rect 529611 48043 529677 48044
rect 526483 47836 526549 47837
rect 526483 47772 526484 47836
rect 526548 47772 526549 47836
rect 526483 47771 526549 47772
rect 520963 47564 521029 47565
rect 520963 47500 520964 47564
rect 521028 47500 521029 47564
rect 520963 47499 521029 47500
rect 518755 42804 518821 42805
rect 518755 42740 518756 42804
rect 518820 42740 518821 42804
rect 518755 42739 518821 42740
rect 520966 42125 521026 47499
rect 522067 47292 522133 47293
rect 522067 47228 522068 47292
rect 522132 47228 522133 47292
rect 522067 47227 522133 47228
rect 522070 42125 522130 47227
rect 526486 42125 526546 47771
rect 529614 42125 529674 48043
rect 515443 42124 515509 42125
rect 515443 42060 515444 42124
rect 515508 42060 515509 42124
rect 515443 42059 515509 42060
rect 520963 42124 521029 42125
rect 520963 42060 520964 42124
rect 521028 42060 521029 42124
rect 520963 42059 521029 42060
rect 522067 42124 522133 42125
rect 522067 42060 522068 42124
rect 522132 42060 522133 42124
rect 522067 42059 522133 42060
rect 526483 42124 526549 42125
rect 526483 42060 526484 42124
rect 526548 42060 526549 42124
rect 526483 42059 526549 42060
rect 529611 42124 529677 42125
rect 529611 42060 529612 42124
rect 529676 42060 529677 42124
rect 529611 42059 529677 42060
rect 464107 41852 464173 41853
rect 464107 41788 464108 41852
rect 464172 41788 464173 41852
rect 464107 41787 464173 41788
rect 141739 40356 141805 40357
rect 141739 40292 141740 40356
rect 141804 40292 141805 40356
rect 141739 40291 141805 40292
<< via4 >>
rect 591902 223412 592138 223498
rect 591902 223348 591988 223412
rect 591988 223348 592052 223412
rect 592052 223348 592138 223412
rect 591902 223262 592138 223348
rect 649494 222582 649730 222818
rect 651886 222582 652122 222818
rect 668078 222582 668314 222818
rect 647102 94062 647338 94298
rect 650230 93382 650466 93618
rect 361902 41852 362138 41938
rect 361902 41788 361988 41852
rect 361988 41788 362052 41852
rect 362052 41788 362138 41852
rect 361902 41702 362138 41788
rect 402566 41702 402802 41938
rect 365582 41022 365818 41258
rect 422162 41702 422398 41938
rect 441390 41702 441626 41938
rect 463654 41702 463890 41938
rect 415446 40342 415682 40578
rect 461262 40342 461498 40578
<< metal5 >>
rect 78610 1018624 90778 1030789
rect 130010 1018624 142178 1030789
rect 181410 1018624 193578 1030789
rect 231810 1018624 243978 1030789
rect 284410 1018624 296578 1030789
rect 334810 1018624 346978 1030789
rect 386210 1018624 398378 1030789
rect 475210 1018624 487378 1030789
rect 526610 1018624 538778 1030789
rect 577010 1018624 589178 1030789
rect 628410 1018624 640578 1030789
rect 6811 956610 18976 968778
rect 698624 953022 710789 965190
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 591860 223498 592180 223540
rect 591860 223262 591902 223498
rect 592138 223262 592180 223498
rect 591860 222860 592180 223262
rect 591860 222818 649772 222860
rect 591860 222582 649494 222818
rect 649730 222582 649772 222818
rect 591860 222540 649772 222582
rect 651844 222818 668356 222860
rect 651844 222582 651886 222818
rect 652122 222582 668078 222818
rect 668314 222582 668356 222818
rect 651844 222540 668356 222582
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 647060 94298 647748 94340
rect 647060 94062 647102 94298
rect 647338 94062 647748 94298
rect 647060 94020 647748 94062
rect 647428 93660 647748 94020
rect 647428 93618 650508 93660
rect 647428 93382 650230 93618
rect 650466 93382 650508 93618
rect 647428 93340 650508 93382
rect 6167 70054 19620 80934
rect 361860 41938 402844 41980
rect 361860 41702 361902 41938
rect 362138 41702 402566 41938
rect 402802 41702 402844 41938
rect 361860 41660 402844 41702
rect 403444 41660 412044 41980
rect 403444 41300 403764 41660
rect 365540 41258 403764 41300
rect 365540 41022 365582 41258
rect 365818 41022 403764 41258
rect 365540 40980 403764 41022
rect 411724 41300 412044 41660
rect 412460 41660 421796 41980
rect 422120 41938 441668 41980
rect 422120 41702 422162 41938
rect 422398 41702 441390 41938
rect 441626 41702 441668 41938
rect 422120 41660 441668 41702
rect 442084 41660 450684 41980
rect 412460 41300 412780 41660
rect 411724 40980 412780 41300
rect 421476 41300 421796 41660
rect 442084 41300 442404 41660
rect 421476 40980 442404 41300
rect 450364 41300 450684 41660
rect 451100 41660 461080 41980
rect 451100 41300 451420 41660
rect 450364 40980 451420 41300
rect 460760 41300 461080 41660
rect 461404 41938 463932 41980
rect 461404 41702 463654 41938
rect 463890 41702 463932 41938
rect 461404 41660 463932 41702
rect 461404 41300 461724 41660
rect 460760 40980 461724 41300
rect 415404 40578 461540 40620
rect 415404 40342 415446 40578
rect 415682 40342 461262 40578
rect 461498 40342 461540 40578
rect 415404 40300 461540 40342
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use caravan_logo  caravan_logo
timestamp 0
transform 1 0 255300 0 1 6032
box 0 0 1 1
use caravan_motto  caravan_motto
timestamp 0
transform 1 0 -54560 0 1 -52
box 0 0 1 1
use copyright_block_a  copyright_block_a
timestamp 0
transform 1 0 149582 0 1 16298
box 0 0 1 1
use open_source  open_source
timestamp 0
transform 1 0 206074 0 1 2336
box 0 0 1 1
use xres_buf  rstb_level
timestamp 1666279203
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use user_id_textblock  user_id_textblock
timestamp 0
transform 1 0 96272 0 1 6890
box 0 0 1 1
use caravel_clocking  clock_ctrl
timestamp 1666279203
transform 1 0 626764 0 1 55284
box 136 496 20000 20000
use buff_flash_clkrst  flash_clkrst_buffers
timestamp 1666279203
transform 1 0 458400 0 1 47600
box 330 0 7699 5000
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1666279203
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1666279203
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1666279203
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use digital_pll  pll
timestamp 1666279203
transform 1 0 628146 0 1 80944
box 0 0 20000 15000
use simple_por  por
timestamp 1666279203
transform 1 0 650146 0 -1 55282
box -14 11 11344 8684
use user_id_programming  user_id_value
timestamp 1666279203
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1666279203
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1666279203
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1666279203
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1666279203
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1666279203
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1666279203
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1666279203
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use spare_logic_block  spare_logic\[2\]
timestamp 1666279203
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1666279203
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1666279203
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1666279203
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use mgmt_protect  mgmt_buffers
timestamp 1666279203
transform 1 0 128180 0 1 232036
box 1066 -400 424400 32400
use spare_logic_block  spare_logic\[0\]
timestamp 1666279203
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1666279203
transform 1 0 108632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1666279203
transform 1 0 578632 0 1 232528
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1666279203
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1666279203
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1666279203
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1666279203
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1666279203
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1666279203
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1666279203
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1666279203
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1666279203
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1666279203
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1666279203
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1666279203
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1666279203
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1666279203
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1666279203
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1666279203
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1666279203
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1666279203
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1666279203
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1666279203
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1666279203
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1666279203
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1666279203
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1666279203
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1666279203
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1666279203
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1666279203
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1666279203
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1666279203
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1666279203
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1666279203
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1666279203
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1666279203
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1666279203
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1666279203
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1666279203
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1666279203
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1666279203
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1666279203
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1666279203
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1666279203
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1666279203
transform -1 0 710203 0 1 884800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1666279203
transform -1 0 709467 0 1 897800
box -38 0 6018 2224
use caravan_power_routing  caravan_power_routing
timestamp 1666279203
transform 1 0 0 0 1 0
box 6022 30806 711814 997678
use caravan_signal_routing  caravan_signal_routing
timestamp 1666279203
transform 1 0 0 0 1 0
box 39764 415548 677806 997846
use user_analog_project_wrapper  mprj
timestamp 1666279203
transform 1 0 65308 0 1 278718
box -800 -800 584800 704800
use chip_io_alt  padframe
timestamp 1666279203
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use gpio_signal_buffering_alt  sigbuf
timestamp 1666279203
transform 1 0 0 0 1 0
box 40023 41960 677583 728321
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698624 953022 710789 965190 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 628410 1018624 640578 1030789 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 526610 1018624 538778 1030789 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 475210 1018624 487378 1030789 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 386210 1018624 398378 1030789 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 284410 1018624 296578 1030789 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 231810 1018624 243978 1030789 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 181410 1018624 193578 1030789 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 130010 1018624 142178 1030789 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 78610 1018624 90778 1030789 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6811 956610 18976 968778 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144150 18309 6 resetb
port 44 nsew signal input
rlabel metal5 s 6167 70054 19620 80934 6 vccd
port 45 nsew signal bidirectional
rlabel metal5 s 697980 909666 711433 920546 6 vccd1
port 46 nsew signal bidirectional
rlabel metal5 s 6167 914054 19620 924934 6 vccd2
port 47 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18976 6 vdda
port 48 nsew signal bidirectional
rlabel metal5 s 698624 819822 710789 831990 6 vdda1
port 49 nsew signal bidirectional
rlabel metal5 s 698624 505222 710789 517390 6 vdda1_2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 484410 18976 496578 6 vdda2
port 51 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio
port 52 nsew signal bidirectional
rlabel metal5 s 6811 871210 18976 883378 6 vddio_2
port 53 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18976 6 vssa
port 54 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1
port 55 nsew signal bidirectional
rlabel metal5 s 698624 417022 710789 429190 6 vssa1_2
port 56 nsew signal bidirectional
rlabel metal5 s 6811 829010 18976 841178 6 vssa2
port 57 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19620 6 vssd
port 58 nsew signal bidirectional
rlabel metal5 s 697980 461866 711433 472746 6 vssd1
port 59 nsew signal bidirectional
rlabel metal5 s 6167 442854 19620 453734 6 vssd2
port 60 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio
port 61 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030789 6 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
