magic
tech sky130A
magscale 1 2
timestamp 1637463856
<< error_p >>
rect 111554 1006757 112632 1006758
rect 111554 1006005 111555 1006757
rect 112631 1006005 112632 1006757
rect 111554 1006004 112632 1006005
rect 162954 1006757 164032 1006758
rect 162954 1006005 162955 1006757
rect 164031 1006005 164032 1006757
rect 162954 1006004 164032 1006005
rect 214354 1006757 215432 1006758
rect 214354 1006005 214355 1006757
rect 215431 1006005 215432 1006757
rect 214354 1006004 215432 1006005
rect 265754 1006757 266832 1006758
rect 265754 1006005 265755 1006757
rect 266831 1006005 266832 1006757
rect 265754 1006004 266832 1006005
rect 317354 1006757 318432 1006758
rect 317354 1006005 317355 1006757
rect 318431 1006005 318432 1006757
rect 317354 1006004 318432 1006005
rect 367754 1006757 368832 1006758
rect 367754 1006005 367755 1006757
rect 368831 1006005 368832 1006757
rect 367754 1006004 368832 1006005
rect 435154 1006757 436232 1006758
rect 435154 1006005 435155 1006757
rect 436231 1006005 436232 1006757
rect 435154 1006004 436232 1006005
rect 512154 1006757 513232 1006758
rect 512154 1006005 512155 1006757
rect 513231 1006005 513232 1006757
rect 512154 1006004 513232 1006005
rect 563554 1006757 564632 1006758
rect 563554 1006005 563555 1006757
rect 564631 1006005 564632 1006757
rect 563554 1006004 564632 1006005
rect 109980 1000219 111064 1000220
rect 109980 999459 109981 1000219
rect 111063 999459 111064 1000219
rect 109980 999458 111064 999459
rect 161380 1000219 162464 1000220
rect 161380 999459 161381 1000219
rect 162463 999459 162464 1000219
rect 161380 999458 162464 999459
rect 212780 1000219 213864 1000220
rect 212780 999459 212781 1000219
rect 213863 999459 213864 1000219
rect 212780 999458 213864 999459
rect 264180 1000219 265264 1000220
rect 264180 999459 264181 1000219
rect 265263 999459 265264 1000219
rect 264180 999458 265264 999459
rect 315780 1000219 316864 1000220
rect 315780 999459 315781 1000219
rect 316863 999459 316864 1000219
rect 315780 999458 316864 999459
rect 366180 1000219 367264 1000220
rect 366180 999459 366181 1000219
rect 367263 999459 367264 1000219
rect 366180 999458 367264 999459
rect 433580 1000219 434664 1000220
rect 433580 999459 433581 1000219
rect 434663 999459 434664 1000219
rect 433580 999458 434664 999459
rect 510580 1000219 511664 1000220
rect 510580 999459 510581 1000219
rect 511663 999459 511664 1000219
rect 510580 999458 511664 999459
rect 561980 1000219 563064 1000220
rect 561980 999459 561981 1000219
rect 563063 999459 563064 1000219
rect 561980 999458 563064 999459
rect 30820 946631 31574 946632
rect 30820 945555 30821 946631
rect 31573 945555 31574 946631
rect 30820 945554 31574 945555
rect 37358 945063 38120 945064
rect 37358 943981 37359 945063
rect 38119 943981 38120 945063
rect 37358 943980 38120 943981
rect 686002 943031 686756 943032
rect 686002 941955 686003 943031
rect 686755 941955 686756 943031
rect 686002 941954 686756 941955
rect 679456 941463 680218 941464
rect 679456 940381 679457 941463
rect 680217 940381 680218 941463
rect 679456 940380 680218 940381
rect 30820 820831 31574 820832
rect 30820 819755 30821 820831
rect 31573 819755 31574 820831
rect 30820 819754 31574 819755
rect 37358 819263 38120 819264
rect 37358 818181 37359 819263
rect 38119 818181 38120 819263
rect 37358 818180 38120 818181
rect 30820 777631 31574 777632
rect 30820 776555 30821 777631
rect 31573 776555 31574 777631
rect 30820 776554 31574 776555
rect 37358 776063 38120 776064
rect 37358 774981 37359 776063
rect 38119 774981 38120 776063
rect 37358 774980 38120 774981
rect 686012 764631 686766 764632
rect 686012 763555 686013 764631
rect 686765 763555 686766 764631
rect 686012 763554 686766 763555
rect 679466 763063 680228 763064
rect 679466 761981 679467 763063
rect 680227 761981 680228 763063
rect 679466 761980 680228 761981
rect 30820 734431 31574 734432
rect 30820 733355 30821 734431
rect 31573 733355 31574 734431
rect 30820 733354 31574 733355
rect 37358 732863 38120 732864
rect 37358 731781 37359 732863
rect 38119 731781 38120 732863
rect 37358 731780 38120 731781
rect 686012 719631 686766 719632
rect 686012 718555 686013 719631
rect 686765 718555 686766 719631
rect 686012 718554 686766 718555
rect 679466 718063 680228 718064
rect 679466 716981 679467 718063
rect 680227 716981 680228 718063
rect 679466 716980 680228 716981
rect 30820 691231 31574 691232
rect 30820 690155 30821 691231
rect 31573 690155 31574 691231
rect 30820 690154 31574 690155
rect 37358 689663 38120 689664
rect 37358 688581 37359 689663
rect 38119 688581 38120 689663
rect 37358 688580 38120 688581
rect 686012 674431 686766 674432
rect 686012 673355 686013 674431
rect 686765 673355 686766 674431
rect 686012 673354 686766 673355
rect 679466 672863 680228 672864
rect 679466 671781 679467 672863
rect 680227 671781 680228 672863
rect 679466 671780 680228 671781
rect 30820 648031 31574 648032
rect 30820 646955 30821 648031
rect 31573 646955 31574 648031
rect 30820 646954 31574 646955
rect 37358 646463 38120 646464
rect 37358 645381 37359 646463
rect 38119 645381 38120 646463
rect 37358 645380 38120 645381
rect 686012 629431 686766 629432
rect 686012 628355 686013 629431
rect 686765 628355 686766 629431
rect 686012 628354 686766 628355
rect 679466 627863 680228 627864
rect 679466 626781 679467 627863
rect 680227 626781 680228 627863
rect 679466 626780 680228 626781
rect 30820 604831 31574 604832
rect 30820 603755 30821 604831
rect 31573 603755 31574 604831
rect 30820 603754 31574 603755
rect 37358 603263 38120 603264
rect 37358 602181 37359 603263
rect 38119 602181 38120 603263
rect 37358 602180 38120 602181
rect 686012 584231 686766 584232
rect 686012 583155 686013 584231
rect 686765 583155 686766 584231
rect 686012 583154 686766 583155
rect 679466 582663 680228 582664
rect 679466 581581 679467 582663
rect 680227 581581 680228 582663
rect 679466 581580 680228 581581
rect 30820 561631 31574 561632
rect 30820 560555 30821 561631
rect 31573 560555 31574 561631
rect 30820 560554 31574 560555
rect 37358 560063 38120 560064
rect 37358 558981 37359 560063
rect 38119 558981 38120 560063
rect 37358 558980 38120 558981
rect 686012 539231 686766 539232
rect 686012 538155 686013 539231
rect 686765 538155 686766 539231
rect 686012 538154 686766 538155
rect 679466 537663 680228 537664
rect 679466 536581 679467 537663
rect 680227 536581 680228 537663
rect 679466 536580 680228 536581
rect 686012 495231 686766 495232
rect 686012 494155 686013 495231
rect 686765 494155 686766 495231
rect 686012 494154 686766 494155
rect 679466 493663 680228 493664
rect 679466 492581 679467 493663
rect 680227 492581 680228 493663
rect 679466 492580 680228 492581
rect 30820 434031 31574 434032
rect 30820 432955 30821 434031
rect 31573 432955 31574 434031
rect 30820 432954 31574 432955
rect 37358 432463 38120 432464
rect 37358 431381 37359 432463
rect 38119 431381 38120 432463
rect 37358 431380 38120 431381
rect 686012 407031 686766 407032
rect 686012 405955 686013 407031
rect 686765 405955 686766 407031
rect 686012 405954 686766 405955
rect 679466 405463 680228 405464
rect 679466 404381 679467 405463
rect 680227 404381 680228 405463
rect 679466 404380 680228 404381
rect 30820 390831 31574 390832
rect 30820 389755 30821 390831
rect 31573 389755 31574 390831
rect 30820 389754 31574 389755
rect 37358 389263 38120 389264
rect 37358 388181 37359 389263
rect 38119 388181 38120 389263
rect 37358 388180 38120 388181
rect 686012 361831 686766 361832
rect 686012 360755 686013 361831
rect 686765 360755 686766 361831
rect 686012 360754 686766 360755
rect 679466 360263 680228 360264
rect 679466 359181 679467 360263
rect 680227 359181 680228 360263
rect 679466 359180 680228 359181
rect 30820 347631 31574 347632
rect 30820 346555 30821 347631
rect 31573 346555 31574 347631
rect 30820 346554 31574 346555
rect 37358 346063 38120 346064
rect 37358 344981 37359 346063
rect 38119 344981 38120 346063
rect 37358 344980 38120 344981
rect 686012 316831 686766 316832
rect 686012 315755 686013 316831
rect 686765 315755 686766 316831
rect 686012 315754 686766 315755
rect 679466 315263 680228 315264
rect 679466 314181 679467 315263
rect 680227 314181 680228 315263
rect 679466 314180 680228 314181
rect 30820 304431 31574 304432
rect 30820 303355 30821 304431
rect 31573 303355 31574 304431
rect 30820 303354 31574 303355
rect 37358 302863 38120 302864
rect 37358 301781 37359 302863
rect 38119 301781 38120 302863
rect 37358 301780 38120 301781
rect 686012 271831 686766 271832
rect 686012 270755 686013 271831
rect 686765 270755 686766 271831
rect 686012 270754 686766 270755
rect 679466 270263 680228 270264
rect 679466 269181 679467 270263
rect 680227 269181 680228 270263
rect 679466 269180 680228 269181
rect 30820 261231 31574 261232
rect 30820 260155 30821 261231
rect 31573 260155 31574 261231
rect 30820 260154 31574 260155
rect 37358 259663 38120 259664
rect 37358 258581 37359 259663
rect 38119 258581 38120 259663
rect 37358 258580 38120 258581
rect 686012 226631 686766 226632
rect 686012 225555 686013 226631
rect 686765 225555 686766 226631
rect 686012 225554 686766 225555
rect 679466 225063 680228 225064
rect 679466 223981 679467 225063
rect 680227 223981 680228 225063
rect 679466 223980 680228 223981
rect 30820 218031 31574 218032
rect 30820 216955 30821 218031
rect 31573 216955 31574 218031
rect 30820 216954 31574 216955
rect 37358 216463 38120 216464
rect 37358 215381 37359 216463
rect 38119 215381 38120 216463
rect 37358 215380 38120 215381
rect 686012 181631 686766 181632
rect 686012 180555 686013 181631
rect 686765 180555 686766 181631
rect 686012 180554 686766 180555
rect 679466 180063 680228 180064
rect 679466 178981 679467 180063
rect 680227 178981 680228 180063
rect 679466 178980 680228 178981
rect 686012 136431 686766 136432
rect 686012 135355 686013 136431
rect 686765 135355 686766 136431
rect 686012 135354 686766 135355
rect 679466 134863 680228 134864
rect 679466 133781 679467 134863
rect 680227 133781 680228 134863
rect 679466 133780 680228 133781
rect 670566 32563 674216 32564
rect 670566 32055 670567 32563
rect 674215 32055 674216 32563
rect 670566 32054 674216 32055
<< metal3 >>
rect 575700 997056 580479 997678
rect 575700 995134 575788 997056
rect 580384 995134 580479 997056
rect 575700 995032 580479 995134
rect 585678 997062 590458 997678
rect 585678 995140 585758 997062
rect 590354 995140 590458 997062
rect 585678 995032 590458 995140
rect 39852 842324 50002 842458
rect 39852 837800 47908 842324
rect 49694 837800 50002 842324
rect 39852 837678 50002 837800
rect 667172 833206 677818 833301
rect 39852 832392 50002 832479
rect 39852 827868 47908 832392
rect 49694 827868 50002 832392
rect 667172 828630 667284 833206
rect 669732 828630 677818 833206
rect 667172 828521 677818 828630
rect 39852 827699 50002 827868
rect 667172 823212 677818 823322
rect 667172 818636 667270 823212
rect 669718 818636 677818 823212
rect 667172 818542 677818 818636
rect 667062 518582 677700 518701
rect 667062 514056 667336 518582
rect 669706 514056 677700 518582
rect 667062 513921 677700 514056
rect 667062 508592 677700 508722
rect 667062 504066 667350 508592
rect 669720 504066 677700 508592
rect 667062 503942 677700 504066
rect 39924 497732 52292 497858
rect 39924 493250 50364 497732
rect 52092 493250 52292 497732
rect 39924 493078 52292 493250
rect 39924 487742 52292 487879
rect 39924 483260 50352 487742
rect 52080 483260 52292 487742
rect 39924 483099 52292 483260
rect 663914 430390 677712 430501
rect 663914 425684 664134 430390
rect 666540 425748 677712 430390
rect 666540 425684 667110 425748
rect 663914 425562 667110 425684
rect 663914 420462 677712 420522
rect 663914 415856 664112 420462
rect 666528 415856 677712 420462
rect 663914 415742 677712 415856
rect 39934 124982 45766 125058
rect 39934 120338 42826 124982
rect 45696 120338 45766 124982
rect 39934 120278 45766 120338
rect 39934 115018 45766 115079
rect 39934 110374 42822 115018
rect 45692 110374 45766 115018
rect 39934 110299 45766 110374
rect 241690 45716 246049 45786
rect 241690 42842 241740 45716
rect 245986 42842 246049 45716
rect 241690 39426 246049 42842
rect 251300 45730 255702 45786
rect 251300 42856 251392 45730
rect 255638 42856 255702 45730
rect 251300 39426 255702 42856
rect 622942 45708 627722 45818
rect 622942 42878 623000 45708
rect 627626 42878 627722 45708
rect 622942 39838 627722 42878
rect 632921 45698 637701 45818
rect 632921 42868 633000 45698
rect 637626 42868 637701 45698
rect 632921 39838 637701 42868
rect 670476 32564 674286 41774
rect 670476 32054 670566 32564
rect 674216 32054 674286 32564
rect 670476 31974 674286 32054
<< via3 >>
rect 575788 995134 580384 997056
rect 585758 995140 590354 997062
rect 47908 837800 49694 842324
rect 47908 827868 49694 832392
rect 667284 828630 669732 833206
rect 667270 818636 669718 823212
rect 667336 514056 669706 518582
rect 667350 504066 669720 508592
rect 50364 493250 52092 497732
rect 50352 483260 52080 487742
rect 664134 425684 666540 430390
rect 664112 415856 666528 420462
rect 42826 120338 45696 124982
rect 42822 110374 45692 115018
rect 241740 42842 245986 45716
rect 251392 42856 255638 45730
rect 623000 42878 627626 45708
rect 633000 42868 637626 45698
rect 670566 32054 674216 32564
<< metal4 >>
rect 575680 997056 580478 997130
rect 575680 995134 575788 997056
rect 580384 995134 580478 997056
rect 575680 993314 580478 995134
rect 575680 990884 575762 993314
rect 580384 990884 580478 993314
rect 575680 990788 580478 990884
rect 585670 997062 590468 997144
rect 585670 995140 585758 997062
rect 590354 995140 590468 997062
rect 585670 993328 590468 995140
rect 585670 990898 585758 993328
rect 590380 990898 590468 993328
rect 585670 990802 590468 990898
rect 47792 842324 49822 842462
rect 47792 837800 47908 842324
rect 49694 837800 49822 842324
rect 47792 837658 49822 837800
rect 667202 833206 669802 833310
rect 47792 832392 49822 832506
rect 47792 827868 47908 832392
rect 49694 827868 49822 832392
rect 667202 828630 667284 833206
rect 669732 828630 669802 833206
rect 667202 828520 669802 828630
rect 47792 827702 49822 827868
rect 667214 823212 669814 823336
rect 667214 818636 667270 823212
rect 669718 818636 669814 823212
rect 667214 818546 669814 818636
rect 667206 518582 669814 518696
rect 667206 514056 667336 518582
rect 669706 514056 669814 518582
rect 667206 513920 669814 514056
rect 667218 508592 669826 508726
rect 667218 504066 667350 508592
rect 669720 504066 669826 508592
rect 667218 503950 669826 504066
rect 50172 497732 52196 497874
rect 50172 493250 50364 497732
rect 52092 493250 52196 497732
rect 50172 493084 52196 493250
rect 50198 487742 52222 487884
rect 50198 483260 50352 487742
rect 52080 483260 52222 487742
rect 50198 483094 52222 483260
rect 664008 430390 666612 430490
rect 664008 425684 664134 430390
rect 666540 425684 666612 430390
rect 664008 425572 666612 425684
rect 664018 420462 666634 420524
rect 664018 415856 664112 420462
rect 666528 415856 666634 420462
rect 664018 415760 666634 415856
rect 42764 124982 45774 125050
rect 42764 120338 42826 124982
rect 45696 120338 45774 124982
rect 42764 120264 45774 120338
rect 42762 115018 45772 115082
rect 42762 110374 42822 115018
rect 45692 110374 45772 115018
rect 42762 110296 45772 110374
rect 241680 45716 246056 45792
rect 241680 42842 241740 45716
rect 245986 42842 246056 45716
rect 241680 42784 246056 42842
rect 251302 45730 255700 45784
rect 251302 42856 251392 45730
rect 255638 42856 255700 45730
rect 251302 42788 255700 42856
rect 622940 45708 627718 45784
rect 622940 42878 623000 45708
rect 627626 42878 627718 45708
rect 622940 42780 627718 42878
rect 632920 45698 637698 45790
rect 632920 42868 633000 45698
rect 637626 42868 637698 45698
rect 632920 42786 637698 42868
<< via4 >>
rect 575762 990884 580384 993314
rect 585758 990898 590380 993328
rect 47908 837800 49694 842324
rect 47908 827868 49694 832392
rect 667284 828630 669732 833206
rect 667270 818636 669718 823212
rect 667336 514056 669706 518582
rect 667350 504066 669720 508592
rect 50364 493250 52092 497732
rect 50352 483260 52080 487742
rect 664134 425684 666540 430390
rect 664112 415856 666528 420462
rect 42826 120338 45696 124982
rect 42822 110374 45692 115018
rect 241740 42842 245986 45716
rect 251392 42856 255638 45730
rect 623000 42878 627626 45708
rect 633000 42868 637626 45698
<< metal5 >>
rect 52598 995502 676620 996702
rect 47798 842324 49798 992152
rect 47798 837800 47908 842324
rect 49694 837800 49798 842324
rect 47798 832392 49798 837800
rect 47798 827868 47908 832392
rect 49694 827868 49798 832392
rect 47798 243300 49798 827868
rect 50198 497732 52198 992152
rect 50198 493250 50364 497732
rect 52092 493250 52198 497732
rect 50198 487742 52198 493250
rect 50198 483260 50352 487742
rect 52080 483260 52198 487742
rect 50198 243300 52198 483260
rect 42768 124982 45768 176144
rect 42768 120338 42826 124982
rect 45696 120338 45768 124982
rect 42768 115018 45768 120338
rect 42768 110374 42822 115018
rect 45692 110374 45768 115018
rect 42768 42872 45768 110374
rect 47836 45444 50836 240850
rect 52598 217742 53798 995502
rect 54198 993902 673420 995102
rect 54198 219342 55398 993902
rect 575640 993328 666620 993396
rect 575640 993314 585758 993328
rect 575640 990884 575762 993314
rect 580384 990898 585758 993314
rect 590380 990898 666620 993328
rect 670820 992696 673420 993902
rect 674020 992696 676620 995502
rect 580384 990884 666620 990898
rect 575640 990796 666620 990884
rect 664020 430390 666620 990796
rect 664020 425684 664134 430390
rect 666540 425684 666620 430390
rect 664020 420462 666620 425684
rect 664020 415856 664112 420462
rect 666528 415856 666620 420462
rect 59154 260466 189024 263466
rect 417154 260466 657074 263466
rect 59154 256466 189024 259466
rect 417154 256466 657074 259466
rect 59154 252466 189024 255466
rect 417154 252466 657074 255466
rect 59154 248466 189024 251466
rect 417154 248466 657074 251466
rect 59154 244466 189024 247466
rect 417154 244466 657074 247466
rect 59154 240466 189024 243466
rect 417154 240466 657074 243466
rect 59154 236466 189024 239466
rect 417154 236466 657074 239466
rect 59154 232466 189024 235466
rect 417154 232466 657074 235466
rect 598374 51222 601374 228738
rect 162222 48222 601374 51222
rect 602390 48502 605390 228790
rect 664020 215484 666620 415856
rect 667220 833206 669820 992690
rect 667220 828630 667284 833206
rect 669732 828630 669820 833206
rect 667220 823212 669820 828630
rect 667220 818636 667270 823212
rect 669718 818636 669820 823212
rect 667220 518582 669820 818636
rect 667220 514056 667336 518582
rect 669706 514056 669820 518582
rect 667220 508592 669820 514056
rect 667220 504066 667350 508592
rect 669720 504066 669820 508592
rect 667220 215428 669820 504066
rect 162222 45444 165222 48222
rect 47836 42444 165222 45444
rect 241654 45730 613240 45788
rect 241654 45716 251392 45730
rect 241654 42842 241740 45716
rect 245986 42856 251392 45716
rect 255638 42856 613240 45730
rect 245986 42842 613240 42856
rect 241654 42788 613240 42842
rect 622918 45708 644430 45788
rect 622918 42878 623000 45708
rect 627626 45698 644430 45708
rect 627626 42878 633000 45698
rect 622918 42868 633000 42878
rect 637626 42868 644430 45698
rect 666426 43548 669426 211904
rect 622918 42788 644430 42868
<< comment >>
rect 0 1037400 717600 1037600
rect 0 200 200 1037400
rect 717400 200 717600 1037400
rect 0 0 717600 200
use gpio_control_power_routing  gpio_control_power_routing_0
timestamp 1637447660
transform 1 0 -10 0 1 0
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_1
timestamp 1637447660
transform 1 0 -10 0 1 43200
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_14
timestamp 1637447660
transform -1 0 717846 0 1 -81600
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_13
timestamp 1637447660
transform -1 0 717846 0 1 -36400
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_12
timestamp 1637447660
transform -1 0 717846 0 1 8600
box 6032 203748 46270 221470
use gpio_control_power_routing  gpio_control_power_routing_2
timestamp 1637447660
transform 1 0 -10 0 1 86400
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_3
timestamp 1637447660
transform 1 0 -10 0 1 129600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_4
timestamp 1637447660
transform 1 0 -10 0 1 172800
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_11
timestamp 1637447660
transform -1 0 717846 0 1 53800
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_10
timestamp 1637447660
transform -1 0 717846 0 1 98800
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_9
timestamp 1637447660
transform -1 0 717846 0 1 143800
box 6032 203748 46270 221470
use gpio_control_power_routing  gpio_control_power_routing_5
timestamp 1637447660
transform 1 0 -10 0 1 216000
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_8
timestamp 1637447660
transform -1 0 717846 0 1 189000
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_7
timestamp 1637447660
transform -1 0 717846 0 1 277200
box 6032 203748 46270 221470
use gpio_control_power_routing  gpio_control_power_routing_6
timestamp 1637447660
transform 1 0 -10 0 1 343600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_7
timestamp 1637447660
transform 1 0 -10 0 1 386800
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_8
timestamp 1637447660
transform 1 0 -10 0 1 430000
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_6
timestamp 1637447660
transform -1 0 717846 0 1 321200
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_5
timestamp 1637447660
transform -1 0 717846 0 1 366200
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_4
timestamp 1637447660
transform -1 0 717846 0 1 411400
box 6032 203748 46270 221470
use gpio_control_power_routing  gpio_control_power_routing_9
timestamp 1637447660
transform 1 0 -10 0 1 473200
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_11
timestamp 1637447660
transform 1 0 -10 0 1 559600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_10
timestamp 1637447660
transform 1 0 -10 0 1 516400
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_3
timestamp 1637447660
transform -1 0 717846 0 1 456400
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_2
timestamp 1637447660
transform -1 0 717846 0 1 501600
box 6032 203748 46270 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_1
timestamp 1637447660
transform -1 0 717846 0 1 546600
box 6032 203748 46270 221470
use gpio_control_power_routing  gpio_control_power_routing_12
timestamp 1637447660
transform 1 0 -10 0 1 602800
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_13
timestamp 1637447660
transform 1 0 -10 0 1 728600
box 6032 203748 55470 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_0
timestamp 1637447660
transform 0 1 -105400 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_1
timestamp 1637447660
transform 0 1 -54000 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_3
timestamp 1637447660
transform 0 1 48800 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_2
timestamp 1637447660
transform 0 1 -2600 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_4
timestamp 1637447660
transform 0 1 100400 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_5
timestamp 1637447660
transform 0 1 150800 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_6
timestamp 1637447660
transform 0 1 218200 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_7
timestamp 1637447660
transform 0 1 295200 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_8
timestamp 1637447660
transform 0 1 346600 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_0
timestamp 1637447660
transform -1 0 717836 0 1 725000
box 6032 203748 46270 221470
<< labels >>
flabel metal5 54316 219436 55324 219998 0 FreeSans 1600 0 0 0 vccd1
flabel metal5 52692 217826 53700 218388 0 FreeSans 1600 0 0 0 vssd1
flabel metal5 664092 215580 666518 216304 0 FreeSans 3200 0 0 0 vssa1
flabel metal5 667280 215542 669706 216266 0 FreeSans 3200 0 0 0 vdda1
flabel metal5 47904 243444 49660 243998 0 FreeSans 3200 0 0 0 vssa2
flabel metal5 50338 243444 52094 243998 0 FreeSans 3200 0 0 0 vdda2
<< end >>
