VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO empty_macro_1
  CLASS BLOCK ;
  FOREIGN empty_macro_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 120.000 BY 200.000 ;
END empty_macro_1
END LIBRARY