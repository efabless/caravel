magic
tech sky130A
magscale 1 2
timestamp 1638030917
<< checkpaint >>
rect -194 -220 7278 7292
<< nwell >>
rect 2304 2369 2397 2389
<< viali >>
rect 4353 5117 4387 5151
rect 5273 5117 5307 5151
rect 2145 4641 2179 4675
rect 3249 4641 3283 4675
rect 3617 4641 3651 4675
rect 4721 4641 4755 4675
rect 1593 4029 1627 4063
rect 2053 4029 2087 4063
rect 4445 4029 4479 4063
rect 4721 4029 4755 4063
rect 5549 4029 5583 4063
rect 1685 3553 1719 3587
rect 1961 3553 1995 3587
rect 2697 3553 2731 3587
rect 3157 3553 3191 3587
rect 3433 3553 3467 3587
rect 4261 3553 4295 3587
rect 4813 3553 4847 3587
rect 5273 3553 5307 3587
rect 1593 2941 1627 2975
rect 4813 2397 4847 2431
rect 5089 2397 5123 2431
rect 1593 1853 1627 1887
rect 2145 1853 2179 1887
rect 2605 1853 2639 1887
rect 2881 1853 2915 1887
rect 3249 1853 3283 1887
rect 4077 1853 4111 1887
rect 5641 1853 5675 1887
rect 1685 1377 1719 1411
rect 2973 1377 3007 1411
rect 4629 1377 4663 1411
<< metal1 >>
rect 1104 6010 5980 6032
rect 1104 5958 2607 6010
rect 2659 5958 2671 6010
rect 2723 5958 2735 6010
rect 2787 5958 2799 6010
rect 2851 5958 4232 6010
rect 4284 5958 4296 6010
rect 4348 5958 4360 6010
rect 4412 5958 4424 6010
rect 4476 5958 5980 6010
rect 1104 5936 5980 5958
rect 1104 5466 5980 5488
rect 1104 5414 1794 5466
rect 1846 5414 1858 5466
rect 1910 5414 1922 5466
rect 1974 5414 1986 5466
rect 2038 5414 3420 5466
rect 3472 5414 3484 5466
rect 3536 5414 3548 5466
rect 3600 5414 3612 5466
rect 3664 5414 5045 5466
rect 5097 5414 5109 5466
rect 5161 5414 5173 5466
rect 5225 5414 5237 5466
rect 5289 5414 5980 5466
rect 1104 5392 5980 5414
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 4157 5148 4215 5157
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 4120 5120 4353 5148
rect 4120 5108 4126 5120
rect 4157 5111 4215 5120
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 4614 5108 4620 5160
rect 4672 5148 4678 5160
rect 5077 5148 5135 5157
rect 5261 5151 5319 5157
rect 5261 5148 5273 5151
rect 4672 5120 5273 5148
rect 4672 5108 4678 5120
rect 5077 5111 5135 5120
rect 5261 5117 5273 5120
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 1104 4922 5980 4944
rect 1104 4870 2607 4922
rect 2659 4870 2671 4922
rect 2723 4870 2735 4922
rect 2787 4870 2799 4922
rect 2851 4870 4232 4922
rect 4284 4870 4296 4922
rect 4348 4870 4360 4922
rect 4412 4870 4424 4922
rect 4476 4870 5980 4922
rect 1104 4848 5980 4870
rect 1949 4672 2007 4681
rect 2133 4675 2191 4681
rect 2133 4672 2145 4675
rect 1949 4644 2145 4672
rect 1949 4635 2007 4644
rect 2133 4641 2145 4644
rect 2179 4672 2191 4675
rect 2958 4672 2964 4684
rect 2179 4644 2964 4672
rect 2179 4641 2191 4644
rect 2133 4635 2191 4641
rect 2958 4632 2964 4644
rect 3016 4632 3022 4684
rect 3050 4672 3114 4684
rect 3234 4672 3240 4684
rect 3050 4644 3240 4672
rect 3050 4632 3114 4644
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 3418 4672 3482 4684
rect 3602 4675 3666 4684
rect 3602 4672 3617 4675
rect 3418 4644 3617 4672
rect 3418 4632 3482 4644
rect 3602 4641 3617 4644
rect 3651 4641 3666 4675
rect 3602 4632 3666 4641
rect 4522 4674 4586 4684
rect 4706 4675 4770 4684
rect 4706 4674 4721 4675
rect 4522 4644 4721 4674
rect 4522 4632 4586 4644
rect 4706 4641 4721 4644
rect 4755 4641 4770 4675
rect 4706 4632 4770 4641
rect 3620 4468 3648 4632
rect 4720 4539 4755 4632
rect 4720 4505 4754 4539
rect 4720 4480 4755 4505
rect 3878 4468 3884 4480
rect 3620 4440 3884 4468
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 4706 4428 4712 4480
rect 4764 4428 4770 4480
rect 1104 4378 5980 4400
rect 1104 4326 1794 4378
rect 1846 4326 1858 4378
rect 1910 4326 1922 4378
rect 1974 4326 1986 4378
rect 2038 4326 3420 4378
rect 3472 4326 3484 4378
rect 3536 4326 3548 4378
rect 3600 4326 3612 4378
rect 3664 4326 5045 4378
rect 5097 4326 5109 4378
rect 5161 4326 5173 4378
rect 5225 4326 5237 4378
rect 5289 4326 5980 4378
rect 1104 4304 5980 4326
rect 3050 4224 3056 4276
rect 3108 4264 3114 4276
rect 3108 4236 4568 4264
rect 3108 4224 3114 4236
rect 1394 4156 1400 4208
rect 1452 4196 1458 4208
rect 1452 4168 1902 4196
rect 1452 4156 1458 4168
rect 1394 4060 1458 4072
rect 1578 4060 1584 4072
rect 1394 4032 1584 4060
rect 1394 4020 1458 4032
rect 1578 4020 1584 4032
rect 1636 4020 1642 4072
rect 1870 4069 1902 4168
rect 2222 4088 2228 4140
rect 2280 4128 2286 4140
rect 2280 4100 3924 4128
rect 2280 4088 2286 4100
rect 1857 4059 1915 4069
rect 2041 4063 2099 4069
rect 2041 4059 2053 4063
rect 1857 4031 2053 4059
rect 1857 4023 1915 4031
rect 2041 4029 2053 4031
rect 2087 4029 2099 4063
rect 2041 4023 2099 4029
rect 3896 3992 3924 4100
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 4540 4069 4568 4236
rect 4249 4060 4307 4069
rect 4433 4063 4491 4069
rect 4433 4060 4445 4063
rect 4120 4032 4445 4060
rect 4120 4020 4126 4032
rect 4249 4023 4307 4032
rect 4433 4029 4445 4032
rect 4479 4029 4491 4063
rect 4433 4023 4491 4029
rect 4525 4060 4583 4069
rect 4709 4063 4767 4069
rect 4709 4060 4721 4063
rect 4525 4032 4721 4060
rect 4525 4023 4583 4032
rect 4709 4029 4721 4032
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 5350 4020 5356 4072
rect 5408 4060 5414 4072
rect 5537 4063 5595 4069
rect 5537 4060 5549 4063
rect 5408 4031 5549 4060
rect 5408 4020 5414 4031
rect 5537 4029 5549 4031
rect 5583 4029 5595 4063
rect 5537 4023 5595 4029
rect 4890 3992 4896 4004
rect 3896 3964 4896 3992
rect 4890 3952 4896 3964
rect 4948 3952 4954 4004
rect 1104 3834 5980 3856
rect 1104 3782 2607 3834
rect 2659 3782 2671 3834
rect 2723 3782 2735 3834
rect 2787 3782 2799 3834
rect 2851 3782 4232 3834
rect 4284 3782 4296 3834
rect 4348 3782 4360 3834
rect 4412 3782 4424 3834
rect 4476 3782 5980 3834
rect 1104 3760 5980 3782
rect 566 3680 572 3732
rect 624 3720 630 3732
rect 4706 3720 4712 3732
rect 624 3692 4712 3720
rect 624 3680 630 3692
rect 4706 3680 4712 3692
rect 4764 3680 4770 3732
rect 5902 3652 5908 3664
rect 1964 3624 5908 3652
rect 1486 3584 1550 3596
rect 1670 3584 1676 3596
rect 1486 3556 1676 3584
rect 1486 3544 1550 3556
rect 1670 3544 1676 3556
rect 1728 3544 1734 3596
rect 1964 3593 1992 3624
rect 5902 3612 5908 3624
rect 5960 3612 5966 3664
rect 1765 3584 1823 3593
rect 1949 3587 2007 3593
rect 1949 3584 1961 3587
rect 1765 3556 1961 3584
rect 1765 3547 1823 3556
rect 1949 3553 1961 3556
rect 1995 3553 2007 3587
rect 1949 3547 2007 3553
rect 2501 3586 2559 3593
rect 2685 3587 2743 3593
rect 2685 3586 2697 3587
rect 2501 3555 2697 3586
rect 2501 3547 2559 3555
rect 2685 3553 2697 3555
rect 2731 3586 2743 3587
rect 2774 3586 2780 3596
rect 2731 3555 2780 3586
rect 2731 3553 2743 3555
rect 2685 3547 2743 3553
rect 2774 3544 2780 3555
rect 2832 3544 2838 3596
rect 2958 3584 3022 3596
rect 3142 3584 3148 3596
rect 2958 3556 3148 3584
rect 2958 3544 3022 3556
rect 3142 3544 3148 3556
rect 3200 3544 3206 3596
rect 3234 3585 3298 3596
rect 3418 3587 3482 3596
rect 3418 3585 3433 3587
rect 3234 3557 3433 3585
rect 3234 3544 3298 3557
rect 3418 3553 3433 3557
rect 3467 3553 3482 3587
rect 3418 3544 3482 3553
rect 4065 3584 4123 3593
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 4065 3556 4261 3584
rect 4065 3547 4123 3556
rect 4249 3553 4261 3556
rect 4295 3584 4307 3587
rect 4522 3584 4528 3596
rect 4295 3556 4528 3584
rect 4295 3553 4307 3556
rect 4249 3547 4307 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 4614 3585 4678 3596
rect 4798 3587 4862 3596
rect 4798 3585 4813 3587
rect 4614 3557 4813 3585
rect 4614 3544 4678 3557
rect 4798 3553 4813 3557
rect 4847 3553 4862 3587
rect 4798 3544 4862 3553
rect 4982 3544 4988 3596
rect 5040 3584 5046 3596
rect 5077 3584 5135 3593
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 5040 3556 5273 3584
rect 5040 3544 5046 3556
rect 5077 3547 5135 3556
rect 5261 3553 5273 3556
rect 5307 3553 5319 3587
rect 5261 3547 5319 3553
rect 2222 3408 2228 3460
rect 2280 3448 2286 3460
rect 3438 3448 3466 3544
rect 4706 3448 4712 3460
rect 2280 3420 3280 3448
rect 3438 3420 4712 3448
rect 2280 3408 2286 3420
rect 3252 3380 3280 3420
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 4814 3380 4842 3544
rect 3252 3352 4842 3380
rect 1104 3290 2150 3312
rect 1104 3238 1794 3290
rect 1846 3238 1858 3290
rect 1910 3238 1922 3290
rect 1974 3238 1986 3290
rect 2038 3238 2150 3290
rect 1104 3216 2150 3238
rect 2181 3290 5902 3312
rect 2181 3238 3420 3290
rect 3472 3238 3484 3290
rect 3536 3238 3548 3290
rect 3600 3238 3612 3290
rect 3664 3238 5045 3290
rect 5097 3238 5109 3290
rect 5161 3238 5173 3290
rect 5225 3238 5237 3290
rect 5289 3238 5902 3290
rect 2181 3216 5902 3238
rect 5966 3216 5980 3312
rect 2773 3131 2779 3183
rect 2831 3174 2837 3183
rect 5902 3174 5908 3188
rect 2831 3143 5908 3174
rect 2831 3131 2837 3143
rect 5902 3136 5908 3143
rect 5960 3136 5966 3188
rect 1397 2972 1455 2981
rect 1581 2975 1639 2981
rect 1581 2972 1593 2975
rect 1397 2944 1593 2972
rect 1397 2935 1455 2944
rect 1581 2941 1593 2944
rect 1627 2972 1639 2975
rect 3050 2972 3056 2984
rect 1627 2944 3056 2972
rect 1627 2941 1639 2944
rect 1581 2935 1639 2941
rect 3050 2932 3056 2944
rect 3108 2932 3114 2984
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 4614 2836 4620 2848
rect 1728 2808 4620 2836
rect 1728 2796 1734 2808
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 1104 2746 5980 2768
rect 1104 2694 2607 2746
rect 2659 2694 2671 2746
rect 2723 2694 2735 2746
rect 2787 2694 2799 2746
rect 2851 2694 4232 2746
rect 4284 2694 4296 2746
rect 4348 2694 4360 2746
rect 4412 2694 4424 2746
rect 4476 2694 5980 2746
rect 1104 2672 5980 2694
rect 5442 2496 5448 2508
rect 4815 2468 5448 2496
rect 4815 2437 4843 2468
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 4617 2429 4675 2437
rect 4801 2431 4859 2437
rect 4801 2429 4813 2431
rect 4617 2401 4813 2429
rect 4617 2391 4675 2401
rect 4801 2397 4813 2401
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 4890 2388 4896 2440
rect 4948 2428 4954 2440
rect 5077 2431 5135 2437
rect 5077 2428 5089 2431
rect 4948 2400 5089 2428
rect 4948 2388 4954 2400
rect 5077 2397 5089 2400
rect 5123 2397 5135 2431
rect 5077 2391 5135 2397
rect 2314 2320 2320 2372
rect 2372 2360 2378 2372
rect 6454 2360 6460 2372
rect 2372 2332 6460 2360
rect 2372 2320 2378 2332
rect 6454 2320 6460 2332
rect 6512 2320 6518 2372
rect 1104 2202 5980 2224
rect 1104 2150 1794 2202
rect 1846 2150 1858 2202
rect 1910 2150 1922 2202
rect 1974 2150 1986 2202
rect 2038 2150 3420 2202
rect 3472 2150 3484 2202
rect 3536 2150 3548 2202
rect 3600 2150 3612 2202
rect 3664 2150 5045 2202
rect 5097 2150 5109 2202
rect 5161 2150 5173 2202
rect 5225 2150 5237 2202
rect 5289 2150 5980 2202
rect 1104 2128 5980 2150
rect 3970 2020 3976 2032
rect 2976 1992 3976 2020
rect 1210 1912 1216 1964
rect 1268 1952 1274 1964
rect 1268 1924 2452 1952
rect 1268 1912 1274 1924
rect 1397 1884 1455 1893
rect 1581 1887 1639 1893
rect 1581 1884 1593 1887
rect 1397 1856 1593 1884
rect 1397 1847 1455 1856
rect 1581 1853 1593 1856
rect 1627 1853 1639 1887
rect 1581 1847 1639 1853
rect 1949 1884 2007 1893
rect 2133 1887 2191 1893
rect 2133 1884 2145 1887
rect 1949 1856 2145 1884
rect 1949 1847 2007 1856
rect 2133 1853 2145 1856
rect 2179 1884 2191 1887
rect 2314 1884 2320 1896
rect 2179 1856 2320 1884
rect 2179 1853 2191 1856
rect 2133 1847 2191 1853
rect 1596 1816 1624 1847
rect 2314 1844 2320 1856
rect 2372 1844 2378 1896
rect 2424 1893 2452 1924
rect 2409 1884 2467 1893
rect 2593 1887 2651 1893
rect 2593 1884 2605 1887
rect 2409 1856 2605 1884
rect 2409 1847 2467 1856
rect 2593 1853 2605 1856
rect 2639 1853 2651 1887
rect 2593 1847 2651 1853
rect 2685 1884 2743 1893
rect 2869 1887 2927 1893
rect 2869 1884 2881 1887
rect 2685 1856 2881 1884
rect 2685 1847 2743 1856
rect 2869 1853 2881 1856
rect 2915 1884 2927 1887
rect 2976 1884 3004 1992
rect 3970 1980 3976 1992
rect 4028 1980 4034 2032
rect 2915 1856 3004 1884
rect 3050 1884 3114 1896
rect 3234 1884 3240 1896
rect 3050 1856 3240 1884
rect 2915 1853 2927 1856
rect 2869 1847 2927 1853
rect 3050 1844 3114 1856
rect 3234 1844 3240 1856
rect 3292 1844 3298 1896
rect 3786 1844 3792 1896
rect 3844 1884 3850 1896
rect 3881 1884 3939 1893
rect 4065 1887 4123 1893
rect 4065 1884 4077 1887
rect 3844 1856 4077 1884
rect 3844 1844 3850 1856
rect 3881 1847 3939 1856
rect 4065 1853 4077 1856
rect 4111 1853 4123 1887
rect 4065 1847 4123 1853
rect 5442 1884 5506 1896
rect 5626 1884 5632 1896
rect 5442 1856 5632 1884
rect 5442 1844 5506 1856
rect 5626 1844 5632 1856
rect 5684 1844 5690 1896
rect 1596 1788 3004 1816
rect 2976 1748 3004 1788
rect 3234 1748 3240 1760
rect 2976 1720 3240 1748
rect 3234 1708 3240 1720
rect 3292 1708 3298 1760
rect 1104 1658 5980 1680
rect 1104 1606 2607 1658
rect 2659 1606 2671 1658
rect 2723 1606 2735 1658
rect 2787 1606 2799 1658
rect 2851 1606 4232 1658
rect 4284 1606 4296 1658
rect 4348 1606 4360 1658
rect 4412 1606 4424 1658
rect 4476 1606 5980 1658
rect 1104 1584 5980 1606
rect 1118 1368 1124 1420
rect 1176 1408 1182 1420
rect 1489 1408 1547 1417
rect 1673 1411 1731 1417
rect 1673 1408 1685 1411
rect 1176 1380 1685 1408
rect 1176 1368 1182 1380
rect 1489 1371 1547 1380
rect 1673 1377 1685 1380
rect 1719 1377 1731 1411
rect 1673 1371 1731 1377
rect 2774 1408 2838 1420
rect 2958 1408 2964 1420
rect 2774 1380 2964 1408
rect 2774 1368 2838 1380
rect 2958 1368 2964 1380
rect 3016 1368 3022 1420
rect 4430 1408 4494 1420
rect 4614 1408 4620 1420
rect 4430 1380 4620 1408
rect 4430 1368 4494 1380
rect 4614 1368 4620 1380
rect 4672 1368 4678 1420
rect 1104 1114 5980 1136
rect 1104 1062 1794 1114
rect 1846 1062 1858 1114
rect 1910 1062 1922 1114
rect 1974 1062 1986 1114
rect 2038 1062 3420 1114
rect 3472 1062 3484 1114
rect 3536 1062 3548 1114
rect 3600 1062 3612 1114
rect 3664 1062 5045 1114
rect 5097 1062 5109 1114
rect 5161 1062 5173 1114
rect 5225 1062 5237 1114
rect 5289 1062 5980 1114
rect 1104 1040 5980 1062
<< via1 >>
rect 2607 5958 2659 6010
rect 2671 5958 2723 6010
rect 2735 5958 2787 6010
rect 2799 5958 2851 6010
rect 4232 5958 4284 6010
rect 4296 5958 4348 6010
rect 4360 5958 4412 6010
rect 4424 5958 4476 6010
rect 1794 5414 1846 5466
rect 1858 5414 1910 5466
rect 1922 5414 1974 5466
rect 1986 5414 2038 5466
rect 3420 5414 3472 5466
rect 3484 5414 3536 5466
rect 3548 5414 3600 5466
rect 3612 5414 3664 5466
rect 5045 5414 5097 5466
rect 5109 5414 5161 5466
rect 5173 5414 5225 5466
rect 5237 5414 5289 5466
rect 4068 5108 4120 5160
rect 4620 5108 4672 5160
rect 2607 4870 2659 4922
rect 2671 4870 2723 4922
rect 2735 4870 2787 4922
rect 2799 4870 2851 4922
rect 4232 4870 4284 4922
rect 4296 4870 4348 4922
rect 4360 4870 4412 4922
rect 4424 4870 4476 4922
rect 2964 4632 3016 4684
rect 3240 4675 3292 4684
rect 3240 4641 3249 4675
rect 3249 4641 3283 4675
rect 3283 4641 3292 4675
rect 3240 4632 3292 4641
rect 3884 4428 3936 4480
rect 4712 4428 4764 4480
rect 1794 4326 1846 4378
rect 1858 4326 1910 4378
rect 1922 4326 1974 4378
rect 1986 4326 2038 4378
rect 3420 4326 3472 4378
rect 3484 4326 3536 4378
rect 3548 4326 3600 4378
rect 3612 4326 3664 4378
rect 5045 4326 5097 4378
rect 5109 4326 5161 4378
rect 5173 4326 5225 4378
rect 5237 4326 5289 4378
rect 3056 4224 3108 4276
rect 1400 4156 1452 4208
rect 1584 4063 1636 4072
rect 1584 4029 1593 4063
rect 1593 4029 1627 4063
rect 1627 4029 1636 4063
rect 1584 4020 1636 4029
rect 2228 4088 2280 4140
rect 4068 4020 4120 4072
rect 5356 4020 5408 4072
rect 4896 3952 4948 4004
rect 2607 3782 2659 3834
rect 2671 3782 2723 3834
rect 2735 3782 2787 3834
rect 2799 3782 2851 3834
rect 4232 3782 4284 3834
rect 4296 3782 4348 3834
rect 4360 3782 4412 3834
rect 4424 3782 4476 3834
rect 572 3680 624 3732
rect 4712 3680 4764 3732
rect 1676 3587 1728 3596
rect 1676 3553 1685 3587
rect 1685 3553 1719 3587
rect 1719 3553 1728 3587
rect 1676 3544 1728 3553
rect 5908 3612 5960 3664
rect 2780 3544 2832 3596
rect 3148 3587 3200 3596
rect 3148 3553 3157 3587
rect 3157 3553 3191 3587
rect 3191 3553 3200 3587
rect 3148 3544 3200 3553
rect 4528 3544 4580 3596
rect 4988 3544 5040 3596
rect 2228 3408 2280 3460
rect 4712 3408 4764 3460
rect 1794 3238 1846 3290
rect 1858 3238 1910 3290
rect 1922 3238 1974 3290
rect 1986 3238 2038 3290
rect 3420 3238 3472 3290
rect 3484 3238 3536 3290
rect 3548 3238 3600 3290
rect 3612 3238 3664 3290
rect 5045 3238 5097 3290
rect 5109 3238 5161 3290
rect 5173 3238 5225 3290
rect 5237 3238 5289 3290
rect 2779 3131 2831 3183
rect 5908 3136 5960 3188
rect 3056 2932 3108 2984
rect 1676 2796 1728 2848
rect 4620 2796 4672 2848
rect 2607 2694 2659 2746
rect 2671 2694 2723 2746
rect 2735 2694 2787 2746
rect 2799 2694 2851 2746
rect 4232 2694 4284 2746
rect 4296 2694 4348 2746
rect 4360 2694 4412 2746
rect 4424 2694 4476 2746
rect 5448 2456 5500 2508
rect 4896 2388 4948 2440
rect 2320 2320 2372 2372
rect 6460 2320 6512 2372
rect 1794 2150 1846 2202
rect 1858 2150 1910 2202
rect 1922 2150 1974 2202
rect 1986 2150 2038 2202
rect 3420 2150 3472 2202
rect 3484 2150 3536 2202
rect 3548 2150 3600 2202
rect 3612 2150 3664 2202
rect 5045 2150 5097 2202
rect 5109 2150 5161 2202
rect 5173 2150 5225 2202
rect 5237 2150 5289 2202
rect 1216 1912 1268 1964
rect 2320 1844 2372 1896
rect 3976 1980 4028 2032
rect 3240 1887 3292 1896
rect 3240 1853 3249 1887
rect 3249 1853 3283 1887
rect 3283 1853 3292 1887
rect 3240 1844 3292 1853
rect 3792 1844 3844 1896
rect 5632 1887 5684 1896
rect 5632 1853 5641 1887
rect 5641 1853 5675 1887
rect 5675 1853 5684 1887
rect 5632 1844 5684 1853
rect 3240 1708 3292 1760
rect 2607 1606 2659 1658
rect 2671 1606 2723 1658
rect 2735 1606 2787 1658
rect 2799 1606 2851 1658
rect 4232 1606 4284 1658
rect 4296 1606 4348 1658
rect 4360 1606 4412 1658
rect 4424 1606 4476 1658
rect 1124 1368 1176 1420
rect 2964 1411 3016 1420
rect 2964 1377 2973 1411
rect 2973 1377 3007 1411
rect 3007 1377 3016 1411
rect 2964 1368 3016 1377
rect 4620 1411 4672 1420
rect 4620 1377 4629 1411
rect 4629 1377 4663 1411
rect 4663 1377 4672 1411
rect 4620 1368 4672 1377
rect 1794 1062 1846 1114
rect 1858 1062 1910 1114
rect 1922 1062 1974 1114
rect 1986 1062 2038 1114
rect 3420 1062 3472 1114
rect 3484 1062 3536 1114
rect 3548 1062 3600 1114
rect 3612 1062 3664 1114
rect 5045 1062 5097 1114
rect 5109 1062 5161 1114
rect 5173 1062 5225 1114
rect 5237 1062 5289 1114
<< metal2 >>
rect 1122 6277 1178 7077
rect 1674 6277 1730 7077
rect 2226 6277 2282 7077
rect 2962 6277 3018 7077
rect 3514 6277 3570 7077
rect 4066 6277 4122 7077
rect 4802 6277 4858 7077
rect 5354 6277 5410 7077
rect 5906 6277 5962 7077
rect 6458 6277 6514 7077
rect 572 3732 624 3738
rect 572 3674 624 3680
rect 584 800 612 3674
rect 1136 1426 1164 6277
rect 1582 4448 1638 4457
rect 1582 4383 1638 4392
rect 1400 4208 1452 4214
rect 1400 4150 1452 4156
rect 1412 2553 1440 4150
rect 1596 4078 1624 4383
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1688 3602 1716 6277
rect 1768 5468 2064 5488
rect 1824 5466 1848 5468
rect 1904 5466 1928 5468
rect 1984 5466 2008 5468
rect 1846 5414 1848 5466
rect 1910 5414 1922 5466
rect 1984 5414 1986 5466
rect 1824 5412 1848 5414
rect 1904 5412 1928 5414
rect 1984 5412 2008 5414
rect 1768 5392 2064 5412
rect 1768 4380 2064 4400
rect 1824 4378 1848 4380
rect 1904 4378 1928 4380
rect 1984 4378 2008 4380
rect 1846 4326 1848 4378
rect 1910 4326 1922 4378
rect 1984 4326 1986 4378
rect 1824 4324 1848 4326
rect 1904 4324 1928 4326
rect 1984 4324 2008 4326
rect 1768 4304 2064 4324
rect 2240 4146 2268 6277
rect 2581 6012 2877 6032
rect 2637 6010 2661 6012
rect 2717 6010 2741 6012
rect 2797 6010 2821 6012
rect 2659 5958 2661 6010
rect 2723 5958 2735 6010
rect 2797 5958 2799 6010
rect 2637 5956 2661 5958
rect 2717 5956 2741 5958
rect 2797 5956 2821 5958
rect 2581 5936 2877 5956
rect 2581 4924 2877 4944
rect 2637 4922 2661 4924
rect 2717 4922 2741 4924
rect 2797 4922 2821 4924
rect 2659 4870 2661 4922
rect 2723 4870 2735 4922
rect 2797 4870 2799 4922
rect 2637 4868 2661 4870
rect 2717 4868 2741 4870
rect 2797 4868 2821 4870
rect 2581 4848 2877 4868
rect 2976 4690 3004 6277
rect 3528 5658 3556 6277
rect 3528 5630 3832 5658
rect 3394 5468 3690 5488
rect 3450 5466 3474 5468
rect 3530 5466 3554 5468
rect 3610 5466 3634 5468
rect 3472 5414 3474 5466
rect 3536 5414 3548 5466
rect 3610 5414 3612 5466
rect 3450 5412 3474 5414
rect 3530 5412 3554 5414
rect 3610 5412 3634 5414
rect 3394 5392 3690 5412
rect 3054 5264 3110 5273
rect 3054 5199 3110 5208
rect 3238 5264 3294 5273
rect 3238 5199 3294 5208
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 3068 4282 3096 5199
rect 3252 4690 3280 5199
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3394 4380 3690 4400
rect 3450 4378 3474 4380
rect 3530 4378 3554 4380
rect 3610 4378 3634 4380
rect 3472 4326 3474 4378
rect 3536 4326 3548 4378
rect 3610 4326 3612 4378
rect 3450 4324 3474 4326
rect 3530 4324 3554 4326
rect 3610 4324 3634 4326
rect 3394 4304 3690 4324
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2581 3836 2877 3856
rect 2637 3834 2661 3836
rect 2717 3834 2741 3836
rect 2797 3834 2821 3836
rect 2659 3782 2661 3834
rect 2723 3782 2735 3834
rect 2797 3782 2799 3834
rect 2637 3780 2661 3782
rect 2717 3780 2741 3782
rect 2797 3780 2821 3782
rect 2581 3760 2877 3780
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 2228 3460 2280 3466
rect 2228 3402 2280 3408
rect 1768 3292 2064 3312
rect 1824 3290 1848 3292
rect 1904 3290 1928 3292
rect 1984 3290 2008 3292
rect 1846 3238 1848 3290
rect 1910 3238 1922 3290
rect 1984 3238 1986 3290
rect 1824 3236 1848 3238
rect 1904 3236 1928 3238
rect 1984 3236 2008 3238
rect 1768 3216 2064 3236
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1398 2544 1454 2553
rect 1398 2479 1454 2488
rect 1216 1964 1268 1970
rect 1216 1906 1268 1912
rect 1124 1420 1176 1426
rect 1124 1362 1176 1368
rect 1228 1034 1256 1906
rect 1136 1006 1256 1034
rect 1136 800 1164 1006
rect 1688 800 1716 2790
rect 1768 2204 2064 2224
rect 1824 2202 1848 2204
rect 1904 2202 1928 2204
rect 1984 2202 2008 2204
rect 1846 2150 1848 2202
rect 1910 2150 1922 2202
rect 1984 2150 1986 2202
rect 1824 2148 1848 2150
rect 1904 2148 1928 2150
rect 1984 2148 2008 2150
rect 1768 2128 2064 2148
rect 1768 1116 2064 1136
rect 1824 1114 1848 1116
rect 1904 1114 1928 1116
rect 1984 1114 2008 1116
rect 1846 1062 1848 1114
rect 1910 1062 1922 1114
rect 1984 1062 1986 1114
rect 1824 1060 1848 1062
rect 1904 1060 1928 1062
rect 1984 1060 2008 1062
rect 1768 1040 2064 1060
rect 2240 800 2268 3402
rect 2792 3189 2820 3538
rect 2779 3183 2831 3189
rect 2779 3125 2831 3131
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 2581 2748 2877 2768
rect 2637 2746 2661 2748
rect 2717 2746 2741 2748
rect 2797 2746 2821 2748
rect 2659 2694 2661 2746
rect 2723 2694 2735 2746
rect 2797 2694 2799 2746
rect 2637 2692 2661 2694
rect 2717 2692 2741 2694
rect 2797 2692 2821 2694
rect 2581 2672 2877 2692
rect 2962 2544 3018 2553
rect 2962 2479 3018 2488
rect 2320 2372 2372 2378
rect 2320 2314 2372 2320
rect 2332 1902 2360 2314
rect 2320 1896 2372 1902
rect 2320 1838 2372 1844
rect 2581 1660 2877 1680
rect 2637 1658 2661 1660
rect 2717 1658 2741 1660
rect 2797 1658 2821 1660
rect 2659 1606 2661 1658
rect 2723 1606 2735 1658
rect 2797 1606 2799 1658
rect 2637 1604 2661 1606
rect 2717 1604 2741 1606
rect 2797 1604 2821 1606
rect 2581 1584 2877 1604
rect 2976 1426 3004 2479
rect 2964 1420 3016 1426
rect 2964 1362 3016 1368
rect 3068 1170 3096 2926
rect 3160 1873 3188 3538
rect 3394 3292 3690 3312
rect 3450 3290 3474 3292
rect 3530 3290 3554 3292
rect 3610 3290 3634 3292
rect 3472 3238 3474 3290
rect 3536 3238 3548 3290
rect 3610 3238 3612 3290
rect 3450 3236 3474 3238
rect 3530 3236 3554 3238
rect 3610 3236 3634 3238
rect 3394 3216 3690 3236
rect 3238 3088 3294 3097
rect 3238 3023 3294 3032
rect 3252 1902 3280 3023
rect 3394 2204 3690 2224
rect 3450 2202 3474 2204
rect 3530 2202 3554 2204
rect 3610 2202 3634 2204
rect 3472 2150 3474 2202
rect 3536 2150 3548 2202
rect 3610 2150 3612 2202
rect 3450 2148 3474 2150
rect 3530 2148 3554 2150
rect 3610 2148 3634 2150
rect 3394 2128 3690 2148
rect 3804 1902 3832 5630
rect 4080 5250 4108 6277
rect 4206 6012 4502 6032
rect 4262 6010 4286 6012
rect 4342 6010 4366 6012
rect 4422 6010 4446 6012
rect 4284 5958 4286 6010
rect 4348 5958 4360 6010
rect 4422 5958 4424 6010
rect 4262 5956 4286 5958
rect 4342 5956 4366 5958
rect 4422 5956 4446 5958
rect 4206 5936 4502 5956
rect 4526 5808 4582 5817
rect 4526 5743 4582 5752
rect 3988 5222 4108 5250
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3240 1896 3292 1902
rect 3146 1864 3202 1873
rect 3240 1838 3292 1844
rect 3792 1896 3844 1902
rect 3792 1838 3844 1844
rect 3146 1799 3202 1808
rect 3240 1760 3292 1766
rect 3240 1702 3292 1708
rect 2976 1142 3096 1170
rect 2976 800 3004 1142
rect 3252 898 3280 1702
rect 3394 1116 3690 1136
rect 3450 1114 3474 1116
rect 3530 1114 3554 1116
rect 3610 1114 3634 1116
rect 3472 1062 3474 1114
rect 3536 1062 3548 1114
rect 3610 1062 3612 1114
rect 3450 1060 3474 1062
rect 3530 1060 3554 1062
rect 3610 1060 3634 1062
rect 3394 1040 3690 1060
rect 3896 921 3924 4422
rect 3988 2038 4016 5222
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4080 4593 4108 5102
rect 4206 4924 4502 4944
rect 4262 4922 4286 4924
rect 4342 4922 4366 4924
rect 4422 4922 4446 4924
rect 4284 4870 4286 4922
rect 4348 4870 4360 4922
rect 4422 4870 4424 4922
rect 4262 4868 4286 4870
rect 4342 4868 4366 4870
rect 4422 4868 4446 4870
rect 4206 4848 4502 4868
rect 4066 4584 4122 4593
rect 4066 4519 4122 4528
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3976 2032 4028 2038
rect 3976 1974 4028 1980
rect 3882 912 3938 921
rect 3252 870 3556 898
rect 3528 800 3556 870
rect 3882 847 3938 856
rect 4080 800 4108 4014
rect 4206 3836 4502 3856
rect 4262 3834 4286 3836
rect 4342 3834 4366 3836
rect 4422 3834 4446 3836
rect 4284 3782 4286 3834
rect 4348 3782 4360 3834
rect 4422 3782 4424 3834
rect 4262 3780 4286 3782
rect 4342 3780 4366 3782
rect 4422 3780 4446 3782
rect 4206 3760 4502 3780
rect 4540 3602 4568 5743
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4632 2854 4660 5102
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4724 3738 4752 4422
rect 4816 4127 4844 6277
rect 5019 5468 5315 5488
rect 5075 5466 5099 5468
rect 5155 5466 5179 5468
rect 5235 5466 5259 5468
rect 5097 5414 5099 5466
rect 5161 5414 5173 5466
rect 5235 5414 5237 5466
rect 5075 5412 5099 5414
rect 5155 5412 5179 5414
rect 5235 5412 5259 5414
rect 5019 5392 5315 5412
rect 5019 4380 5315 4400
rect 5075 4378 5099 4380
rect 5155 4378 5179 4380
rect 5235 4378 5259 4380
rect 5097 4326 5099 4378
rect 5161 4326 5173 4378
rect 5235 4326 5237 4378
rect 5075 4324 5099 4326
rect 5155 4324 5179 4326
rect 5235 4324 5259 4326
rect 5019 4304 5315 4324
rect 5368 4298 5396 6277
rect 5368 4270 5488 4298
rect 4816 4099 5028 4127
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4712 3732 4764 3738
rect 4712 3674 4764 3680
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4206 2748 4502 2768
rect 4262 2746 4286 2748
rect 4342 2746 4366 2748
rect 4422 2746 4446 2748
rect 4284 2694 4286 2746
rect 4348 2694 4360 2746
rect 4422 2694 4424 2746
rect 4262 2692 4286 2694
rect 4342 2692 4366 2694
rect 4422 2692 4446 2694
rect 4206 2672 4502 2692
rect 4618 1728 4674 1737
rect 4206 1660 4502 1680
rect 4724 1714 4752 3402
rect 4908 2446 4936 3946
rect 5000 3602 5028 4099
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 5019 3292 5315 3312
rect 5075 3290 5099 3292
rect 5155 3290 5179 3292
rect 5235 3290 5259 3292
rect 5097 3238 5099 3290
rect 5161 3238 5173 3290
rect 5235 3238 5237 3290
rect 5075 3236 5099 3238
rect 5155 3236 5179 3238
rect 5235 3236 5259 3238
rect 5019 3216 5315 3236
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5019 2204 5315 2224
rect 5075 2202 5099 2204
rect 5155 2202 5179 2204
rect 5235 2202 5259 2204
rect 5097 2150 5099 2202
rect 5161 2150 5173 2202
rect 5235 2150 5237 2202
rect 5075 2148 5099 2150
rect 5155 2148 5179 2150
rect 5235 2148 5259 2150
rect 5019 2128 5315 2148
rect 4724 1686 4844 1714
rect 4618 1663 4674 1672
rect 4262 1658 4286 1660
rect 4342 1658 4366 1660
rect 4422 1658 4446 1660
rect 4284 1606 4286 1658
rect 4348 1606 4360 1658
rect 4422 1606 4424 1658
rect 4262 1604 4286 1606
rect 4342 1604 4366 1606
rect 4422 1604 4446 1606
rect 4206 1584 4502 1604
rect 4632 1426 4660 1663
rect 4620 1420 4672 1426
rect 4620 1362 4672 1368
rect 4816 800 4844 1686
rect 5019 1116 5315 1136
rect 5075 1114 5099 1116
rect 5155 1114 5179 1116
rect 5235 1114 5259 1116
rect 5097 1062 5099 1114
rect 5161 1062 5173 1114
rect 5235 1062 5237 1114
rect 5075 1060 5099 1062
rect 5155 1060 5179 1062
rect 5235 1060 5259 1062
rect 5019 1040 5315 1060
rect 5368 800 5396 4014
rect 5460 2514 5488 4270
rect 5920 3670 5948 6277
rect 5908 3664 5960 3670
rect 5630 3632 5686 3641
rect 5908 3606 5960 3612
rect 5630 3567 5686 3576
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5644 1902 5672 3567
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5632 1896 5684 1902
rect 5632 1838 5684 1844
rect 5920 800 5948 3130
rect 6472 2378 6500 6277
rect 6460 2372 6512 2378
rect 6460 2314 6512 2320
rect 570 0 626 800
rect 1122 0 1178 800
rect 1674 0 1730 800
rect 2226 0 2282 800
rect 2962 0 3018 800
rect 3514 0 3570 800
rect 4066 0 4122 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
<< via2 >>
rect 1582 4392 1638 4448
rect 1768 5466 1824 5468
rect 1848 5466 1904 5468
rect 1928 5466 1984 5468
rect 2008 5466 2064 5468
rect 1768 5414 1794 5466
rect 1794 5414 1824 5466
rect 1848 5414 1858 5466
rect 1858 5414 1904 5466
rect 1928 5414 1974 5466
rect 1974 5414 1984 5466
rect 2008 5414 2038 5466
rect 2038 5414 2064 5466
rect 1768 5412 1824 5414
rect 1848 5412 1904 5414
rect 1928 5412 1984 5414
rect 2008 5412 2064 5414
rect 1768 4378 1824 4380
rect 1848 4378 1904 4380
rect 1928 4378 1984 4380
rect 2008 4378 2064 4380
rect 1768 4326 1794 4378
rect 1794 4326 1824 4378
rect 1848 4326 1858 4378
rect 1858 4326 1904 4378
rect 1928 4326 1974 4378
rect 1974 4326 1984 4378
rect 2008 4326 2038 4378
rect 2038 4326 2064 4378
rect 1768 4324 1824 4326
rect 1848 4324 1904 4326
rect 1928 4324 1984 4326
rect 2008 4324 2064 4326
rect 2581 6010 2637 6012
rect 2661 6010 2717 6012
rect 2741 6010 2797 6012
rect 2821 6010 2877 6012
rect 2581 5958 2607 6010
rect 2607 5958 2637 6010
rect 2661 5958 2671 6010
rect 2671 5958 2717 6010
rect 2741 5958 2787 6010
rect 2787 5958 2797 6010
rect 2821 5958 2851 6010
rect 2851 5958 2877 6010
rect 2581 5956 2637 5958
rect 2661 5956 2717 5958
rect 2741 5956 2797 5958
rect 2821 5956 2877 5958
rect 2581 4922 2637 4924
rect 2661 4922 2717 4924
rect 2741 4922 2797 4924
rect 2821 4922 2877 4924
rect 2581 4870 2607 4922
rect 2607 4870 2637 4922
rect 2661 4870 2671 4922
rect 2671 4870 2717 4922
rect 2741 4870 2787 4922
rect 2787 4870 2797 4922
rect 2821 4870 2851 4922
rect 2851 4870 2877 4922
rect 2581 4868 2637 4870
rect 2661 4868 2717 4870
rect 2741 4868 2797 4870
rect 2821 4868 2877 4870
rect 3394 5466 3450 5468
rect 3474 5466 3530 5468
rect 3554 5466 3610 5468
rect 3634 5466 3690 5468
rect 3394 5414 3420 5466
rect 3420 5414 3450 5466
rect 3474 5414 3484 5466
rect 3484 5414 3530 5466
rect 3554 5414 3600 5466
rect 3600 5414 3610 5466
rect 3634 5414 3664 5466
rect 3664 5414 3690 5466
rect 3394 5412 3450 5414
rect 3474 5412 3530 5414
rect 3554 5412 3610 5414
rect 3634 5412 3690 5414
rect 3054 5208 3110 5264
rect 3238 5208 3294 5264
rect 3394 4378 3450 4380
rect 3474 4378 3530 4380
rect 3554 4378 3610 4380
rect 3634 4378 3690 4380
rect 3394 4326 3420 4378
rect 3420 4326 3450 4378
rect 3474 4326 3484 4378
rect 3484 4326 3530 4378
rect 3554 4326 3600 4378
rect 3600 4326 3610 4378
rect 3634 4326 3664 4378
rect 3664 4326 3690 4378
rect 3394 4324 3450 4326
rect 3474 4324 3530 4326
rect 3554 4324 3610 4326
rect 3634 4324 3690 4326
rect 2581 3834 2637 3836
rect 2661 3834 2717 3836
rect 2741 3834 2797 3836
rect 2821 3834 2877 3836
rect 2581 3782 2607 3834
rect 2607 3782 2637 3834
rect 2661 3782 2671 3834
rect 2671 3782 2717 3834
rect 2741 3782 2787 3834
rect 2787 3782 2797 3834
rect 2821 3782 2851 3834
rect 2851 3782 2877 3834
rect 2581 3780 2637 3782
rect 2661 3780 2717 3782
rect 2741 3780 2797 3782
rect 2821 3780 2877 3782
rect 1768 3290 1824 3292
rect 1848 3290 1904 3292
rect 1928 3290 1984 3292
rect 2008 3290 2064 3292
rect 1768 3238 1794 3290
rect 1794 3238 1824 3290
rect 1848 3238 1858 3290
rect 1858 3238 1904 3290
rect 1928 3238 1974 3290
rect 1974 3238 1984 3290
rect 2008 3238 2038 3290
rect 2038 3238 2064 3290
rect 1768 3236 1824 3238
rect 1848 3236 1904 3238
rect 1928 3236 1984 3238
rect 2008 3236 2064 3238
rect 1398 2488 1454 2544
rect 1768 2202 1824 2204
rect 1848 2202 1904 2204
rect 1928 2202 1984 2204
rect 2008 2202 2064 2204
rect 1768 2150 1794 2202
rect 1794 2150 1824 2202
rect 1848 2150 1858 2202
rect 1858 2150 1904 2202
rect 1928 2150 1974 2202
rect 1974 2150 1984 2202
rect 2008 2150 2038 2202
rect 2038 2150 2064 2202
rect 1768 2148 1824 2150
rect 1848 2148 1904 2150
rect 1928 2148 1984 2150
rect 2008 2148 2064 2150
rect 1768 1114 1824 1116
rect 1848 1114 1904 1116
rect 1928 1114 1984 1116
rect 2008 1114 2064 1116
rect 1768 1062 1794 1114
rect 1794 1062 1824 1114
rect 1848 1062 1858 1114
rect 1858 1062 1904 1114
rect 1928 1062 1974 1114
rect 1974 1062 1984 1114
rect 2008 1062 2038 1114
rect 2038 1062 2064 1114
rect 1768 1060 1824 1062
rect 1848 1060 1904 1062
rect 1928 1060 1984 1062
rect 2008 1060 2064 1062
rect 2581 2746 2637 2748
rect 2661 2746 2717 2748
rect 2741 2746 2797 2748
rect 2821 2746 2877 2748
rect 2581 2694 2607 2746
rect 2607 2694 2637 2746
rect 2661 2694 2671 2746
rect 2671 2694 2717 2746
rect 2741 2694 2787 2746
rect 2787 2694 2797 2746
rect 2821 2694 2851 2746
rect 2851 2694 2877 2746
rect 2581 2692 2637 2694
rect 2661 2692 2717 2694
rect 2741 2692 2797 2694
rect 2821 2692 2877 2694
rect 2962 2488 3018 2544
rect 2581 1658 2637 1660
rect 2661 1658 2717 1660
rect 2741 1658 2797 1660
rect 2821 1658 2877 1660
rect 2581 1606 2607 1658
rect 2607 1606 2637 1658
rect 2661 1606 2671 1658
rect 2671 1606 2717 1658
rect 2741 1606 2787 1658
rect 2787 1606 2797 1658
rect 2821 1606 2851 1658
rect 2851 1606 2877 1658
rect 2581 1604 2637 1606
rect 2661 1604 2717 1606
rect 2741 1604 2797 1606
rect 2821 1604 2877 1606
rect 3394 3290 3450 3292
rect 3474 3290 3530 3292
rect 3554 3290 3610 3292
rect 3634 3290 3690 3292
rect 3394 3238 3420 3290
rect 3420 3238 3450 3290
rect 3474 3238 3484 3290
rect 3484 3238 3530 3290
rect 3554 3238 3600 3290
rect 3600 3238 3610 3290
rect 3634 3238 3664 3290
rect 3664 3238 3690 3290
rect 3394 3236 3450 3238
rect 3474 3236 3530 3238
rect 3554 3236 3610 3238
rect 3634 3236 3690 3238
rect 3238 3032 3294 3088
rect 3394 2202 3450 2204
rect 3474 2202 3530 2204
rect 3554 2202 3610 2204
rect 3634 2202 3690 2204
rect 3394 2150 3420 2202
rect 3420 2150 3450 2202
rect 3474 2150 3484 2202
rect 3484 2150 3530 2202
rect 3554 2150 3600 2202
rect 3600 2150 3610 2202
rect 3634 2150 3664 2202
rect 3664 2150 3690 2202
rect 3394 2148 3450 2150
rect 3474 2148 3530 2150
rect 3554 2148 3610 2150
rect 3634 2148 3690 2150
rect 4206 6010 4262 6012
rect 4286 6010 4342 6012
rect 4366 6010 4422 6012
rect 4446 6010 4502 6012
rect 4206 5958 4232 6010
rect 4232 5958 4262 6010
rect 4286 5958 4296 6010
rect 4296 5958 4342 6010
rect 4366 5958 4412 6010
rect 4412 5958 4422 6010
rect 4446 5958 4476 6010
rect 4476 5958 4502 6010
rect 4206 5956 4262 5958
rect 4286 5956 4342 5958
rect 4366 5956 4422 5958
rect 4446 5956 4502 5958
rect 4526 5752 4582 5808
rect 3146 1808 3202 1864
rect 3394 1114 3450 1116
rect 3474 1114 3530 1116
rect 3554 1114 3610 1116
rect 3634 1114 3690 1116
rect 3394 1062 3420 1114
rect 3420 1062 3450 1114
rect 3474 1062 3484 1114
rect 3484 1062 3530 1114
rect 3554 1062 3600 1114
rect 3600 1062 3610 1114
rect 3634 1062 3664 1114
rect 3664 1062 3690 1114
rect 3394 1060 3450 1062
rect 3474 1060 3530 1062
rect 3554 1060 3610 1062
rect 3634 1060 3690 1062
rect 4206 4922 4262 4924
rect 4286 4922 4342 4924
rect 4366 4922 4422 4924
rect 4446 4922 4502 4924
rect 4206 4870 4232 4922
rect 4232 4870 4262 4922
rect 4286 4870 4296 4922
rect 4296 4870 4342 4922
rect 4366 4870 4412 4922
rect 4412 4870 4422 4922
rect 4446 4870 4476 4922
rect 4476 4870 4502 4922
rect 4206 4868 4262 4870
rect 4286 4868 4342 4870
rect 4366 4868 4422 4870
rect 4446 4868 4502 4870
rect 4066 4528 4122 4584
rect 3882 856 3938 912
rect 4206 3834 4262 3836
rect 4286 3834 4342 3836
rect 4366 3834 4422 3836
rect 4446 3834 4502 3836
rect 4206 3782 4232 3834
rect 4232 3782 4262 3834
rect 4286 3782 4296 3834
rect 4296 3782 4342 3834
rect 4366 3782 4412 3834
rect 4412 3782 4422 3834
rect 4446 3782 4476 3834
rect 4476 3782 4502 3834
rect 4206 3780 4262 3782
rect 4286 3780 4342 3782
rect 4366 3780 4422 3782
rect 4446 3780 4502 3782
rect 5019 5466 5075 5468
rect 5099 5466 5155 5468
rect 5179 5466 5235 5468
rect 5259 5466 5315 5468
rect 5019 5414 5045 5466
rect 5045 5414 5075 5466
rect 5099 5414 5109 5466
rect 5109 5414 5155 5466
rect 5179 5414 5225 5466
rect 5225 5414 5235 5466
rect 5259 5414 5289 5466
rect 5289 5414 5315 5466
rect 5019 5412 5075 5414
rect 5099 5412 5155 5414
rect 5179 5412 5235 5414
rect 5259 5412 5315 5414
rect 5019 4378 5075 4380
rect 5099 4378 5155 4380
rect 5179 4378 5235 4380
rect 5259 4378 5315 4380
rect 5019 4326 5045 4378
rect 5045 4326 5075 4378
rect 5099 4326 5109 4378
rect 5109 4326 5155 4378
rect 5179 4326 5225 4378
rect 5225 4326 5235 4378
rect 5259 4326 5289 4378
rect 5289 4326 5315 4378
rect 5019 4324 5075 4326
rect 5099 4324 5155 4326
rect 5179 4324 5235 4326
rect 5259 4324 5315 4326
rect 4206 2746 4262 2748
rect 4286 2746 4342 2748
rect 4366 2746 4422 2748
rect 4446 2746 4502 2748
rect 4206 2694 4232 2746
rect 4232 2694 4262 2746
rect 4286 2694 4296 2746
rect 4296 2694 4342 2746
rect 4366 2694 4412 2746
rect 4412 2694 4422 2746
rect 4446 2694 4476 2746
rect 4476 2694 4502 2746
rect 4206 2692 4262 2694
rect 4286 2692 4342 2694
rect 4366 2692 4422 2694
rect 4446 2692 4502 2694
rect 4618 1672 4674 1728
rect 5019 3290 5075 3292
rect 5099 3290 5155 3292
rect 5179 3290 5235 3292
rect 5259 3290 5315 3292
rect 5019 3238 5045 3290
rect 5045 3238 5075 3290
rect 5099 3238 5109 3290
rect 5109 3238 5155 3290
rect 5179 3238 5225 3290
rect 5225 3238 5235 3290
rect 5259 3238 5289 3290
rect 5289 3238 5315 3290
rect 5019 3236 5075 3238
rect 5099 3236 5155 3238
rect 5179 3236 5235 3238
rect 5259 3236 5315 3238
rect 5019 2202 5075 2204
rect 5099 2202 5155 2204
rect 5179 2202 5235 2204
rect 5259 2202 5315 2204
rect 5019 2150 5045 2202
rect 5045 2150 5075 2202
rect 5099 2150 5109 2202
rect 5109 2150 5155 2202
rect 5179 2150 5225 2202
rect 5225 2150 5235 2202
rect 5259 2150 5289 2202
rect 5289 2150 5315 2202
rect 5019 2148 5075 2150
rect 5099 2148 5155 2150
rect 5179 2148 5235 2150
rect 5259 2148 5315 2150
rect 4206 1658 4262 1660
rect 4286 1658 4342 1660
rect 4366 1658 4422 1660
rect 4446 1658 4502 1660
rect 4206 1606 4232 1658
rect 4232 1606 4262 1658
rect 4286 1606 4296 1658
rect 4296 1606 4342 1658
rect 4366 1606 4412 1658
rect 4412 1606 4422 1658
rect 4446 1606 4476 1658
rect 4476 1606 4502 1658
rect 4206 1604 4262 1606
rect 4286 1604 4342 1606
rect 4366 1604 4422 1606
rect 4446 1604 4502 1606
rect 5019 1114 5075 1116
rect 5099 1114 5155 1116
rect 5179 1114 5235 1116
rect 5259 1114 5315 1116
rect 5019 1062 5045 1114
rect 5045 1062 5075 1114
rect 5099 1062 5109 1114
rect 5109 1062 5155 1114
rect 5179 1062 5225 1114
rect 5225 1062 5235 1114
rect 5259 1062 5289 1114
rect 5289 1062 5315 1114
rect 5019 1060 5075 1062
rect 5099 1060 5155 1062
rect 5179 1060 5235 1062
rect 5259 1060 5315 1062
rect 5630 3576 5686 3632
<< metal3 >>
rect 0 6082 800 6112
rect 0 6022 2330 6082
rect 0 5992 800 6022
rect 2270 5810 2330 6022
rect 2569 6016 2889 6017
rect 2569 5952 2577 6016
rect 2641 5952 2657 6016
rect 2721 5952 2737 6016
rect 2801 5952 2817 6016
rect 2881 5952 2889 6016
rect 2569 5951 2889 5952
rect 4194 6016 4514 6017
rect 4194 5952 4202 6016
rect 4266 5952 4282 6016
rect 4346 5952 4362 6016
rect 4426 5952 4442 6016
rect 4506 5952 4514 6016
rect 4194 5951 4514 5952
rect 4521 5810 4587 5813
rect 2270 5808 4587 5810
rect 2270 5752 4526 5808
rect 4582 5752 4587 5808
rect 2270 5750 4587 5752
rect 4521 5747 4587 5750
rect 1756 5472 2076 5473
rect 1756 5408 1764 5472
rect 1828 5408 1844 5472
rect 1908 5408 1924 5472
rect 1988 5408 2004 5472
rect 2068 5408 2076 5472
rect 1756 5407 2076 5408
rect 3382 5472 3702 5473
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 5407 3702 5408
rect 5007 5472 5327 5473
rect 5007 5408 5015 5472
rect 5079 5408 5095 5472
rect 5159 5408 5175 5472
rect 5239 5408 5255 5472
rect 5319 5408 5327 5472
rect 5007 5407 5327 5408
rect 0 5266 800 5296
rect 3049 5266 3115 5269
rect 0 5264 3115 5266
rect 0 5208 3054 5264
rect 3110 5208 3115 5264
rect 0 5206 3115 5208
rect 0 5176 800 5206
rect 3049 5203 3115 5206
rect 3233 5266 3299 5269
rect 6309 5266 7109 5296
rect 3233 5264 7109 5266
rect 3233 5208 3238 5264
rect 3294 5208 7109 5264
rect 3233 5206 7109 5208
rect 3233 5203 3299 5206
rect 6309 5176 7109 5206
rect 2569 4928 2889 4929
rect 2569 4864 2577 4928
rect 2641 4864 2657 4928
rect 2721 4864 2737 4928
rect 2801 4864 2817 4928
rect 2881 4864 2889 4928
rect 2569 4863 2889 4864
rect 4194 4928 4514 4929
rect 4194 4864 4202 4928
rect 4266 4864 4282 4928
rect 4346 4864 4362 4928
rect 4426 4864 4442 4928
rect 4506 4864 4514 4928
rect 4194 4863 4514 4864
rect 4061 4586 4127 4589
rect 4061 4584 5458 4586
rect 4061 4528 4066 4584
rect 4122 4528 5458 4584
rect 4061 4526 5458 4528
rect 4061 4523 4127 4526
rect 0 4450 800 4480
rect 1577 4450 1643 4453
rect 0 4448 1643 4450
rect 0 4392 1582 4448
rect 1638 4392 1643 4448
rect 0 4390 1643 4392
rect 5398 4450 5458 4526
rect 6309 4450 7109 4480
rect 5398 4390 7109 4450
rect 0 4360 800 4390
rect 1577 4387 1643 4390
rect 1756 4384 2076 4385
rect 1756 4320 1764 4384
rect 1828 4320 1844 4384
rect 1908 4320 1924 4384
rect 1988 4320 2004 4384
rect 2068 4320 2076 4384
rect 1756 4319 2076 4320
rect 3382 4384 3702 4385
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 4319 3702 4320
rect 5007 4384 5327 4385
rect 5007 4320 5015 4384
rect 5079 4320 5095 4384
rect 5159 4320 5175 4384
rect 5239 4320 5255 4384
rect 5319 4320 5327 4384
rect 6309 4360 7109 4390
rect 5007 4319 5327 4320
rect 2569 3840 2889 3841
rect 2569 3776 2577 3840
rect 2641 3776 2657 3840
rect 2721 3776 2737 3840
rect 2801 3776 2817 3840
rect 2881 3776 2889 3840
rect 2569 3775 2889 3776
rect 4194 3840 4514 3841
rect 4194 3776 4202 3840
rect 4266 3776 4282 3840
rect 4346 3776 4362 3840
rect 4426 3776 4442 3840
rect 4506 3776 4514 3840
rect 4194 3775 4514 3776
rect 5625 3634 5691 3637
rect 6309 3634 7109 3664
rect 5625 3632 7109 3634
rect 5625 3576 5630 3632
rect 5686 3576 7109 3632
rect 5625 3574 7109 3576
rect 5625 3571 5691 3574
rect 6309 3544 7109 3574
rect 0 3362 800 3392
rect 0 3302 1594 3362
rect 0 3272 800 3302
rect 1534 3090 1594 3302
rect 1756 3296 2076 3297
rect 1756 3232 1764 3296
rect 1828 3232 1844 3296
rect 1908 3232 1924 3296
rect 1988 3232 2004 3296
rect 2068 3232 2076 3296
rect 1756 3231 2076 3232
rect 3382 3296 3702 3297
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 3231 3702 3232
rect 5007 3296 5327 3297
rect 5007 3232 5015 3296
rect 5079 3232 5095 3296
rect 5159 3232 5175 3296
rect 5239 3232 5255 3296
rect 5319 3232 5327 3296
rect 5007 3231 5327 3232
rect 3233 3090 3299 3093
rect 1534 3088 3299 3090
rect 1534 3032 3238 3088
rect 3294 3032 3299 3088
rect 1534 3030 3299 3032
rect 3233 3027 3299 3030
rect 2569 2752 2889 2753
rect 2569 2688 2577 2752
rect 2641 2688 2657 2752
rect 2721 2688 2737 2752
rect 2801 2688 2817 2752
rect 2881 2688 2889 2752
rect 2569 2687 2889 2688
rect 4194 2752 4514 2753
rect 4194 2688 4202 2752
rect 4266 2688 4282 2752
rect 4346 2688 4362 2752
rect 4426 2688 4442 2752
rect 4506 2688 4514 2752
rect 4194 2687 4514 2688
rect 0 2546 800 2576
rect 1393 2546 1459 2549
rect 0 2544 1459 2546
rect 0 2488 1398 2544
rect 1454 2488 1459 2544
rect 0 2486 1459 2488
rect 0 2456 800 2486
rect 1393 2483 1459 2486
rect 2957 2546 3023 2549
rect 6309 2546 7109 2576
rect 2957 2544 7109 2546
rect 2957 2488 2962 2544
rect 3018 2488 7109 2544
rect 2957 2486 7109 2488
rect 2957 2483 3023 2486
rect 6309 2456 7109 2486
rect 1756 2208 2076 2209
rect 1756 2144 1764 2208
rect 1828 2144 1844 2208
rect 1908 2144 1924 2208
rect 1988 2144 2004 2208
rect 2068 2144 2076 2208
rect 1756 2143 2076 2144
rect 3382 2208 3702 2209
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 2143 3702 2144
rect 5007 2208 5327 2209
rect 5007 2144 5015 2208
rect 5079 2144 5095 2208
rect 5159 2144 5175 2208
rect 5239 2144 5255 2208
rect 5319 2144 5327 2208
rect 5007 2143 5327 2144
rect 3141 1866 3207 1869
rect 1534 1864 3207 1866
rect 1534 1808 3146 1864
rect 3202 1808 3207 1864
rect 1534 1806 3207 1808
rect 0 1730 800 1760
rect 1534 1730 1594 1806
rect 3141 1803 3207 1806
rect 0 1670 1594 1730
rect 4613 1730 4679 1733
rect 6309 1730 7109 1760
rect 4613 1728 7109 1730
rect 4613 1672 4618 1728
rect 4674 1672 7109 1728
rect 4613 1670 7109 1672
rect 0 1640 800 1670
rect 4613 1667 4679 1670
rect 2569 1664 2889 1665
rect 2569 1600 2577 1664
rect 2641 1600 2657 1664
rect 2721 1600 2737 1664
rect 2801 1600 2817 1664
rect 2881 1600 2889 1664
rect 2569 1599 2889 1600
rect 4194 1664 4514 1665
rect 4194 1600 4202 1664
rect 4266 1600 4282 1664
rect 4346 1600 4362 1664
rect 4426 1600 4442 1664
rect 4506 1600 4514 1664
rect 6309 1640 7109 1670
rect 4194 1599 4514 1600
rect 1756 1120 2076 1121
rect 1756 1056 1764 1120
rect 1828 1056 1844 1120
rect 1908 1056 1924 1120
rect 1988 1056 2004 1120
rect 2068 1056 2076 1120
rect 1756 1055 2076 1056
rect 3382 1120 3702 1121
rect 3382 1056 3390 1120
rect 3454 1056 3470 1120
rect 3534 1056 3550 1120
rect 3614 1056 3630 1120
rect 3694 1056 3702 1120
rect 3382 1055 3702 1056
rect 5007 1120 5327 1121
rect 5007 1056 5015 1120
rect 5079 1056 5095 1120
rect 5159 1056 5175 1120
rect 5239 1056 5255 1120
rect 5319 1056 5327 1120
rect 5007 1055 5327 1056
rect 3877 914 3943 917
rect 6309 914 7109 944
rect 3877 912 7109 914
rect 3877 856 3882 912
rect 3938 856 7109 912
rect 3877 854 7109 856
rect 3877 851 3943 854
rect 6309 824 7109 854
<< via3 >>
rect 2577 6012 2641 6016
rect 2577 5956 2581 6012
rect 2581 5956 2637 6012
rect 2637 5956 2641 6012
rect 2577 5952 2641 5956
rect 2657 6012 2721 6016
rect 2657 5956 2661 6012
rect 2661 5956 2717 6012
rect 2717 5956 2721 6012
rect 2657 5952 2721 5956
rect 2737 6012 2801 6016
rect 2737 5956 2741 6012
rect 2741 5956 2797 6012
rect 2797 5956 2801 6012
rect 2737 5952 2801 5956
rect 2817 6012 2881 6016
rect 2817 5956 2821 6012
rect 2821 5956 2877 6012
rect 2877 5956 2881 6012
rect 2817 5952 2881 5956
rect 4202 6012 4266 6016
rect 4202 5956 4206 6012
rect 4206 5956 4262 6012
rect 4262 5956 4266 6012
rect 4202 5952 4266 5956
rect 4282 6012 4346 6016
rect 4282 5956 4286 6012
rect 4286 5956 4342 6012
rect 4342 5956 4346 6012
rect 4282 5952 4346 5956
rect 4362 6012 4426 6016
rect 4362 5956 4366 6012
rect 4366 5956 4422 6012
rect 4422 5956 4426 6012
rect 4362 5952 4426 5956
rect 4442 6012 4506 6016
rect 4442 5956 4446 6012
rect 4446 5956 4502 6012
rect 4502 5956 4506 6012
rect 4442 5952 4506 5956
rect 1764 5468 1828 5472
rect 1764 5412 1768 5468
rect 1768 5412 1824 5468
rect 1824 5412 1828 5468
rect 1764 5408 1828 5412
rect 1844 5468 1908 5472
rect 1844 5412 1848 5468
rect 1848 5412 1904 5468
rect 1904 5412 1908 5468
rect 1844 5408 1908 5412
rect 1924 5468 1988 5472
rect 1924 5412 1928 5468
rect 1928 5412 1984 5468
rect 1984 5412 1988 5468
rect 1924 5408 1988 5412
rect 2004 5468 2068 5472
rect 2004 5412 2008 5468
rect 2008 5412 2064 5468
rect 2064 5412 2068 5468
rect 2004 5408 2068 5412
rect 3390 5468 3454 5472
rect 3390 5412 3394 5468
rect 3394 5412 3450 5468
rect 3450 5412 3454 5468
rect 3390 5408 3454 5412
rect 3470 5468 3534 5472
rect 3470 5412 3474 5468
rect 3474 5412 3530 5468
rect 3530 5412 3534 5468
rect 3470 5408 3534 5412
rect 3550 5468 3614 5472
rect 3550 5412 3554 5468
rect 3554 5412 3610 5468
rect 3610 5412 3614 5468
rect 3550 5408 3614 5412
rect 3630 5468 3694 5472
rect 3630 5412 3634 5468
rect 3634 5412 3690 5468
rect 3690 5412 3694 5468
rect 3630 5408 3694 5412
rect 5015 5468 5079 5472
rect 5015 5412 5019 5468
rect 5019 5412 5075 5468
rect 5075 5412 5079 5468
rect 5015 5408 5079 5412
rect 5095 5468 5159 5472
rect 5095 5412 5099 5468
rect 5099 5412 5155 5468
rect 5155 5412 5159 5468
rect 5095 5408 5159 5412
rect 5175 5468 5239 5472
rect 5175 5412 5179 5468
rect 5179 5412 5235 5468
rect 5235 5412 5239 5468
rect 5175 5408 5239 5412
rect 5255 5468 5319 5472
rect 5255 5412 5259 5468
rect 5259 5412 5315 5468
rect 5315 5412 5319 5468
rect 5255 5408 5319 5412
rect 2577 4924 2641 4928
rect 2577 4868 2581 4924
rect 2581 4868 2637 4924
rect 2637 4868 2641 4924
rect 2577 4864 2641 4868
rect 2657 4924 2721 4928
rect 2657 4868 2661 4924
rect 2661 4868 2717 4924
rect 2717 4868 2721 4924
rect 2657 4864 2721 4868
rect 2737 4924 2801 4928
rect 2737 4868 2741 4924
rect 2741 4868 2797 4924
rect 2797 4868 2801 4924
rect 2737 4864 2801 4868
rect 2817 4924 2881 4928
rect 2817 4868 2821 4924
rect 2821 4868 2877 4924
rect 2877 4868 2881 4924
rect 2817 4864 2881 4868
rect 4202 4924 4266 4928
rect 4202 4868 4206 4924
rect 4206 4868 4262 4924
rect 4262 4868 4266 4924
rect 4202 4864 4266 4868
rect 4282 4924 4346 4928
rect 4282 4868 4286 4924
rect 4286 4868 4342 4924
rect 4342 4868 4346 4924
rect 4282 4864 4346 4868
rect 4362 4924 4426 4928
rect 4362 4868 4366 4924
rect 4366 4868 4422 4924
rect 4422 4868 4426 4924
rect 4362 4864 4426 4868
rect 4442 4924 4506 4928
rect 4442 4868 4446 4924
rect 4446 4868 4502 4924
rect 4502 4868 4506 4924
rect 4442 4864 4506 4868
rect 1764 4380 1828 4384
rect 1764 4324 1768 4380
rect 1768 4324 1824 4380
rect 1824 4324 1828 4380
rect 1764 4320 1828 4324
rect 1844 4380 1908 4384
rect 1844 4324 1848 4380
rect 1848 4324 1904 4380
rect 1904 4324 1908 4380
rect 1844 4320 1908 4324
rect 1924 4380 1988 4384
rect 1924 4324 1928 4380
rect 1928 4324 1984 4380
rect 1984 4324 1988 4380
rect 1924 4320 1988 4324
rect 2004 4380 2068 4384
rect 2004 4324 2008 4380
rect 2008 4324 2064 4380
rect 2064 4324 2068 4380
rect 2004 4320 2068 4324
rect 3390 4380 3454 4384
rect 3390 4324 3394 4380
rect 3394 4324 3450 4380
rect 3450 4324 3454 4380
rect 3390 4320 3454 4324
rect 3470 4380 3534 4384
rect 3470 4324 3474 4380
rect 3474 4324 3530 4380
rect 3530 4324 3534 4380
rect 3470 4320 3534 4324
rect 3550 4380 3614 4384
rect 3550 4324 3554 4380
rect 3554 4324 3610 4380
rect 3610 4324 3614 4380
rect 3550 4320 3614 4324
rect 3630 4380 3694 4384
rect 3630 4324 3634 4380
rect 3634 4324 3690 4380
rect 3690 4324 3694 4380
rect 3630 4320 3694 4324
rect 5015 4380 5079 4384
rect 5015 4324 5019 4380
rect 5019 4324 5075 4380
rect 5075 4324 5079 4380
rect 5015 4320 5079 4324
rect 5095 4380 5159 4384
rect 5095 4324 5099 4380
rect 5099 4324 5155 4380
rect 5155 4324 5159 4380
rect 5095 4320 5159 4324
rect 5175 4380 5239 4384
rect 5175 4324 5179 4380
rect 5179 4324 5235 4380
rect 5235 4324 5239 4380
rect 5175 4320 5239 4324
rect 5255 4380 5319 4384
rect 5255 4324 5259 4380
rect 5259 4324 5315 4380
rect 5315 4324 5319 4380
rect 5255 4320 5319 4324
rect 2577 3836 2641 3840
rect 2577 3780 2581 3836
rect 2581 3780 2637 3836
rect 2637 3780 2641 3836
rect 2577 3776 2641 3780
rect 2657 3836 2721 3840
rect 2657 3780 2661 3836
rect 2661 3780 2717 3836
rect 2717 3780 2721 3836
rect 2657 3776 2721 3780
rect 2737 3836 2801 3840
rect 2737 3780 2741 3836
rect 2741 3780 2797 3836
rect 2797 3780 2801 3836
rect 2737 3776 2801 3780
rect 2817 3836 2881 3840
rect 2817 3780 2821 3836
rect 2821 3780 2877 3836
rect 2877 3780 2881 3836
rect 2817 3776 2881 3780
rect 4202 3836 4266 3840
rect 4202 3780 4206 3836
rect 4206 3780 4262 3836
rect 4262 3780 4266 3836
rect 4202 3776 4266 3780
rect 4282 3836 4346 3840
rect 4282 3780 4286 3836
rect 4286 3780 4342 3836
rect 4342 3780 4346 3836
rect 4282 3776 4346 3780
rect 4362 3836 4426 3840
rect 4362 3780 4366 3836
rect 4366 3780 4422 3836
rect 4422 3780 4426 3836
rect 4362 3776 4426 3780
rect 4442 3836 4506 3840
rect 4442 3780 4446 3836
rect 4446 3780 4502 3836
rect 4502 3780 4506 3836
rect 4442 3776 4506 3780
rect 1764 3292 1828 3296
rect 1764 3236 1768 3292
rect 1768 3236 1824 3292
rect 1824 3236 1828 3292
rect 1764 3232 1828 3236
rect 1844 3292 1908 3296
rect 1844 3236 1848 3292
rect 1848 3236 1904 3292
rect 1904 3236 1908 3292
rect 1844 3232 1908 3236
rect 1924 3292 1988 3296
rect 1924 3236 1928 3292
rect 1928 3236 1984 3292
rect 1984 3236 1988 3292
rect 1924 3232 1988 3236
rect 2004 3292 2068 3296
rect 2004 3236 2008 3292
rect 2008 3236 2064 3292
rect 2064 3236 2068 3292
rect 2004 3232 2068 3236
rect 3390 3292 3454 3296
rect 3390 3236 3394 3292
rect 3394 3236 3450 3292
rect 3450 3236 3454 3292
rect 3390 3232 3454 3236
rect 3470 3292 3534 3296
rect 3470 3236 3474 3292
rect 3474 3236 3530 3292
rect 3530 3236 3534 3292
rect 3470 3232 3534 3236
rect 3550 3292 3614 3296
rect 3550 3236 3554 3292
rect 3554 3236 3610 3292
rect 3610 3236 3614 3292
rect 3550 3232 3614 3236
rect 3630 3292 3694 3296
rect 3630 3236 3634 3292
rect 3634 3236 3690 3292
rect 3690 3236 3694 3292
rect 3630 3232 3694 3236
rect 5015 3292 5079 3296
rect 5015 3236 5019 3292
rect 5019 3236 5075 3292
rect 5075 3236 5079 3292
rect 5015 3232 5079 3236
rect 5095 3292 5159 3296
rect 5095 3236 5099 3292
rect 5099 3236 5155 3292
rect 5155 3236 5159 3292
rect 5095 3232 5159 3236
rect 5175 3292 5239 3296
rect 5175 3236 5179 3292
rect 5179 3236 5235 3292
rect 5235 3236 5239 3292
rect 5175 3232 5239 3236
rect 5255 3292 5319 3296
rect 5255 3236 5259 3292
rect 5259 3236 5315 3292
rect 5315 3236 5319 3292
rect 5255 3232 5319 3236
rect 2577 2748 2641 2752
rect 2577 2692 2581 2748
rect 2581 2692 2637 2748
rect 2637 2692 2641 2748
rect 2577 2688 2641 2692
rect 2657 2748 2721 2752
rect 2657 2692 2661 2748
rect 2661 2692 2717 2748
rect 2717 2692 2721 2748
rect 2657 2688 2721 2692
rect 2737 2748 2801 2752
rect 2737 2692 2741 2748
rect 2741 2692 2797 2748
rect 2797 2692 2801 2748
rect 2737 2688 2801 2692
rect 2817 2748 2881 2752
rect 2817 2692 2821 2748
rect 2821 2692 2877 2748
rect 2877 2692 2881 2748
rect 2817 2688 2881 2692
rect 4202 2748 4266 2752
rect 4202 2692 4206 2748
rect 4206 2692 4262 2748
rect 4262 2692 4266 2748
rect 4202 2688 4266 2692
rect 4282 2748 4346 2752
rect 4282 2692 4286 2748
rect 4286 2692 4342 2748
rect 4342 2692 4346 2748
rect 4282 2688 4346 2692
rect 4362 2748 4426 2752
rect 4362 2692 4366 2748
rect 4366 2692 4422 2748
rect 4422 2692 4426 2748
rect 4362 2688 4426 2692
rect 4442 2748 4506 2752
rect 4442 2692 4446 2748
rect 4446 2692 4502 2748
rect 4502 2692 4506 2748
rect 4442 2688 4506 2692
rect 1764 2204 1828 2208
rect 1764 2148 1768 2204
rect 1768 2148 1824 2204
rect 1824 2148 1828 2204
rect 1764 2144 1828 2148
rect 1844 2204 1908 2208
rect 1844 2148 1848 2204
rect 1848 2148 1904 2204
rect 1904 2148 1908 2204
rect 1844 2144 1908 2148
rect 1924 2204 1988 2208
rect 1924 2148 1928 2204
rect 1928 2148 1984 2204
rect 1984 2148 1988 2204
rect 1924 2144 1988 2148
rect 2004 2204 2068 2208
rect 2004 2148 2008 2204
rect 2008 2148 2064 2204
rect 2064 2148 2068 2204
rect 2004 2144 2068 2148
rect 3390 2204 3454 2208
rect 3390 2148 3394 2204
rect 3394 2148 3450 2204
rect 3450 2148 3454 2204
rect 3390 2144 3454 2148
rect 3470 2204 3534 2208
rect 3470 2148 3474 2204
rect 3474 2148 3530 2204
rect 3530 2148 3534 2204
rect 3470 2144 3534 2148
rect 3550 2204 3614 2208
rect 3550 2148 3554 2204
rect 3554 2148 3610 2204
rect 3610 2148 3614 2204
rect 3550 2144 3614 2148
rect 3630 2204 3694 2208
rect 3630 2148 3634 2204
rect 3634 2148 3690 2204
rect 3690 2148 3694 2204
rect 3630 2144 3694 2148
rect 5015 2204 5079 2208
rect 5015 2148 5019 2204
rect 5019 2148 5075 2204
rect 5075 2148 5079 2204
rect 5015 2144 5079 2148
rect 5095 2204 5159 2208
rect 5095 2148 5099 2204
rect 5099 2148 5155 2204
rect 5155 2148 5159 2204
rect 5095 2144 5159 2148
rect 5175 2204 5239 2208
rect 5175 2148 5179 2204
rect 5179 2148 5235 2204
rect 5235 2148 5239 2204
rect 5175 2144 5239 2148
rect 5255 2204 5319 2208
rect 5255 2148 5259 2204
rect 5259 2148 5315 2204
rect 5315 2148 5319 2204
rect 5255 2144 5319 2148
rect 2577 1660 2641 1664
rect 2577 1604 2581 1660
rect 2581 1604 2637 1660
rect 2637 1604 2641 1660
rect 2577 1600 2641 1604
rect 2657 1660 2721 1664
rect 2657 1604 2661 1660
rect 2661 1604 2717 1660
rect 2717 1604 2721 1660
rect 2657 1600 2721 1604
rect 2737 1660 2801 1664
rect 2737 1604 2741 1660
rect 2741 1604 2797 1660
rect 2797 1604 2801 1660
rect 2737 1600 2801 1604
rect 2817 1660 2881 1664
rect 2817 1604 2821 1660
rect 2821 1604 2877 1660
rect 2877 1604 2881 1660
rect 2817 1600 2881 1604
rect 4202 1660 4266 1664
rect 4202 1604 4206 1660
rect 4206 1604 4262 1660
rect 4262 1604 4266 1660
rect 4202 1600 4266 1604
rect 4282 1660 4346 1664
rect 4282 1604 4286 1660
rect 4286 1604 4342 1660
rect 4342 1604 4346 1660
rect 4282 1600 4346 1604
rect 4362 1660 4426 1664
rect 4362 1604 4366 1660
rect 4366 1604 4422 1660
rect 4422 1604 4426 1660
rect 4362 1600 4426 1604
rect 4442 1660 4506 1664
rect 4442 1604 4446 1660
rect 4446 1604 4502 1660
rect 4502 1604 4506 1660
rect 4442 1600 4506 1604
rect 1764 1116 1828 1120
rect 1764 1060 1768 1116
rect 1768 1060 1824 1116
rect 1824 1060 1828 1116
rect 1764 1056 1828 1060
rect 1844 1116 1908 1120
rect 1844 1060 1848 1116
rect 1848 1060 1904 1116
rect 1904 1060 1908 1116
rect 1844 1056 1908 1060
rect 1924 1116 1988 1120
rect 1924 1060 1928 1116
rect 1928 1060 1984 1116
rect 1984 1060 1988 1116
rect 1924 1056 1988 1060
rect 2004 1116 2068 1120
rect 2004 1060 2008 1116
rect 2008 1060 2064 1116
rect 2064 1060 2068 1116
rect 2004 1056 2068 1060
rect 3390 1116 3454 1120
rect 3390 1060 3394 1116
rect 3394 1060 3450 1116
rect 3450 1060 3454 1116
rect 3390 1056 3454 1060
rect 3470 1116 3534 1120
rect 3470 1060 3474 1116
rect 3474 1060 3530 1116
rect 3530 1060 3534 1116
rect 3470 1056 3534 1060
rect 3550 1116 3614 1120
rect 3550 1060 3554 1116
rect 3554 1060 3610 1116
rect 3610 1060 3614 1116
rect 3550 1056 3614 1060
rect 3630 1116 3694 1120
rect 3630 1060 3634 1116
rect 3634 1060 3690 1116
rect 3690 1060 3694 1116
rect 3630 1056 3694 1060
rect 5015 1116 5079 1120
rect 5015 1060 5019 1116
rect 5019 1060 5075 1116
rect 5075 1060 5079 1116
rect 5015 1056 5079 1060
rect 5095 1116 5159 1120
rect 5095 1060 5099 1116
rect 5099 1060 5155 1116
rect 5155 1060 5159 1116
rect 5095 1056 5159 1060
rect 5175 1116 5239 1120
rect 5175 1060 5179 1116
rect 5179 1060 5235 1116
rect 5235 1060 5239 1116
rect 5175 1056 5239 1060
rect 5255 1116 5319 1120
rect 5255 1060 5259 1116
rect 5259 1060 5315 1116
rect 5315 1060 5319 1116
rect 5255 1056 5319 1060
<< metal4 >>
rect 1756 5472 2076 6032
rect 1756 5408 1764 5472
rect 1828 5408 1844 5472
rect 1908 5408 1924 5472
rect 1988 5408 2004 5472
rect 2068 5408 2076 5472
rect 1756 5238 2076 5408
rect 1756 5002 1798 5238
rect 2034 5002 2076 5238
rect 1756 4384 2076 5002
rect 1756 4320 1764 4384
rect 1828 4320 1844 4384
rect 1908 4320 1924 4384
rect 1988 4320 2004 4384
rect 2068 4320 2076 4384
rect 1756 3606 2076 4320
rect 1756 3370 1798 3606
rect 2034 3370 2076 3606
rect 1756 3296 2076 3370
rect 1756 3232 1764 3296
rect 1828 3232 1844 3296
rect 1908 3232 1924 3296
rect 1988 3232 2004 3296
rect 2068 3232 2076 3296
rect 1756 2208 2076 3232
rect 1756 2144 1764 2208
rect 1828 2144 1844 2208
rect 1908 2144 1924 2208
rect 1988 2144 2004 2208
rect 2068 2144 2076 2208
rect 1756 1974 2076 2144
rect 1756 1738 1798 1974
rect 2034 1738 2076 1974
rect 1756 1120 2076 1738
rect 1756 1056 1764 1120
rect 1828 1056 1844 1120
rect 1908 1056 1924 1120
rect 1988 1056 2004 1120
rect 2068 1056 2076 1120
rect 1756 1040 2076 1056
rect 2569 6016 2889 6032
rect 2569 5952 2577 6016
rect 2641 5952 2657 6016
rect 2721 5952 2737 6016
rect 2801 5952 2817 6016
rect 2881 5952 2889 6016
rect 2569 4928 2889 5952
rect 2569 4864 2577 4928
rect 2641 4864 2657 4928
rect 2721 4864 2737 4928
rect 2801 4864 2817 4928
rect 2881 4864 2889 4928
rect 2569 4422 2889 4864
rect 2569 4186 2611 4422
rect 2847 4186 2889 4422
rect 2569 3840 2889 4186
rect 2569 3776 2577 3840
rect 2641 3776 2657 3840
rect 2721 3776 2737 3840
rect 2801 3776 2817 3840
rect 2881 3776 2889 3840
rect 2569 2790 2889 3776
rect 2569 2752 2611 2790
rect 2847 2752 2889 2790
rect 2569 2688 2577 2752
rect 2881 2688 2889 2752
rect 2569 2554 2611 2688
rect 2847 2554 2889 2688
rect 2569 1664 2889 2554
rect 2569 1600 2577 1664
rect 2641 1600 2657 1664
rect 2721 1600 2737 1664
rect 2801 1600 2817 1664
rect 2881 1600 2889 1664
rect 2569 1040 2889 1600
rect 3382 5472 3702 6032
rect 3382 5408 3390 5472
rect 3454 5408 3470 5472
rect 3534 5408 3550 5472
rect 3614 5408 3630 5472
rect 3694 5408 3702 5472
rect 3382 5238 3702 5408
rect 3382 5002 3424 5238
rect 3660 5002 3702 5238
rect 3382 4384 3702 5002
rect 3382 4320 3390 4384
rect 3454 4320 3470 4384
rect 3534 4320 3550 4384
rect 3614 4320 3630 4384
rect 3694 4320 3702 4384
rect 3382 3606 3702 4320
rect 3382 3370 3424 3606
rect 3660 3370 3702 3606
rect 3382 3296 3702 3370
rect 3382 3232 3390 3296
rect 3454 3232 3470 3296
rect 3534 3232 3550 3296
rect 3614 3232 3630 3296
rect 3694 3232 3702 3296
rect 3382 2208 3702 3232
rect 3382 2144 3390 2208
rect 3454 2144 3470 2208
rect 3534 2144 3550 2208
rect 3614 2144 3630 2208
rect 3694 2144 3702 2208
rect 3382 1974 3702 2144
rect 3382 1738 3424 1974
rect 3660 1738 3702 1974
rect 3382 1120 3702 1738
rect 3382 1056 3390 1120
rect 3454 1056 3470 1120
rect 3534 1056 3550 1120
rect 3614 1056 3630 1120
rect 3694 1056 3702 1120
rect 3382 1040 3702 1056
rect 4194 6016 4514 6032
rect 4194 5952 4202 6016
rect 4266 5952 4282 6016
rect 4346 5952 4362 6016
rect 4426 5952 4442 6016
rect 4506 5952 4514 6016
rect 4194 4928 4514 5952
rect 4194 4864 4202 4928
rect 4266 4864 4282 4928
rect 4346 4864 4362 4928
rect 4426 4864 4442 4928
rect 4506 4864 4514 4928
rect 4194 4422 4514 4864
rect 4194 4186 4236 4422
rect 4472 4186 4514 4422
rect 4194 3840 4514 4186
rect 4194 3776 4202 3840
rect 4266 3776 4282 3840
rect 4346 3776 4362 3840
rect 4426 3776 4442 3840
rect 4506 3776 4514 3840
rect 4194 2790 4514 3776
rect 4194 2752 4236 2790
rect 4472 2752 4514 2790
rect 4194 2688 4202 2752
rect 4506 2688 4514 2752
rect 4194 2554 4236 2688
rect 4472 2554 4514 2688
rect 4194 1664 4514 2554
rect 4194 1600 4202 1664
rect 4266 1600 4282 1664
rect 4346 1600 4362 1664
rect 4426 1600 4442 1664
rect 4506 1600 4514 1664
rect 4194 1040 4514 1600
rect 5007 5472 5327 6032
rect 5007 5408 5015 5472
rect 5079 5408 5095 5472
rect 5159 5408 5175 5472
rect 5239 5408 5255 5472
rect 5319 5408 5327 5472
rect 5007 5238 5327 5408
rect 5007 5002 5049 5238
rect 5285 5002 5327 5238
rect 5007 4384 5327 5002
rect 5007 4320 5015 4384
rect 5079 4320 5095 4384
rect 5159 4320 5175 4384
rect 5239 4320 5255 4384
rect 5319 4320 5327 4384
rect 5007 3606 5327 4320
rect 5007 3370 5049 3606
rect 5285 3370 5327 3606
rect 5007 3296 5327 3370
rect 5007 3232 5015 3296
rect 5079 3232 5095 3296
rect 5159 3232 5175 3296
rect 5239 3232 5255 3296
rect 5319 3232 5327 3296
rect 5007 2208 5327 3232
rect 5007 2144 5015 2208
rect 5079 2144 5095 2208
rect 5159 2144 5175 2208
rect 5239 2144 5255 2208
rect 5319 2144 5327 2208
rect 5007 1974 5327 2144
rect 5007 1738 5049 1974
rect 5285 1738 5327 1974
rect 5007 1120 5327 1738
rect 5007 1056 5015 1120
rect 5079 1056 5095 1120
rect 5159 1056 5175 1120
rect 5239 1056 5255 1120
rect 5319 1056 5327 1120
rect 5007 1040 5327 1056
<< via4 >>
rect 1798 5002 2034 5238
rect 1798 3370 2034 3606
rect 1798 1738 2034 1974
rect 2611 4186 2847 4422
rect 2611 2752 2847 2790
rect 2611 2688 2641 2752
rect 2641 2688 2657 2752
rect 2657 2688 2721 2752
rect 2721 2688 2737 2752
rect 2737 2688 2801 2752
rect 2801 2688 2817 2752
rect 2817 2688 2847 2752
rect 2611 2554 2847 2688
rect 3424 5002 3660 5238
rect 3424 3370 3660 3606
rect 3424 1738 3660 1974
rect 4236 4186 4472 4422
rect 4236 2752 4472 2790
rect 4236 2688 4266 2752
rect 4266 2688 4282 2752
rect 4282 2688 4346 2752
rect 4346 2688 4362 2752
rect 4362 2688 4426 2752
rect 4426 2688 4442 2752
rect 4442 2688 4472 2752
rect 4236 2554 4472 2688
rect 5049 5002 5285 5238
rect 5049 3370 5285 3606
rect 5049 1738 5285 1974
<< metal5 >>
rect 1104 5238 5980 5280
rect 1104 5002 1798 5238
rect 2034 5002 3424 5238
rect 3660 5002 5049 5238
rect 5285 5002 5980 5238
rect 1104 4960 5980 5002
rect 1104 4422 5980 4464
rect 1104 4186 2611 4422
rect 2847 4186 4236 4422
rect 4472 4186 5980 4422
rect 1104 4144 5980 4186
rect 1104 3606 5980 3648
rect 1104 3370 1798 3606
rect 2034 3370 3424 3606
rect 3660 3370 5049 3606
rect 5285 3370 5980 3606
rect 1104 3328 5980 3370
rect 1104 2790 5980 2832
rect 1104 2554 2611 2790
rect 2847 2554 4236 2790
rect 4472 2554 5980 2790
rect 1104 2512 5980 2554
rect 1104 1974 5980 2016
rect 1104 1738 1798 1974
rect 2034 1738 3424 1974
rect 3660 1738 5049 1974
rect 5285 1738 5980 1974
rect 1104 1696 5980 1738
use sky130_fd_sc_hd__decap_8  FILLER_0_7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 1748 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21
timestamp 1641350499
transform 1 0 3036 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39
timestamp 1641350499
transform 1 0 4692 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_42
timestamp 1641350499
transform 1 0 4968 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_23
timestamp 1641350499
transform 1 0 3220 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_12
timestamp 1641350499
transform 1 0 2208 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_40
timestamp 1641350499
transform 1 0 4784 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 3312 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_32
timestamp 1641350499
transform 1 0 4048 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_44
timestamp 1641350499
transform 1 0 5152 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_40
timestamp 1641350499
transform 1 0 4784 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1641350499
transform 1 0 1380 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_36
timestamp 1641350499
transform 1 0 4416 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_27
timestamp 1641350499
transform 1 0 3588 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_44
timestamp 1641350499
transform 1 0 5152 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[3\] $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 1380 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[28\]
timestamp 1641350499
transform 1 0 1932 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[27\]
timestamp 1641350499
transform 1 0 1472 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[20\]
timestamp 1641350499
transform 1 0 2760 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[1\]
timestamp 1641350499
transform 1 0 3036 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[11\]
timestamp 1641350499
transform 1 0 2668 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[0\]
timestamp 1641350499
transform 1 0 2392 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[7\]
timestamp 1641350499
transform 1 0 3864 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[15\]
timestamp 1641350499
transform 1 0 4416 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[4\]
timestamp 1641350499
transform 1 0 5428 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[13\]
timestamp 1641350499
transform 1 0 4600 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[9\]
timestamp 1641350499
transform 1 0 4876 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[31\]
timestamp 1641350499
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[24\]
timestamp 1641350499
transform 1 0 1748 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[17\]
timestamp 1641350499
transform 1 0 1472 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[8\]
timestamp 1641350499
transform 1 0 3220 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[25\]
timestamp 1641350499
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[14\]
timestamp 1641350499
transform 1 0 2484 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[22\]
timestamp 1641350499
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[16\]
timestamp 1641350499
transform 1 0 4600 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[26\]
timestamp 1641350499
transform 1 0 5060 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[6\]
timestamp 1641350499
transform 1 0 1380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[2\]
timestamp 1641350499
transform 1 0 1840 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[18\]
timestamp 1641350499
transform 1 0 4508 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[10\]
timestamp 1641350499
transform 1 0 4232 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[29\]
timestamp 1641350499
transform 1 0 5336 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[19\]
timestamp 1641350499
transform 1 0 1932 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[30\]
timestamp 1641350499
transform 1 0 3036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[21\]
timestamp 1641350499
transform 1 0 3404 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[5\]
timestamp 1641350499
transform 1 0 4140 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[12\]
timestamp 1641350499
transform 1 0 4508 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  mask_rev_value\[23\]
timestamp 1641350499
transform 1 0 5060 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 2208 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1641350499
transform 1 0 3772 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_45
timestamp 1641350499
transform 1 0 5244 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_18
timestamp 1641350499
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 1641350499
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_6
timestamp 1641350499
transform 1 0 1656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1641350499
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 4140 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1641350499
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1641350499
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_6
timestamp 1641350499
transform 1 0 1656 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_18
timestamp 1641350499
transform 1 0 2760 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_30
timestamp 1641350499
transform 1 0 3864 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_11
timestamp 1641350499
transform 1 0 2116 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1641350499
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1641350499
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1641350499
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1641350499
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1641350499
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 1380 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_20
timestamp 1641350499
transform 1 0 2944 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1641350499
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_14
timestamp 1641350499
transform 1 0 2392 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_30
timestamp 1641350499
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_49
timestamp 1641350499
transform 1 0 5612 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_24
timestamp 1641350499
transform 1 0 3312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_20
timestamp 1641350499
transform 1 0 2944 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 1641350499
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_42
timestamp 1641350499
transform 1 0 4968 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 1656 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1641350499
transform 1 0 1104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1641350499
transform 1 0 1104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15
timestamp 1641350499
transform 1 0 2484 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47
timestamp 1641350499
transform 1 0 5428 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1641350499
transform -1 0 5980 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1641350499
transform -1 0 5980 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1641350499
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1641350499
transform -1 0 5980 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1641350499
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1641350499
transform -1 0 5980 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1641350499
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_35
timestamp 1641350499
transform 1 0 4324 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1641350499
transform -1 0 5980 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1641350499
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_31
timestamp 1641350499
transform 1 0 3956 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1641350499
transform -1 0 5980 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1641350499
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1641350499
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_28
timestamp 1641350499
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1641350499
transform -1 0 5980 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1641350499
transform -1 0 5980 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1641350499
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1641350499
transform -1 0 5980 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 3956 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_19
timestamp 1641350499
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_20
timestamp 1641350499
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_21
timestamp 1641350499
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_22
timestamp 1641350499
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1641350499
transform 1 0 4048 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1641350499
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1641350499
transform 1 0 2024 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_26
timestamp 1641350499
transform 1 0 3496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_46
timestamp 1641350499
transform 1 0 5336 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1641350499
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_46
timestamp 1641350499
transform 1 0 5336 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1641350499
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
<< labels >>
rlabel metal2 s 4066 6277 4122 7077 4 mask_rev[0]
port 1 nsew
rlabel metal2 s 4066 0 4122 800 4 mask_rev[10]
port 2 nsew
rlabel metal2 s 1122 0 1178 800 4 mask_rev[11]
port 3 nsew
rlabel metal2 s 570 0 626 800 4 mask_rev[12]
port 4 nsew
rlabel metal2 s 5354 6277 5410 7077 4 mask_rev[13]
port 5 nsew
rlabel metal2 s 5906 0 5962 800 4 mask_rev[14]
port 6 nsew
rlabel metal3 s 6309 1640 7109 1760 4 mask_rev[15]
port 7 nsew
rlabel metal2 s 2226 0 2282 800 4 mask_rev[16]
port 8 nsew
rlabel metal2 s 1674 6277 1730 7077 4 mask_rev[17]
port 9 nsew
rlabel metal3 s 0 5176 800 5296 4 mask_rev[18]
port 10 nsew
rlabel metal2 s 2962 6277 3018 7077 4 mask_rev[19]
port 11 nsew
rlabel metal3 s 0 3272 800 3392 4 mask_rev[1]
port 12 nsew
rlabel metal3 s 6309 2456 7109 2576 4 mask_rev[20]
port 13 nsew
rlabel metal3 s 6309 824 7109 944 4 mask_rev[21]
port 14 nsew
rlabel metal3 s 0 5992 800 6112 4 mask_rev[22]
port 15 nsew
rlabel metal2 s 1674 0 1730 800 4 mask_rev[23]
port 16 nsew
rlabel metal2 s 5906 6277 5962 7077 4 mask_rev[24]
port 17 nsew
rlabel metal3 s 0 1640 800 1760 4 mask_rev[25]
port 18 nsew
rlabel metal2 s 4802 6277 4858 7077 4 mask_rev[26]
port 19 nsew
rlabel metal2 s 1122 6277 1178 7077 4 mask_rev[27]
port 20 nsew
rlabel metal2 s 6458 6277 6514 7077 4 mask_rev[28]
port 21 nsew
rlabel metal2 s 5354 0 5410 800 4 mask_rev[29]
port 22 nsew
rlabel metal3 s 0 2456 800 2576 4 mask_rev[2]
port 23 nsew
rlabel metal3 s 6309 5176 7109 5296 4 mask_rev[30]
port 24 nsew
rlabel metal2 s 2962 0 3018 800 4 mask_rev[31]
port 25 nsew
rlabel metal2 s 3514 0 3570 800 4 mask_rev[3]
port 26 nsew
rlabel metal3 s 6309 3544 7109 3664 4 mask_rev[4]
port 27 nsew
rlabel metal3 s 6309 4360 7109 4480 4 mask_rev[5]
port 28 nsew
rlabel metal3 s 0 4360 800 4480 4 mask_rev[6]
port 29 nsew
rlabel metal2 s 3514 6277 3570 7077 4 mask_rev[7]
port 30 nsew
rlabel metal2 s 4802 0 4858 800 4 mask_rev[8]
port 31 nsew
rlabel metal2 s 2226 6277 2282 7077 4 mask_rev[9]
port 32 nsew
rlabel metal5 s 1104 1696 5980 2016 4 VPWR
port 33 nsew
rlabel metal5 s 1104 2512 5980 2832 4 VGND
port 34 nsew
<< properties >>
string FIXED_BBOX 0 0 7109 7077
string GDS_FILE ../gds/user_id_programming.gds
string GDS_START 0
<< end >>
