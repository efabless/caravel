magic
tech sky130A
magscale 1 2
timestamp 1666198072
<< metal1 >>
rect 132494 1001920 132500 1001972
rect 132552 1001960 132558 1001972
rect 133690 1001960 133696 1001972
rect 132552 1001932 133696 1001960
rect 132552 1001920 132558 1001932
rect 133690 1001920 133696 1001932
rect 133748 1001920 133754 1001972
rect 401686 992196 401692 992248
rect 401744 992236 401750 992248
rect 404354 992236 404360 992248
rect 401744 992208 404360 992236
rect 401744 992196 401750 992208
rect 404354 992196 404360 992208
rect 404412 992196 404418 992248
rect 396074 990836 396080 990888
rect 396132 990876 396138 990888
rect 400214 990876 400220 990888
rect 396132 990848 400220 990876
rect 396132 990836 396138 990848
rect 400214 990836 400220 990848
rect 400272 990836 400278 990888
rect 242250 989068 242256 989120
rect 242308 989108 242314 989120
rect 245654 989108 245660 989120
rect 242308 989080 245660 989108
rect 242308 989068 242314 989080
rect 245654 989068 245660 989080
rect 245712 989068 245718 989120
rect 293954 988184 293960 988236
rect 294012 988224 294018 988236
rect 298094 988224 298100 988236
rect 294012 988196 298100 988224
rect 294012 988184 294018 988196
rect 298094 988184 298100 988196
rect 298152 988184 298158 988236
rect 389174 987504 389180 987556
rect 389232 987544 389238 987556
rect 391934 987544 391940 987556
rect 389232 987516 391940 987544
rect 389232 987504 389238 987516
rect 391934 987504 391940 987516
rect 391992 987504 391998 987556
rect 399754 986348 399760 986400
rect 399812 986388 399818 986400
rect 401686 986388 401692 986400
rect 399812 986360 401692 986388
rect 399812 986348 399818 986360
rect 401686 986348 401692 986360
rect 401744 986348 401750 986400
rect 238662 985940 238668 985992
rect 238720 985980 238726 985992
rect 242250 985980 242256 985992
rect 238720 985952 242256 985980
rect 238720 985940 238726 985952
rect 242250 985940 242256 985952
rect 242308 985940 242314 985992
rect 289722 985396 289728 985448
rect 289780 985436 289786 985448
rect 293954 985436 293960 985448
rect 289780 985408 293960 985436
rect 289780 985396 289786 985408
rect 293954 985396 293960 985408
rect 294012 985396 294018 985448
rect 394418 983492 394424 983544
rect 394476 983532 394482 983544
rect 396074 983532 396080 983544
rect 394476 983504 396080 983532
rect 394476 983492 394482 983504
rect 396074 983492 396080 983504
rect 396132 983492 396138 983544
rect 483014 982472 483020 982524
rect 483072 982512 483078 982524
rect 483842 982512 483848 982524
rect 483072 982484 483848 982512
rect 483072 982472 483078 982484
rect 483842 982472 483848 982484
rect 483900 982472 483906 982524
rect 651374 959080 651380 959132
rect 651432 959120 651438 959132
rect 677410 959120 677416 959132
rect 651432 959092 677416 959120
rect 651432 959080 651438 959092
rect 677410 959080 677416 959092
rect 677468 959080 677474 959132
rect 30098 954932 30104 954984
rect 30156 954972 30162 954984
rect 63402 954972 63408 954984
rect 30156 954944 63408 954972
rect 30156 954932 30162 954944
rect 63402 954932 63408 954944
rect 63460 954932 63466 954984
rect 676030 897104 676036 897116
rect 663766 897076 676036 897104
rect 656158 896996 656164 897048
rect 656216 897036 656222 897048
rect 663766 897036 663794 897076
rect 676030 897064 676036 897076
rect 676088 897064 676094 897116
rect 656216 897008 663794 897036
rect 656216 896996 656222 897008
rect 672718 895772 672724 895824
rect 672776 895812 672782 895824
rect 676030 895812 676036 895824
rect 672776 895784 676036 895812
rect 672776 895772 672782 895784
rect 676030 895772 676036 895784
rect 676088 895772 676094 895824
rect 654778 895636 654784 895688
rect 654836 895676 654842 895688
rect 675846 895676 675852 895688
rect 654836 895648 675852 895676
rect 654836 895636 654842 895648
rect 675846 895636 675852 895648
rect 675904 895636 675910 895688
rect 671890 894412 671896 894464
rect 671948 894452 671954 894464
rect 676030 894452 676036 894464
rect 671948 894424 676036 894452
rect 671948 894412 671954 894424
rect 676030 894412 676036 894424
rect 676088 894412 676094 894464
rect 671062 894276 671068 894328
rect 671120 894316 671126 894328
rect 675846 894316 675852 894328
rect 671120 894288 675852 894316
rect 671120 894276 671126 894288
rect 675846 894276 675852 894288
rect 675904 894276 675910 894328
rect 673270 892984 673276 893036
rect 673328 893024 673334 893036
rect 675846 893024 675852 893036
rect 673328 892996 675852 893024
rect 673328 892984 673334 892996
rect 675846 892984 675852 892996
rect 675904 892984 675910 893036
rect 672258 892848 672264 892900
rect 672316 892888 672322 892900
rect 676030 892888 676036 892900
rect 672316 892860 676036 892888
rect 672316 892848 672322 892860
rect 676030 892848 676036 892860
rect 676088 892848 676094 892900
rect 674834 890332 674840 890384
rect 674892 890372 674898 890384
rect 676030 890372 676036 890384
rect 674892 890344 676036 890372
rect 674892 890332 674898 890344
rect 676030 890332 676036 890344
rect 676088 890332 676094 890384
rect 676214 890128 676220 890180
rect 676272 890168 676278 890180
rect 676858 890168 676864 890180
rect 676272 890140 676864 890168
rect 676272 890128 676278 890140
rect 676858 890128 676864 890140
rect 676916 890128 676922 890180
rect 674374 888904 674380 888956
rect 674432 888944 674438 888956
rect 676030 888944 676036 888956
rect 674432 888916 676036 888944
rect 674432 888904 674438 888916
rect 676030 888904 676036 888916
rect 676088 888904 676094 888956
rect 675018 888700 675024 888752
rect 675076 888740 675082 888752
rect 675846 888740 675852 888752
rect 675076 888712 675852 888740
rect 675076 888700 675082 888712
rect 675846 888700 675852 888712
rect 675904 888700 675910 888752
rect 676214 888700 676220 888752
rect 676272 888740 676278 888752
rect 677042 888740 677048 888752
rect 676272 888712 677048 888740
rect 676272 888700 676278 888712
rect 677042 888700 677048 888712
rect 677100 888700 677106 888752
rect 674650 888496 674656 888548
rect 674708 888536 674714 888548
rect 676030 888536 676036 888548
rect 674708 888508 676036 888536
rect 674708 888496 674714 888508
rect 676030 888496 676036 888508
rect 676088 888496 676094 888548
rect 674190 887272 674196 887324
rect 674248 887312 674254 887324
rect 676030 887312 676036 887324
rect 674248 887284 676036 887312
rect 674248 887272 674254 887284
rect 676030 887272 676036 887284
rect 676088 887272 676094 887324
rect 670878 886864 670884 886916
rect 670936 886904 670942 886916
rect 676030 886904 676036 886916
rect 670936 886876 676036 886904
rect 670936 886864 670942 886876
rect 676030 886864 676036 886876
rect 676088 886864 676094 886916
rect 675570 886592 675576 886644
rect 675628 886632 675634 886644
rect 676398 886632 676404 886644
rect 675628 886604 676404 886632
rect 675628 886592 675634 886604
rect 676398 886592 676404 886604
rect 676456 886592 676462 886644
rect 653398 880472 653404 880524
rect 653456 880512 653462 880524
rect 667290 880512 667296 880524
rect 653456 880484 667296 880512
rect 653456 880472 653462 880484
rect 667290 880472 667296 880484
rect 667348 880472 667354 880524
rect 679618 880444 679624 880456
rect 676186 880416 679624 880444
rect 675386 880336 675392 880388
rect 675444 880376 675450 880388
rect 676186 880376 676214 880416
rect 679618 880404 679624 880416
rect 679676 880404 679682 880456
rect 675444 880348 676214 880376
rect 675444 880336 675450 880348
rect 667290 879588 667296 879640
rect 667348 879628 667354 879640
rect 675570 879628 675576 879640
rect 667348 879600 675576 879628
rect 667348 879588 667354 879600
rect 675570 879588 675576 879600
rect 675628 879588 675634 879640
rect 675754 879316 675760 879368
rect 675812 879356 675818 879368
rect 676858 879356 676864 879368
rect 675812 879328 676864 879356
rect 675812 879316 675818 879328
rect 676858 879316 676864 879328
rect 676916 879316 676922 879368
rect 675938 879180 675944 879232
rect 675996 879220 676002 879232
rect 678238 879220 678244 879232
rect 675996 879192 678244 879220
rect 675996 879180 676002 879192
rect 678238 879180 678244 879192
rect 678296 879180 678302 879232
rect 677042 879084 677048 879096
rect 675128 879056 677048 879084
rect 674006 878976 674012 879028
rect 674064 879016 674070 879028
rect 675128 879016 675156 879056
rect 677042 879044 677048 879056
rect 677100 879044 677106 879096
rect 674064 878988 675156 879016
rect 674064 878976 674070 878988
rect 675754 878364 675760 878416
rect 675812 878364 675818 878416
rect 675772 878200 675800 878364
rect 675588 878172 675800 878200
rect 675588 877384 675616 878172
rect 675496 877356 675616 877384
rect 675496 877260 675524 877356
rect 675478 877208 675484 877260
rect 675536 877208 675542 877260
rect 674834 874896 674840 874948
rect 674892 874936 674898 874948
rect 675386 874936 675392 874948
rect 674892 874908 675392 874936
rect 674892 874896 674898 874908
rect 675386 874896 675392 874908
rect 675444 874896 675450 874948
rect 674006 873672 674012 873724
rect 674064 873712 674070 873724
rect 675386 873712 675392 873724
rect 674064 873684 675392 873712
rect 674064 873672 674070 873684
rect 675386 873672 675392 873684
rect 675444 873672 675450 873724
rect 674190 871972 674196 872024
rect 674248 872012 674254 872024
rect 674650 872012 674656 872024
rect 674248 871984 674656 872012
rect 674248 871972 674254 871984
rect 674650 871972 674656 871984
rect 674708 871972 674714 872024
rect 657538 869388 657544 869440
rect 657596 869428 657602 869440
rect 674650 869428 674656 869440
rect 657596 869400 674656 869428
rect 657596 869388 657602 869400
rect 674650 869388 674656 869400
rect 674708 869388 674714 869440
rect 651466 868844 651472 868896
rect 651524 868884 651530 868896
rect 654778 868884 654784 868896
rect 651524 868856 654784 868884
rect 651524 868844 651530 868856
rect 654778 868844 654784 868856
rect 654836 868844 654842 868896
rect 654134 868028 654140 868080
rect 654192 868068 654198 868080
rect 674834 868068 674840 868080
rect 654192 868040 674840 868068
rect 654192 868028 654198 868040
rect 674834 868028 674840 868040
rect 674892 868028 674898 868080
rect 651466 867892 651472 867944
rect 651524 867932 651530 867944
rect 656158 867932 656164 867944
rect 651524 867904 656164 867932
rect 651524 867892 651530 867904
rect 656158 867892 656164 867904
rect 656216 867892 656222 867944
rect 674650 867892 674656 867944
rect 674708 867932 674714 867944
rect 675202 867932 675208 867944
rect 674708 867904 675208 867932
rect 674708 867892 674714 867904
rect 675202 867892 675208 867904
rect 675260 867892 675266 867944
rect 651466 866600 651472 866652
rect 651524 866640 651530 866652
rect 672718 866640 672724 866652
rect 651524 866612 672724 866640
rect 651524 866600 651530 866612
rect 672718 866600 672724 866612
rect 672776 866600 672782 866652
rect 651374 865172 651380 865224
rect 651432 865212 651438 865224
rect 653398 865212 653404 865224
rect 651432 865184 653404 865212
rect 651432 865172 651438 865184
rect 653398 865172 653404 865184
rect 653456 865172 653462 865224
rect 651466 863812 651472 863864
rect 651524 863852 651530 863864
rect 657538 863852 657544 863864
rect 651524 863824 657544 863852
rect 651524 863812 651530 863824
rect 657538 863812 657544 863824
rect 657596 863812 657602 863864
rect 651466 862452 651472 862504
rect 651524 862492 651530 862504
rect 654134 862492 654140 862504
rect 651524 862464 654140 862492
rect 651524 862452 651530 862464
rect 654134 862452 654140 862464
rect 654192 862452 654198 862504
rect 35802 816960 35808 817012
rect 35860 817000 35866 817012
rect 58618 817000 58624 817012
rect 35860 816972 58624 817000
rect 35860 816960 35866 816972
rect 58618 816960 58624 816972
rect 58676 816960 58682 817012
rect 35802 815736 35808 815788
rect 35860 815776 35866 815788
rect 43438 815776 43444 815788
rect 35860 815748 43444 815776
rect 35860 815736 35866 815748
rect 43438 815736 43444 815748
rect 43496 815736 43502 815788
rect 35618 815600 35624 815652
rect 35676 815640 35682 815652
rect 61378 815640 61384 815652
rect 35676 815612 61384 815640
rect 35676 815600 35682 815612
rect 61378 815600 61384 815612
rect 61436 815600 61442 815652
rect 35434 814852 35440 814904
rect 35492 814892 35498 814904
rect 62758 814892 62764 814904
rect 35492 814864 62764 814892
rect 35492 814852 35498 814864
rect 62758 814852 62764 814864
rect 62816 814852 62822 814904
rect 35618 814376 35624 814428
rect 35676 814416 35682 814428
rect 42886 814416 42892 814428
rect 35676 814388 42892 814416
rect 35676 814376 35682 814388
rect 42886 814376 42892 814388
rect 42944 814376 42950 814428
rect 35802 814240 35808 814292
rect 35860 814280 35866 814292
rect 44726 814280 44732 814292
rect 35860 814252 44732 814280
rect 35860 814240 35866 814252
rect 44726 814240 44732 814252
rect 44784 814240 44790 814292
rect 41322 812812 41328 812864
rect 41380 812852 41386 812864
rect 44174 812852 44180 812864
rect 41380 812824 44180 812852
rect 41380 812812 41386 812824
rect 44174 812812 44180 812824
rect 44232 812812 44238 812864
rect 41322 811724 41328 811776
rect 41380 811764 41386 811776
rect 43070 811764 43076 811776
rect 41380 811736 43076 811764
rect 41380 811724 41386 811736
rect 43070 811724 43076 811736
rect 43128 811724 43134 811776
rect 40954 810704 40960 810756
rect 41012 810744 41018 810756
rect 42610 810744 42616 810756
rect 41012 810716 42616 810744
rect 41012 810704 41018 810716
rect 42610 810704 42616 810716
rect 42668 810704 42674 810756
rect 41322 808596 41328 808648
rect 41380 808636 41386 808648
rect 42242 808636 42248 808648
rect 41380 808608 42248 808636
rect 41380 808596 41386 808608
rect 42242 808596 42248 808608
rect 42300 808596 42306 808648
rect 41322 807440 41328 807492
rect 41380 807480 41386 807492
rect 43254 807480 43260 807492
rect 41380 807452 43260 807480
rect 41380 807440 41386 807452
rect 43254 807440 43260 807452
rect 43312 807440 43318 807492
rect 41138 807304 41144 807356
rect 41196 807344 41202 807356
rect 44358 807344 44364 807356
rect 41196 807316 44364 807344
rect 41196 807304 41202 807316
rect 44358 807304 44364 807316
rect 44416 807304 44422 807356
rect 41322 806080 41328 806132
rect 41380 806120 41386 806132
rect 50338 806120 50344 806132
rect 41380 806092 50344 806120
rect 41380 806080 41386 806092
rect 50338 806080 50344 806092
rect 50396 806080 50402 806132
rect 41138 805944 41144 805996
rect 41196 805984 41202 805996
rect 64138 805984 64144 805996
rect 41196 805956 64144 805984
rect 41196 805944 41202 805956
rect 64138 805944 64144 805956
rect 64196 805944 64202 805996
rect 34514 802408 34520 802460
rect 34572 802448 34578 802460
rect 42150 802448 42156 802460
rect 34572 802420 42156 802448
rect 34572 802408 34578 802420
rect 42150 802408 42156 802420
rect 42208 802408 42214 802460
rect 37918 801728 37924 801780
rect 37976 801768 37982 801780
rect 41966 801768 41972 801780
rect 37976 801740 41972 801768
rect 37976 801728 37982 801740
rect 41966 801728 41972 801740
rect 42024 801728 42030 801780
rect 36538 801252 36544 801304
rect 36596 801292 36602 801304
rect 42610 801292 42616 801304
rect 36596 801264 42616 801292
rect 36596 801252 36602 801264
rect 42610 801252 42616 801264
rect 42668 801252 42674 801304
rect 41966 801116 41972 801168
rect 42024 801156 42030 801168
rect 42702 801156 42708 801168
rect 42024 801128 42708 801156
rect 42024 801116 42030 801128
rect 42702 801116 42708 801128
rect 42760 801116 42766 801168
rect 31018 801048 31024 801100
rect 31076 801088 31082 801100
rect 31076 801060 41414 801088
rect 31076 801048 31082 801060
rect 41386 801020 41414 801060
rect 42794 801020 42800 801032
rect 41386 800992 42800 801020
rect 42794 800980 42800 800992
rect 42852 800980 42858 801032
rect 43622 799076 43628 799128
rect 43680 799116 43686 799128
rect 53098 799116 53104 799128
rect 43680 799088 53104 799116
rect 43680 799076 43686 799088
rect 53098 799076 53104 799088
rect 53156 799076 53162 799128
rect 43806 797648 43812 797700
rect 43864 797688 43870 797700
rect 62942 797688 62948 797700
rect 43864 797660 62948 797688
rect 43864 797648 43870 797660
rect 62942 797648 62948 797660
rect 63000 797648 63006 797700
rect 42242 795608 42248 795660
rect 42300 795648 42306 795660
rect 43806 795648 43812 795660
rect 42300 795620 43812 795648
rect 42300 795608 42306 795620
rect 43806 795608 43812 795620
rect 43864 795608 43870 795660
rect 44358 794900 44364 794912
rect 42352 794872 44364 794900
rect 42352 794368 42380 794872
rect 44358 794860 44364 794872
rect 44416 794860 44422 794912
rect 42334 794316 42340 794368
rect 42392 794316 42398 794368
rect 653398 790780 653404 790832
rect 653456 790820 653462 790832
rect 675386 790820 675392 790832
rect 653456 790792 675392 790820
rect 653456 790780 653462 790792
rect 675386 790780 675392 790792
rect 675444 790780 675450 790832
rect 53098 790712 53104 790764
rect 53156 790752 53162 790764
rect 62206 790752 62212 790764
rect 53156 790724 62212 790752
rect 53156 790712 53162 790724
rect 62206 790712 62212 790724
rect 62264 790712 62270 790764
rect 42150 790100 42156 790152
rect 42208 790140 42214 790152
rect 42702 790140 42708 790152
rect 42208 790112 42708 790140
rect 42208 790100 42214 790112
rect 42702 790100 42708 790112
rect 42760 790100 42766 790152
rect 61378 788604 61384 788656
rect 61436 788644 61442 788656
rect 62942 788644 62948 788656
rect 61436 788616 62948 788644
rect 61436 788604 61442 788616
rect 62942 788604 62948 788616
rect 63000 788604 63006 788656
rect 42610 787992 42616 788044
rect 42668 788032 42674 788044
rect 43070 788032 43076 788044
rect 42668 788004 43076 788032
rect 42668 787992 42674 788004
rect 43070 787992 43076 788004
rect 43128 787992 43134 788044
rect 42702 786632 42708 786684
rect 42760 786672 42766 786684
rect 62114 786672 62120 786684
rect 42760 786644 62120 786672
rect 42760 786632 42766 786644
rect 62114 786632 62120 786644
rect 62172 786632 62178 786684
rect 58618 786496 58624 786548
rect 58676 786536 58682 786548
rect 62114 786536 62120 786548
rect 58676 786508 62120 786536
rect 58676 786496 58682 786508
rect 62114 786496 62120 786508
rect 62172 786496 62178 786548
rect 670602 784252 670608 784304
rect 670660 784292 670666 784304
rect 675110 784292 675116 784304
rect 670660 784264 675116 784292
rect 670660 784252 670666 784264
rect 675110 784252 675116 784264
rect 675168 784252 675174 784304
rect 669222 784116 669228 784168
rect 669280 784156 669286 784168
rect 675386 784156 675392 784168
rect 669280 784128 675392 784156
rect 669280 784116 669286 784128
rect 675386 784116 675392 784128
rect 675444 784116 675450 784168
rect 673914 782620 673920 782672
rect 673972 782660 673978 782672
rect 675110 782660 675116 782672
rect 673972 782632 675116 782660
rect 673972 782620 673978 782632
rect 675110 782620 675116 782632
rect 675168 782620 675174 782672
rect 669038 782484 669044 782536
rect 669096 782524 669102 782536
rect 675294 782524 675300 782536
rect 669096 782496 675300 782524
rect 669096 782484 669102 782496
rect 675294 782484 675300 782496
rect 675352 782484 675358 782536
rect 655514 781056 655520 781108
rect 655572 781096 655578 781108
rect 675202 781096 675208 781108
rect 655572 781068 675208 781096
rect 655572 781056 655578 781068
rect 675202 781056 675208 781068
rect 675260 781056 675266 781108
rect 655054 778336 655060 778388
rect 655112 778376 655118 778388
rect 674926 778376 674932 778388
rect 655112 778348 674932 778376
rect 655112 778336 655118 778348
rect 674926 778336 674932 778348
rect 674984 778336 674990 778388
rect 651466 777588 651472 777640
rect 651524 777628 651530 777640
rect 660298 777628 660304 777640
rect 651524 777600 660304 777628
rect 651524 777588 651530 777600
rect 660298 777588 660304 777600
rect 660356 777588 660362 777640
rect 670418 776976 670424 777028
rect 670476 777016 670482 777028
rect 675294 777016 675300 777028
rect 670476 776988 675300 777016
rect 670476 776976 670482 776988
rect 675294 776976 675300 776988
rect 675352 776976 675358 777028
rect 672718 775616 672724 775668
rect 672776 775656 672782 775668
rect 674926 775656 674932 775668
rect 672776 775628 674932 775656
rect 672776 775616 672782 775628
rect 674926 775616 674932 775628
rect 674984 775616 674990 775668
rect 651466 775548 651472 775600
rect 651524 775588 651530 775600
rect 669958 775588 669964 775600
rect 651524 775560 669964 775588
rect 651524 775548 651530 775560
rect 669958 775548 669964 775560
rect 670016 775548 670022 775600
rect 651374 775276 651380 775328
rect 651432 775316 651438 775328
rect 653398 775316 653404 775328
rect 651432 775288 653404 775316
rect 651432 775276 651438 775288
rect 653398 775276 653404 775288
rect 653456 775276 653462 775328
rect 35802 774188 35808 774240
rect 35860 774228 35866 774240
rect 41690 774228 41696 774240
rect 35860 774200 41696 774228
rect 35860 774188 35866 774200
rect 41690 774188 41696 774200
rect 41748 774188 41754 774240
rect 42058 774188 42064 774240
rect 42116 774228 42122 774240
rect 58618 774228 58624 774240
rect 42116 774200 58624 774228
rect 42116 774188 42122 774200
rect 58618 774188 58624 774200
rect 58676 774188 58682 774240
rect 651466 774120 651472 774172
rect 651524 774160 651530 774172
rect 655514 774160 655520 774172
rect 651524 774132 655520 774160
rect 651524 774120 651530 774132
rect 655514 774120 655520 774132
rect 655572 774120 655578 774172
rect 651466 773780 651472 773832
rect 651524 773820 651530 773832
rect 655054 773820 655060 773832
rect 651524 773792 655060 773820
rect 651524 773780 651530 773792
rect 655054 773780 655060 773792
rect 655112 773780 655118 773832
rect 671430 773372 671436 773424
rect 671488 773412 671494 773424
rect 675294 773412 675300 773424
rect 671488 773384 675300 773412
rect 671488 773372 671494 773384
rect 675294 773372 675300 773384
rect 675352 773372 675358 773424
rect 35802 773304 35808 773356
rect 35860 773344 35866 773356
rect 40310 773344 40316 773356
rect 35860 773316 40316 773344
rect 35860 773304 35866 773316
rect 40310 773304 40316 773316
rect 40368 773304 40374 773356
rect 35802 773100 35808 773152
rect 35860 773140 35866 773152
rect 39574 773140 39580 773152
rect 35860 773112 39580 773140
rect 35860 773100 35866 773112
rect 39574 773100 39580 773112
rect 39632 773100 39638 773152
rect 35618 772964 35624 773016
rect 35676 773004 35682 773016
rect 41690 773004 41696 773016
rect 35676 772976 41696 773004
rect 35676 772964 35682 772976
rect 41690 772964 41696 772976
rect 41748 772964 41754 773016
rect 42058 772964 42064 773016
rect 42116 773004 42122 773016
rect 44542 773004 44548 773016
rect 42116 772976 44548 773004
rect 42116 772964 42122 772976
rect 44542 772964 44548 772976
rect 44600 772964 44606 773016
rect 35434 772828 35440 772880
rect 35492 772868 35498 772880
rect 41690 772868 41696 772880
rect 35492 772840 41696 772868
rect 35492 772828 35498 772840
rect 41690 772828 41696 772840
rect 41748 772828 41754 772880
rect 42058 772828 42064 772880
rect 42116 772868 42122 772880
rect 61378 772868 61384 772880
rect 42116 772840 61384 772868
rect 42116 772828 42122 772840
rect 61378 772828 61384 772840
rect 61436 772828 61442 772880
rect 35618 771808 35624 771860
rect 35676 771848 35682 771860
rect 40770 771848 40776 771860
rect 35676 771820 40776 771848
rect 35676 771808 35682 771820
rect 40770 771808 40776 771820
rect 40828 771808 40834 771860
rect 41690 771644 41696 771656
rect 41386 771616 41696 771644
rect 35802 771536 35808 771588
rect 35860 771576 35866 771588
rect 41386 771576 41414 771616
rect 41690 771604 41696 771616
rect 41748 771604 41754 771656
rect 42058 771604 42064 771656
rect 42116 771644 42122 771656
rect 44726 771644 44732 771656
rect 42116 771616 44732 771644
rect 42116 771604 42122 771616
rect 44726 771604 44732 771616
rect 44784 771604 44790 771656
rect 35860 771548 41414 771576
rect 35860 771536 35866 771548
rect 35434 771400 35440 771452
rect 35492 771440 35498 771452
rect 41690 771440 41696 771452
rect 35492 771412 41696 771440
rect 35492 771400 35498 771412
rect 41690 771400 41696 771412
rect 41748 771400 41754 771452
rect 42058 771400 42064 771452
rect 42116 771440 42122 771452
rect 44358 771440 44364 771452
rect 42116 771412 44364 771440
rect 42116 771400 42122 771412
rect 44358 771400 44364 771412
rect 44416 771400 44422 771452
rect 35802 770448 35808 770500
rect 35860 770488 35866 770500
rect 40494 770488 40500 770500
rect 35860 770460 40500 770488
rect 35860 770448 35866 770460
rect 40494 770448 40500 770460
rect 40552 770448 40558 770500
rect 39942 770284 39948 770296
rect 36004 770256 39948 770284
rect 35434 770176 35440 770228
rect 35492 770216 35498 770228
rect 36004 770216 36032 770256
rect 39942 770244 39948 770256
rect 40000 770244 40006 770296
rect 35492 770188 36032 770216
rect 35492 770176 35498 770188
rect 35618 770040 35624 770092
rect 35676 770080 35682 770092
rect 41690 770080 41696 770092
rect 35676 770052 41696 770080
rect 35676 770040 35682 770052
rect 41690 770040 41696 770052
rect 41748 770040 41754 770092
rect 42058 770040 42064 770092
rect 42116 770080 42122 770092
rect 44174 770080 44180 770092
rect 42116 770052 44180 770080
rect 42116 770040 42122 770052
rect 44174 770040 44180 770052
rect 44232 770040 44238 770092
rect 652018 768884 652024 768936
rect 652076 768924 652082 768936
rect 656158 768924 656164 768936
rect 652076 768896 656164 768924
rect 652076 768884 652082 768896
rect 656158 768884 656164 768896
rect 656216 768884 656222 768936
rect 35618 768816 35624 768868
rect 35676 768856 35682 768868
rect 41690 768856 41696 768868
rect 35676 768828 41696 768856
rect 35676 768816 35682 768828
rect 41690 768816 41696 768828
rect 41748 768816 41754 768868
rect 35802 768680 35808 768732
rect 35860 768720 35866 768732
rect 40034 768720 40040 768732
rect 35860 768692 40040 768720
rect 35860 768680 35866 768692
rect 40034 768680 40040 768692
rect 40092 768680 40098 768732
rect 35802 767592 35808 767644
rect 35860 767632 35866 767644
rect 36538 767632 36544 767644
rect 35860 767604 36544 767632
rect 35860 767592 35866 767604
rect 36538 767592 36544 767604
rect 36596 767592 36602 767644
rect 35802 765892 35808 765944
rect 35860 765932 35866 765944
rect 39758 765932 39764 765944
rect 35860 765904 39764 765932
rect 35860 765892 35866 765904
rect 39758 765892 39764 765904
rect 39816 765892 39822 765944
rect 40034 765280 40040 765332
rect 40092 765320 40098 765332
rect 41690 765320 41696 765332
rect 40092 765292 41696 765320
rect 40092 765280 40098 765292
rect 41690 765280 41696 765292
rect 41748 765280 41754 765332
rect 42058 765144 42064 765196
rect 42116 765184 42122 765196
rect 42518 765184 42524 765196
rect 42116 765156 42524 765184
rect 42116 765144 42122 765156
rect 42518 765144 42524 765156
rect 42576 765144 42582 765196
rect 35802 764804 35808 764856
rect 35860 764844 35866 764856
rect 39206 764844 39212 764856
rect 35860 764816 39212 764844
rect 35860 764804 35866 764816
rect 39206 764804 39212 764816
rect 39264 764804 39270 764856
rect 35802 764532 35808 764584
rect 35860 764572 35866 764584
rect 39758 764572 39764 764584
rect 35860 764544 39764 764572
rect 35860 764532 35866 764544
rect 39758 764532 39764 764544
rect 39816 764532 39822 764584
rect 35618 763444 35624 763496
rect 35676 763484 35682 763496
rect 41690 763484 41696 763496
rect 35676 763456 41696 763484
rect 35676 763444 35682 763456
rect 41690 763444 41696 763456
rect 41748 763444 41754 763496
rect 40696 763252 41736 763280
rect 35802 763172 35808 763224
rect 35860 763212 35866 763224
rect 40696 763212 40724 763252
rect 35860 763184 40724 763212
rect 35860 763172 35866 763184
rect 41708 763156 41736 763252
rect 57238 763212 57244 763224
rect 41984 763184 57244 763212
rect 41690 763104 41696 763156
rect 41748 763104 41754 763156
rect 41984 763076 42012 763184
rect 57238 763172 57244 763184
rect 57296 763172 57302 763224
rect 42610 763076 42616 763088
rect 41984 763048 42616 763076
rect 42610 763036 42616 763048
rect 42668 763036 42674 763088
rect 42058 761880 42064 761932
rect 42116 761920 42122 761932
rect 48958 761920 48964 761932
rect 42116 761892 48964 761920
rect 42116 761880 42122 761892
rect 48958 761880 48964 761892
rect 49016 761880 49022 761932
rect 35802 761812 35808 761864
rect 35860 761852 35866 761864
rect 41690 761852 41696 761864
rect 35860 761824 41696 761852
rect 35860 761812 35866 761824
rect 41690 761812 41696 761824
rect 41748 761812 41754 761864
rect 35158 759772 35164 759824
rect 35216 759812 35222 759824
rect 41690 759812 41696 759824
rect 35216 759784 41696 759812
rect 35216 759772 35222 759784
rect 41690 759772 41696 759784
rect 41748 759772 41754 759824
rect 32398 759636 32404 759688
rect 32456 759676 32462 759688
rect 41598 759676 41604 759688
rect 32456 759648 41604 759676
rect 32456 759636 32462 759648
rect 41598 759636 41604 759648
rect 41656 759636 41662 759688
rect 33778 758276 33784 758328
rect 33836 758316 33842 758328
rect 39298 758316 39304 758328
rect 33836 758288 39304 758316
rect 33836 758276 33842 758288
rect 39298 758276 39304 758288
rect 39356 758276 39362 758328
rect 42426 758072 42432 758124
rect 42484 758112 42490 758124
rect 42794 758112 42800 758124
rect 42484 758084 42800 758112
rect 42484 758072 42490 758084
rect 42794 758072 42800 758084
rect 42852 758072 42858 758124
rect 42058 757936 42064 757988
rect 42116 757976 42122 757988
rect 42426 757976 42432 757988
rect 42116 757948 42432 757976
rect 42116 757936 42122 757948
rect 42426 757936 42432 757948
rect 42484 757936 42490 757988
rect 45094 755488 45100 755540
rect 45152 755528 45158 755540
rect 62758 755528 62764 755540
rect 45152 755500 62764 755528
rect 45152 755488 45158 755500
rect 62758 755488 62764 755500
rect 62816 755488 62822 755540
rect 42886 754876 42892 754928
rect 42944 754916 42950 754928
rect 44726 754916 44732 754928
rect 42944 754888 44732 754916
rect 42944 754876 42950 754888
rect 44726 754876 44732 754888
rect 44784 754876 44790 754928
rect 42242 754264 42248 754316
rect 42300 754304 42306 754316
rect 45094 754304 45100 754316
rect 42300 754276 45100 754304
rect 42300 754264 42306 754276
rect 45094 754264 45100 754276
rect 45152 754264 45158 754316
rect 44174 753556 44180 753568
rect 42260 753528 44180 753556
rect 42260 753432 42288 753528
rect 44174 753516 44180 753528
rect 44232 753516 44238 753568
rect 42242 753380 42248 753432
rect 42300 753380 42306 753432
rect 42334 749980 42340 750032
rect 42392 749980 42398 750032
rect 42352 749352 42380 749980
rect 42334 749300 42340 749352
rect 42392 749300 42398 749352
rect 61378 747124 61384 747176
rect 61436 747164 61442 747176
rect 63034 747164 63040 747176
rect 61436 747136 63040 747164
rect 61436 747124 61442 747136
rect 63034 747124 63040 747136
rect 63092 747124 63098 747176
rect 653398 746580 653404 746632
rect 653456 746620 653462 746632
rect 675386 746620 675392 746632
rect 653456 746592 675392 746620
rect 653456 746580 653462 746592
rect 675386 746580 675392 746592
rect 675444 746580 675450 746632
rect 45094 746512 45100 746564
rect 45152 746552 45158 746564
rect 62114 746552 62120 746564
rect 45152 746524 62120 746552
rect 45152 746512 45158 746524
rect 62114 746512 62120 746524
rect 62172 746512 62178 746564
rect 42150 745424 42156 745476
rect 42208 745464 42214 745476
rect 42702 745464 42708 745476
rect 42208 745436 42708 745464
rect 42208 745424 42214 745436
rect 42702 745424 42708 745436
rect 42760 745424 42766 745476
rect 42794 744064 42800 744116
rect 42852 744104 42858 744116
rect 42852 744076 45554 744104
rect 42852 744064 42858 744076
rect 45526 743900 45554 744076
rect 62114 743900 62120 743912
rect 45526 743872 62120 743900
rect 62114 743860 62120 743872
rect 62172 743860 62178 743912
rect 671706 743860 671712 743912
rect 671764 743900 671770 743912
rect 675110 743900 675116 743912
rect 671764 743872 675116 743900
rect 671764 743860 671770 743872
rect 675110 743860 675116 743872
rect 675168 743860 675174 743912
rect 46198 743724 46204 743776
rect 46256 743764 46262 743776
rect 62114 743764 62120 743776
rect 46256 743736 62120 743764
rect 46256 743724 46262 743736
rect 62114 743724 62120 743736
rect 62172 743724 62178 743776
rect 58618 742364 58624 742416
rect 58676 742404 58682 742416
rect 62114 742404 62120 742416
rect 58676 742376 62120 742404
rect 58676 742364 58682 742376
rect 62114 742364 62120 742376
rect 62172 742364 62178 742416
rect 671798 742160 671804 742212
rect 671856 742200 671862 742212
rect 675478 742200 675484 742212
rect 671856 742172 675484 742200
rect 671856 742160 671862 742172
rect 675478 742160 675484 742172
rect 675536 742160 675542 742212
rect 674834 739780 674840 739832
rect 674892 739820 674898 739832
rect 675386 739820 675392 739832
rect 674892 739792 675392 739820
rect 674892 739780 674898 739792
rect 675386 739780 675392 739792
rect 675444 739780 675450 739832
rect 672442 739100 672448 739152
rect 672500 739140 672506 739152
rect 675294 739140 675300 739152
rect 672500 739112 675300 739140
rect 672500 739100 672506 739112
rect 675294 739100 675300 739112
rect 675352 739100 675358 739152
rect 673454 738624 673460 738676
rect 673512 738664 673518 738676
rect 675386 738664 675392 738676
rect 673512 738636 675392 738664
rect 673512 738624 673518 738636
rect 675386 738624 675392 738636
rect 675444 738624 675450 738676
rect 669590 738284 669596 738336
rect 669648 738324 669654 738336
rect 669648 738296 675340 738324
rect 669648 738284 669654 738296
rect 675312 737996 675340 738296
rect 675294 737944 675300 737996
rect 675352 737944 675358 737996
rect 675202 735740 675208 735752
rect 663766 735712 675208 735740
rect 657538 735564 657544 735616
rect 657596 735604 657602 735616
rect 663766 735604 663794 735712
rect 675202 735700 675208 735712
rect 675260 735700 675266 735752
rect 657596 735576 663794 735604
rect 657596 735564 657602 735576
rect 654778 734136 654784 734188
rect 654836 734176 654842 734188
rect 675294 734176 675300 734188
rect 654836 734148 675300 734176
rect 654836 734136 654842 734148
rect 675294 734136 675300 734148
rect 675352 734136 675358 734188
rect 675294 733660 675300 733712
rect 675352 733660 675358 733712
rect 651466 733388 651472 733440
rect 651524 733428 651530 733440
rect 668578 733428 668584 733440
rect 651524 733400 668584 733428
rect 651524 733388 651530 733400
rect 668578 733388 668584 733400
rect 668636 733388 668642 733440
rect 675312 733372 675340 733660
rect 675294 733320 675300 733372
rect 675352 733320 675358 733372
rect 651466 731416 651472 731468
rect 651524 731456 651530 731468
rect 658918 731456 658924 731468
rect 651524 731428 658924 731456
rect 651524 731416 651530 731428
rect 658918 731416 658924 731428
rect 658976 731416 658982 731468
rect 651374 731076 651380 731128
rect 651432 731116 651438 731128
rect 653398 731116 653404 731128
rect 651432 731088 653404 731116
rect 651432 731076 651438 731088
rect 653398 731076 653404 731088
rect 653456 731076 653462 731128
rect 652662 730668 652668 730720
rect 652720 730708 652726 730720
rect 661678 730708 661684 730720
rect 652720 730680 661684 730708
rect 652720 730668 652726 730680
rect 661678 730668 661684 730680
rect 661736 730668 661742 730720
rect 673822 730464 673828 730516
rect 673880 730504 673886 730516
rect 674650 730504 674656 730516
rect 673880 730476 674656 730504
rect 673880 730464 673886 730476
rect 674650 730464 674656 730476
rect 674708 730464 674714 730516
rect 675294 730464 675300 730516
rect 675352 730464 675358 730516
rect 43622 730328 43628 730380
rect 43680 730368 43686 730380
rect 58618 730368 58624 730380
rect 43680 730340 58624 730368
rect 43680 730328 43686 730340
rect 58618 730328 58624 730340
rect 58676 730328 58682 730380
rect 651466 729988 651472 730040
rect 651524 730028 651530 730040
rect 657538 730028 657544 730040
rect 651524 730000 657544 730028
rect 651524 729988 651530 730000
rect 657538 729988 657544 730000
rect 657596 729988 657602 730040
rect 675018 729852 675024 729904
rect 675076 729892 675082 729904
rect 675312 729892 675340 730464
rect 675076 729864 675340 729892
rect 675076 729852 675082 729864
rect 42426 729308 42432 729360
rect 42484 729348 42490 729360
rect 62758 729348 62764 729360
rect 42484 729320 62764 729348
rect 42484 729308 42490 729320
rect 62758 729308 62764 729320
rect 62816 729308 62822 729360
rect 41322 728764 41328 728816
rect 41380 728804 41386 728816
rect 41690 728804 41696 728816
rect 41380 728776 41696 728804
rect 41380 728764 41386 728776
rect 41690 728764 41696 728776
rect 41748 728764 41754 728816
rect 42058 728764 42064 728816
rect 42116 728804 42122 728816
rect 44358 728804 44364 728816
rect 42116 728776 44364 728804
rect 42116 728764 42122 728776
rect 44358 728764 44364 728776
rect 44416 728764 44422 728816
rect 41322 728628 41328 728680
rect 41380 728668 41386 728680
rect 41690 728668 41696 728680
rect 41380 728640 41696 728668
rect 41380 728628 41386 728640
rect 41690 728628 41696 728640
rect 41748 728628 41754 728680
rect 42058 728628 42064 728680
rect 42116 728668 42122 728680
rect 44542 728668 44548 728680
rect 42116 728640 44548 728668
rect 42116 728628 42122 728640
rect 44542 728628 44548 728640
rect 44600 728628 44606 728680
rect 651466 728492 651472 728544
rect 651524 728532 651530 728544
rect 654778 728532 654784 728544
rect 651524 728504 654784 728532
rect 651524 728492 651530 728504
rect 654778 728492 654784 728504
rect 654836 728492 654842 728544
rect 673086 728288 673092 728340
rect 673144 728328 673150 728340
rect 673144 728300 674176 728328
rect 673144 728288 673150 728300
rect 670878 728084 670884 728136
rect 670936 728124 670942 728136
rect 670936 728096 674058 728124
rect 670936 728084 670942 728096
rect 40678 727404 40684 727456
rect 40736 727444 40742 727456
rect 41690 727444 41696 727456
rect 40736 727416 41696 727444
rect 40736 727404 40742 727416
rect 41690 727404 41696 727416
rect 41748 727404 41754 727456
rect 42058 727404 42064 727456
rect 42116 727444 42122 727456
rect 43438 727444 43444 727456
rect 42116 727416 43444 727444
rect 42116 727404 42122 727416
rect 43438 727404 43444 727416
rect 43496 727404 43502 727456
rect 40862 727268 40868 727320
rect 40920 727308 40926 727320
rect 41690 727308 41696 727320
rect 40920 727280 41696 727308
rect 40920 727268 40926 727280
rect 41690 727268 41696 727280
rect 41748 727268 41754 727320
rect 42058 727268 42064 727320
rect 42116 727308 42122 727320
rect 43438 727308 43444 727320
rect 42116 727280 43444 727308
rect 42116 727268 42122 727280
rect 43438 727268 43444 727280
rect 43496 727268 43502 727320
rect 674742 727200 674748 727252
rect 674800 727240 674806 727252
rect 680998 727240 681004 727252
rect 674800 727212 681004 727240
rect 674800 727200 674806 727212
rect 680998 727200 681004 727212
rect 681056 727200 681062 727252
rect 674466 726656 674472 726708
rect 674524 726696 674530 726708
rect 684126 726696 684132 726708
rect 674524 726668 684132 726696
rect 674524 726656 674530 726668
rect 684126 726656 684132 726668
rect 684184 726656 684190 726708
rect 674282 726452 674288 726504
rect 674340 726492 674346 726504
rect 674340 726464 674834 726492
rect 674340 726452 674346 726464
rect 674806 726424 674834 726464
rect 683482 726424 683488 726436
rect 674806 726396 683488 726424
rect 683482 726384 683488 726396
rect 683540 726384 683546 726436
rect 41138 726044 41144 726096
rect 41196 726084 41202 726096
rect 41598 726084 41604 726096
rect 41196 726056 41604 726084
rect 41196 726044 41202 726056
rect 41598 726044 41604 726056
rect 41656 726044 41662 726096
rect 40954 725908 40960 725960
rect 41012 725948 41018 725960
rect 41414 725948 41420 725960
rect 41012 725920 41420 725948
rect 41012 725908 41018 725920
rect 41414 725908 41420 725920
rect 41472 725908 41478 725960
rect 673822 724384 673828 724396
rect 673380 724356 673828 724384
rect 673380 724260 673408 724356
rect 673822 724344 673828 724356
rect 673880 724344 673886 724396
rect 673362 724208 673368 724260
rect 673420 724208 673426 724260
rect 675294 721692 675300 721744
rect 675352 721692 675358 721744
rect 675312 721268 675340 721692
rect 675294 721216 675300 721268
rect 675352 721216 675358 721268
rect 675294 720808 675300 720860
rect 675352 720808 675358 720860
rect 675312 720520 675340 720808
rect 675294 720468 675300 720520
rect 675352 720468 675358 720520
rect 42794 718972 42800 719024
rect 42852 719012 42858 719024
rect 61378 719012 61384 719024
rect 42852 718984 61384 719012
rect 42852 718972 42858 718984
rect 61378 718972 61384 718984
rect 61436 718972 61442 719024
rect 32398 716864 32404 716916
rect 32456 716904 32462 716916
rect 40218 716904 40224 716916
rect 32456 716876 40224 716904
rect 32456 716864 32462 716876
rect 40218 716864 40224 716876
rect 40276 716864 40282 716916
rect 674282 716456 674288 716508
rect 674340 716496 674346 716508
rect 676030 716496 676036 716508
rect 674340 716468 676036 716496
rect 674340 716456 674346 716468
rect 676030 716456 676036 716468
rect 676088 716456 676094 716508
rect 656158 716252 656164 716304
rect 656216 716292 656222 716304
rect 674006 716292 674012 716304
rect 656216 716264 674012 716292
rect 656216 716252 656222 716264
rect 674006 716252 674012 716264
rect 674064 716252 674070 716304
rect 669958 715708 669964 715760
rect 670016 715748 670022 715760
rect 674006 715748 674012 715760
rect 670016 715720 674012 715748
rect 670016 715708 670022 715720
rect 674006 715708 674012 715720
rect 674064 715708 674070 715760
rect 35158 715640 35164 715692
rect 35216 715680 35222 715692
rect 41506 715680 41512 715692
rect 35216 715652 41512 715680
rect 35216 715640 35222 715652
rect 41506 715640 41512 715652
rect 41564 715640 41570 715692
rect 31662 715504 31668 715556
rect 31720 715544 31726 715556
rect 40586 715544 40592 715556
rect 31720 715516 40592 715544
rect 31720 715504 31726 715516
rect 40586 715504 40592 715516
rect 40644 715504 40650 715556
rect 671062 715436 671068 715488
rect 671120 715476 671126 715488
rect 674006 715476 674012 715488
rect 671120 715448 674012 715476
rect 671120 715436 671126 715448
rect 674006 715436 674012 715448
rect 674064 715436 674070 715488
rect 674282 715436 674288 715488
rect 674340 715476 674346 715488
rect 675846 715476 675852 715488
rect 674340 715448 675852 715476
rect 674340 715436 674346 715448
rect 675846 715436 675852 715448
rect 675904 715436 675910 715488
rect 674282 715300 674288 715352
rect 674340 715340 674346 715352
rect 676030 715340 676036 715352
rect 674340 715312 676036 715340
rect 674340 715300 674346 715312
rect 676030 715300 676036 715312
rect 676088 715300 676094 715352
rect 42058 715028 42064 715080
rect 42116 715068 42122 715080
rect 42426 715068 42432 715080
rect 42116 715040 42432 715068
rect 42116 715028 42122 715040
rect 42426 715028 42432 715040
rect 42484 715028 42490 715080
rect 674006 714932 674012 714944
rect 663766 714904 674012 714932
rect 660298 714824 660304 714876
rect 660356 714864 660362 714876
rect 663766 714864 663794 714904
rect 674006 714892 674012 714904
rect 674064 714892 674070 714944
rect 660356 714836 663794 714864
rect 660356 714824 660362 714836
rect 39298 714756 39304 714808
rect 39356 714796 39362 714808
rect 41690 714796 41696 714808
rect 39356 714768 41696 714796
rect 39356 714756 39362 714768
rect 41690 714756 41696 714768
rect 41748 714756 41754 714808
rect 671890 714484 671896 714536
rect 671948 714524 671954 714536
rect 674006 714524 674012 714536
rect 671948 714496 674012 714524
rect 671948 714484 671954 714496
rect 674006 714484 674012 714496
rect 674064 714484 674070 714536
rect 671062 713192 671068 713244
rect 671120 713232 671126 713244
rect 674006 713232 674012 713244
rect 671120 713204 674012 713232
rect 671120 713192 671126 713204
rect 674006 713192 674012 713204
rect 674064 713192 674070 713244
rect 672258 712852 672264 712904
rect 672316 712892 672322 712904
rect 674006 712892 674012 712904
rect 672316 712864 674012 712892
rect 672316 712852 672322 712864
rect 674006 712852 674012 712864
rect 674064 712852 674070 712904
rect 671890 712376 671896 712428
rect 671948 712416 671954 712428
rect 674006 712416 674012 712428
rect 671948 712388 674012 712416
rect 671948 712376 671954 712388
rect 674006 712376 674012 712388
rect 674064 712376 674070 712428
rect 43806 712240 43812 712292
rect 43864 712280 43870 712292
rect 51718 712280 51724 712292
rect 43864 712252 51724 712280
rect 43864 712240 43870 712252
rect 51718 712240 51724 712252
rect 51776 712240 51782 712292
rect 42334 711084 42340 711136
rect 42392 711124 42398 711136
rect 43806 711124 43812 711136
rect 42392 711096 43812 711124
rect 42392 711084 42398 711096
rect 43806 711084 43812 711096
rect 43864 711084 43870 711136
rect 43806 710948 43812 711000
rect 43864 710988 43870 711000
rect 44726 710988 44732 711000
rect 43864 710960 44732 710988
rect 43864 710948 43870 710960
rect 44726 710948 44732 710960
rect 44784 710948 44790 711000
rect 42334 710404 42340 710456
rect 42392 710444 42398 710456
rect 42794 710444 42800 710456
rect 42392 710416 42800 710444
rect 42392 710404 42398 710416
rect 42794 710404 42800 710416
rect 42852 710404 42858 710456
rect 671430 709996 671436 710048
rect 671488 710036 671494 710048
rect 674006 710036 674012 710048
rect 671488 710008 674012 710036
rect 671488 709996 671494 710008
rect 674006 709996 674012 710008
rect 674064 709996 674070 710048
rect 674282 709452 674288 709504
rect 674340 709492 674346 709504
rect 676030 709492 676036 709504
rect 674340 709464 676036 709492
rect 674340 709452 674346 709464
rect 676030 709452 676036 709464
rect 676088 709452 676094 709504
rect 669038 709316 669044 709368
rect 669096 709356 669102 709368
rect 674006 709356 674012 709368
rect 669096 709328 674012 709356
rect 669096 709316 669102 709328
rect 674006 709316 674012 709328
rect 674064 709316 674070 709368
rect 670602 709180 670608 709232
rect 670660 709220 670666 709232
rect 674006 709220 674012 709232
rect 670660 709192 674012 709220
rect 670660 709180 670666 709192
rect 674006 709180 674012 709192
rect 674064 709180 674070 709232
rect 674650 707548 674656 707600
rect 674708 707588 674714 707600
rect 676030 707588 676036 707600
rect 674708 707560 676036 707588
rect 674708 707548 674714 707560
rect 676030 707548 676036 707560
rect 676088 707548 676094 707600
rect 670418 705916 670424 705968
rect 670476 705956 670482 705968
rect 674006 705956 674012 705968
rect 670476 705928 674012 705956
rect 670476 705916 670482 705928
rect 674006 705916 674012 705928
rect 674064 705916 674070 705968
rect 674282 705780 674288 705832
rect 674340 705820 674346 705832
rect 676030 705820 676036 705832
rect 674340 705792 676036 705820
rect 674340 705780 674346 705792
rect 676030 705780 676036 705792
rect 676088 705780 676094 705832
rect 674466 705304 674472 705356
rect 674524 705344 674530 705356
rect 683114 705344 683120 705356
rect 674524 705316 683120 705344
rect 674524 705304 674530 705316
rect 683114 705304 683120 705316
rect 683172 705304 683178 705356
rect 669222 705168 669228 705220
rect 669280 705208 669286 705220
rect 674006 705208 674012 705220
rect 669280 705180 674012 705208
rect 669280 705168 669286 705180
rect 674006 705168 674012 705180
rect 674064 705168 674070 705220
rect 51718 705100 51724 705152
rect 51776 705140 51782 705152
rect 62114 705140 62120 705152
rect 51776 705112 62120 705140
rect 51776 705100 51782 705112
rect 62114 705100 62120 705112
rect 62172 705100 62178 705152
rect 674282 704012 674288 704064
rect 674340 704052 674346 704064
rect 676030 704052 676036 704064
rect 674340 704024 676036 704052
rect 674340 704012 674346 704024
rect 676030 704012 676036 704024
rect 676088 704012 676094 704064
rect 667842 703808 667848 703860
rect 667900 703848 667906 703860
rect 674006 703848 674012 703860
rect 667900 703820 674012 703848
rect 667900 703808 667906 703820
rect 674006 703808 674012 703820
rect 674064 703808 674070 703860
rect 44726 703740 44732 703792
rect 44784 703780 44790 703792
rect 62114 703780 62120 703792
rect 44784 703752 62120 703780
rect 44784 703740 44790 703752
rect 62114 703740 62120 703752
rect 62172 703740 62178 703792
rect 654778 701156 654784 701208
rect 654836 701196 654842 701208
rect 674006 701196 674012 701208
rect 654836 701168 674012 701196
rect 654836 701156 654842 701168
rect 674006 701156 674012 701168
rect 674064 701156 674070 701208
rect 674282 701088 674288 701140
rect 674340 701128 674346 701140
rect 675386 701128 675392 701140
rect 674340 701100 675392 701128
rect 674340 701088 674346 701100
rect 675386 701088 675392 701100
rect 675444 701088 675450 701140
rect 42794 701020 42800 701072
rect 42852 701060 42858 701072
rect 62206 701060 62212 701072
rect 42852 701032 62212 701060
rect 42852 701020 42858 701032
rect 62206 701020 62212 701032
rect 62264 701020 62270 701072
rect 666462 701020 666468 701072
rect 666520 701060 666526 701072
rect 674006 701060 674012 701072
rect 666520 701032 674012 701060
rect 666520 701020 666526 701032
rect 674006 701020 674012 701032
rect 674064 701020 674070 701072
rect 46198 700272 46204 700324
rect 46256 700312 46262 700324
rect 62114 700312 62120 700324
rect 46256 700284 62120 700312
rect 46256 700272 46262 700284
rect 62114 700272 62120 700284
rect 62172 700272 62178 700324
rect 58618 699524 58624 699576
rect 58676 699564 58682 699576
rect 62298 699564 62304 699576
rect 58676 699536 62304 699564
rect 58676 699524 58682 699536
rect 62298 699524 62304 699536
rect 62356 699524 62362 699576
rect 666278 696940 666284 696992
rect 666336 696980 666342 696992
rect 674006 696980 674012 696992
rect 666336 696952 674012 696980
rect 666336 696940 666342 696952
rect 674006 696940 674012 696952
rect 674064 696940 674070 696992
rect 674282 696940 674288 696992
rect 674340 696980 674346 696992
rect 675110 696980 675116 696992
rect 674340 696952 675116 696980
rect 674340 696940 674346 696952
rect 675110 696940 675116 696952
rect 675168 696940 675174 696992
rect 674282 693132 674288 693184
rect 674340 693172 674346 693184
rect 675110 693172 675116 693184
rect 674340 693144 675116 693172
rect 674340 693132 674346 693144
rect 675110 693132 675116 693144
rect 675168 693132 675174 693184
rect 668946 693064 668952 693116
rect 669004 693104 669010 693116
rect 674006 693104 674012 693116
rect 669004 693076 674012 693104
rect 669004 693064 669010 693076
rect 674006 693064 674012 693076
rect 674064 693064 674070 693116
rect 674282 692996 674288 693048
rect 674340 693036 674346 693048
rect 675386 693036 675392 693048
rect 674340 693008 675392 693036
rect 674340 692996 674346 693008
rect 675386 692996 675392 693008
rect 675444 692996 675450 693048
rect 656434 690072 656440 690124
rect 656492 690112 656498 690124
rect 674006 690112 674012 690124
rect 656492 690084 674012 690112
rect 656492 690072 656498 690084
rect 674006 690072 674012 690084
rect 674064 690072 674070 690124
rect 674466 690004 674472 690056
rect 674524 690044 674530 690056
rect 675110 690044 675116 690056
rect 674524 690016 675116 690044
rect 674524 690004 674530 690016
rect 675110 690004 675116 690016
rect 675168 690004 675174 690056
rect 674742 688984 674748 689036
rect 674800 689024 674806 689036
rect 675202 689024 675208 689036
rect 674800 688996 675208 689024
rect 674800 688984 674806 688996
rect 675202 688984 675208 688996
rect 675260 688984 675266 689036
rect 652754 688780 652760 688832
rect 652812 688820 652818 688832
rect 674006 688820 674012 688832
rect 652812 688792 674012 688820
rect 652812 688780 652818 688792
rect 674006 688780 674012 688792
rect 674064 688780 674070 688832
rect 651466 688644 651472 688696
rect 651524 688684 651530 688696
rect 657538 688684 657544 688696
rect 651524 688656 657544 688684
rect 651524 688644 651530 688656
rect 657538 688644 657544 688656
rect 657596 688644 657602 688696
rect 35802 687488 35808 687540
rect 35860 687528 35866 687540
rect 41690 687528 41696 687540
rect 35860 687500 41696 687528
rect 35860 687488 35866 687500
rect 41690 687488 41696 687500
rect 41748 687488 41754 687540
rect 35434 687216 35440 687268
rect 35492 687256 35498 687268
rect 35492 687228 38654 687256
rect 35492 687216 35498 687228
rect 38626 687188 38654 687228
rect 651466 687216 651472 687268
rect 651524 687256 651530 687268
rect 669958 687256 669964 687268
rect 651524 687228 669964 687256
rect 651524 687216 651530 687228
rect 669958 687216 669964 687228
rect 670016 687216 670022 687268
rect 41690 687188 41696 687200
rect 38626 687160 41696 687188
rect 41690 687148 41696 687160
rect 41748 687148 41754 687200
rect 651466 687012 651472 687064
rect 651524 687052 651530 687064
rect 654778 687052 654784 687064
rect 651524 687024 654784 687052
rect 651524 687012 651530 687024
rect 654778 687012 654784 687024
rect 654836 687012 654842 687064
rect 42058 686468 42064 686520
rect 42116 686508 42122 686520
rect 63402 686508 63408 686520
rect 42116 686480 63408 686508
rect 42116 686468 42122 686480
rect 63402 686468 63408 686480
rect 63460 686468 63466 686520
rect 651650 686468 651656 686520
rect 651708 686508 651714 686520
rect 667198 686508 667204 686520
rect 651708 686480 667204 686508
rect 651708 686468 651714 686480
rect 667198 686468 667204 686480
rect 667256 686468 667262 686520
rect 35618 686400 35624 686452
rect 35676 686440 35682 686452
rect 41690 686440 41696 686452
rect 35676 686412 41696 686440
rect 35676 686400 35682 686412
rect 41690 686400 41696 686412
rect 41748 686400 41754 686452
rect 35802 686264 35808 686316
rect 35860 686304 35866 686316
rect 41690 686304 41696 686316
rect 35860 686276 41696 686304
rect 35860 686264 35866 686276
rect 41690 686264 41696 686276
rect 41748 686264 41754 686316
rect 42058 686264 42064 686316
rect 42116 686304 42122 686316
rect 43806 686304 43812 686316
rect 42116 686276 43812 686304
rect 42116 686264 42122 686276
rect 43806 686264 43812 686276
rect 43864 686264 43870 686316
rect 42058 686060 42064 686112
rect 42116 686100 42122 686112
rect 44542 686100 44548 686112
rect 42116 686072 44548 686100
rect 42116 686060 42122 686072
rect 44542 686060 44548 686072
rect 44600 686060 44606 686112
rect 35802 685992 35808 686044
rect 35860 686032 35866 686044
rect 41690 686032 41696 686044
rect 35860 686004 41696 686032
rect 35860 685992 35866 686004
rect 41690 685992 41696 686004
rect 41748 685992 41754 686044
rect 670878 685924 670884 685976
rect 670936 685964 670942 685976
rect 672994 685964 673000 685976
rect 670936 685936 673000 685964
rect 670936 685924 670942 685936
rect 672994 685924 673000 685936
rect 673052 685924 673058 685976
rect 35434 685856 35440 685908
rect 35492 685896 35498 685908
rect 41690 685896 41696 685908
rect 35492 685868 41696 685896
rect 35492 685856 35498 685868
rect 41690 685856 41696 685868
rect 41748 685856 41754 685908
rect 42058 685856 42064 685908
rect 42116 685896 42122 685908
rect 44266 685896 44272 685908
rect 42116 685868 44272 685896
rect 42116 685856 42122 685868
rect 44266 685856 44272 685868
rect 44324 685856 44330 685908
rect 651466 685516 651472 685568
rect 651524 685556 651530 685568
rect 656434 685556 656440 685568
rect 651524 685528 656440 685556
rect 651524 685516 651530 685528
rect 656434 685516 656440 685528
rect 656492 685516 656498 685568
rect 35802 684972 35808 685024
rect 35860 685012 35866 685024
rect 35860 684972 35894 685012
rect 35866 684808 35894 684972
rect 42058 684904 42064 684956
rect 42116 684944 42122 684956
rect 45094 684944 45100 684956
rect 42116 684916 45100 684944
rect 42116 684904 42122 684916
rect 45094 684904 45100 684916
rect 45152 684904 45158 684956
rect 41322 684808 41328 684820
rect 35866 684780 41328 684808
rect 41322 684768 41328 684780
rect 41380 684768 41386 684820
rect 35618 684632 35624 684684
rect 35676 684672 35682 684684
rect 41506 684672 41512 684684
rect 35676 684644 41512 684672
rect 35676 684632 35682 684644
rect 41506 684632 41512 684644
rect 41564 684632 41570 684684
rect 35802 684496 35808 684548
rect 35860 684536 35866 684548
rect 41690 684536 41696 684548
rect 35860 684508 41696 684536
rect 35860 684496 35866 684508
rect 41690 684496 41696 684508
rect 41748 684496 41754 684548
rect 35802 683408 35808 683460
rect 35860 683448 35866 683460
rect 41690 683448 41696 683460
rect 35860 683420 41696 683448
rect 35860 683408 35866 683420
rect 41690 683408 41696 683420
rect 41748 683408 41754 683460
rect 35618 683272 35624 683324
rect 35676 683312 35682 683324
rect 41506 683312 41512 683324
rect 35676 683284 41512 683312
rect 35676 683272 35682 683284
rect 41506 683272 41512 683284
rect 41564 683272 41570 683324
rect 35434 683136 35440 683188
rect 35492 683176 35498 683188
rect 41690 683176 41696 683188
rect 35492 683148 41696 683176
rect 35492 683136 35498 683148
rect 41690 683136 41696 683148
rect 41748 683136 41754 683188
rect 42058 683136 42064 683188
rect 42116 683176 42122 683188
rect 44358 683176 44364 683188
rect 42116 683148 44364 683176
rect 42116 683136 42122 683148
rect 44358 683136 44364 683148
rect 44416 683136 44422 683188
rect 674834 682524 674840 682576
rect 674892 682564 674898 682576
rect 683206 682564 683212 682576
rect 674892 682536 683212 682564
rect 674892 682524 674898 682536
rect 683206 682524 683212 682536
rect 683264 682524 683270 682576
rect 674834 682388 674840 682440
rect 674892 682428 674898 682440
rect 683482 682428 683488 682440
rect 674892 682400 683488 682428
rect 674892 682388 674898 682400
rect 683482 682388 683488 682400
rect 683540 682388 683546 682440
rect 35618 681844 35624 681896
rect 35676 681884 35682 681896
rect 41598 681884 41604 681896
rect 35676 681856 41604 681884
rect 35676 681844 35682 681856
rect 41598 681844 41604 681856
rect 41656 681844 41662 681896
rect 35802 681708 35808 681760
rect 35860 681748 35866 681760
rect 41414 681748 41420 681760
rect 35860 681720 41420 681748
rect 35860 681708 35866 681720
rect 41414 681708 41420 681720
rect 41472 681708 41478 681760
rect 42058 681708 42064 681760
rect 42116 681748 42122 681760
rect 42610 681748 42616 681760
rect 42116 681720 42616 681748
rect 42116 681708 42122 681720
rect 42610 681708 42616 681720
rect 42668 681708 42674 681760
rect 35802 680620 35808 680672
rect 35860 680660 35866 680672
rect 41690 680660 41696 680672
rect 35860 680632 41696 680660
rect 35860 680620 35866 680632
rect 41690 680620 41696 680632
rect 41748 680620 41754 680672
rect 35802 679396 35808 679448
rect 35860 679436 35866 679448
rect 41690 679436 41696 679448
rect 35860 679408 41696 679436
rect 35860 679396 35866 679408
rect 41690 679396 41696 679408
rect 41748 679396 41754 679448
rect 41690 679232 41696 679244
rect 41386 679204 41696 679232
rect 35618 679124 35624 679176
rect 35676 679164 35682 679176
rect 41386 679164 41414 679204
rect 41690 679192 41696 679204
rect 41748 679192 41754 679244
rect 42058 679192 42064 679244
rect 42116 679232 42122 679244
rect 44174 679232 44180 679244
rect 42116 679204 44180 679232
rect 42116 679192 42122 679204
rect 44174 679192 44180 679204
rect 44232 679192 44238 679244
rect 35676 679136 41414 679164
rect 35676 679124 35682 679136
rect 35434 678988 35440 679040
rect 35492 679028 35498 679040
rect 41690 679028 41696 679040
rect 35492 679000 41696 679028
rect 35492 678988 35498 679000
rect 41690 678988 41696 679000
rect 41748 678988 41754 679040
rect 42058 678988 42064 679040
rect 42116 679028 42122 679040
rect 44634 679028 44640 679040
rect 42116 679000 44640 679028
rect 42116 678988 42122 679000
rect 44634 678988 44640 679000
rect 44692 678988 44698 679040
rect 40770 677696 40776 677748
rect 40828 677736 40834 677748
rect 41598 677736 41604 677748
rect 40828 677708 41604 677736
rect 40828 677696 40834 677708
rect 41598 677696 41604 677708
rect 41656 677696 41662 677748
rect 42794 676200 42800 676252
rect 42852 676240 42858 676252
rect 55858 676240 55864 676252
rect 42852 676212 55864 676240
rect 42852 676200 42858 676212
rect 55858 676200 55864 676212
rect 55916 676200 55922 676252
rect 33042 674092 33048 674144
rect 33100 674132 33106 674144
rect 41506 674132 41512 674144
rect 33100 674104 41512 674132
rect 33100 674092 33106 674104
rect 41506 674092 41512 674104
rect 41564 674092 41570 674144
rect 35158 672868 35164 672920
rect 35216 672908 35222 672920
rect 39574 672908 39580 672920
rect 35216 672880 39580 672908
rect 35216 672868 35222 672880
rect 39574 672868 39580 672880
rect 39632 672868 39638 672920
rect 31018 672732 31024 672784
rect 31076 672772 31082 672784
rect 31076 672744 41414 672772
rect 31076 672732 31082 672744
rect 41386 672636 41414 672744
rect 41690 672636 41696 672648
rect 41386 672608 41696 672636
rect 41690 672596 41696 672608
rect 41748 672596 41754 672648
rect 42058 672528 42064 672580
rect 42116 672568 42122 672580
rect 42794 672568 42800 672580
rect 42116 672540 42800 672568
rect 42116 672528 42122 672540
rect 42794 672528 42800 672540
rect 42852 672528 42858 672580
rect 42610 672392 42616 672444
rect 42668 672432 42674 672444
rect 42668 672404 42840 672432
rect 42668 672392 42674 672404
rect 42812 672240 42840 672404
rect 42794 672188 42800 672240
rect 42852 672188 42858 672240
rect 673730 671304 673736 671356
rect 673788 671344 673794 671356
rect 673788 671316 673960 671344
rect 673788 671304 673794 671316
rect 668578 671100 668584 671152
rect 668636 671140 668642 671152
rect 673730 671140 673736 671152
rect 668636 671112 673736 671140
rect 668636 671100 668642 671112
rect 673730 671100 673736 671112
rect 673788 671100 673794 671152
rect 661678 670692 661684 670744
rect 661736 670732 661742 670744
rect 673932 670732 673960 671316
rect 661736 670704 673960 670732
rect 661736 670692 661742 670704
rect 674834 669808 674840 669860
rect 674892 669848 674898 669860
rect 676490 669848 676496 669860
rect 674892 669820 676496 669848
rect 674892 669808 674898 669820
rect 676490 669808 676496 669820
rect 676548 669808 676554 669860
rect 658918 669468 658924 669520
rect 658976 669508 658982 669520
rect 673730 669508 673736 669520
rect 658976 669480 673736 669508
rect 658976 669468 658982 669480
rect 673730 669468 673736 669480
rect 673788 669468 673794 669520
rect 45830 669400 45836 669452
rect 45888 669440 45894 669452
rect 45888 669412 51074 669440
rect 45888 669400 45894 669412
rect 51046 669372 51074 669412
rect 53098 669372 53104 669384
rect 51046 669344 53104 669372
rect 53098 669332 53104 669344
rect 53156 669332 53162 669384
rect 670234 669332 670240 669384
rect 670292 669372 670298 669384
rect 673362 669372 673368 669384
rect 670292 669344 673368 669372
rect 670292 669332 670298 669344
rect 673362 669332 673368 669344
rect 673420 669332 673426 669384
rect 673730 668652 673736 668704
rect 673788 668692 673794 668704
rect 673788 668664 673960 668692
rect 673788 668652 673794 668664
rect 671062 668516 671068 668568
rect 671120 668556 671126 668568
rect 673730 668556 673736 668568
rect 671120 668528 673736 668556
rect 671120 668516 671126 668528
rect 673730 668516 673736 668528
rect 673788 668516 673794 668568
rect 671430 668176 671436 668228
rect 671488 668216 671494 668228
rect 673932 668216 673960 668664
rect 671488 668188 673960 668216
rect 671488 668176 671494 668188
rect 45646 667904 45652 667956
rect 45704 667944 45710 667956
rect 58618 667944 58624 667956
rect 45704 667916 58624 667944
rect 45704 667904 45710 667916
rect 58618 667904 58624 667916
rect 58676 667904 58682 667956
rect 671062 667904 671068 667956
rect 671120 667944 671126 667956
rect 673730 667944 673736 667956
rect 671120 667916 673736 667944
rect 671120 667904 671126 667916
rect 673730 667904 673736 667916
rect 673788 667904 673794 667956
rect 673730 667292 673736 667344
rect 673788 667332 673794 667344
rect 673788 667304 673960 667332
rect 673788 667292 673794 667304
rect 671614 667156 671620 667208
rect 671672 667196 671678 667208
rect 673730 667196 673736 667208
rect 671672 667168 673736 667196
rect 671672 667156 671678 667168
rect 673730 667156 673736 667168
rect 673788 667156 673794 667208
rect 42242 666884 42248 666936
rect 42300 666924 42306 666936
rect 44174 666924 44180 666936
rect 42300 666896 44180 666924
rect 42300 666884 42306 666896
rect 44174 666884 44180 666896
rect 44232 666884 44238 666936
rect 671890 666884 671896 666936
rect 671948 666924 671954 666936
rect 673932 666924 673960 667304
rect 671948 666896 673960 666924
rect 671948 666884 671954 666896
rect 44634 666584 44640 666596
rect 42352 666556 44640 666584
rect 42352 665712 42380 666556
rect 44634 666544 44640 666556
rect 44692 666544 44698 666596
rect 671890 666544 671896 666596
rect 671948 666584 671954 666596
rect 673730 666584 673736 666596
rect 671948 666556 673736 666584
rect 671948 666544 671954 666556
rect 673730 666544 673736 666556
rect 673788 666544 673794 666596
rect 42334 665660 42340 665712
rect 42392 665660 42398 665712
rect 669590 665252 669596 665304
rect 669648 665292 669654 665304
rect 673730 665292 673736 665304
rect 669648 665264 673736 665292
rect 669648 665252 669654 665264
rect 673730 665252 673736 665264
rect 673788 665252 673794 665304
rect 672442 665116 672448 665168
rect 672500 665156 672506 665168
rect 673362 665156 673368 665168
rect 672500 665128 673368 665156
rect 672500 665116 672506 665128
rect 673362 665116 673368 665128
rect 673420 665116 673426 665168
rect 671706 664368 671712 664420
rect 671764 664408 671770 664420
rect 673730 664408 673736 664420
rect 671764 664380 673736 664408
rect 671764 664368 671770 664380
rect 673730 664368 673736 664380
rect 673788 664368 673794 664420
rect 669406 663892 669412 663944
rect 669464 663932 669470 663944
rect 673730 663932 673736 663944
rect 669464 663904 673736 663932
rect 669464 663892 669470 663904
rect 673730 663892 673736 663904
rect 673788 663892 673794 663944
rect 674834 663756 674840 663808
rect 674892 663796 674898 663808
rect 676030 663796 676036 663808
rect 674892 663768 676036 663796
rect 674892 663756 674898 663768
rect 676030 663756 676036 663768
rect 676088 663756 676094 663808
rect 672074 663416 672080 663468
rect 672132 663456 672138 663468
rect 673362 663456 673368 663468
rect 672132 663428 673368 663456
rect 672132 663416 672138 663428
rect 673362 663416 673368 663428
rect 673420 663416 673426 663468
rect 42242 663008 42248 663060
rect 42300 663048 42306 663060
rect 43990 663048 43996 663060
rect 42300 663020 43996 663048
rect 42300 663008 42306 663020
rect 43990 663008 43996 663020
rect 44048 663008 44054 663060
rect 42426 662872 42432 662924
rect 42484 662912 42490 662924
rect 45554 662912 45560 662924
rect 42484 662884 45560 662912
rect 42484 662872 42490 662884
rect 45554 662872 45560 662884
rect 45612 662872 45618 662924
rect 671246 661580 671252 661632
rect 671304 661620 671310 661632
rect 673730 661620 673736 661632
rect 671304 661592 673736 661620
rect 671304 661580 671310 661592
rect 673730 661580 673736 661592
rect 673788 661580 673794 661632
rect 668210 661104 668216 661156
rect 668268 661144 668274 661156
rect 673730 661144 673736 661156
rect 668268 661116 673736 661144
rect 668268 661104 668274 661116
rect 673730 661104 673736 661116
rect 673788 661104 673794 661156
rect 53098 660900 53104 660952
rect 53156 660940 53162 660952
rect 62114 660940 62120 660952
rect 53156 660912 62120 660940
rect 53156 660900 53162 660912
rect 62114 660900 62120 660912
rect 62172 660900 62178 660952
rect 668762 660084 668768 660136
rect 668820 660124 668826 660136
rect 673730 660124 673736 660136
rect 668820 660096 673736 660124
rect 668820 660084 668826 660096
rect 673730 660084 673736 660096
rect 673788 660084 673794 660136
rect 674834 659812 674840 659864
rect 674892 659852 674898 659864
rect 683114 659852 683120 659864
rect 674892 659824 683120 659852
rect 674892 659812 674898 659824
rect 683114 659812 683120 659824
rect 683172 659812 683178 659864
rect 58618 659540 58624 659592
rect 58676 659580 58682 659592
rect 62114 659580 62120 659592
rect 58676 659552 62120 659580
rect 58676 659540 58682 659552
rect 62114 659540 62120 659552
rect 62172 659540 62178 659592
rect 45370 658928 45376 658980
rect 45428 658968 45434 658980
rect 62298 658968 62304 658980
rect 45428 658940 62304 658968
rect 45428 658928 45434 658940
rect 62298 658928 62304 658940
rect 62356 658928 62362 658980
rect 42518 657500 42524 657552
rect 42576 657540 42582 657552
rect 62114 657540 62120 657552
rect 42576 657512 62120 657540
rect 42576 657500 42582 657512
rect 62114 657500 62120 657512
rect 62172 657500 62178 657552
rect 46198 656820 46204 656872
rect 46256 656860 46262 656872
rect 62114 656860 62120 656872
rect 46256 656832 62120 656860
rect 46256 656820 46262 656832
rect 62114 656820 62120 656832
rect 62172 656820 62178 656872
rect 653398 655528 653404 655580
rect 653456 655568 653462 655580
rect 673730 655568 673736 655580
rect 653456 655540 673736 655568
rect 653456 655528 653462 655540
rect 673730 655528 673736 655540
rect 673788 655528 673794 655580
rect 655514 645872 655520 645924
rect 655572 645912 655578 645924
rect 673730 645912 673736 645924
rect 655572 645884 673736 645912
rect 655572 645872 655578 645884
rect 673730 645872 673736 645884
rect 673788 645872 673794 645924
rect 35802 644444 35808 644496
rect 35860 644484 35866 644496
rect 39758 644484 39764 644496
rect 35860 644456 39764 644484
rect 35860 644444 35866 644456
rect 39758 644444 39764 644456
rect 39816 644444 39822 644496
rect 35802 643492 35808 643544
rect 35860 643532 35866 643544
rect 40218 643532 40224 643544
rect 35860 643504 40224 643532
rect 35860 643492 35866 643504
rect 40218 643492 40224 643504
rect 40276 643492 40282 643544
rect 41690 643328 41696 643340
rect 41386 643300 41696 643328
rect 35526 643220 35532 643272
rect 35584 643260 35590 643272
rect 41386 643260 41414 643300
rect 41690 643288 41696 643300
rect 41748 643288 41754 643340
rect 42058 643288 42064 643340
rect 42116 643328 42122 643340
rect 43806 643328 43812 643340
rect 42116 643300 43812 643328
rect 42116 643288 42122 643300
rect 43806 643288 43812 643300
rect 43864 643288 43870 643340
rect 35584 643232 41414 643260
rect 35584 643220 35590 643232
rect 35342 643084 35348 643136
rect 35400 643124 35406 643136
rect 41690 643124 41696 643136
rect 35400 643096 41696 643124
rect 35400 643084 35406 643096
rect 41690 643084 41696 643096
rect 41748 643084 41754 643136
rect 42058 643084 42064 643136
rect 42116 643124 42122 643136
rect 58618 643124 58624 643136
rect 42116 643096 58624 643124
rect 42116 643084 42122 643096
rect 58618 643084 58624 643096
rect 58676 643084 58682 643136
rect 655330 643084 655336 643136
rect 655388 643124 655394 643136
rect 673730 643124 673736 643136
rect 655388 643096 673736 643124
rect 655388 643084 655394 643096
rect 673730 643084 673736 643096
rect 673788 643084 673794 643136
rect 38562 642472 38568 642524
rect 38620 642512 38626 642524
rect 41690 642512 41696 642524
rect 38620 642484 41696 642512
rect 38620 642472 38626 642484
rect 41690 642472 41696 642484
rect 41748 642472 41754 642524
rect 42058 642336 42064 642388
rect 42116 642376 42122 642388
rect 62942 642376 62948 642388
rect 42116 642348 62948 642376
rect 42116 642336 42122 642348
rect 62942 642336 62948 642348
rect 63000 642336 63006 642388
rect 651466 642336 651472 642388
rect 651524 642376 651530 642388
rect 660298 642376 660304 642388
rect 651524 642348 660304 642376
rect 651524 642336 651530 642348
rect 660298 642336 660304 642348
rect 660356 642336 660362 642388
rect 35802 642132 35808 642184
rect 35860 642172 35866 642184
rect 39574 642172 39580 642184
rect 35860 642144 39580 642172
rect 35860 642132 35866 642144
rect 39574 642132 39580 642144
rect 39632 642132 39638 642184
rect 40770 642036 40776 642048
rect 36004 642008 40776 642036
rect 35802 641860 35808 641912
rect 35860 641900 35866 641912
rect 36004 641900 36032 642008
rect 40770 641996 40776 642008
rect 40828 641996 40834 642048
rect 35860 641872 36032 641900
rect 35860 641860 35866 641872
rect 35618 641724 35624 641776
rect 35676 641764 35682 641776
rect 41690 641764 41696 641776
rect 35676 641736 41696 641764
rect 35676 641724 35682 641736
rect 41690 641724 41696 641736
rect 41748 641724 41754 641776
rect 42058 641724 42064 641776
rect 42116 641764 42122 641776
rect 45278 641764 45284 641776
rect 42116 641736 45284 641764
rect 42116 641724 42122 641736
rect 45278 641724 45284 641736
rect 45336 641724 45342 641776
rect 35802 640772 35808 640824
rect 35860 640812 35866 640824
rect 35860 640772 35894 640812
rect 35866 640744 35894 640772
rect 39298 640744 39304 640756
rect 35866 640716 39304 640744
rect 39298 640704 39304 640716
rect 39356 640704 39362 640756
rect 40402 640540 40408 640552
rect 36004 640512 40408 640540
rect 35802 640432 35808 640484
rect 35860 640472 35866 640484
rect 36004 640472 36032 640512
rect 40402 640500 40408 640512
rect 40460 640500 40466 640552
rect 35860 640444 36032 640472
rect 35860 640432 35866 640444
rect 674834 640364 674840 640416
rect 674892 640364 674898 640416
rect 35618 640296 35624 640348
rect 35676 640336 35682 640348
rect 40862 640336 40868 640348
rect 35676 640308 40868 640336
rect 35676 640296 35682 640308
rect 40862 640296 40868 640308
rect 40920 640296 40926 640348
rect 651466 640296 651472 640348
rect 651524 640336 651530 640348
rect 668578 640336 668584 640348
rect 651524 640308 668584 640336
rect 651524 640296 651530 640308
rect 668578 640296 668584 640308
rect 668636 640296 668642 640348
rect 674852 640268 674880 640364
rect 675294 640268 675300 640280
rect 674852 640240 675300 640268
rect 675294 640228 675300 640240
rect 675352 640228 675358 640280
rect 651374 640092 651380 640144
rect 651432 640132 651438 640144
rect 653398 640132 653404 640144
rect 651432 640104 653404 640132
rect 651432 640092 651438 640104
rect 653398 640092 653404 640104
rect 653456 640092 653462 640144
rect 35802 639208 35808 639260
rect 35860 639248 35866 639260
rect 41690 639248 41696 639260
rect 35860 639220 41696 639248
rect 35860 639208 35866 639220
rect 41690 639208 41696 639220
rect 41748 639208 41754 639260
rect 35526 638936 35532 638988
rect 35584 638976 35590 638988
rect 39298 638976 39304 638988
rect 35584 638948 39304 638976
rect 35584 638936 35590 638948
rect 39298 638936 39304 638948
rect 39356 638936 39362 638988
rect 651650 638868 651656 638920
rect 651708 638908 651714 638920
rect 655330 638908 655336 638920
rect 651708 638880 655336 638908
rect 651708 638868 651714 638880
rect 655330 638868 655336 638880
rect 655388 638868 655394 638920
rect 651466 638732 651472 638784
rect 651524 638772 651530 638784
rect 655514 638772 655520 638784
rect 651524 638744 655520 638772
rect 651524 638732 651530 638744
rect 655514 638732 655520 638744
rect 655572 638732 655578 638784
rect 34422 638188 34428 638240
rect 34480 638228 34486 638240
rect 41690 638228 41696 638240
rect 34480 638200 41696 638228
rect 34480 638188 34486 638200
rect 41690 638188 41696 638200
rect 41748 638188 41754 638240
rect 35802 637848 35808 637900
rect 35860 637888 35866 637900
rect 36538 637888 36544 637900
rect 35860 637860 36544 637888
rect 35860 637848 35866 637860
rect 36538 637848 36544 637860
rect 36596 637848 36602 637900
rect 674466 636964 674472 637016
rect 674524 637004 674530 637016
rect 683206 637004 683212 637016
rect 674524 636976 683212 637004
rect 674524 636964 674530 636976
rect 683206 636964 683212 636976
rect 683264 636964 683270 637016
rect 35618 636896 35624 636948
rect 35676 636936 35682 636948
rect 40586 636936 40592 636948
rect 35676 636908 40592 636936
rect 35676 636896 35682 636908
rect 40586 636896 40592 636908
rect 40644 636896 40650 636948
rect 674282 636828 674288 636880
rect 674340 636868 674346 636880
rect 683390 636868 683396 636880
rect 674340 636840 683396 636868
rect 674340 636828 674346 636840
rect 683390 636828 683396 636840
rect 683448 636828 683454 636880
rect 35802 636692 35808 636744
rect 35860 636732 35866 636744
rect 35860 636692 35894 636732
rect 35866 636664 35894 636692
rect 40126 636664 40132 636676
rect 35866 636636 40132 636664
rect 40126 636624 40132 636636
rect 40184 636624 40190 636676
rect 40770 636460 40776 636472
rect 36004 636432 40776 636460
rect 35802 636352 35808 636404
rect 35860 636392 35866 636404
rect 36004 636392 36032 636432
rect 40770 636420 40776 636432
rect 40828 636420 40834 636472
rect 35860 636364 36032 636392
rect 35860 636352 35866 636364
rect 35526 636216 35532 636268
rect 35584 636256 35590 636268
rect 40586 636256 40592 636268
rect 35584 636228 40592 636256
rect 35584 636216 35590 636228
rect 40586 636216 40592 636228
rect 40644 636216 40650 636268
rect 671982 636148 671988 636200
rect 672040 636188 672046 636200
rect 672166 636188 672172 636200
rect 672040 636160 672172 636188
rect 672040 636148 672046 636160
rect 672166 636148 672172 636160
rect 672224 636148 672230 636200
rect 651834 635468 651840 635520
rect 651892 635508 651898 635520
rect 661678 635508 661684 635520
rect 651892 635480 661684 635508
rect 651892 635468 651898 635480
rect 661678 635468 661684 635480
rect 661736 635468 661742 635520
rect 674926 635468 674932 635520
rect 674984 635508 674990 635520
rect 675662 635508 675668 635520
rect 674984 635480 675668 635508
rect 674984 635468 674990 635480
rect 675662 635468 675668 635480
rect 675720 635468 675726 635520
rect 35802 634788 35808 634840
rect 35860 634828 35866 634840
rect 39942 634828 39948 634840
rect 35860 634800 39948 634828
rect 35860 634788 35866 634800
rect 39942 634788 39948 634800
rect 40000 634788 40006 634840
rect 35802 633836 35808 633888
rect 35860 633876 35866 633888
rect 35860 633836 35894 633876
rect 35866 633740 35894 633836
rect 40494 633740 40500 633752
rect 35866 633712 40500 633740
rect 40494 633700 40500 633712
rect 40552 633700 40558 633752
rect 35802 633428 35808 633480
rect 35860 633468 35866 633480
rect 41506 633468 41512 633480
rect 35860 633440 41512 633468
rect 35860 633428 35866 633440
rect 41506 633428 41512 633440
rect 41564 633428 41570 633480
rect 42150 633428 42156 633480
rect 42208 633468 42214 633480
rect 63402 633468 63408 633480
rect 42208 633440 63408 633468
rect 42208 633428 42214 633440
rect 63402 633428 63408 633440
rect 63460 633428 63466 633480
rect 671522 632952 671528 633004
rect 671580 632952 671586 633004
rect 671338 632924 671344 632936
rect 671172 632896 671344 632924
rect 671172 632652 671200 632896
rect 671338 632884 671344 632896
rect 671396 632884 671402 632936
rect 671338 632748 671344 632800
rect 671396 632788 671402 632800
rect 671540 632788 671568 632952
rect 671396 632760 671568 632788
rect 671396 632748 671402 632760
rect 671522 632652 671528 632664
rect 671172 632624 671528 632652
rect 671522 632612 671528 632624
rect 671580 632612 671586 632664
rect 36538 630572 36544 630624
rect 36596 630612 36602 630624
rect 36596 630584 41414 630612
rect 36596 630572 36602 630584
rect 41386 630544 41414 630584
rect 41598 630544 41604 630556
rect 41386 630516 41604 630544
rect 41598 630504 41604 630516
rect 41656 630504 41662 630556
rect 671890 630028 671896 630080
rect 671948 630068 671954 630080
rect 671948 630040 672120 630068
rect 671948 630028 671954 630040
rect 672092 629400 672120 630040
rect 672074 629348 672080 629400
rect 672132 629348 672138 629400
rect 35158 628532 35164 628584
rect 35216 628572 35222 628584
rect 39666 628572 39672 628584
rect 35216 628544 39672 628572
rect 35216 628532 35222 628544
rect 39666 628532 39672 628544
rect 39724 628532 39730 628584
rect 667198 626084 667204 626136
rect 667256 626124 667262 626136
rect 672810 626124 672816 626136
rect 667256 626096 672816 626124
rect 667256 626084 667262 626096
rect 672810 626084 672816 626096
rect 672868 626084 672874 626136
rect 44174 625812 44180 625864
rect 44232 625852 44238 625864
rect 63126 625852 63132 625864
rect 44232 625824 63132 625852
rect 44232 625812 44238 625824
rect 63126 625812 63132 625824
rect 63184 625812 63190 625864
rect 669958 625540 669964 625592
rect 670016 625580 670022 625592
rect 672166 625580 672172 625592
rect 670016 625552 672172 625580
rect 670016 625540 670022 625552
rect 672166 625540 672172 625552
rect 672224 625540 672230 625592
rect 42334 625132 42340 625184
rect 42392 625172 42398 625184
rect 44358 625172 44364 625184
rect 42392 625144 44364 625172
rect 42392 625132 42398 625144
rect 44358 625132 44364 625144
rect 44416 625132 44422 625184
rect 657538 625132 657544 625184
rect 657596 625172 657602 625184
rect 672810 625172 672816 625184
rect 657596 625144 672816 625172
rect 657596 625132 657602 625144
rect 672810 625132 672816 625144
rect 672868 625132 672874 625184
rect 670234 624996 670240 625048
rect 670292 625036 670298 625048
rect 672810 625036 672816 625048
rect 670292 625008 672816 625036
rect 670292 624996 670298 625008
rect 672810 624996 672816 625008
rect 672868 624996 672874 625048
rect 670418 624656 670424 624708
rect 670476 624696 670482 624708
rect 672810 624696 672816 624708
rect 670476 624668 672816 624696
rect 670476 624656 670482 624668
rect 672810 624656 672816 624668
rect 672868 624656 672874 624708
rect 671430 624316 671436 624368
rect 671488 624356 671494 624368
rect 672810 624356 672816 624368
rect 671488 624328 672816 624356
rect 671488 624316 671494 624328
rect 672810 624316 672816 624328
rect 672868 624316 672874 624368
rect 670234 623840 670240 623892
rect 670292 623880 670298 623892
rect 672810 623880 672816 623892
rect 670292 623852 672816 623880
rect 670292 623840 670298 623852
rect 672810 623840 672816 623852
rect 672868 623840 672874 623892
rect 44082 623812 44088 623824
rect 42352 623784 44088 623812
rect 42352 623416 42380 623784
rect 44082 623772 44088 623784
rect 44140 623772 44146 623824
rect 671062 623500 671068 623552
rect 671120 623540 671126 623552
rect 672810 623540 672816 623552
rect 671120 623512 672816 623540
rect 671120 623500 671126 623512
rect 672810 623500 672816 623512
rect 672868 623500 672874 623552
rect 42334 623364 42340 623416
rect 42392 623364 42398 623416
rect 669406 623024 669412 623076
rect 669464 623064 669470 623076
rect 672810 623064 672816 623076
rect 669464 623036 672816 623064
rect 669464 623024 669470 623036
rect 672810 623024 672816 623036
rect 672868 623024 672874 623076
rect 674650 623024 674656 623076
rect 674708 623064 674714 623076
rect 683390 623064 683396 623076
rect 674708 623036 683396 623064
rect 674708 623024 674714 623036
rect 683390 623024 683396 623036
rect 683448 623024 683454 623076
rect 42426 621460 42432 621512
rect 42484 621500 42490 621512
rect 42484 621472 42656 621500
rect 42484 621460 42490 621472
rect 42628 621240 42656 621472
rect 42610 621188 42616 621240
rect 42668 621188 42674 621240
rect 666462 621052 666468 621104
rect 666520 621092 666526 621104
rect 672810 621092 672816 621104
rect 666520 621064 672816 621092
rect 666520 621052 666526 621064
rect 672810 621052 672816 621064
rect 672868 621052 672874 621104
rect 674282 620984 674288 621036
rect 674340 621024 674346 621036
rect 676214 621024 676220 621036
rect 674340 620996 676220 621024
rect 674340 620984 674346 620996
rect 676214 620984 676220 620996
rect 676272 620984 676278 621036
rect 668946 620236 668952 620288
rect 669004 620276 669010 620288
rect 672810 620276 672816 620288
rect 669004 620248 672816 620276
rect 669004 620236 669010 620248
rect 672810 620236 672816 620248
rect 672868 620236 672874 620288
rect 670878 619964 670884 620016
rect 670936 620004 670942 620016
rect 672810 620004 672816 620016
rect 670936 619976 672816 620004
rect 670936 619964 670942 619976
rect 672810 619964 672816 619976
rect 672868 619964 672874 620016
rect 666278 619692 666284 619744
rect 666336 619732 666342 619744
rect 672810 619732 672816 619744
rect 666336 619704 672816 619732
rect 666336 619692 666342 619704
rect 672810 619692 672816 619704
rect 672868 619692 672874 619744
rect 674374 619692 674380 619744
rect 674432 619732 674438 619744
rect 676030 619732 676036 619744
rect 674432 619704 676036 619732
rect 674432 619692 674438 619704
rect 676030 619692 676036 619704
rect 676088 619692 676094 619744
rect 42242 619624 42248 619676
rect 42300 619664 42306 619676
rect 42886 619664 42892 619676
rect 42300 619636 42892 619664
rect 42300 619624 42306 619636
rect 42886 619624 42892 619636
rect 42944 619624 42950 619676
rect 42702 618876 42708 618928
rect 42760 618916 42766 618928
rect 43898 618916 43904 618928
rect 42760 618888 43904 618916
rect 42760 618876 42766 618888
rect 43898 618876 43904 618888
rect 43956 618876 43962 618928
rect 674282 618468 674288 618520
rect 674340 618508 674346 618520
rect 676214 618508 676220 618520
rect 674340 618480 676220 618508
rect 674340 618468 674346 618480
rect 676214 618468 676220 618480
rect 676272 618468 676278 618520
rect 674282 617992 674288 618044
rect 674340 618032 674346 618044
rect 676490 618032 676496 618044
rect 674340 618004 676496 618032
rect 674340 617992 674346 618004
rect 676490 617992 676496 618004
rect 676548 617992 676554 618044
rect 674282 617856 674288 617908
rect 674340 617896 674346 617908
rect 676214 617896 676220 617908
rect 674340 617868 676220 617896
rect 674340 617856 674346 617868
rect 676214 617856 676220 617868
rect 676272 617856 676278 617908
rect 670602 617448 670608 617500
rect 670660 617488 670666 617500
rect 674006 617488 674012 617500
rect 670660 617460 674012 617488
rect 670660 617448 670666 617460
rect 674006 617448 674012 617460
rect 674064 617448 674070 617500
rect 674282 617448 674288 617500
rect 674340 617488 674346 617500
rect 676214 617488 676220 617500
rect 674340 617460 676220 617488
rect 674340 617448 674346 617460
rect 676214 617448 676220 617460
rect 676272 617448 676278 617500
rect 42150 617108 42156 617160
rect 42208 617148 42214 617160
rect 42702 617148 42708 617160
rect 42208 617120 42708 617148
rect 42208 617108 42214 617120
rect 42702 617108 42708 617120
rect 42760 617108 42766 617160
rect 668394 616836 668400 616888
rect 668452 616876 668458 616888
rect 674006 616876 674012 616888
rect 668452 616848 674012 616876
rect 668452 616836 668458 616848
rect 674006 616836 674012 616848
rect 674064 616836 674070 616888
rect 44174 616768 44180 616820
rect 44232 616808 44238 616820
rect 62114 616808 62120 616820
rect 44232 616780 62120 616808
rect 44232 616768 44238 616780
rect 62114 616768 62120 616780
rect 62172 616768 62178 616820
rect 669774 615612 669780 615664
rect 669832 615652 669838 615664
rect 674006 615652 674012 615664
rect 669832 615624 674012 615652
rect 669832 615612 669838 615624
rect 674006 615612 674012 615624
rect 674064 615612 674070 615664
rect 674282 615476 674288 615528
rect 674340 615516 674346 615528
rect 683114 615516 683120 615528
rect 674340 615488 683120 615516
rect 674340 615476 674346 615488
rect 683114 615476 683120 615488
rect 683172 615476 683178 615528
rect 674282 614592 674288 614644
rect 674340 614632 674346 614644
rect 676214 614632 676220 614644
rect 674340 614604 676220 614632
rect 674340 614592 674346 614604
rect 676214 614592 676220 614604
rect 676272 614592 676278 614644
rect 42794 614116 42800 614168
rect 42852 614156 42858 614168
rect 62114 614156 62120 614168
rect 42852 614128 62120 614156
rect 42852 614116 42858 614128
rect 62114 614116 62120 614128
rect 62172 614116 62178 614168
rect 670602 614116 670608 614168
rect 670660 614156 670666 614168
rect 674006 614156 674012 614168
rect 670660 614128 674012 614156
rect 670660 614116 670666 614128
rect 674006 614116 674012 614128
rect 674064 614116 674070 614168
rect 58618 613980 58624 614032
rect 58676 614020 58682 614032
rect 62114 614020 62120 614032
rect 58676 613992 62120 614020
rect 58676 613980 58682 613992
rect 62114 613980 62120 613992
rect 62172 613980 62178 614032
rect 46198 613368 46204 613420
rect 46256 613408 46262 613420
rect 62114 613408 62120 613420
rect 46256 613380 62120 613408
rect 46256 613368 46262 613380
rect 62114 613368 62120 613380
rect 62172 613368 62178 613420
rect 43070 612824 43076 612876
rect 43128 612864 43134 612876
rect 43128 612836 43760 612864
rect 43128 612824 43134 612836
rect 43732 612728 43760 612836
rect 43898 612728 43904 612740
rect 43732 612700 43904 612728
rect 43898 612688 43904 612700
rect 43956 612688 43962 612740
rect 43254 612620 43260 612672
rect 43312 612660 43318 612672
rect 43312 612632 43691 612660
rect 43312 612620 43318 612632
rect 42242 612348 42248 612400
rect 42300 612388 42306 612400
rect 42300 612360 43562 612388
rect 42300 612348 42306 612360
rect 43663 612306 43691 612632
rect 53098 612592 53104 612604
rect 43778 612564 53104 612592
rect 43778 612170 43806 612564
rect 53098 612552 53104 612564
rect 53156 612552 53162 612604
rect 44910 611980 44916 611992
rect 43901 611952 44916 611980
rect 44910 611940 44916 611952
rect 44968 611940 44974 611992
rect 46198 611708 46204 611720
rect 44022 611680 46204 611708
rect 46198 611668 46204 611680
rect 46256 611668 46262 611720
rect 44088 611584 44140 611590
rect 44088 611526 44140 611532
rect 653398 611328 653404 611380
rect 653456 611368 653462 611380
rect 674006 611368 674012 611380
rect 653456 611340 674012 611368
rect 653456 611328 653462 611340
rect 674006 611328 674012 611340
rect 674064 611328 674070 611380
rect 674282 611328 674288 611380
rect 674340 611368 674346 611380
rect 675386 611368 675392 611380
rect 674340 611340 675392 611368
rect 674340 611328 674346 611340
rect 675386 611328 675392 611340
rect 675444 611328 675450 611380
rect 50154 611300 50160 611312
rect 44237 611272 50160 611300
rect 50154 611260 50160 611272
rect 50212 611260 50218 611312
rect 44312 611124 44318 611176
rect 44370 611124 44376 611176
rect 44461 610864 45554 610892
rect 44726 610756 44732 610768
rect 44574 610728 44732 610756
rect 44726 610716 44732 610728
rect 44784 610716 44790 610768
rect 45526 610008 45554 610864
rect 50154 610104 50160 610156
rect 50212 610144 50218 610156
rect 58618 610144 58624 610156
rect 50212 610116 58624 610144
rect 50212 610104 50218 610116
rect 58618 610104 58624 610116
rect 58676 610104 58682 610156
rect 64322 610008 64328 610020
rect 45526 609980 64328 610008
rect 64322 609968 64328 609980
rect 64380 609968 64386 610020
rect 669038 608608 669044 608660
rect 669096 608648 669102 608660
rect 674006 608648 674012 608660
rect 669096 608620 674012 608648
rect 669096 608608 669102 608620
rect 674006 608608 674012 608620
rect 674064 608608 674070 608660
rect 674282 608608 674288 608660
rect 674340 608648 674346 608660
rect 675110 608648 675116 608660
rect 674340 608620 675116 608648
rect 674340 608608 674346 608620
rect 675110 608608 675116 608620
rect 675168 608608 675174 608660
rect 673546 607248 673552 607300
rect 673604 607248 673610 607300
rect 673564 607096 673592 607248
rect 673546 607044 673552 607096
rect 673604 607044 673610 607096
rect 673270 603508 673276 603560
rect 673328 603548 673334 603560
rect 674006 603548 674012 603560
rect 673328 603520 674012 603548
rect 673328 603508 673334 603520
rect 674006 603508 674012 603520
rect 674064 603508 674070 603560
rect 674282 603236 674288 603288
rect 674340 603276 674346 603288
rect 675110 603276 675116 603288
rect 674340 603248 675116 603276
rect 674340 603236 674346 603248
rect 675110 603236 675116 603248
rect 675168 603236 675174 603288
rect 657538 600312 657544 600364
rect 657596 600352 657602 600364
rect 674006 600352 674012 600364
rect 657596 600324 674012 600352
rect 657596 600312 657602 600324
rect 674006 600312 674012 600324
rect 674064 600312 674070 600364
rect 674006 599400 674012 599412
rect 663766 599372 674012 599400
rect 654778 598952 654784 599004
rect 654836 598992 654842 599004
rect 663766 598992 663794 599372
rect 674006 599360 674012 599372
rect 674064 599360 674070 599412
rect 654836 598964 663794 598992
rect 654836 598952 654842 598964
rect 674558 598952 674564 599004
rect 674616 598992 674622 599004
rect 675294 598992 675300 599004
rect 674616 598964 675300 598992
rect 674616 598952 674622 598964
rect 675294 598952 675300 598964
rect 675352 598952 675358 599004
rect 674466 598340 674472 598392
rect 674524 598380 674530 598392
rect 675294 598380 675300 598392
rect 674524 598352 675300 598380
rect 674524 598340 674530 598352
rect 675294 598340 675300 598352
rect 675352 598340 675358 598392
rect 651466 597524 651472 597576
rect 651524 597564 651530 597576
rect 669958 597564 669964 597576
rect 651524 597536 669964 597564
rect 651524 597524 651530 597536
rect 669958 597524 669964 597536
rect 670016 597524 670022 597576
rect 43070 597388 43076 597440
rect 43128 597388 43134 597440
rect 43088 597032 43116 597388
rect 43070 596980 43076 597032
rect 43128 596980 43134 597032
rect 651466 596164 651472 596216
rect 651524 596204 651530 596216
rect 667198 596204 667204 596216
rect 651524 596176 667204 596204
rect 651524 596164 651530 596176
rect 667198 596164 667204 596176
rect 667256 596164 667262 596216
rect 40126 595756 40132 595808
rect 40184 595796 40190 595808
rect 41690 595796 41696 595808
rect 40184 595768 41696 595796
rect 40184 595756 40190 595768
rect 41690 595756 41696 595768
rect 41748 595756 41754 595808
rect 651650 595484 651656 595536
rect 651708 595524 651714 595536
rect 653398 595524 653404 595536
rect 651708 595496 653404 595524
rect 651708 595484 651714 595496
rect 653398 595484 653404 595496
rect 653456 595484 653462 595536
rect 41322 594804 41328 594856
rect 41380 594844 41386 594856
rect 41690 594844 41696 594856
rect 41380 594816 41696 594844
rect 41380 594804 41386 594816
rect 41690 594804 41696 594816
rect 41748 594804 41754 594856
rect 651466 594804 651472 594856
rect 651524 594844 651530 594856
rect 658918 594844 658924 594856
rect 651524 594816 658924 594844
rect 651524 594804 651530 594816
rect 658918 594804 658924 594816
rect 658976 594804 658982 594856
rect 39942 594668 39948 594720
rect 40000 594708 40006 594720
rect 41690 594708 41696 594720
rect 40000 594680 41696 594708
rect 40000 594668 40006 594680
rect 41690 594668 41696 594680
rect 41748 594668 41754 594720
rect 651466 594668 651472 594720
rect 651524 594708 651530 594720
rect 657538 594708 657544 594720
rect 651524 594680 657544 594708
rect 651524 594668 651530 594680
rect 657538 594668 657544 594680
rect 657596 594668 657602 594720
rect 651466 593240 651472 593292
rect 651524 593280 651530 593292
rect 654778 593280 654784 593292
rect 651524 593252 654784 593280
rect 651524 593240 651530 593252
rect 654778 593240 654784 593252
rect 654836 593240 654842 593292
rect 683390 592668 683396 592680
rect 678946 592640 683396 592668
rect 674742 592560 674748 592612
rect 674800 592600 674806 592612
rect 678946 592600 678974 592640
rect 683390 592628 683396 592640
rect 683448 592628 683454 592680
rect 674800 592572 678974 592600
rect 674800 592560 674806 592572
rect 39298 591404 39304 591456
rect 39356 591444 39362 591456
rect 41414 591444 41420 591456
rect 39356 591416 41420 591444
rect 39356 591404 39362 591416
rect 41414 591404 41420 591416
rect 41472 591404 41478 591456
rect 35802 590928 35808 590980
rect 35860 590968 35866 590980
rect 40770 590968 40776 590980
rect 35860 590940 40776 590968
rect 35860 590928 35866 590940
rect 40770 590928 40776 590940
rect 40828 590928 40834 590980
rect 41690 590764 41696 590776
rect 36004 590736 41696 590764
rect 35618 590656 35624 590708
rect 35676 590696 35682 590708
rect 36004 590696 36032 590736
rect 41690 590724 41696 590736
rect 41748 590724 41754 590776
rect 35676 590668 36032 590696
rect 35676 590656 35682 590668
rect 42058 590656 42064 590708
rect 42116 590696 42122 590708
rect 43254 590696 43260 590708
rect 42116 590668 43260 590696
rect 42116 590656 42122 590668
rect 43254 590656 43260 590668
rect 43312 590656 43318 590708
rect 674834 590588 674840 590640
rect 674892 590628 674898 590640
rect 682378 590628 682384 590640
rect 674892 590600 682384 590628
rect 674892 590588 674898 590600
rect 682378 590588 682384 590600
rect 682436 590588 682442 590640
rect 675294 590424 675300 590436
rect 675128 590396 675300 590424
rect 675128 590232 675156 590396
rect 675294 590384 675300 590396
rect 675352 590384 675358 590436
rect 675110 590180 675116 590232
rect 675168 590180 675174 590232
rect 674466 588548 674472 588600
rect 674524 588588 674530 588600
rect 684034 588588 684040 588600
rect 674524 588560 684040 588588
rect 674524 588548 674530 588560
rect 684034 588548 684040 588560
rect 684092 588548 684098 588600
rect 33042 587120 33048 587172
rect 33100 587160 33106 587172
rect 41506 587160 41512 587172
rect 33100 587132 41512 587160
rect 33100 587120 33106 587132
rect 41506 587120 41512 587132
rect 41564 587120 41570 587172
rect 37918 585828 37924 585880
rect 37976 585868 37982 585880
rect 41690 585868 41696 585880
rect 37976 585840 41696 585868
rect 37976 585828 37982 585840
rect 41690 585828 41696 585840
rect 41748 585828 41754 585880
rect 42058 585828 42064 585880
rect 42116 585868 42122 585880
rect 42610 585868 42616 585880
rect 42116 585840 42616 585868
rect 42116 585828 42122 585840
rect 42610 585828 42616 585840
rect 42668 585828 42674 585880
rect 31018 585692 31024 585744
rect 31076 585732 31082 585744
rect 41690 585732 41696 585744
rect 31076 585704 41696 585732
rect 31076 585692 31082 585704
rect 41690 585692 41696 585704
rect 41748 585692 41754 585744
rect 42058 585624 42064 585676
rect 42116 585664 42122 585676
rect 42702 585664 42708 585676
rect 42116 585636 42708 585664
rect 42116 585624 42122 585636
rect 42702 585624 42708 585636
rect 42760 585624 42766 585676
rect 672258 584400 672264 584452
rect 672316 584440 672322 584452
rect 672626 584440 672632 584452
rect 672316 584412 672632 584440
rect 672316 584400 672322 584412
rect 672626 584400 672632 584412
rect 672684 584400 672690 584452
rect 42426 582428 42432 582480
rect 42484 582428 42490 582480
rect 42242 582088 42248 582140
rect 42300 582128 42306 582140
rect 42444 582128 42472 582428
rect 42300 582100 42472 582128
rect 42300 582088 42306 582100
rect 661678 581000 661684 581052
rect 661736 581040 661742 581052
rect 673638 581040 673644 581052
rect 661736 581012 673644 581040
rect 661736 581000 661742 581012
rect 673638 581000 673644 581012
rect 673696 581000 673702 581052
rect 42426 580592 42432 580644
rect 42484 580632 42490 580644
rect 43254 580632 43260 580644
rect 42484 580604 43260 580632
rect 42484 580592 42490 580604
rect 43254 580592 43260 580604
rect 43312 580592 43318 580644
rect 668578 580252 668584 580304
rect 668636 580292 668642 580304
rect 673638 580292 673644 580304
rect 668636 580264 673644 580292
rect 668636 580252 668642 580264
rect 673638 580252 673644 580264
rect 673696 580252 673702 580304
rect 42242 580048 42248 580100
rect 42300 580048 42306 580100
rect 42260 579964 42288 580048
rect 42242 579912 42248 579964
rect 42300 579912 42306 579964
rect 670418 579844 670424 579896
rect 670476 579884 670482 579896
rect 673638 579884 673644 579896
rect 670476 579856 673644 579884
rect 670476 579844 670482 579856
rect 673638 579844 673644 579856
rect 673696 579844 673702 579896
rect 660298 579640 660304 579692
rect 660356 579680 660362 579692
rect 673086 579680 673092 579692
rect 660356 579652 673092 579680
rect 660356 579640 660362 579652
rect 673086 579640 673092 579652
rect 673144 579640 673150 579692
rect 670786 579368 670792 579420
rect 670844 579408 670850 579420
rect 673638 579408 673644 579420
rect 670844 579380 673644 579408
rect 670844 579368 670850 579380
rect 673638 579368 673644 579380
rect 673696 579368 673702 579420
rect 670234 579028 670240 579080
rect 670292 579068 670298 579080
rect 673638 579068 673644 579080
rect 670292 579040 673644 579068
rect 670292 579028 670298 579040
rect 673638 579028 673644 579040
rect 673696 579028 673702 579080
rect 671154 578552 671160 578604
rect 671212 578592 671218 578604
rect 673638 578592 673644 578604
rect 671212 578564 673644 578592
rect 671212 578552 671218 578564
rect 673638 578552 673644 578564
rect 673696 578552 673702 578604
rect 669406 578144 669412 578196
rect 669464 578184 669470 578196
rect 673638 578184 673644 578196
rect 669464 578156 673644 578184
rect 669464 578144 669470 578156
rect 673638 578144 673644 578156
rect 673696 578144 673702 578196
rect 670234 577736 670240 577788
rect 670292 577776 670298 577788
rect 673638 577776 673644 577788
rect 670292 577748 673644 577776
rect 670292 577736 670298 577748
rect 673638 577736 673644 577748
rect 673696 577736 673702 577788
rect 671430 577396 671436 577448
rect 671488 577436 671494 577448
rect 673638 577436 673644 577448
rect 671488 577408 673644 577436
rect 671488 577396 671494 577408
rect 673638 577396 673644 577408
rect 673696 577396 673702 577448
rect 669406 576920 669412 576972
rect 669464 576960 669470 576972
rect 673638 576960 673644 576972
rect 669464 576932 673644 576960
rect 669464 576920 669470 576932
rect 673638 576920 673644 576932
rect 673696 576920 673702 576972
rect 45094 575424 45100 575476
rect 45152 575464 45158 575476
rect 62114 575464 62120 575476
rect 45152 575436 62120 575464
rect 45152 575424 45158 575436
rect 62114 575424 62120 575436
rect 62172 575424 62178 575476
rect 671614 574540 671620 574592
rect 671672 574580 671678 574592
rect 673638 574580 673644 574592
rect 671672 574552 673644 574580
rect 671672 574540 671678 574552
rect 673638 574540 673644 574552
rect 673696 574540 673702 574592
rect 671982 574132 671988 574184
rect 672040 574172 672046 574184
rect 673638 574172 673644 574184
rect 672040 574144 673644 574172
rect 672040 574132 672046 574144
rect 673638 574132 673644 574144
rect 673696 574132 673702 574184
rect 51718 573996 51724 574048
rect 51776 574036 51782 574048
rect 62114 574036 62120 574048
rect 51776 574008 62120 574036
rect 51776 573996 51782 574008
rect 62114 573996 62120 574008
rect 62172 573996 62178 574048
rect 672258 573996 672264 574048
rect 672316 574036 672322 574048
rect 673086 574036 673092 574048
rect 672316 574008 673092 574036
rect 672316 573996 672322 574008
rect 673086 573996 673092 574008
rect 673144 573996 673150 574048
rect 42242 573452 42248 573504
rect 42300 573492 42306 573504
rect 42702 573492 42708 573504
rect 42300 573464 42708 573492
rect 42300 573452 42306 573464
rect 42702 573452 42708 573464
rect 42760 573452 42766 573504
rect 669590 572228 669596 572280
rect 669648 572268 669654 572280
rect 673638 572268 673644 572280
rect 669648 572240 673644 572268
rect 669648 572228 669654 572240
rect 673638 572228 673644 572240
rect 673696 572228 673702 572280
rect 674466 571548 674472 571600
rect 674524 571588 674530 571600
rect 676214 571588 676220 571600
rect 674524 571560 676220 571588
rect 674524 571548 674530 571560
rect 676214 571548 676220 571560
rect 676272 571548 676278 571600
rect 671798 571412 671804 571464
rect 671856 571452 671862 571464
rect 673638 571452 673644 571464
rect 671856 571424 673644 571452
rect 671856 571412 671862 571424
rect 673638 571412 673644 571424
rect 673696 571412 673702 571464
rect 42058 570936 42064 570988
rect 42116 570976 42122 570988
rect 42610 570976 42616 570988
rect 42116 570948 42616 570976
rect 42116 570936 42122 570948
rect 42610 570936 42616 570948
rect 42668 570936 42674 570988
rect 674834 570460 674840 570512
rect 674892 570500 674898 570512
rect 675478 570500 675484 570512
rect 674892 570472 675484 570500
rect 674892 570460 674898 570472
rect 675478 570460 675484 570472
rect 675536 570500 675542 570512
rect 683114 570500 683120 570512
rect 675536 570472 683120 570500
rect 675536 570460 675542 570472
rect 683114 570460 683120 570472
rect 683172 570460 683178 570512
rect 671338 570392 671344 570444
rect 671396 570432 671402 570444
rect 671396 570404 673868 570432
rect 671396 570392 671402 570404
rect 671982 570120 671988 570172
rect 672040 570160 672046 570172
rect 673638 570160 673644 570172
rect 672040 570132 673644 570160
rect 672040 570120 672046 570132
rect 673638 570120 673644 570132
rect 673696 570120 673702 570172
rect 673638 569916 673644 569968
rect 673696 569956 673702 569968
rect 673840 569956 673868 570404
rect 673696 569928 673868 569956
rect 673696 569916 673702 569928
rect 669774 568556 669780 568608
rect 669832 568596 669838 568608
rect 673638 568596 673644 568608
rect 669832 568568 673644 568596
rect 669832 568556 669838 568568
rect 673638 568556 673644 568568
rect 673696 568556 673702 568608
rect 653398 565836 653404 565888
rect 653456 565876 653462 565888
rect 673638 565876 673644 565888
rect 653456 565848 673644 565876
rect 653456 565836 653462 565848
rect 673638 565836 673644 565848
rect 673696 565836 673702 565888
rect 665082 564544 665088 564596
rect 665140 564584 665146 564596
rect 673638 564584 673644 564596
rect 665140 564556 673644 564584
rect 665140 564544 665146 564556
rect 673638 564544 673644 564556
rect 673696 564544 673702 564596
rect 661034 554752 661040 554804
rect 661092 554792 661098 554804
rect 673638 554792 673644 554804
rect 661092 554764 673644 554792
rect 661092 554752 661098 554764
rect 673638 554752 673644 554764
rect 673696 554752 673702 554804
rect 655146 553392 655152 553444
rect 655204 553432 655210 553444
rect 673638 553432 673644 553444
rect 655204 553404 673644 553432
rect 655204 553392 655210 553404
rect 673638 553392 673644 553404
rect 673696 553392 673702 553444
rect 651466 552644 651472 552696
rect 651524 552684 651530 552696
rect 665818 552684 665824 552696
rect 651524 552656 665824 552684
rect 651524 552644 651530 552656
rect 665818 552644 665824 552656
rect 665876 552644 665882 552696
rect 675202 552576 675208 552628
rect 675260 552576 675266 552628
rect 675220 552356 675248 552576
rect 675202 552304 675208 552356
rect 675260 552304 675266 552356
rect 674650 550604 674656 550656
rect 674708 550644 674714 550656
rect 674834 550644 674840 550656
rect 674708 550616 674840 550644
rect 674708 550604 674714 550616
rect 674834 550604 674840 550616
rect 674892 550604 674898 550656
rect 40954 550468 40960 550520
rect 41012 550508 41018 550520
rect 41690 550508 41696 550520
rect 41012 550480 41696 550508
rect 41012 550468 41018 550480
rect 41690 550468 41696 550480
rect 41748 550468 41754 550520
rect 675202 550468 675208 550520
rect 675260 550468 675266 550520
rect 651650 550332 651656 550384
rect 651708 550372 651714 550384
rect 653398 550372 653404 550384
rect 651708 550344 653404 550372
rect 651708 550332 651714 550344
rect 653398 550332 653404 550344
rect 653456 550332 653462 550384
rect 675220 549964 675248 550468
rect 675220 549936 675340 549964
rect 651466 549856 651472 549908
rect 651524 549896 651530 549908
rect 664438 549896 664444 549908
rect 651524 549868 664444 549896
rect 651524 549856 651530 549868
rect 664438 549856 664444 549868
rect 664496 549856 664502 549908
rect 675312 549840 675340 549936
rect 675294 549788 675300 549840
rect 675352 549788 675358 549840
rect 651466 549176 651472 549228
rect 651524 549216 651530 549228
rect 661034 549216 661040 549228
rect 651524 549188 661040 549216
rect 651524 549176 651530 549188
rect 661034 549176 661040 549188
rect 661092 549176 661098 549228
rect 651466 548836 651472 548888
rect 651524 548876 651530 548888
rect 655146 548876 655152 548888
rect 651524 548848 655152 548876
rect 651524 548836 651530 548848
rect 655146 548836 655152 548848
rect 655204 548836 655210 548888
rect 41322 547952 41328 548004
rect 41380 547992 41386 548004
rect 41380 547952 41414 547992
rect 41386 547924 41414 547952
rect 41690 547924 41696 547936
rect 41386 547896 41696 547924
rect 41690 547884 41696 547896
rect 41748 547884 41754 547936
rect 42058 547884 42064 547936
rect 42116 547924 42122 547936
rect 43254 547924 43260 547936
rect 42116 547896 43260 547924
rect 42116 547884 42122 547896
rect 43254 547884 43260 547896
rect 43312 547884 43318 547936
rect 29638 547136 29644 547188
rect 29696 547176 29702 547188
rect 41690 547176 41696 547188
rect 29696 547148 41696 547176
rect 29696 547136 29702 547148
rect 41690 547136 41696 547148
rect 41748 547136 41754 547188
rect 675570 547136 675576 547188
rect 675628 547176 675634 547188
rect 683206 547176 683212 547188
rect 675628 547148 683212 547176
rect 675628 547136 675634 547148
rect 683206 547136 683212 547148
rect 683264 547136 683270 547188
rect 674834 545980 674840 546032
rect 674892 545980 674898 546032
rect 674852 545884 674880 545980
rect 682378 545884 682384 545896
rect 674852 545856 682384 545884
rect 682378 545844 682384 545856
rect 682436 545844 682442 545896
rect 667198 535916 667204 535968
rect 667256 535956 667262 535968
rect 672626 535956 672632 535968
rect 667256 535928 672632 535956
rect 667256 535916 667262 535928
rect 672626 535916 672632 535928
rect 672684 535916 672690 535968
rect 669958 535644 669964 535696
rect 670016 535684 670022 535696
rect 672626 535684 672632 535696
rect 670016 535656 672632 535684
rect 670016 535644 670022 535656
rect 672626 535644 672632 535656
rect 672684 535644 672690 535696
rect 670786 534828 670792 534880
rect 670844 534868 670850 534880
rect 672626 534868 672632 534880
rect 670844 534840 672632 534868
rect 670844 534828 670850 534840
rect 672626 534828 672632 534840
rect 672684 534828 672690 534880
rect 671154 534556 671160 534608
rect 671212 534596 671218 534608
rect 672626 534596 672632 534608
rect 671212 534568 672632 534596
rect 671212 534556 671218 534568
rect 672626 534556 672632 534568
rect 672684 534556 672690 534608
rect 658918 534216 658924 534268
rect 658976 534256 658982 534268
rect 672626 534256 672632 534268
rect 658976 534228 672632 534256
rect 658976 534216 658982 534228
rect 672626 534216 672632 534228
rect 672684 534216 672690 534268
rect 674282 534080 674288 534132
rect 674340 534120 674346 534132
rect 676030 534120 676036 534132
rect 674340 534092 676036 534120
rect 674340 534080 674346 534092
rect 676030 534080 676036 534092
rect 676088 534080 676094 534132
rect 670234 533332 670240 533384
rect 670292 533372 670298 533384
rect 672442 533372 672448 533384
rect 670292 533344 672448 533372
rect 670292 533332 670298 533344
rect 672442 533332 672448 533344
rect 672500 533332 672506 533384
rect 674282 533332 674288 533384
rect 674340 533372 674346 533384
rect 683574 533372 683580 533384
rect 674340 533344 683580 533372
rect 674340 533332 674346 533344
rect 683574 533332 683580 533344
rect 683632 533332 683638 533384
rect 42426 532720 42432 532772
rect 42484 532760 42490 532772
rect 43070 532760 43076 532772
rect 42484 532732 43076 532760
rect 42484 532720 42490 532732
rect 43070 532720 43076 532732
rect 43128 532720 43134 532772
rect 669406 532516 669412 532568
rect 669464 532556 669470 532568
rect 672442 532556 672448 532568
rect 669464 532528 672448 532556
rect 669464 532516 669470 532528
rect 672442 532516 672448 532528
rect 672500 532516 672506 532568
rect 673822 532176 673828 532228
rect 673880 532176 673886 532228
rect 673840 531820 673868 532176
rect 675478 531972 675484 532024
rect 675536 532012 675542 532024
rect 676214 532012 676220 532024
rect 675536 531984 676220 532012
rect 675536 531972 675542 531984
rect 676214 531972 676220 531984
rect 676272 531972 676278 532024
rect 673822 531768 673828 531820
rect 673880 531768 673886 531820
rect 51718 531224 51724 531276
rect 51776 531264 51782 531276
rect 62114 531264 62120 531276
rect 51776 531236 62120 531264
rect 51776 531224 51782 531236
rect 62114 531224 62120 531236
rect 62172 531224 62178 531276
rect 45278 531088 45284 531140
rect 45336 531128 45342 531140
rect 62114 531128 62120 531140
rect 45336 531100 62120 531128
rect 45336 531088 45342 531100
rect 62114 531088 62120 531100
rect 62172 531088 62178 531140
rect 673270 530884 673276 530936
rect 673328 530924 673334 530936
rect 674006 530924 674012 530936
rect 673328 530896 674012 530924
rect 673328 530884 673334 530896
rect 674006 530884 674012 530896
rect 674064 530884 674070 530936
rect 674282 530816 674288 530868
rect 674340 530856 674346 530868
rect 676030 530856 676036 530868
rect 674340 530828 676036 530856
rect 674340 530816 674346 530828
rect 676030 530816 676036 530828
rect 676088 530816 676094 530868
rect 667382 529932 667388 529984
rect 667440 529972 667446 529984
rect 674006 529972 674012 529984
rect 667440 529944 674012 529972
rect 667440 529932 667446 529944
rect 674006 529932 674012 529944
rect 674064 529932 674070 529984
rect 674282 529932 674288 529984
rect 674340 529972 674346 529984
rect 676030 529972 676036 529984
rect 674340 529944 676036 529972
rect 674340 529932 674346 529944
rect 676030 529932 676036 529944
rect 676088 529932 676094 529984
rect 42150 529456 42156 529508
rect 42208 529496 42214 529508
rect 42610 529496 42616 529508
rect 42208 529468 42616 529496
rect 42208 529456 42214 529468
rect 42610 529456 42616 529468
rect 42668 529456 42674 529508
rect 670970 529252 670976 529304
rect 671028 529292 671034 529304
rect 674006 529292 674012 529304
rect 671028 529264 674012 529292
rect 671028 529252 671034 529264
rect 674006 529252 674012 529264
rect 674064 529252 674070 529304
rect 674282 529184 674288 529236
rect 674340 529224 674346 529236
rect 676030 529224 676036 529236
rect 674340 529196 676036 529224
rect 674340 529184 674346 529196
rect 676030 529184 676036 529196
rect 676088 529184 676094 529236
rect 674282 528980 674288 529032
rect 674340 529020 674346 529032
rect 676214 529020 676220 529032
rect 674340 528992 676220 529020
rect 674340 528980 674346 528992
rect 676214 528980 676220 528992
rect 676272 528980 676278 529032
rect 45278 528572 45284 528624
rect 45336 528612 45342 528624
rect 62114 528612 62120 528624
rect 45336 528584 62120 528612
rect 45336 528572 45342 528584
rect 62114 528572 62120 528584
rect 62172 528572 62178 528624
rect 668854 528572 668860 528624
rect 668912 528612 668918 528624
rect 674006 528612 674012 528624
rect 668912 528584 674012 528612
rect 668912 528572 668918 528584
rect 674006 528572 674012 528584
rect 674064 528572 674070 528624
rect 54478 527076 54484 527128
rect 54536 527116 54542 527128
rect 62114 527116 62120 527128
rect 54536 527088 62120 527116
rect 54536 527076 54542 527088
rect 62114 527076 62120 527088
rect 62172 527076 62178 527128
rect 42058 527008 42064 527060
rect 42116 527048 42122 527060
rect 42610 527048 42616 527060
rect 42116 527020 42616 527048
rect 42116 527008 42122 527020
rect 42610 527008 42616 527020
rect 42668 527008 42674 527060
rect 674650 526736 674656 526788
rect 674708 526776 674714 526788
rect 676030 526776 676036 526788
rect 674708 526748 676036 526776
rect 674708 526736 674714 526748
rect 676030 526736 676036 526748
rect 676088 526736 676094 526788
rect 674282 526328 674288 526380
rect 674340 526368 674346 526380
rect 676030 526368 676036 526380
rect 674340 526340 676036 526368
rect 674340 526328 674346 526340
rect 676030 526328 676036 526340
rect 676088 526328 676094 526380
rect 667566 524424 667572 524476
rect 667624 524464 667630 524476
rect 674006 524464 674012 524476
rect 667624 524436 674012 524464
rect 667624 524424 667630 524436
rect 674006 524424 674012 524436
rect 674064 524424 674070 524476
rect 674282 524424 674288 524476
rect 674340 524464 674346 524476
rect 683114 524464 683120 524476
rect 674340 524436 683120 524464
rect 674340 524424 674346 524436
rect 683114 524424 683120 524436
rect 683172 524424 683178 524476
rect 663794 521568 663800 521620
rect 663852 521608 663858 521620
rect 667566 521608 667572 521620
rect 663852 521580 667572 521608
rect 663852 521568 663858 521580
rect 667566 521568 667572 521580
rect 667624 521568 667630 521620
rect 675478 520208 675484 520260
rect 675536 520248 675542 520260
rect 678974 520248 678980 520260
rect 675536 520220 678980 520248
rect 675536 520208 675542 520220
rect 678974 520208 678980 520220
rect 679032 520208 679038 520260
rect 675662 518780 675668 518832
rect 675720 518820 675726 518832
rect 677870 518820 677876 518832
rect 675720 518792 677876 518820
rect 675720 518780 675726 518792
rect 677870 518780 677876 518792
rect 677928 518780 677934 518832
rect 656342 514020 656348 514072
rect 656400 514060 656406 514072
rect 663794 514060 663800 514072
rect 656400 514032 663800 514060
rect 656400 514020 656406 514032
rect 663794 514020 663800 514032
rect 663852 514020 663858 514072
rect 653398 510620 653404 510672
rect 653456 510660 653462 510672
rect 656342 510660 656348 510672
rect 653456 510632 656348 510660
rect 653456 510620 653462 510632
rect 656342 510620 656348 510632
rect 656400 510620 656406 510672
rect 675110 503616 675116 503668
rect 675168 503656 675174 503668
rect 679618 503656 679624 503668
rect 675168 503628 679624 503656
rect 675168 503616 675174 503628
rect 679618 503616 679624 503628
rect 679676 503616 679682 503668
rect 675294 503480 675300 503532
rect 675352 503520 675358 503532
rect 680998 503520 681004 503532
rect 675352 503492 681004 503520
rect 675352 503480 675358 503492
rect 680998 503480 681004 503492
rect 681056 503480 681062 503532
rect 674834 500896 674840 500948
rect 674892 500936 674898 500948
rect 681182 500936 681188 500948
rect 674892 500908 681188 500936
rect 674892 500896 674898 500908
rect 681182 500896 681188 500908
rect 681240 500896 681246 500948
rect 652018 500216 652024 500268
rect 652076 500256 652082 500268
rect 669958 500256 669964 500268
rect 652076 500228 669964 500256
rect 652076 500216 652082 500228
rect 669958 500216 669964 500228
rect 670016 500216 670022 500268
rect 650638 494708 650644 494760
rect 650696 494748 650702 494760
rect 653398 494748 653404 494760
rect 650696 494720 653404 494748
rect 650696 494708 650702 494720
rect 653398 494708 653404 494720
rect 653456 494708 653462 494760
rect 674282 491988 674288 492040
rect 674340 492028 674346 492040
rect 674650 492028 674656 492040
rect 674340 492000 674656 492028
rect 674340 491988 674346 492000
rect 674650 491988 674656 492000
rect 674708 491988 674714 492040
rect 669958 491852 669964 491904
rect 670016 491892 670022 491904
rect 674006 491892 674012 491904
rect 670016 491864 674012 491892
rect 670016 491852 670022 491864
rect 674006 491852 674012 491864
rect 674064 491852 674070 491904
rect 674282 491784 674288 491836
rect 674340 491824 674346 491836
rect 675846 491824 675852 491836
rect 674340 491796 675852 491824
rect 674340 491784 674346 491796
rect 675846 491784 675852 491796
rect 675904 491784 675910 491836
rect 674282 491648 674288 491700
rect 674340 491688 674346 491700
rect 676030 491688 676036 491700
rect 674340 491660 676036 491688
rect 674340 491648 674346 491660
rect 676030 491648 676036 491660
rect 676088 491648 676094 491700
rect 665818 491444 665824 491496
rect 665876 491484 665882 491496
rect 674006 491484 674012 491496
rect 665876 491456 674012 491484
rect 665876 491444 665882 491456
rect 674006 491444 674012 491456
rect 674064 491444 674070 491496
rect 664438 491308 664444 491360
rect 664496 491348 664502 491360
rect 673822 491348 673828 491360
rect 664496 491320 673828 491348
rect 664496 491308 664502 491320
rect 673822 491308 673828 491320
rect 673880 491308 673886 491360
rect 670786 490900 670792 490952
rect 670844 490940 670850 490952
rect 674006 490940 674012 490952
rect 670844 490912 674012 490940
rect 670844 490900 670850 490912
rect 674006 490900 674012 490912
rect 674064 490900 674070 490952
rect 672442 490424 672448 490476
rect 672500 490464 672506 490476
rect 674006 490464 674012 490476
rect 672500 490436 674012 490464
rect 672500 490424 672506 490436
rect 674006 490424 674012 490436
rect 674064 490424 674070 490476
rect 672626 490084 672632 490136
rect 672684 490124 672690 490136
rect 674006 490124 674012 490136
rect 672684 490096 674012 490124
rect 672684 490084 672690 490096
rect 674006 490084 674012 490096
rect 674064 490084 674070 490136
rect 672626 489608 672632 489660
rect 672684 489648 672690 489660
rect 674006 489648 674012 489660
rect 672684 489620 674012 489648
rect 672684 489608 672690 489620
rect 674006 489608 674012 489620
rect 674064 489608 674070 489660
rect 671614 489268 671620 489320
rect 671672 489308 671678 489320
rect 674006 489308 674012 489320
rect 671672 489280 674012 489308
rect 671672 489268 671678 489280
rect 674006 489268 674012 489280
rect 674064 489268 674070 489320
rect 671154 488452 671160 488504
rect 671212 488492 671218 488504
rect 674006 488492 674012 488504
rect 671212 488464 674012 488492
rect 671212 488452 671218 488464
rect 674006 488452 674012 488464
rect 674064 488452 674070 488504
rect 674282 486140 674288 486192
rect 674340 486180 674346 486192
rect 676030 486180 676036 486192
rect 674340 486152 676036 486180
rect 674340 486140 674346 486152
rect 676030 486140 676036 486152
rect 676088 486140 676094 486192
rect 672258 486004 672264 486056
rect 672316 486044 672322 486056
rect 673822 486044 673828 486056
rect 672316 486016 673828 486044
rect 672316 486004 672322 486016
rect 673822 486004 673828 486016
rect 673880 486004 673886 486056
rect 665082 485800 665088 485852
rect 665140 485840 665146 485852
rect 674006 485840 674012 485852
rect 665140 485812 674012 485840
rect 665140 485800 665146 485812
rect 674006 485800 674012 485812
rect 674064 485800 674070 485852
rect 674282 485120 674288 485172
rect 674340 485160 674346 485172
rect 676030 485160 676036 485172
rect 674340 485132 676036 485160
rect 674340 485120 674346 485132
rect 676030 485120 676036 485132
rect 676088 485120 676094 485172
rect 667014 484372 667020 484424
rect 667072 484412 667078 484424
rect 674006 484412 674012 484424
rect 667072 484384 674012 484412
rect 667072 484372 667078 484384
rect 674006 484372 674012 484384
rect 674064 484372 674070 484424
rect 674466 483964 674472 484016
rect 674524 484004 674530 484016
rect 676030 484004 676036 484016
rect 674524 483976 676036 484004
rect 674524 483964 674530 483976
rect 676030 483964 676036 483976
rect 676088 483964 676094 484016
rect 671798 483148 671804 483200
rect 671856 483188 671862 483200
rect 674006 483188 674012 483200
rect 671856 483160 674012 483188
rect 671856 483148 671862 483160
rect 674006 483148 674012 483160
rect 674064 483148 674070 483200
rect 676214 482944 676220 482996
rect 676272 482984 676278 482996
rect 677410 482984 677416 482996
rect 676272 482956 677416 482984
rect 676272 482944 676278 482956
rect 677410 482944 677416 482956
rect 677468 482944 677474 482996
rect 669958 480700 669964 480752
rect 670016 480740 670022 480752
rect 670418 480740 670424 480752
rect 670016 480712 670424 480740
rect 670016 480700 670022 480712
rect 670418 480700 670424 480712
rect 670476 480740 670482 480752
rect 674006 480740 674012 480752
rect 670476 480712 674012 480740
rect 670476 480700 670482 480712
rect 674006 480700 674012 480712
rect 674064 480700 674070 480752
rect 674282 480360 674288 480412
rect 674340 480400 674346 480412
rect 683114 480400 683120 480412
rect 674340 480372 683120 480400
rect 674340 480360 674346 480372
rect 683114 480360 683120 480372
rect 683172 480360 683178 480412
rect 676030 476076 676036 476128
rect 676088 476116 676094 476128
rect 680354 476116 680360 476128
rect 676088 476088 680360 476116
rect 676088 476076 676094 476088
rect 680354 476076 680360 476088
rect 680412 476076 680418 476128
rect 657538 467100 657544 467152
rect 657596 467140 657602 467152
rect 669958 467140 669964 467152
rect 657596 467112 669964 467140
rect 657596 467100 657602 467112
rect 669958 467100 669964 467112
rect 670016 467100 670022 467152
rect 653398 460164 653404 460216
rect 653456 460204 653462 460216
rect 657538 460204 657544 460216
rect 653456 460176 657544 460204
rect 653456 460164 653462 460176
rect 657538 460164 657544 460176
rect 657596 460164 657602 460216
rect 667842 456560 667848 456612
rect 667900 456600 667906 456612
rect 667900 456572 673988 456600
rect 667900 456560 667906 456572
rect 673960 456246 673988 456572
rect 669222 455948 669228 456000
rect 669280 455988 669286 456000
rect 669280 455960 673854 455988
rect 669280 455948 669286 455960
rect 673362 455812 673368 455864
rect 673420 455852 673426 455864
rect 673420 455824 673762 455852
rect 673420 455812 673426 455824
rect 668210 455608 668216 455660
rect 668268 455648 668274 455660
rect 668268 455620 673624 455648
rect 668268 455608 668274 455620
rect 673270 455336 673276 455388
rect 673328 455336 673334 455388
rect 673288 455022 673316 455336
rect 673388 455252 673440 455258
rect 673388 455194 673440 455200
rect 673506 455252 673558 455258
rect 673506 455194 673558 455200
rect 674282 454860 674288 454912
rect 674340 454900 674346 454912
rect 675846 454900 675852 454912
rect 674340 454872 675852 454900
rect 674340 454860 674346 454872
rect 675846 454860 675852 454872
rect 675904 454860 675910 454912
rect 672074 454792 672080 454844
rect 672132 454832 672138 454844
rect 672132 454804 673190 454832
rect 672132 454792 672138 454804
rect 673046 454640 673098 454646
rect 674282 454588 674288 454640
rect 674340 454628 674346 454640
rect 675478 454628 675484 454640
rect 674340 454600 675484 454628
rect 674340 454588 674346 454600
rect 675478 454588 675484 454600
rect 675536 454588 675542 454640
rect 673046 454582 673098 454588
rect 672810 454452 672816 454504
rect 672868 454452 672874 454504
rect 672828 454206 672856 454452
rect 672954 454368 673006 454374
rect 674282 454316 674288 454368
rect 674340 454356 674346 454368
rect 675662 454356 675668 454368
rect 674340 454328 675668 454356
rect 674340 454316 674346 454328
rect 675662 454316 675668 454328
rect 675720 454316 675726 454368
rect 672954 454310 673006 454316
rect 672258 453908 672264 453960
rect 672316 453948 672322 453960
rect 672316 453920 672750 453948
rect 672316 453908 672322 453920
rect 674282 453908 674288 453960
rect 674340 453948 674346 453960
rect 676030 453948 676036 453960
rect 674340 453920 676036 453948
rect 674340 453908 674346 453920
rect 676030 453908 676036 453920
rect 676088 453908 676094 453960
rect 44818 451392 44824 451444
rect 44876 451432 44882 451444
rect 47762 451432 47768 451444
rect 44876 451404 47768 451432
rect 44876 451392 44882 451404
rect 47762 451392 47768 451404
rect 47820 451392 47826 451444
rect 35802 429156 35808 429208
rect 35860 429196 35866 429208
rect 41322 429196 41328 429208
rect 35860 429168 41328 429196
rect 35860 429156 35866 429168
rect 41322 429156 41328 429168
rect 41380 429156 41386 429208
rect 35802 427932 35808 427984
rect 35860 427972 35866 427984
rect 41598 427972 41604 427984
rect 35860 427944 41604 427972
rect 35860 427932 35866 427944
rect 41598 427932 41604 427944
rect 41656 427932 41662 427984
rect 41138 424328 41144 424380
rect 41196 424368 41202 424380
rect 41690 424368 41696 424380
rect 41196 424340 41696 424368
rect 41196 424328 41202 424340
rect 41690 424328 41696 424340
rect 41748 424328 41754 424380
rect 33042 417392 33048 417444
rect 33100 417432 33106 417444
rect 41690 417432 41696 417444
rect 33100 417404 41696 417432
rect 33100 417392 33106 417404
rect 41690 417392 41696 417404
rect 41748 417392 41754 417444
rect 42058 417256 42064 417308
rect 42116 417296 42122 417308
rect 42518 417296 42524 417308
rect 42116 417268 42524 417296
rect 42116 417256 42122 417268
rect 42518 417256 42524 417268
rect 42576 417256 42582 417308
rect 34514 416032 34520 416084
rect 34572 416072 34578 416084
rect 41598 416072 41604 416084
rect 34572 416044 41604 416072
rect 34572 416032 34578 416044
rect 41598 416032 41604 416044
rect 41656 416032 41662 416084
rect 42242 409776 42248 409828
rect 42300 409816 42306 409828
rect 42702 409816 42708 409828
rect 42300 409788 42708 409816
rect 42300 409776 42306 409788
rect 42702 409776 42708 409788
rect 42760 409776 42766 409828
rect 42242 407668 42248 407720
rect 42300 407708 42306 407720
rect 42610 407708 42616 407720
rect 42300 407680 42616 407708
rect 42300 407668 42306 407680
rect 42610 407668 42616 407680
rect 42668 407668 42674 407720
rect 51074 404268 51080 404320
rect 51132 404308 51138 404320
rect 62114 404308 62120 404320
rect 51132 404280 62120 404308
rect 51132 404268 51138 404280
rect 62114 404268 62120 404280
rect 62172 404268 62178 404320
rect 674558 403248 674564 403300
rect 674616 403288 674622 403300
rect 676214 403288 676220 403300
rect 674616 403260 676220 403288
rect 674616 403248 674622 403260
rect 676214 403248 676220 403260
rect 676272 403248 676278 403300
rect 51442 402908 51448 402960
rect 51500 402948 51506 402960
rect 62114 402948 62120 402960
rect 51500 402920 62120 402948
rect 51500 402908 51506 402920
rect 62114 402908 62120 402920
rect 62172 402908 62178 402960
rect 51074 400188 51080 400240
rect 51132 400228 51138 400240
rect 62114 400228 62120 400240
rect 51132 400200 62120 400228
rect 51132 400188 51138 400200
rect 62114 400188 62120 400200
rect 62172 400188 62178 400240
rect 44818 400052 44824 400104
rect 44876 400092 44882 400104
rect 62114 400092 62120 400104
rect 44876 400064 62120 400092
rect 44876 400052 44882 400064
rect 62114 400052 62120 400064
rect 62172 400052 62178 400104
rect 674926 398828 674932 398880
rect 674984 398868 674990 398880
rect 676030 398868 676036 398880
rect 674984 398840 676036 398868
rect 674984 398828 674990 398840
rect 676030 398828 676036 398840
rect 676088 398828 676094 398880
rect 54478 398760 54484 398812
rect 54536 398800 54542 398812
rect 62114 398800 62120 398812
rect 54536 398772 62120 398800
rect 54536 398760 54542 398772
rect 62114 398760 62120 398772
rect 62172 398760 62178 398812
rect 675018 395700 675024 395752
rect 675076 395740 675082 395752
rect 676214 395740 676220 395752
rect 675076 395712 676220 395740
rect 675076 395700 675082 395712
rect 676214 395700 676220 395712
rect 676272 395700 676278 395752
rect 674374 395496 674380 395548
rect 674432 395536 674438 395548
rect 676214 395536 676220 395548
rect 674432 395508 676220 395536
rect 674432 395496 674438 395508
rect 676214 395496 676220 395508
rect 676272 395496 676278 395548
rect 674466 394272 674472 394324
rect 674524 394312 674530 394324
rect 676214 394312 676220 394324
rect 674524 394284 676220 394312
rect 674524 394272 674530 394284
rect 676214 394272 676220 394284
rect 676272 394272 676278 394324
rect 679618 386764 679624 386776
rect 675588 386736 679624 386764
rect 41322 386384 41328 386436
rect 41380 386424 41386 386436
rect 41598 386424 41604 386436
rect 41380 386396 41604 386424
rect 41380 386384 41386 386396
rect 41598 386384 41604 386396
rect 41656 386384 41662 386436
rect 675588 386424 675616 386736
rect 679618 386724 679624 386736
rect 679676 386724 679682 386776
rect 675496 386396 675616 386424
rect 674834 386112 674840 386164
rect 674892 386152 674898 386164
rect 675294 386152 675300 386164
rect 674892 386124 675300 386152
rect 674892 386112 674898 386124
rect 675294 386112 675300 386124
rect 675352 386112 675358 386164
rect 675496 386028 675524 386396
rect 675478 385976 675484 386028
rect 675536 385976 675542 386028
rect 41322 382508 41328 382560
rect 41380 382548 41386 382560
rect 41598 382548 41604 382560
rect 41380 382520 41604 382548
rect 41380 382508 41386 382520
rect 41598 382508 41604 382520
rect 41656 382508 41662 382560
rect 35802 379516 35808 379568
rect 35860 379556 35866 379568
rect 40402 379556 40408 379568
rect 35860 379528 40408 379556
rect 35860 379516 35866 379528
rect 40402 379516 40408 379528
rect 40460 379516 40466 379568
rect 674466 378088 674472 378140
rect 674524 378128 674530 378140
rect 675110 378128 675116 378140
rect 674524 378100 675116 378128
rect 674524 378088 674530 378100
rect 675110 378088 675116 378100
rect 675168 378088 675174 378140
rect 35802 376728 35808 376780
rect 35860 376768 35866 376780
rect 41690 376768 41696 376780
rect 35860 376740 41696 376768
rect 35860 376728 35866 376740
rect 41690 376728 41696 376740
rect 41748 376728 41754 376780
rect 674374 375300 674380 375352
rect 674432 375340 674438 375352
rect 675110 375340 675116 375352
rect 674432 375312 675116 375340
rect 674432 375300 674438 375312
rect 675110 375300 675116 375312
rect 675168 375300 675174 375352
rect 651466 373940 651472 373992
rect 651524 373980 651530 373992
rect 663058 373980 663064 373992
rect 651524 373952 663064 373980
rect 651524 373940 651530 373952
rect 663058 373940 663064 373952
rect 663116 373940 663122 373992
rect 33962 373260 33968 373312
rect 34020 373300 34026 373312
rect 41690 373300 41696 373312
rect 34020 373272 41696 373300
rect 34020 373260 34026 373272
rect 41690 373260 41696 373272
rect 41748 373260 41754 373312
rect 39298 371628 39304 371680
rect 39356 371668 39362 371680
rect 41690 371668 41696 371680
rect 39356 371640 41696 371668
rect 39356 371628 39362 371640
rect 41690 371628 41696 371640
rect 41748 371628 41754 371680
rect 42058 371560 42064 371612
rect 42116 371600 42122 371612
rect 42518 371600 42524 371612
rect 42116 371572 42524 371600
rect 42116 371560 42122 371572
rect 42518 371560 42524 371572
rect 42576 371560 42582 371612
rect 651466 370948 651472 371000
rect 651524 370988 651530 371000
rect 654778 370988 654784 371000
rect 651524 370960 654784 370988
rect 651524 370948 651530 370960
rect 654778 370948 654784 370960
rect 654836 370948 654842 371000
rect 42242 365304 42248 365356
rect 42300 365344 42306 365356
rect 43070 365344 43076 365356
rect 42300 365316 43076 365344
rect 42300 365304 42306 365316
rect 43070 365304 43076 365316
rect 43128 365304 43134 365356
rect 662414 364352 662420 364404
rect 662472 364392 662478 364404
rect 666462 364392 666468 364404
rect 662472 364364 666468 364392
rect 662472 364352 662478 364364
rect 666462 364352 666468 364364
rect 666520 364352 666526 364404
rect 42242 362856 42248 362908
rect 42300 362856 42306 362908
rect 42260 362636 42288 362856
rect 42242 362584 42248 362636
rect 42300 362584 42306 362636
rect 44726 361496 44732 361548
rect 44784 361536 44790 361548
rect 62114 361536 62120 361548
rect 44784 361508 62120 361536
rect 44784 361496 44790 361508
rect 62114 361496 62120 361508
rect 62172 361496 62178 361548
rect 657538 360204 657544 360256
rect 657596 360244 657602 360256
rect 662414 360244 662420 360256
rect 657596 360216 662420 360244
rect 657596 360204 657602 360216
rect 662414 360204 662420 360216
rect 662472 360204 662478 360256
rect 51074 360136 51080 360188
rect 51132 360176 51138 360188
rect 62114 360176 62120 360188
rect 51132 360148 62120 360176
rect 51132 360136 51138 360148
rect 62114 360136 62120 360148
rect 62172 360136 62178 360188
rect 42150 359932 42156 359984
rect 42208 359972 42214 359984
rect 42886 359972 42892 359984
rect 42208 359944 42892 359972
rect 42208 359932 42214 359944
rect 42886 359932 42892 359944
rect 42944 359932 42950 359984
rect 54478 356668 54484 356720
rect 54536 356708 54542 356720
rect 62114 356708 62120 356720
rect 54536 356680 62120 356708
rect 54536 356668 54542 356680
rect 62114 356668 62120 356680
rect 62172 356668 62178 356720
rect 44634 354968 44640 355020
rect 44692 355008 44698 355020
rect 44692 354980 45002 355008
rect 44692 354968 44698 354980
rect 44634 354832 44640 354884
rect 44692 354872 44698 354884
rect 44692 354844 44895 354872
rect 44692 354832 44698 354844
rect 44640 354544 44692 354550
rect 44640 354486 44692 354492
rect 44732 354408 44784 354414
rect 44732 354350 44784 354356
rect 44867 354314 44895 354844
rect 44974 354110 45002 354980
rect 45646 353852 45652 353864
rect 45105 353824 45652 353852
rect 45646 353812 45652 353824
rect 45704 353812 45710 353864
rect 45830 353716 45836 353728
rect 45218 353688 45836 353716
rect 45830 353676 45836 353688
rect 45888 353676 45894 353728
rect 45646 353444 45652 353456
rect 45329 353416 45652 353444
rect 45646 353404 45652 353416
rect 45704 353404 45710 353456
rect 46014 353240 46020 353252
rect 45448 353212 46020 353240
rect 46014 353200 46020 353212
rect 46072 353200 46078 353252
rect 652018 348372 652024 348424
rect 652076 348412 652082 348424
rect 657538 348412 657544 348424
rect 652076 348384 657544 348412
rect 652076 348372 652082 348384
rect 657538 348372 657544 348384
rect 657596 348372 657602 348424
rect 35802 343748 35808 343800
rect 35860 343788 35866 343800
rect 40218 343788 40224 343800
rect 35860 343760 40224 343788
rect 35860 343748 35866 343760
rect 40218 343748 40224 343760
rect 40276 343748 40282 343800
rect 35526 343612 35532 343664
rect 35584 343652 35590 343664
rect 40034 343652 40040 343664
rect 35584 343624 40040 343652
rect 35584 343612 35590 343624
rect 40034 343612 40040 343624
rect 40092 343612 40098 343664
rect 35802 341300 35808 341352
rect 35860 341340 35866 341352
rect 39850 341340 39856 341352
rect 35860 341312 39856 341340
rect 35860 341300 35866 341312
rect 39850 341300 39856 341312
rect 39908 341300 39914 341352
rect 35802 341164 35808 341216
rect 35860 341204 35866 341216
rect 40218 341204 40224 341216
rect 35860 341176 40224 341204
rect 35860 341164 35866 341176
rect 40218 341164 40224 341176
rect 40276 341164 40282 341216
rect 35526 341028 35532 341080
rect 35584 341068 35590 341080
rect 40034 341068 40040 341080
rect 35584 341040 40040 341068
rect 35584 341028 35590 341040
rect 40034 341028 40040 341040
rect 40092 341028 40098 341080
rect 35802 339600 35808 339652
rect 35860 339640 35866 339652
rect 37918 339640 37924 339652
rect 35860 339612 37924 339640
rect 35860 339600 35866 339612
rect 37918 339600 37924 339612
rect 37976 339600 37982 339652
rect 35526 339464 35532 339516
rect 35584 339504 35590 339516
rect 38930 339504 38936 339516
rect 35584 339476 38936 339504
rect 35584 339464 35590 339476
rect 38930 339464 38936 339476
rect 38988 339464 38994 339516
rect 35802 335316 35808 335368
rect 35860 335356 35866 335368
rect 40218 335356 40224 335368
rect 35860 335328 40224 335356
rect 35860 335316 35866 335328
rect 40218 335316 40224 335328
rect 40276 335316 40282 335368
rect 35802 334092 35808 334144
rect 35860 334132 35866 334144
rect 39758 334132 39764 334144
rect 35860 334104 39764 334132
rect 35860 334092 35866 334104
rect 39758 334092 39764 334104
rect 39816 334092 39822 334144
rect 674466 331032 674472 331084
rect 674524 331072 674530 331084
rect 675110 331072 675116 331084
rect 674524 331044 675116 331072
rect 674524 331032 674530 331044
rect 675110 331032 675116 331044
rect 675168 331032 675174 331084
rect 651466 328244 651472 328296
rect 651524 328284 651530 328296
rect 654778 328284 654784 328296
rect 651524 328256 654784 328284
rect 651524 328244 651530 328256
rect 654778 328244 654784 328256
rect 654836 328244 654842 328296
rect 651742 325592 651748 325644
rect 651800 325632 651806 325644
rect 653582 325632 653588 325644
rect 651800 325604 653588 325632
rect 651800 325592 651806 325604
rect 653582 325592 653588 325604
rect 653640 325592 653646 325644
rect 650822 322940 650828 322992
rect 650880 322980 650886 322992
rect 653398 322980 653404 322992
rect 650880 322952 653404 322980
rect 650880 322940 650886 322952
rect 653398 322940 653404 322952
rect 653456 322940 653462 322992
rect 42242 320220 42248 320272
rect 42300 320220 42306 320272
rect 42260 320124 42288 320220
rect 42260 320096 42656 320124
rect 42628 320000 42656 320096
rect 42610 319948 42616 320000
rect 42668 319948 42674 320000
rect 53834 317364 53840 317416
rect 53892 317404 53898 317416
rect 62114 317404 62120 317416
rect 53892 317376 62120 317404
rect 53892 317364 53898 317376
rect 62114 317364 62120 317376
rect 62172 317364 62178 317416
rect 53834 314712 53840 314764
rect 53892 314752 53898 314764
rect 62114 314752 62120 314764
rect 53892 314724 62120 314752
rect 53892 314712 53898 314724
rect 62114 314712 62120 314724
rect 62172 314712 62178 314764
rect 674374 311992 674380 312044
rect 674432 312032 674438 312044
rect 675478 312032 675484 312044
rect 674432 312004 675484 312032
rect 674432 311992 674438 312004
rect 675478 311992 675484 312004
rect 675536 311992 675542 312044
rect 676214 306348 676220 306400
rect 676272 306388 676278 306400
rect 676858 306388 676864 306400
rect 676272 306360 676864 306388
rect 676272 306348 676278 306360
rect 676858 306348 676864 306360
rect 676916 306348 676922 306400
rect 50522 305600 50528 305652
rect 50580 305640 50586 305652
rect 58802 305640 58808 305652
rect 50580 305612 58808 305640
rect 50580 305600 50586 305612
rect 58802 305600 58808 305612
rect 58860 305600 58866 305652
rect 675846 304852 675852 304904
rect 675904 304892 675910 304904
rect 676398 304892 676404 304904
rect 675904 304864 676404 304892
rect 675904 304852 675910 304864
rect 676398 304852 676404 304864
rect 676456 304852 676462 304904
rect 651374 303356 651380 303408
rect 651432 303396 651438 303408
rect 653398 303396 653404 303408
rect 651432 303368 653404 303396
rect 651432 303356 651438 303368
rect 653398 303356 653404 303368
rect 653456 303356 653462 303408
rect 651466 300772 651472 300824
rect 651524 300812 651530 300824
rect 658918 300812 658924 300824
rect 651524 300784 658924 300812
rect 651524 300772 651530 300784
rect 658918 300772 658924 300784
rect 658976 300772 658982 300824
rect 41138 299072 41144 299124
rect 41196 299112 41202 299124
rect 41690 299112 41696 299124
rect 41196 299084 41696 299112
rect 41196 299072 41202 299084
rect 41690 299072 41696 299084
rect 41748 299072 41754 299124
rect 651466 298120 651472 298172
rect 651524 298160 651530 298172
rect 660574 298160 660580 298172
rect 651524 298132 660580 298160
rect 651524 298120 651530 298132
rect 660574 298120 660580 298132
rect 660632 298120 660638 298172
rect 675846 298052 675852 298104
rect 675904 298092 675910 298104
rect 678238 298092 678244 298104
rect 675904 298064 678244 298092
rect 675904 298052 675910 298064
rect 678238 298052 678244 298064
rect 678296 298052 678302 298104
rect 651650 296760 651656 296812
rect 651708 296800 651714 296812
rect 651708 296772 654134 296800
rect 651708 296760 651714 296772
rect 654106 296732 654134 296772
rect 658918 296732 658924 296744
rect 654106 296704 658924 296732
rect 658918 296692 658924 296704
rect 658976 296692 658982 296744
rect 675478 296352 675484 296404
rect 675536 296352 675542 296404
rect 675294 296148 675300 296200
rect 675352 296148 675358 296200
rect 675312 295452 675340 296148
rect 675294 295400 675300 295452
rect 675352 295400 675358 295452
rect 675496 295248 675524 296352
rect 675478 295196 675484 295248
rect 675536 295196 675542 295248
rect 41322 294584 41328 294636
rect 41380 294624 41386 294636
rect 41690 294624 41696 294636
rect 41380 294596 41696 294624
rect 41380 294584 41386 294596
rect 41690 294584 41696 294596
rect 41748 294584 41754 294636
rect 42058 294448 42064 294500
rect 42116 294488 42122 294500
rect 42518 294488 42524 294500
rect 42116 294460 42524 294488
rect 42116 294448 42122 294460
rect 42518 294448 42524 294460
rect 42576 294448 42582 294500
rect 57422 294040 57428 294092
rect 57480 294080 57486 294092
rect 62114 294080 62120 294092
rect 57480 294052 62120 294080
rect 57480 294040 57486 294052
rect 62114 294040 62120 294052
rect 62172 294040 62178 294092
rect 651466 293972 651472 294024
rect 651524 294012 651530 294024
rect 664438 294012 664444 294024
rect 651524 293984 664444 294012
rect 651524 293972 651530 293984
rect 664438 293972 664444 293984
rect 664496 293972 664502 294024
rect 47578 293904 47584 293956
rect 47636 293944 47642 293956
rect 50522 293944 50528 293956
rect 47636 293916 50528 293944
rect 47636 293904 47642 293916
rect 50522 293904 50528 293916
rect 50580 293904 50586 293956
rect 40586 292544 40592 292596
rect 40644 292584 40650 292596
rect 41598 292584 41604 292596
rect 40644 292556 41604 292584
rect 40644 292544 40650 292556
rect 41598 292544 41604 292556
rect 41656 292544 41662 292596
rect 56042 292544 56048 292596
rect 56100 292584 56106 292596
rect 62758 292584 62764 292596
rect 56100 292556 62764 292584
rect 56100 292544 56106 292556
rect 62758 292544 62764 292556
rect 62816 292544 62822 292596
rect 651466 292544 651472 292596
rect 651524 292584 651530 292596
rect 660298 292584 660304 292596
rect 651524 292556 660304 292584
rect 651524 292544 651530 292556
rect 660298 292544 660304 292556
rect 660356 292544 660362 292596
rect 54478 292408 54484 292460
rect 54536 292448 54542 292460
rect 62114 292448 62120 292460
rect 54536 292420 62120 292448
rect 54536 292408 54542 292420
rect 62114 292408 62120 292420
rect 62172 292408 62178 292460
rect 35802 291320 35808 291372
rect 35860 291360 35866 291372
rect 41598 291360 41604 291372
rect 35860 291332 41604 291360
rect 35860 291320 35866 291332
rect 41598 291320 41604 291332
rect 41656 291320 41662 291372
rect 51718 291116 51724 291168
rect 51776 291156 51782 291168
rect 62114 291156 62120 291168
rect 51776 291128 62120 291156
rect 51776 291116 51782 291128
rect 62114 291116 62120 291128
rect 62172 291116 62178 291168
rect 649258 290776 649264 290828
rect 649316 290816 649322 290828
rect 651742 290816 651748 290828
rect 649316 290788 651748 290816
rect 649316 290776 649322 290788
rect 651742 290776 651748 290788
rect 651800 290776 651806 290828
rect 651466 289824 651472 289876
rect 651524 289864 651530 289876
rect 663058 289864 663064 289876
rect 651524 289836 663064 289864
rect 651524 289824 651530 289836
rect 663058 289824 663064 289836
rect 663116 289824 663122 289876
rect 51718 288464 51724 288516
rect 51776 288504 51782 288516
rect 62114 288504 62120 288516
rect 51776 288476 62120 288504
rect 51776 288464 51782 288476
rect 62114 288464 62120 288476
rect 62172 288464 62178 288516
rect 651466 288396 651472 288448
rect 651524 288436 651530 288448
rect 672166 288436 672172 288448
rect 651524 288408 672172 288436
rect 651524 288396 651530 288408
rect 672166 288396 672172 288408
rect 672224 288396 672230 288448
rect 33042 287648 33048 287700
rect 33100 287688 33106 287700
rect 41506 287688 41512 287700
rect 33100 287660 41512 287688
rect 33100 287648 33106 287660
rect 41506 287648 41512 287660
rect 41564 287648 41570 287700
rect 651466 287036 651472 287088
rect 651524 287076 651530 287088
rect 667750 287076 667756 287088
rect 651524 287048 667756 287076
rect 651524 287036 651530 287048
rect 667750 287036 667756 287048
rect 667808 287036 667814 287088
rect 674374 286628 674380 286680
rect 674432 286668 674438 286680
rect 675294 286668 675300 286680
rect 674432 286640 675300 286668
rect 674432 286628 674438 286640
rect 675294 286628 675300 286640
rect 675352 286628 675358 286680
rect 35158 286288 35164 286340
rect 35216 286328 35222 286340
rect 41690 286328 41696 286340
rect 35216 286300 41696 286328
rect 35216 286288 35222 286300
rect 41690 286288 41696 286300
rect 41748 286288 41754 286340
rect 42242 286288 42248 286340
rect 42300 286328 42306 286340
rect 42610 286328 42616 286340
rect 42300 286300 42616 286328
rect 42300 286288 42306 286300
rect 42610 286288 42616 286300
rect 42668 286288 42674 286340
rect 46382 285676 46388 285728
rect 46440 285716 46446 285728
rect 62114 285716 62120 285728
rect 46440 285688 62120 285716
rect 46440 285676 46446 285688
rect 62114 285676 62120 285688
rect 62172 285676 62178 285728
rect 651466 285676 651472 285728
rect 651524 285716 651530 285728
rect 667566 285716 667572 285728
rect 651524 285688 667572 285716
rect 651524 285676 651530 285688
rect 667566 285676 667572 285688
rect 667624 285676 667630 285728
rect 47762 284928 47768 284980
rect 47820 284968 47826 284980
rect 59998 284968 60004 284980
rect 47820 284940 60004 284968
rect 47820 284928 47826 284940
rect 59998 284928 60004 284940
rect 60056 284928 60062 284980
rect 45554 284316 45560 284368
rect 45612 284356 45618 284368
rect 62942 284356 62948 284368
rect 45612 284328 62948 284356
rect 45612 284316 45618 284328
rect 62942 284316 62948 284328
rect 63000 284316 63006 284368
rect 651466 284316 651472 284368
rect 651524 284356 651530 284368
rect 672350 284356 672356 284368
rect 651524 284328 672356 284356
rect 651524 284316 651530 284328
rect 672350 284316 672356 284328
rect 672408 284316 672414 284368
rect 651466 282888 651472 282940
rect 651524 282928 651530 282940
rect 667198 282928 667204 282940
rect 651524 282900 667204 282928
rect 651524 282888 651530 282900
rect 667198 282888 667204 282900
rect 667256 282888 667262 282940
rect 54478 280372 54484 280424
rect 54536 280412 54542 280424
rect 62114 280412 62120 280424
rect 54536 280384 62120 280412
rect 54536 280372 54542 280384
rect 62114 280372 62120 280384
rect 62172 280372 62178 280424
rect 53282 280168 53288 280220
rect 53340 280208 53346 280220
rect 62298 280208 62304 280220
rect 53340 280180 62304 280208
rect 53340 280168 53346 280180
rect 62298 280168 62304 280180
rect 62356 280168 62362 280220
rect 651466 280168 651472 280220
rect 651524 280208 651530 280220
rect 667382 280208 667388 280220
rect 651524 280180 667388 280208
rect 651524 280168 651530 280180
rect 667382 280168 667388 280180
rect 667440 280168 667446 280220
rect 62574 278672 62580 278724
rect 62632 278712 62638 278724
rect 671338 278712 671344 278724
rect 62632 278684 671344 278712
rect 62632 278672 62638 278684
rect 671338 278672 671344 278684
rect 671396 278672 671402 278724
rect 63310 278536 63316 278588
rect 63368 278576 63374 278588
rect 63368 278548 669314 278576
rect 63368 278536 63374 278548
rect 669286 278508 669314 278548
rect 671706 278508 671712 278520
rect 669286 278480 671712 278508
rect 671706 278468 671712 278480
rect 671764 278468 671770 278520
rect 58802 278400 58808 278452
rect 58860 278440 58866 278452
rect 650822 278440 650828 278452
rect 58860 278412 650828 278440
rect 58860 278400 58866 278412
rect 650822 278400 650828 278412
rect 650880 278400 650886 278452
rect 50522 278264 50528 278316
rect 50580 278304 50586 278316
rect 69198 278304 69204 278316
rect 50580 278276 69204 278304
rect 50580 278264 50586 278276
rect 69198 278264 69204 278276
rect 69256 278264 69262 278316
rect 649258 278304 649264 278316
rect 69676 278276 649264 278304
rect 59998 278128 60004 278180
rect 60056 278168 60062 278180
rect 69676 278168 69704 278276
rect 649258 278264 649264 278276
rect 649316 278264 649322 278316
rect 650638 278168 650644 278180
rect 60056 278140 69704 278168
rect 74506 278140 650644 278168
rect 60056 278128 60062 278140
rect 69198 277992 69204 278044
rect 69256 278032 69262 278044
rect 74506 278032 74534 278140
rect 650638 278128 650644 278140
rect 650696 278128 650702 278180
rect 69256 278004 74534 278032
rect 69256 277992 69262 278004
rect 45462 277380 45468 277432
rect 45520 277420 45526 277432
rect 637850 277420 637856 277432
rect 45520 277392 637856 277420
rect 45520 277380 45526 277392
rect 637850 277380 637856 277392
rect 637908 277380 637914 277432
rect 42242 277312 42248 277364
rect 42300 277352 42306 277364
rect 43346 277352 43352 277364
rect 42300 277324 43352 277352
rect 42300 277312 42306 277324
rect 43346 277312 43352 277324
rect 43404 277312 43410 277364
rect 487982 277176 487988 277228
rect 488040 277216 488046 277228
rect 565814 277216 565820 277228
rect 488040 277188 565820 277216
rect 488040 277176 488046 277188
rect 565814 277176 565820 277188
rect 565872 277176 565878 277228
rect 497918 277040 497924 277092
rect 497976 277080 497982 277092
rect 579982 277080 579988 277092
rect 497976 277052 579988 277080
rect 497976 277040 497982 277052
rect 579982 277040 579988 277052
rect 580040 277040 580046 277092
rect 511626 276904 511632 276956
rect 511684 276944 511690 276956
rect 600130 276944 600136 276956
rect 511684 276916 600136 276944
rect 511684 276904 511690 276916
rect 600130 276904 600136 276916
rect 600188 276904 600194 276956
rect 42242 276768 42248 276820
rect 42300 276808 42306 276820
rect 42610 276808 42616 276820
rect 42300 276780 42616 276808
rect 42300 276768 42306 276780
rect 42610 276768 42616 276780
rect 42668 276768 42674 276820
rect 514478 276768 514484 276820
rect 514536 276808 514542 276820
rect 603626 276808 603632 276820
rect 514536 276780 603632 276808
rect 514536 276768 514542 276780
rect 603626 276768 603632 276780
rect 603684 276768 603690 276820
rect 518342 276632 518348 276684
rect 518400 276672 518406 276684
rect 609606 276672 609612 276684
rect 518400 276644 609612 276672
rect 518400 276632 518406 276644
rect 609606 276632 609612 276644
rect 609664 276632 609670 276684
rect 479978 276496 479984 276548
rect 480036 276536 480042 276548
rect 555234 276536 555240 276548
rect 480036 276508 555240 276536
rect 480036 276496 480042 276508
rect 555234 276496 555240 276508
rect 555292 276496 555298 276548
rect 482830 276360 482836 276412
rect 482888 276400 482894 276412
rect 557534 276400 557540 276412
rect 482888 276372 557540 276400
rect 482888 276360 482894 276372
rect 557534 276360 557540 276372
rect 557592 276360 557598 276412
rect 477034 276224 477040 276276
rect 477092 276264 477098 276276
rect 550450 276264 550456 276276
rect 477092 276236 550456 276264
rect 477092 276224 477098 276236
rect 550450 276224 550456 276236
rect 550508 276224 550514 276276
rect 471606 276088 471612 276140
rect 471664 276128 471670 276140
rect 543366 276128 543372 276140
rect 471664 276100 543372 276128
rect 471664 276088 471670 276100
rect 543366 276088 543372 276100
rect 543424 276088 543430 276140
rect 107194 275952 107200 276004
rect 107252 275992 107258 276004
rect 163498 275992 163504 276004
rect 107252 275964 163504 275992
rect 107252 275952 107258 275964
rect 163498 275952 163504 275964
rect 163556 275952 163562 276004
rect 167546 275952 167552 276004
rect 167604 275992 167610 276004
rect 178678 275992 178684 276004
rect 167604 275964 178684 275992
rect 167604 275952 167610 275964
rect 178678 275952 178684 275964
rect 178736 275952 178742 276004
rect 185210 275952 185216 276004
rect 185268 275992 185274 276004
rect 221274 275992 221280 276004
rect 185268 275964 221280 275992
rect 185268 275952 185274 275964
rect 221274 275952 221280 275964
rect 221332 275952 221338 276004
rect 232498 275952 232504 276004
rect 232556 275992 232562 276004
rect 240042 275992 240048 276004
rect 232556 275964 240048 275992
rect 232556 275952 232562 275964
rect 240042 275952 240048 275964
rect 240100 275952 240106 276004
rect 410794 275952 410800 276004
rect 410852 275992 410858 276004
rect 455874 275992 455880 276004
rect 410852 275964 455880 275992
rect 410852 275952 410858 275964
rect 455874 275952 455880 275964
rect 455932 275952 455938 276004
rect 456058 275952 456064 276004
rect 456116 275992 456122 276004
rect 509050 275992 509056 276004
rect 456116 275964 509056 275992
rect 456116 275952 456122 275964
rect 509050 275952 509056 275964
rect 509108 275952 509114 276004
rect 513190 275952 513196 276004
rect 513248 275992 513254 276004
rect 601326 275992 601332 276004
rect 513248 275964 601332 275992
rect 513248 275952 513254 275964
rect 601326 275952 601332 275964
rect 601384 275952 601390 276004
rect 139118 275816 139124 275868
rect 139176 275856 139182 275868
rect 174262 275856 174268 275868
rect 139176 275828 174268 275856
rect 139176 275816 139182 275828
rect 174262 275816 174268 275828
rect 174320 275816 174326 275868
rect 178126 275816 178132 275868
rect 178184 275856 178190 275868
rect 216674 275856 216680 275868
rect 178184 275828 216680 275856
rect 178184 275816 178190 275828
rect 216674 275816 216680 275828
rect 216732 275816 216738 275868
rect 224218 275816 224224 275868
rect 224276 275856 224282 275868
rect 232682 275856 232688 275868
rect 224276 275828 232688 275856
rect 224276 275816 224282 275828
rect 232682 275816 232688 275828
rect 232740 275816 232746 275868
rect 236086 275816 236092 275868
rect 236144 275856 236150 275868
rect 250438 275856 250444 275868
rect 236144 275828 250444 275856
rect 236144 275816 236150 275828
rect 250438 275816 250444 275828
rect 250496 275816 250502 275868
rect 284570 275816 284576 275868
rect 284628 275856 284634 275868
rect 290090 275856 290096 275868
rect 284628 275828 290096 275856
rect 284628 275816 284634 275828
rect 290090 275816 290096 275828
rect 290148 275816 290154 275868
rect 430206 275816 430212 275868
rect 430264 275856 430270 275868
rect 484302 275856 484308 275868
rect 430264 275828 484308 275856
rect 430264 275816 430270 275828
rect 484302 275816 484308 275828
rect 484360 275816 484366 275868
rect 490558 275816 490564 275868
rect 490616 275856 490622 275868
rect 505554 275856 505560 275868
rect 490616 275828 505560 275856
rect 490616 275816 490622 275828
rect 505554 275816 505560 275828
rect 505612 275816 505618 275868
rect 522758 275816 522764 275868
rect 522816 275856 522822 275868
rect 615494 275856 615500 275868
rect 522816 275828 615500 275856
rect 522816 275816 522822 275828
rect 615494 275816 615500 275828
rect 615552 275816 615558 275868
rect 260926 275748 260932 275800
rect 260984 275788 260990 275800
rect 266354 275788 266360 275800
rect 260984 275760 266360 275788
rect 260984 275748 260990 275760
rect 266354 275748 266360 275760
rect 266412 275748 266418 275800
rect 93026 275680 93032 275732
rect 93084 275720 93090 275732
rect 152826 275720 152832 275732
rect 93084 275692 152832 275720
rect 93084 275680 93090 275692
rect 152826 275680 152832 275692
rect 152884 275680 152890 275732
rect 160462 275680 160468 275732
rect 160520 275720 160526 275732
rect 199562 275720 199568 275732
rect 160520 275692 199568 275720
rect 160520 275680 160526 275692
rect 199562 275680 199568 275692
rect 199620 275680 199626 275732
rect 217134 275680 217140 275732
rect 217192 275720 217198 275732
rect 224218 275720 224224 275732
rect 217192 275692 224224 275720
rect 217192 275680 217198 275692
rect 224218 275680 224224 275692
rect 224276 275680 224282 275732
rect 229002 275680 229008 275732
rect 229060 275720 229066 275732
rect 243722 275720 243728 275732
rect 229060 275692 243728 275720
rect 229060 275680 229066 275692
rect 243722 275680 243728 275692
rect 243780 275680 243786 275732
rect 250254 275680 250260 275732
rect 250312 275720 250318 275732
rect 259362 275720 259368 275732
rect 250312 275692 259368 275720
rect 250312 275680 250318 275692
rect 259362 275680 259368 275692
rect 259420 275680 259426 275732
rect 286870 275680 286876 275732
rect 286928 275720 286934 275732
rect 291838 275720 291844 275732
rect 286928 275692 291844 275720
rect 286928 275680 286934 275692
rect 291838 275680 291844 275692
rect 291896 275680 291902 275732
rect 445018 275680 445024 275732
rect 445076 275720 445082 275732
rect 498470 275720 498476 275732
rect 445076 275692 498476 275720
rect 445076 275680 445082 275692
rect 498470 275680 498476 275692
rect 498528 275680 498534 275732
rect 498838 275680 498844 275732
rect 498896 275720 498902 275732
rect 512638 275720 512644 275732
rect 498896 275692 512644 275720
rect 498896 275680 498902 275692
rect 512638 275680 512644 275692
rect 512696 275680 512702 275732
rect 528186 275680 528192 275732
rect 528244 275720 528250 275732
rect 622578 275720 622584 275732
rect 528244 275692 622584 275720
rect 528244 275680 528250 275692
rect 622578 275680 622584 275692
rect 622636 275680 622642 275732
rect 76466 275544 76472 275596
rect 76524 275584 76530 275596
rect 86218 275584 86224 275596
rect 76524 275556 86224 275584
rect 76524 275544 76530 275556
rect 86218 275544 86224 275556
rect 86276 275544 86282 275596
rect 90726 275544 90732 275596
rect 90784 275584 90790 275596
rect 154758 275584 154764 275596
rect 90784 275556 154764 275584
rect 90784 275544 90790 275556
rect 154758 275544 154764 275556
rect 154816 275544 154822 275596
rect 171042 275544 171048 275596
rect 171100 275584 171106 275596
rect 211430 275584 211436 275596
rect 171100 275556 211436 275584
rect 171100 275544 171106 275556
rect 211430 275544 211436 275556
rect 211488 275544 211494 275596
rect 218330 275544 218336 275596
rect 218388 275584 218394 275596
rect 233878 275584 233884 275596
rect 218388 275556 233884 275584
rect 218388 275544 218394 275556
rect 233878 275544 233884 275556
rect 233936 275544 233942 275596
rect 239582 275544 239588 275596
rect 239640 275584 239646 275596
rect 255958 275584 255964 275596
rect 239640 275556 255964 275584
rect 239640 275544 239646 275556
rect 255958 275544 255964 275556
rect 256016 275544 256022 275596
rect 257338 275544 257344 275596
rect 257396 275584 257402 275596
rect 262306 275584 262312 275596
rect 257396 275556 262312 275584
rect 257396 275544 257402 275556
rect 262306 275544 262312 275556
rect 262364 275544 262370 275596
rect 266814 275544 266820 275596
rect 266872 275584 266878 275596
rect 276474 275584 276480 275596
rect 266872 275556 276480 275584
rect 266872 275544 266878 275556
rect 276474 275544 276480 275556
rect 276532 275544 276538 275596
rect 363874 275544 363880 275596
rect 363932 275584 363938 275596
rect 388530 275584 388536 275596
rect 363932 275556 388536 275584
rect 363932 275544 363938 275556
rect 388530 275544 388536 275556
rect 388588 275544 388594 275596
rect 416406 275544 416412 275596
rect 416464 275584 416470 275596
rect 462958 275584 462964 275596
rect 416464 275556 462964 275584
rect 416464 275544 416470 275556
rect 462958 275544 462964 275556
rect 463016 275544 463022 275596
rect 463142 275544 463148 275596
rect 463200 275584 463206 275596
rect 516226 275584 516232 275596
rect 463200 275556 516232 275584
rect 463200 275544 463206 275556
rect 516226 275544 516232 275556
rect 516284 275544 516290 275596
rect 516778 275544 516784 275596
rect 516836 275584 516842 275596
rect 526806 275584 526812 275596
rect 516836 275556 526812 275584
rect 516836 275544 516842 275556
rect 526806 275544 526812 275556
rect 526864 275544 526870 275596
rect 532326 275544 532332 275596
rect 532384 275584 532390 275596
rect 629662 275584 629668 275596
rect 532384 275556 629668 275584
rect 532384 275544 532390 275556
rect 629662 275544 629668 275556
rect 629720 275544 629726 275596
rect 277486 275476 277492 275528
rect 277544 275516 277550 275528
rect 285122 275516 285128 275528
rect 277544 275488 285128 275516
rect 277544 275476 277550 275488
rect 285122 275476 285128 275488
rect 285180 275476 285186 275528
rect 100110 275408 100116 275460
rect 100168 275448 100174 275460
rect 100168 275420 142154 275448
rect 100168 275408 100174 275420
rect 71774 275272 71780 275324
rect 71832 275312 71838 275324
rect 141050 275312 141056 275324
rect 71832 275284 141056 275312
rect 71832 275272 71838 275284
rect 141050 275272 141056 275284
rect 141108 275272 141114 275324
rect 142126 275312 142154 275420
rect 156874 275408 156880 275460
rect 156932 275448 156938 275460
rect 156932 275420 161474 275448
rect 156932 275408 156938 275420
rect 159450 275312 159456 275324
rect 142126 275284 159456 275312
rect 159450 275272 159456 275284
rect 159508 275272 159514 275324
rect 161446 275312 161474 275420
rect 163958 275408 163964 275460
rect 164016 275448 164022 275460
rect 206370 275448 206376 275460
rect 164016 275420 206376 275448
rect 164016 275408 164022 275420
rect 206370 275408 206376 275420
rect 206428 275408 206434 275460
rect 221918 275408 221924 275460
rect 221976 275448 221982 275460
rect 243538 275448 243544 275460
rect 221976 275420 243544 275448
rect 221976 275408 221982 275420
rect 243538 275408 243544 275420
rect 243596 275408 243602 275460
rect 256142 275408 256148 275460
rect 256200 275448 256206 275460
rect 270126 275448 270132 275460
rect 256200 275420 270132 275448
rect 256200 275408 256206 275420
rect 270126 275408 270132 275420
rect 270184 275408 270190 275460
rect 358630 275408 358636 275460
rect 358688 275448 358694 275460
rect 381446 275448 381452 275460
rect 358688 275420 381452 275448
rect 358688 275408 358694 275420
rect 381446 275408 381452 275420
rect 381504 275408 381510 275460
rect 386046 275408 386052 275460
rect 386104 275448 386110 275460
rect 420454 275448 420460 275460
rect 386104 275420 420460 275448
rect 386104 275408 386110 275420
rect 420454 275408 420460 275420
rect 420512 275408 420518 275460
rect 435634 275408 435640 275460
rect 435692 275448 435698 275460
rect 481726 275448 481732 275460
rect 435692 275420 481732 275448
rect 435692 275408 435698 275420
rect 481726 275408 481732 275420
rect 481784 275408 481790 275460
rect 483658 275408 483664 275460
rect 483716 275448 483722 275460
rect 530394 275448 530400 275460
rect 483716 275420 530400 275448
rect 483716 275408 483722 275420
rect 530394 275408 530400 275420
rect 530452 275408 530458 275460
rect 537662 275408 537668 275460
rect 537720 275448 537726 275460
rect 636746 275448 636752 275460
rect 537720 275420 636752 275448
rect 537720 275408 537726 275420
rect 636746 275408 636752 275420
rect 636804 275408 636810 275460
rect 297542 275340 297548 275392
rect 297600 275380 297606 275392
rect 299566 275380 299572 275392
rect 297600 275352 299572 275380
rect 297600 275340 297606 275352
rect 299566 275340 299572 275352
rect 299624 275340 299630 275392
rect 299934 275340 299940 275392
rect 299992 275380 299998 275392
rect 301130 275380 301136 275392
rect 299992 275352 301136 275380
rect 299992 275340 299998 275352
rect 301130 275340 301136 275352
rect 301188 275340 301194 275392
rect 201034 275312 201040 275324
rect 161446 275284 201040 275312
rect 201034 275272 201040 275284
rect 201092 275272 201098 275324
rect 214834 275272 214840 275324
rect 214892 275312 214898 275324
rect 239398 275312 239404 275324
rect 214892 275284 239404 275312
rect 214892 275272 214898 275284
rect 239398 275272 239404 275284
rect 239456 275272 239462 275324
rect 243170 275272 243176 275324
rect 243228 275312 243234 275324
rect 256694 275312 256700 275324
rect 243228 275284 256700 275312
rect 243228 275272 243234 275284
rect 256694 275272 256700 275284
rect 256752 275272 256758 275324
rect 263226 275272 263232 275324
rect 263284 275312 263290 275324
rect 273254 275312 273260 275324
rect 263284 275284 273260 275312
rect 263284 275272 263290 275284
rect 273254 275272 273260 275284
rect 273312 275272 273318 275324
rect 276290 275272 276296 275324
rect 276348 275312 276354 275324
rect 283098 275312 283104 275324
rect 276348 275284 283104 275312
rect 276348 275272 276354 275284
rect 283098 275272 283104 275284
rect 283156 275272 283162 275324
rect 285674 275272 285680 275324
rect 285732 275312 285738 275324
rect 291286 275312 291292 275324
rect 285732 275284 291292 275312
rect 285732 275272 285738 275284
rect 291286 275272 291292 275284
rect 291344 275272 291350 275324
rect 291654 275272 291660 275324
rect 291712 275312 291718 275324
rect 295334 275312 295340 275324
rect 291712 275284 295340 275312
rect 291712 275272 291718 275284
rect 295334 275272 295340 275284
rect 295392 275272 295398 275324
rect 326430 275272 326436 275324
rect 326488 275312 326494 275324
rect 335354 275312 335360 275324
rect 326488 275284 335360 275312
rect 326488 275272 326494 275284
rect 335354 275272 335360 275284
rect 335412 275272 335418 275324
rect 371050 275272 371056 275324
rect 371108 275312 371114 275324
rect 399202 275312 399208 275324
rect 371108 275284 399208 275312
rect 371108 275272 371114 275284
rect 399202 275272 399208 275284
rect 399260 275272 399266 275324
rect 418798 275272 418804 275324
rect 418856 275312 418862 275324
rect 466546 275312 466552 275324
rect 418856 275284 466552 275312
rect 418856 275272 418862 275284
rect 466546 275272 466552 275284
rect 466604 275272 466610 275324
rect 467558 275272 467564 275324
rect 467616 275312 467622 275324
rect 537478 275312 537484 275324
rect 467616 275284 537484 275312
rect 467616 275272 467622 275284
rect 537478 275272 537484 275284
rect 537536 275272 537542 275324
rect 542262 275272 542268 275324
rect 542320 275312 542326 275324
rect 643830 275312 643836 275324
rect 542320 275284 643836 275312
rect 542320 275272 542326 275284
rect 643830 275272 643836 275284
rect 643888 275272 643894 275324
rect 298738 275204 298744 275256
rect 298796 275244 298802 275256
rect 300026 275244 300032 275256
rect 298796 275216 300032 275244
rect 298796 275204 298802 275216
rect 300026 275204 300032 275216
rect 300084 275204 300090 275256
rect 96614 275136 96620 275188
rect 96672 275176 96678 275188
rect 149606 275176 149612 275188
rect 96672 275148 149612 275176
rect 96672 275136 96678 275148
rect 149606 275136 149612 275148
rect 149664 275136 149670 275188
rect 153378 275136 153384 275188
rect 153436 275176 153442 275188
rect 169018 275176 169024 275188
rect 153436 275148 169024 275176
rect 153436 275136 153442 275148
rect 169018 275136 169024 275148
rect 169076 275136 169082 275188
rect 189994 275136 190000 275188
rect 190052 275176 190058 275188
rect 222930 275176 222936 275188
rect 190052 275148 222936 275176
rect 190052 275136 190058 275148
rect 222930 275136 222936 275148
rect 222988 275136 222994 275188
rect 292850 275136 292856 275188
rect 292908 275176 292914 275188
rect 295794 275176 295800 275188
rect 292908 275148 295800 275176
rect 292908 275136 292914 275148
rect 295794 275136 295800 275148
rect 295852 275136 295858 275188
rect 427078 275136 427084 275188
rect 427136 275176 427142 275188
rect 477218 275176 477224 275188
rect 427136 275148 477224 275176
rect 427136 275136 427142 275148
rect 477218 275136 477224 275148
rect 477276 275136 477282 275188
rect 481726 275136 481732 275188
rect 481784 275176 481790 275188
rect 491386 275176 491392 275188
rect 481784 275148 491392 275176
rect 481784 275136 481790 275148
rect 491386 275136 491392 275148
rect 491444 275136 491450 275188
rect 507486 275136 507492 275188
rect 507544 275176 507550 275188
rect 594242 275176 594248 275188
rect 507544 275148 594248 275176
rect 507544 275136 507550 275148
rect 594242 275136 594248 275148
rect 594300 275136 594306 275188
rect 269206 275068 269212 275120
rect 269264 275108 269270 275120
rect 274634 275108 274640 275120
rect 269264 275080 274640 275108
rect 269264 275068 269270 275080
rect 274634 275068 274640 275080
rect 274692 275068 274698 275120
rect 136818 275000 136824 275052
rect 136876 275040 136882 275052
rect 137646 275040 137652 275052
rect 136876 275012 137652 275040
rect 136876 275000 136882 275012
rect 137646 275000 137652 275012
rect 137704 275000 137710 275052
rect 146202 275000 146208 275052
rect 146260 275040 146266 275052
rect 185302 275040 185308 275052
rect 146260 275012 185308 275040
rect 146260 275000 146266 275012
rect 185302 275000 185308 275012
rect 185360 275000 185366 275052
rect 288066 275000 288072 275052
rect 288124 275040 288130 275052
rect 292850 275040 292856 275052
rect 288124 275012 292856 275040
rect 288124 275000 288130 275012
rect 292850 275000 292856 275012
rect 292908 275000 292914 275052
rect 420546 275000 420552 275052
rect 420604 275040 420610 275052
rect 470134 275040 470140 275052
rect 420604 275012 470140 275040
rect 420604 275000 420610 275012
rect 470134 275000 470140 275012
rect 470192 275000 470198 275052
rect 503438 275000 503444 275052
rect 503496 275040 503502 275052
rect 587066 275040 587072 275052
rect 503496 275012 587072 275040
rect 503496 275000 503502 275012
rect 587066 275000 587072 275012
rect 587124 275000 587130 275052
rect 81250 274932 81256 274984
rect 81308 274972 81314 274984
rect 81308 274944 84194 274972
rect 81308 274932 81314 274944
rect 84166 274904 84194 274944
rect 293954 274932 293960 274984
rect 294012 274972 294018 274984
rect 296806 274972 296812 274984
rect 294012 274944 296812 274972
rect 294012 274932 294018 274944
rect 296806 274932 296812 274944
rect 296864 274932 296870 274984
rect 145282 274904 145288 274916
rect 84166 274876 145288 274904
rect 145282 274864 145288 274876
rect 145340 274864 145346 274916
rect 149790 274864 149796 274916
rect 149848 274904 149854 274916
rect 189074 274904 189080 274916
rect 149848 274876 189080 274904
rect 149848 274864 149854 274876
rect 189074 274864 189080 274876
rect 189132 274864 189138 274916
rect 289262 274864 289268 274916
rect 289320 274904 289326 274916
rect 292666 274904 292672 274916
rect 289320 274876 292672 274904
rect 289320 274864 289326 274876
rect 292666 274864 292672 274876
rect 292724 274864 292730 274916
rect 473078 274864 473084 274916
rect 473136 274904 473142 274916
rect 544562 274904 544568 274916
rect 473136 274876 544568 274904
rect 473136 274864 473142 274876
rect 544562 274864 544568 274876
rect 544620 274864 544626 274916
rect 295150 274796 295156 274848
rect 295208 274836 295214 274848
rect 297450 274836 297456 274848
rect 295208 274808 297456 274836
rect 295208 274796 295214 274808
rect 297450 274796 297456 274808
rect 297508 274796 297514 274848
rect 128538 274728 128544 274780
rect 128596 274768 128602 274780
rect 168282 274768 168288 274780
rect 128596 274740 168288 274768
rect 128596 274728 128602 274740
rect 168282 274728 168288 274740
rect 168340 274728 168346 274780
rect 207750 274728 207756 274780
rect 207808 274768 207814 274780
rect 210694 274768 210700 274780
rect 207808 274740 210700 274768
rect 207808 274728 207814 274740
rect 210694 274728 210700 274740
rect 210752 274728 210758 274780
rect 476758 274728 476764 274780
rect 476816 274768 476822 274780
rect 523310 274768 523316 274780
rect 476816 274740 523316 274768
rect 476816 274728 476822 274740
rect 523310 274728 523316 274740
rect 523368 274728 523374 274780
rect 523678 274728 523684 274780
rect 523736 274768 523742 274780
rect 533890 274768 533896 274780
rect 523736 274740 533896 274768
rect 523736 274728 523742 274740
rect 533890 274728 533896 274740
rect 533948 274728 533954 274780
rect 534718 274728 534724 274780
rect 534776 274768 534782 274780
rect 540974 274768 540980 274780
rect 534776 274740 540980 274768
rect 534776 274728 534782 274740
rect 540974 274728 540980 274740
rect 541032 274728 541038 274780
rect 74166 274660 74172 274712
rect 74224 274700 74230 274712
rect 76834 274700 76840 274712
rect 74224 274672 76840 274700
rect 74224 274660 74230 274672
rect 76834 274660 76840 274672
rect 76892 274660 76898 274712
rect 85942 274660 85948 274712
rect 86000 274700 86006 274712
rect 90358 274700 90364 274712
rect 86000 274672 90364 274700
rect 86000 274660 86006 274672
rect 90358 274660 90364 274672
rect 90416 274660 90422 274712
rect 103698 274660 103704 274712
rect 103756 274700 103762 274712
rect 104802 274700 104808 274712
rect 103756 274672 104808 274700
rect 103756 274660 103762 274672
rect 104802 274660 104808 274672
rect 104860 274660 104866 274712
rect 110782 274660 110788 274712
rect 110840 274700 110846 274712
rect 111702 274700 111708 274712
rect 110840 274672 111708 274700
rect 110840 274660 110846 274672
rect 111702 274660 111708 274672
rect 111760 274660 111766 274712
rect 253842 274660 253848 274712
rect 253900 274700 253906 274712
rect 256878 274700 256884 274712
rect 253900 274672 256884 274700
rect 253900 274660 253906 274672
rect 256878 274660 256884 274672
rect 256936 274660 256942 274712
rect 275094 274660 275100 274712
rect 275152 274700 275158 274712
rect 278038 274700 278044 274712
rect 275152 274672 278044 274700
rect 275152 274660 275158 274672
rect 278038 274660 278044 274672
rect 278096 274660 278102 274712
rect 283374 274660 283380 274712
rect 283432 274700 283438 274712
rect 289170 274700 289176 274712
rect 283432 274672 289176 274700
rect 283432 274660 283438 274672
rect 289170 274660 289176 274672
rect 289228 274660 289234 274712
rect 290458 274660 290464 274712
rect 290516 274700 290522 274712
rect 294138 274700 294144 274712
rect 290516 274672 294144 274700
rect 290516 274660 290522 274672
rect 294138 274660 294144 274672
rect 294196 274660 294202 274712
rect 296346 274660 296352 274712
rect 296404 274700 296410 274712
rect 298370 274700 298376 274712
rect 296404 274672 298376 274700
rect 296404 274660 296410 274672
rect 298370 274660 298376 274672
rect 298428 274660 298434 274712
rect 303430 274660 303436 274712
rect 303488 274700 303494 274712
rect 303982 274700 303988 274712
rect 303488 274672 303988 274700
rect 303488 274660 303494 274672
rect 303982 274660 303988 274672
rect 304040 274660 304046 274712
rect 321186 274660 321192 274712
rect 321244 274700 321250 274712
rect 328270 274700 328276 274712
rect 321244 274672 328276 274700
rect 321244 274660 321250 274672
rect 328270 274660 328276 274672
rect 328328 274660 328334 274712
rect 114370 274592 114376 274644
rect 114428 274632 114434 274644
rect 171594 274632 171600 274644
rect 114428 274604 171600 274632
rect 114428 274592 114434 274604
rect 171594 274592 171600 274604
rect 171652 274592 171658 274644
rect 179322 274592 179328 274644
rect 179380 274632 179386 274644
rect 214558 274632 214564 274644
rect 179380 274604 214564 274632
rect 179380 274592 179386 274604
rect 214558 274592 214564 274604
rect 214616 274592 214622 274644
rect 409782 274592 409788 274644
rect 409840 274632 409846 274644
rect 453574 274632 453580 274644
rect 409840 274604 453580 274632
rect 409840 274592 409846 274604
rect 453574 274592 453580 274604
rect 453632 274592 453638 274644
rect 457438 274592 457444 274644
rect 457496 274632 457502 274644
rect 480714 274632 480720 274644
rect 457496 274604 480720 274632
rect 457496 274592 457502 274604
rect 480714 274592 480720 274604
rect 480772 274592 480778 274644
rect 486786 274592 486792 274644
rect 486844 274632 486850 274644
rect 563422 274632 563428 274644
rect 486844 274604 563428 274632
rect 486844 274592 486850 274604
rect 563422 274592 563428 274604
rect 563480 274592 563486 274644
rect 101306 274456 101312 274508
rect 101364 274496 101370 274508
rect 160922 274496 160928 274508
rect 101364 274468 160928 274496
rect 101364 274456 101370 274468
rect 160922 274456 160928 274468
rect 160980 274456 160986 274508
rect 168742 274456 168748 274508
rect 168800 274496 168806 274508
rect 208394 274496 208400 274508
rect 168800 274468 208400 274496
rect 168800 274456 168806 274468
rect 208394 274456 208400 274468
rect 208452 274456 208458 274508
rect 381538 274456 381544 274508
rect 381596 274496 381602 274508
rect 392118 274496 392124 274508
rect 381596 274468 392124 274496
rect 381596 274456 381602 274468
rect 392118 274456 392124 274468
rect 392176 274456 392182 274508
rect 413830 274456 413836 274508
rect 413888 274496 413894 274508
rect 460658 274496 460664 274508
rect 413888 274468 460664 274496
rect 413888 274456 413894 274468
rect 460658 274456 460664 274468
rect 460716 274456 460722 274508
rect 463234 274456 463240 274508
rect 463292 274496 463298 274508
rect 483658 274496 483664 274508
rect 463292 274468 483664 274496
rect 463292 274456 463298 274468
rect 483658 274456 483664 274468
rect 483716 274456 483722 274508
rect 488350 274456 488356 274508
rect 488408 274496 488414 274508
rect 567010 274496 567016 274508
rect 488408 274468 567016 274496
rect 488408 274456 488414 274468
rect 567010 274456 567016 274468
rect 567068 274456 567074 274508
rect 95418 274320 95424 274372
rect 95476 274360 95482 274372
rect 157610 274360 157616 274372
rect 95476 274332 157616 274360
rect 95476 274320 95482 274332
rect 157610 274320 157616 274332
rect 157668 274320 157674 274372
rect 159266 274320 159272 274372
rect 159324 274360 159330 274372
rect 202322 274360 202328 274372
rect 159324 274332 202328 274360
rect 159324 274320 159330 274332
rect 202322 274320 202328 274332
rect 202380 274320 202386 274372
rect 223114 274320 223120 274372
rect 223172 274360 223178 274372
rect 247218 274360 247224 274372
rect 223172 274332 247224 274360
rect 223172 274320 223178 274332
rect 247218 274320 247224 274332
rect 247276 274320 247282 274372
rect 369118 274320 369124 274372
rect 369176 274360 369182 274372
rect 387334 274360 387340 274372
rect 369176 274332 387340 274360
rect 369176 274320 369182 274332
rect 387334 274320 387340 274332
rect 387392 274320 387398 274372
rect 419074 274320 419080 274372
rect 419132 274360 419138 274372
rect 467742 274360 467748 274372
rect 419132 274332 467748 274360
rect 419132 274320 419138 274332
rect 467742 274320 467748 274332
rect 467800 274320 467806 274372
rect 506198 274320 506204 274372
rect 506256 274360 506262 274372
rect 591850 274360 591856 274372
rect 506256 274332 591856 274360
rect 506256 274320 506262 274332
rect 591850 274320 591856 274332
rect 591908 274320 591914 274372
rect 331950 274252 331956 274304
rect 332008 274292 332014 274304
rect 337746 274292 337752 274304
rect 332008 274264 337752 274292
rect 332008 274252 332014 274264
rect 337746 274252 337752 274264
rect 337804 274252 337810 274304
rect 67082 274184 67088 274236
rect 67140 274224 67146 274236
rect 130378 274224 130384 274236
rect 67140 274196 130384 274224
rect 67140 274184 67146 274196
rect 130378 274184 130384 274196
rect 130436 274184 130442 274236
rect 130838 274184 130844 274236
rect 130896 274224 130902 274236
rect 182450 274224 182456 274236
rect 130896 274196 182456 274224
rect 130896 274184 130902 274196
rect 182450 274184 182456 274196
rect 182508 274184 182514 274236
rect 192386 274184 192392 274236
rect 192444 274224 192450 274236
rect 224954 274224 224960 274236
rect 192444 274196 224960 274224
rect 192444 274184 192450 274196
rect 224954 274184 224960 274196
rect 225012 274184 225018 274236
rect 240042 274184 240048 274236
rect 240100 274224 240106 274236
rect 253934 274224 253940 274236
rect 240100 274196 253940 274224
rect 240100 274184 240106 274196
rect 253934 274184 253940 274196
rect 253992 274184 253998 274236
rect 359458 274184 359464 274236
rect 359516 274224 359522 274236
rect 380250 274224 380256 274236
rect 359516 274196 380256 274224
rect 359516 274184 359522 274196
rect 380250 274184 380256 274196
rect 380308 274184 380314 274236
rect 388990 274184 388996 274236
rect 389048 274224 389054 274236
rect 425146 274224 425152 274236
rect 389048 274196 425152 274224
rect 389048 274184 389054 274196
rect 425146 274184 425152 274196
rect 425204 274184 425210 274236
rect 425698 274184 425704 274236
rect 425756 274224 425762 274236
rect 474826 274224 474832 274236
rect 425756 274196 474832 274224
rect 425756 274184 425762 274196
rect 474826 274184 474832 274196
rect 474884 274184 474890 274236
rect 511810 274184 511816 274236
rect 511868 274224 511874 274236
rect 598934 274224 598940 274236
rect 511868 274196 598940 274224
rect 511868 274184 511874 274196
rect 598934 274184 598940 274196
rect 598992 274184 598998 274236
rect 77662 274048 77668 274100
rect 77720 274088 77726 274100
rect 144914 274088 144920 274100
rect 77720 274060 144920 274088
rect 77720 274048 77726 274060
rect 144914 274048 144920 274060
rect 144972 274048 144978 274100
rect 154482 274048 154488 274100
rect 154540 274088 154546 274100
rect 198090 274088 198096 274100
rect 154540 274060 198096 274088
rect 154540 274048 154546 274060
rect 198090 274048 198096 274060
rect 198148 274048 198154 274100
rect 210050 274048 210056 274100
rect 210108 274088 210114 274100
rect 237834 274088 237840 274100
rect 210108 274060 237840 274088
rect 210108 274048 210114 274060
rect 237834 274048 237840 274060
rect 237892 274048 237898 274100
rect 249058 274048 249064 274100
rect 249116 274088 249122 274100
rect 265250 274088 265256 274100
rect 249116 274060 265256 274088
rect 249116 274048 249122 274060
rect 265250 274048 265256 274060
rect 265308 274048 265314 274100
rect 266354 274048 266360 274100
rect 266412 274088 266418 274100
rect 273530 274088 273536 274100
rect 266412 274060 273536 274088
rect 266412 274048 266418 274060
rect 273530 274048 273536 274060
rect 273588 274048 273594 274100
rect 278590 274048 278596 274100
rect 278648 274088 278654 274100
rect 285858 274088 285864 274100
rect 278648 274060 285864 274088
rect 278648 274048 278654 274060
rect 285858 274048 285864 274060
rect 285916 274048 285922 274100
rect 337746 274048 337752 274100
rect 337804 274088 337810 274100
rect 351914 274088 351920 274100
rect 337804 274060 351920 274088
rect 337804 274048 337810 274060
rect 351914 274048 351920 274060
rect 351972 274048 351978 274100
rect 353938 274048 353944 274100
rect 353996 274088 354002 274100
rect 369578 274088 369584 274100
rect 353996 274060 369584 274088
rect 353996 274048 354002 274060
rect 369578 274048 369584 274060
rect 369636 274048 369642 274100
rect 373258 274048 373264 274100
rect 373316 274088 373322 274100
rect 400306 274088 400312 274100
rect 373316 274060 400312 274088
rect 373316 274048 373322 274060
rect 400306 274048 400312 274060
rect 400364 274048 400370 274100
rect 401502 274048 401508 274100
rect 401560 274088 401566 274100
rect 442902 274088 442908 274100
rect 401560 274060 442908 274088
rect 401560 274048 401566 274060
rect 442902 274048 442908 274060
rect 442960 274048 442966 274100
rect 451182 274048 451188 274100
rect 451240 274088 451246 274100
rect 513834 274088 513840 274100
rect 451240 274060 513840 274088
rect 451240 274048 451246 274060
rect 513834 274048 513840 274060
rect 513892 274048 513898 274100
rect 536742 274048 536748 274100
rect 536800 274088 536806 274100
rect 634354 274088 634360 274100
rect 536800 274060 634360 274088
rect 536800 274048 536806 274060
rect 634354 274048 634360 274060
rect 634412 274048 634418 274100
rect 69382 273912 69388 273964
rect 69440 273952 69446 273964
rect 139394 273952 139400 273964
rect 69440 273924 139400 273952
rect 69440 273912 69446 273924
rect 139394 273912 139400 273924
rect 139452 273912 139458 273964
rect 148594 273912 148600 273964
rect 148652 273952 148658 273964
rect 194778 273952 194784 273964
rect 148652 273924 194784 273952
rect 148652 273912 148658 273924
rect 194778 273912 194784 273924
rect 194836 273912 194842 273964
rect 208854 273912 208860 273964
rect 208912 273952 208918 273964
rect 237466 273952 237472 273964
rect 208912 273924 237472 273952
rect 208912 273912 208918 273924
rect 237466 273912 237472 273924
rect 237524 273912 237530 273964
rect 238478 273912 238484 273964
rect 238536 273952 238542 273964
rect 238536 273924 238754 273952
rect 238536 273912 238542 273924
rect 88334 273776 88340 273828
rect 88392 273816 88398 273828
rect 119338 273816 119344 273828
rect 88392 273788 119344 273816
rect 88392 273776 88398 273788
rect 119338 273776 119344 273788
rect 119396 273776 119402 273828
rect 120258 273776 120264 273828
rect 120316 273816 120322 273828
rect 175274 273816 175280 273828
rect 120316 273788 175280 273816
rect 120316 273776 120322 273788
rect 175274 273776 175280 273788
rect 175332 273776 175338 273828
rect 193490 273776 193496 273828
rect 193548 273816 193554 273828
rect 226426 273816 226432 273828
rect 193548 273788 226432 273816
rect 193548 273776 193554 273788
rect 226426 273776 226432 273788
rect 226484 273776 226490 273828
rect 238726 273816 238754 273924
rect 271506 273912 271512 273964
rect 271564 273952 271570 273964
rect 280338 273952 280344 273964
rect 271564 273924 280344 273952
rect 271564 273912 271570 273924
rect 280338 273912 280344 273924
rect 280396 273912 280402 273964
rect 322750 273912 322756 273964
rect 322808 273952 322814 273964
rect 330570 273952 330576 273964
rect 322808 273924 330576 273952
rect 322808 273912 322814 273924
rect 330570 273912 330576 273924
rect 330628 273912 330634 273964
rect 335262 273912 335268 273964
rect 335320 273952 335326 273964
rect 348326 273952 348332 273964
rect 335320 273924 348332 273952
rect 335320 273912 335326 273924
rect 348326 273912 348332 273924
rect 348384 273912 348390 273964
rect 350350 273912 350356 273964
rect 350408 273952 350414 273964
rect 368474 273952 368480 273964
rect 350408 273924 368480 273952
rect 350408 273912 350414 273924
rect 368474 273912 368480 273924
rect 368532 273912 368538 273964
rect 377674 273912 377680 273964
rect 377732 273952 377738 273964
rect 408586 273952 408592 273964
rect 377732 273924 408592 273952
rect 377732 273912 377738 273924
rect 408586 273912 408592 273924
rect 408644 273912 408650 273964
rect 422110 273912 422116 273964
rect 422168 273952 422174 273964
rect 472434 273952 472440 273964
rect 422168 273924 472440 273952
rect 422168 273912 422174 273924
rect 472434 273912 472440 273924
rect 472492 273912 472498 273964
rect 474642 273912 474648 273964
rect 474700 273952 474706 273964
rect 545758 273952 545764 273964
rect 474700 273924 545764 273952
rect 474700 273912 474706 273924
rect 545758 273912 545764 273924
rect 545816 273912 545822 273964
rect 545942 273912 545948 273964
rect 546000 273952 546006 273964
rect 639138 273952 639144 273964
rect 546000 273924 639144 273952
rect 546000 273912 546006 273924
rect 639138 273912 639144 273924
rect 639196 273912 639202 273964
rect 258074 273816 258080 273828
rect 238726 273788 258080 273816
rect 258074 273776 258080 273788
rect 258132 273776 258138 273828
rect 396994 273776 397000 273828
rect 397052 273816 397058 273828
rect 435818 273816 435824 273828
rect 397052 273788 435824 273816
rect 397052 273776 397058 273788
rect 435818 273776 435824 273788
rect 435876 273776 435882 273828
rect 438118 273776 438124 273828
rect 438176 273816 438182 273828
rect 473630 273816 473636 273828
rect 438176 273788 473636 273816
rect 438176 273776 438182 273788
rect 473630 273776 473636 273788
rect 473688 273776 473694 273828
rect 481358 273776 481364 273828
rect 481416 273816 481422 273828
rect 556338 273816 556344 273828
rect 481416 273788 556344 273816
rect 481416 273776 481422 273788
rect 556338 273776 556344 273788
rect 556396 273776 556402 273828
rect 556798 273776 556804 273828
rect 556856 273816 556862 273828
rect 590654 273816 590660 273828
rect 556856 273788 590660 273816
rect 556856 273776 556862 273788
rect 590654 273776 590660 273788
rect 590712 273776 590718 273828
rect 119062 273640 119068 273692
rect 119120 273680 119126 273692
rect 173250 273680 173256 273692
rect 119120 273652 173256 273680
rect 119120 273640 119126 273652
rect 173250 273640 173256 273652
rect 173308 273640 173314 273692
rect 447778 273640 447784 273692
rect 447836 273680 447842 273692
rect 481910 273680 481916 273692
rect 447836 273652 481916 273680
rect 447836 273640 447842 273652
rect 481910 273640 481916 273652
rect 481968 273640 481974 273692
rect 484210 273640 484216 273692
rect 484268 273680 484274 273692
rect 559926 273680 559932 273692
rect 484268 273652 559932 273680
rect 484268 273640 484274 273652
rect 559926 273640 559932 273652
rect 559984 273640 559990 273692
rect 132034 273504 132040 273556
rect 132092 273544 132098 273556
rect 153838 273544 153844 273556
rect 132092 273516 153844 273544
rect 132092 273504 132098 273516
rect 153838 273504 153844 273516
rect 153896 273504 153902 273556
rect 259362 273504 259368 273556
rect 259420 273544 259426 273556
rect 266354 273544 266360 273556
rect 259420 273516 266360 273544
rect 259420 273504 259426 273516
rect 266354 273504 266360 273516
rect 266412 273504 266418 273556
rect 440878 273504 440884 273556
rect 440936 273544 440942 273556
rect 471238 273544 471244 273556
rect 440936 273516 471244 273544
rect 440936 273504 440942 273516
rect 471238 273504 471244 273516
rect 471296 273504 471302 273556
rect 478690 273504 478696 273556
rect 478748 273544 478754 273556
rect 552842 273544 552848 273556
rect 478748 273516 552848 273544
rect 478748 273504 478754 273516
rect 552842 273504 552848 273516
rect 552900 273504 552906 273556
rect 145282 273368 145288 273420
rect 145340 273408 145346 273420
rect 147858 273408 147864 273420
rect 145340 273380 147864 273408
rect 145340 273368 145346 273380
rect 147858 273368 147864 273380
rect 147916 273368 147922 273420
rect 476022 273368 476028 273420
rect 476080 273408 476086 273420
rect 549254 273408 549260 273420
rect 476080 273380 549260 273408
rect 476080 273368 476086 273380
rect 549254 273368 549260 273380
rect 549312 273368 549318 273420
rect 549898 273368 549904 273420
rect 549956 273408 549962 273420
rect 583570 273408 583576 273420
rect 549956 273380 583576 273408
rect 549956 273368 549962 273380
rect 583570 273368 583576 273380
rect 583628 273368 583634 273420
rect 460014 273300 460020 273352
rect 460072 273340 460078 273352
rect 461394 273340 461400 273352
rect 460072 273312 461400 273340
rect 460072 273300 460078 273312
rect 461394 273300 461400 273312
rect 461452 273300 461458 273352
rect 327718 273232 327724 273284
rect 327776 273272 327782 273284
rect 329466 273272 329472 273284
rect 327776 273244 329472 273272
rect 327776 273232 327782 273244
rect 329466 273232 329472 273244
rect 329524 273232 329530 273284
rect 42426 273164 42432 273216
rect 42484 273204 42490 273216
rect 42978 273204 42984 273216
rect 42484 273176 42984 273204
rect 42484 273164 42490 273176
rect 42978 273164 42984 273176
rect 43036 273164 43042 273216
rect 108390 273164 108396 273216
rect 108448 273204 108454 273216
rect 165890 273204 165896 273216
rect 108448 273176 165896 273204
rect 108448 273164 108454 273176
rect 165890 273164 165896 273176
rect 165948 273164 165954 273216
rect 186406 273164 186412 273216
rect 186464 273204 186470 273216
rect 218698 273204 218704 273216
rect 186464 273176 218704 273204
rect 186464 273164 186470 273176
rect 218698 273164 218704 273176
rect 218756 273164 218762 273216
rect 362770 273164 362776 273216
rect 362828 273204 362834 273216
rect 385862 273204 385868 273216
rect 362828 273176 385868 273204
rect 362828 273164 362834 273176
rect 385862 273164 385868 273176
rect 385920 273164 385926 273216
rect 400030 273164 400036 273216
rect 400088 273204 400094 273216
rect 439314 273204 439320 273216
rect 400088 273176 439320 273204
rect 400088 273164 400094 273176
rect 439314 273164 439320 273176
rect 439372 273164 439378 273216
rect 444006 273164 444012 273216
rect 444064 273204 444070 273216
rect 503162 273204 503168 273216
rect 444064 273176 503168 273204
rect 444064 273164 444070 273176
rect 503162 273164 503168 273176
rect 503220 273164 503226 273216
rect 504174 273164 504180 273216
rect 504232 273204 504238 273216
rect 511442 273204 511448 273216
rect 504232 273176 511448 273204
rect 504232 273164 504238 273176
rect 511442 273164 511448 273176
rect 511500 273164 511506 273216
rect 515398 273164 515404 273216
rect 515456 273204 515462 273216
rect 519722 273204 519728 273216
rect 515456 273176 519728 273204
rect 515456 273164 515462 273176
rect 519722 273164 519728 273176
rect 519780 273164 519786 273216
rect 521470 273164 521476 273216
rect 521528 273204 521534 273216
rect 614298 273204 614304 273216
rect 521528 273176 614304 273204
rect 521528 273164 521534 273176
rect 614298 273164 614304 273176
rect 614356 273164 614362 273216
rect 102502 273028 102508 273080
rect 102560 273068 102566 273080
rect 162854 273068 162860 273080
rect 102560 273040 162860 273068
rect 102560 273028 102566 273040
rect 162854 273028 162860 273040
rect 162912 273028 162918 273080
rect 172238 273028 172244 273080
rect 172296 273068 172302 273080
rect 209774 273068 209780 273080
rect 172296 273040 209780 273068
rect 172296 273028 172302 273040
rect 209774 273028 209780 273040
rect 209832 273028 209838 273080
rect 219526 273028 219532 273080
rect 219584 273068 219590 273080
rect 244550 273068 244556 273080
rect 219584 273040 244556 273068
rect 219584 273028 219590 273040
rect 244550 273028 244556 273040
rect 244608 273028 244614 273080
rect 280982 273028 280988 273080
rect 281040 273068 281046 273080
rect 286318 273068 286324 273080
rect 281040 273040 286324 273068
rect 281040 273028 281046 273040
rect 286318 273028 286324 273040
rect 286376 273028 286382 273080
rect 361206 273028 361212 273080
rect 361264 273068 361270 273080
rect 384942 273068 384948 273080
rect 361264 273040 384948 273068
rect 361264 273028 361270 273040
rect 384942 273028 384948 273040
rect 385000 273028 385006 273080
rect 385678 273028 385684 273080
rect 385736 273068 385742 273080
rect 395614 273068 395620 273080
rect 385736 273040 395620 273068
rect 385736 273028 385742 273040
rect 395614 273028 395620 273040
rect 395672 273028 395678 273080
rect 404170 273028 404176 273080
rect 404228 273068 404234 273080
rect 446490 273068 446496 273080
rect 404228 273040 446496 273068
rect 404228 273028 404234 273040
rect 446490 273028 446496 273040
rect 446548 273028 446554 273080
rect 446858 273028 446864 273080
rect 446916 273068 446922 273080
rect 507946 273068 507952 273080
rect 446916 273040 507952 273068
rect 446916 273028 446922 273040
rect 507946 273028 507952 273040
rect 508004 273028 508010 273080
rect 518526 273068 518532 273080
rect 509206 273040 518532 273068
rect 94222 272892 94228 272944
rect 94280 272932 94286 272944
rect 155954 272932 155960 272944
rect 94280 272904 155960 272932
rect 94280 272892 94286 272904
rect 155954 272892 155960 272904
rect 156012 272892 156018 272944
rect 166350 272892 166356 272944
rect 166408 272932 166414 272944
rect 207290 272932 207296 272944
rect 166408 272904 207296 272932
rect 166408 272892 166414 272904
rect 207290 272892 207296 272904
rect 207348 272892 207354 272944
rect 211246 272892 211252 272944
rect 211304 272932 211310 272944
rect 220078 272932 220084 272944
rect 211304 272904 220084 272932
rect 211304 272892 211310 272904
rect 220078 272892 220084 272904
rect 220136 272892 220142 272944
rect 220722 272892 220728 272944
rect 220780 272932 220786 272944
rect 245746 272932 245752 272944
rect 220780 272904 245752 272932
rect 220780 272892 220786 272904
rect 245746 272892 245752 272904
rect 245804 272892 245810 272944
rect 247862 272892 247868 272944
rect 247920 272932 247926 272944
rect 264238 272932 264244 272944
rect 247920 272904 264244 272932
rect 247920 272892 247926 272904
rect 264238 272892 264244 272904
rect 264296 272892 264302 272944
rect 333790 272892 333796 272944
rect 333848 272932 333854 272944
rect 345934 272932 345940 272944
rect 333848 272904 345940 272932
rect 333848 272892 333854 272904
rect 345934 272892 345940 272904
rect 345992 272892 345998 272944
rect 348418 272892 348424 272944
rect 348476 272932 348482 272944
rect 362494 272932 362500 272944
rect 348476 272904 362500 272932
rect 348476 272892 348482 272904
rect 362494 272892 362500 272904
rect 362552 272892 362558 272944
rect 365438 272892 365444 272944
rect 365496 272932 365502 272944
rect 390922 272932 390928 272944
rect 365496 272904 390928 272932
rect 365496 272892 365502 272904
rect 390922 272892 390928 272904
rect 390980 272892 390986 272944
rect 405550 272892 405556 272944
rect 405608 272932 405614 272944
rect 448790 272932 448796 272944
rect 405608 272904 448796 272932
rect 405608 272892 405614 272904
rect 448790 272892 448796 272904
rect 448848 272892 448854 272944
rect 455322 272892 455328 272944
rect 455380 272932 455386 272944
rect 457254 272932 457260 272944
rect 455380 272904 457260 272932
rect 455380 272892 455386 272904
rect 457254 272892 457260 272904
rect 457312 272892 457318 272944
rect 457990 272892 457996 272944
rect 458048 272932 458054 272944
rect 465902 272932 465908 272944
rect 458048 272904 465908 272932
rect 458048 272892 458054 272904
rect 465902 272892 465908 272904
rect 465960 272892 465966 272944
rect 466086 272892 466092 272944
rect 466144 272932 466150 272944
rect 509206 272932 509234 273040
rect 518526 273028 518532 273040
rect 518584 273028 518590 273080
rect 518710 273028 518716 273080
rect 518768 273068 518774 273080
rect 569402 273068 569408 273080
rect 518768 273040 569408 273068
rect 518768 273028 518774 273040
rect 569402 273028 569408 273040
rect 569460 273028 569466 273080
rect 515030 272932 515036 272944
rect 466144 272904 509234 272932
rect 512104 272904 515036 272932
rect 466144 272892 466150 272904
rect 82446 272756 82452 272808
rect 82504 272796 82510 272808
rect 148410 272796 148416 272808
rect 82504 272768 148416 272796
rect 82504 272756 82510 272768
rect 148410 272756 148416 272768
rect 148468 272756 148474 272808
rect 155678 272756 155684 272808
rect 155736 272796 155742 272808
rect 200114 272796 200120 272808
rect 155736 272768 200120 272796
rect 155736 272756 155742 272768
rect 200114 272756 200120 272768
rect 200172 272756 200178 272808
rect 205358 272756 205364 272808
rect 205416 272796 205422 272808
rect 234798 272796 234804 272808
rect 205416 272768 234804 272796
rect 205416 272756 205422 272768
rect 234798 272756 234804 272768
rect 234856 272756 234862 272808
rect 245378 272756 245384 272808
rect 245436 272796 245442 272808
rect 245436 272768 258074 272796
rect 245436 272756 245442 272768
rect 72970 272620 72976 272672
rect 73028 272660 73034 272672
rect 142154 272660 142160 272672
rect 73028 272632 142160 272660
rect 73028 272620 73034 272632
rect 142154 272620 142160 272632
rect 142212 272620 142218 272672
rect 142706 272620 142712 272672
rect 142764 272660 142770 272672
rect 145558 272660 145564 272672
rect 142764 272632 145564 272660
rect 142764 272620 142770 272632
rect 145558 272620 145564 272632
rect 145616 272620 145622 272672
rect 147398 272620 147404 272672
rect 147456 272660 147462 272672
rect 193214 272660 193220 272672
rect 147456 272632 193220 272660
rect 147456 272620 147462 272632
rect 193214 272620 193220 272632
rect 193272 272620 193278 272672
rect 197078 272620 197084 272672
rect 197136 272660 197142 272672
rect 229094 272660 229100 272672
rect 197136 272632 229100 272660
rect 197136 272620 197142 272632
rect 229094 272620 229100 272632
rect 229152 272620 229158 272672
rect 233694 272620 233700 272672
rect 233752 272660 233758 272672
rect 254394 272660 254400 272672
rect 233752 272632 254400 272660
rect 233752 272620 233758 272632
rect 254394 272620 254400 272632
rect 254452 272620 254458 272672
rect 258046 272660 258074 272768
rect 262306 272756 262312 272808
rect 262364 272796 262370 272808
rect 270954 272796 270960 272808
rect 262364 272768 270960 272796
rect 262364 272756 262370 272768
rect 270954 272756 270960 272768
rect 271012 272756 271018 272808
rect 273898 272756 273904 272808
rect 273956 272796 273962 272808
rect 282914 272796 282920 272808
rect 273956 272768 282920 272796
rect 273956 272756 273962 272768
rect 282914 272756 282920 272768
rect 282972 272756 282978 272808
rect 325326 272756 325332 272808
rect 325384 272796 325390 272808
rect 332962 272796 332968 272808
rect 325384 272768 332968 272796
rect 325384 272756 325390 272768
rect 332962 272756 332968 272768
rect 333020 272756 333026 272808
rect 344646 272756 344652 272808
rect 344704 272796 344710 272808
rect 361390 272796 361396 272808
rect 344704 272768 361396 272796
rect 344704 272756 344710 272768
rect 361390 272756 361396 272768
rect 361448 272756 361454 272808
rect 362218 272756 362224 272808
rect 362276 272796 362282 272808
rect 370314 272796 370320 272808
rect 362276 272768 370320 272796
rect 362276 272756 362282 272768
rect 370314 272756 370320 272768
rect 370372 272756 370378 272808
rect 370498 272756 370504 272808
rect 370556 272796 370562 272808
rect 396810 272796 396816 272808
rect 370556 272768 396816 272796
rect 370556 272756 370562 272768
rect 396810 272756 396816 272768
rect 396868 272756 396874 272808
rect 406838 272756 406844 272808
rect 406896 272796 406902 272808
rect 449986 272796 449992 272808
rect 406896 272768 449992 272796
rect 406896 272756 406902 272768
rect 449986 272756 449992 272768
rect 450044 272756 450050 272808
rect 452286 272756 452292 272808
rect 452344 272796 452350 272808
rect 512104 272796 512132 272904
rect 515030 272892 515036 272904
rect 515088 272892 515094 272944
rect 532510 272892 532516 272944
rect 532568 272932 532574 272944
rect 532568 272904 538904 272932
rect 532568 272892 532574 272904
rect 452344 272768 512132 272796
rect 452344 272756 452350 272768
rect 513742 272756 513748 272808
rect 513800 272796 513806 272808
rect 525610 272796 525616 272808
rect 513800 272768 525616 272796
rect 513800 272756 513806 272768
rect 525610 272756 525616 272768
rect 525668 272756 525674 272808
rect 529842 272756 529848 272808
rect 529900 272796 529906 272808
rect 532878 272796 532884 272808
rect 529900 272768 532884 272796
rect 529900 272756 529906 272768
rect 532878 272756 532884 272768
rect 532936 272756 532942 272808
rect 533706 272756 533712 272808
rect 533764 272796 533770 272808
rect 538674 272796 538680 272808
rect 533764 272768 538680 272796
rect 533764 272756 533770 272768
rect 538674 272756 538680 272768
rect 538732 272756 538738 272808
rect 538876 272796 538904 272904
rect 539042 272892 539048 272944
rect 539100 272932 539106 272944
rect 624970 272932 624976 272944
rect 539100 272904 624976 272932
rect 539100 272892 539106 272904
rect 624970 272892 624976 272904
rect 625028 272892 625034 272944
rect 632054 272932 632060 272944
rect 628668 272904 632060 272932
rect 628466 272796 628472 272808
rect 538876 272768 628472 272796
rect 628466 272756 628472 272768
rect 628524 272756 628530 272808
rect 262674 272660 262680 272672
rect 258046 272632 262680 272660
rect 262674 272620 262680 272632
rect 262732 272620 262738 272672
rect 264422 272620 264428 272672
rect 264480 272660 264486 272672
rect 276014 272660 276020 272672
rect 264480 272632 276020 272660
rect 264480 272620 264486 272632
rect 276014 272620 276020 272632
rect 276072 272620 276078 272672
rect 324038 272620 324044 272672
rect 324096 272660 324102 272672
rect 331766 272660 331772 272672
rect 324096 272632 331772 272660
rect 324096 272620 324102 272632
rect 331766 272620 331772 272632
rect 331824 272620 331830 272672
rect 332318 272620 332324 272672
rect 332376 272660 332382 272672
rect 343634 272660 343640 272672
rect 332376 272632 343640 272660
rect 332376 272620 332382 272632
rect 343634 272620 343640 272632
rect 343692 272620 343698 272672
rect 346210 272620 346216 272672
rect 346268 272660 346274 272672
rect 363690 272660 363696 272672
rect 346268 272632 363696 272660
rect 346268 272620 346274 272632
rect 363690 272620 363696 272632
rect 363748 272620 363754 272672
rect 376110 272620 376116 272672
rect 376168 272660 376174 272672
rect 406286 272660 406292 272672
rect 376168 272632 406292 272660
rect 376168 272620 376174 272632
rect 406286 272620 406292 272632
rect 406344 272620 406350 272672
rect 412266 272620 412272 272672
rect 412324 272660 412330 272672
rect 457070 272660 457076 272672
rect 412324 272632 457076 272660
rect 412324 272620 412330 272632
rect 457070 272620 457076 272632
rect 457128 272620 457134 272672
rect 457254 272620 457260 272672
rect 457312 272660 457318 272672
rect 460014 272660 460020 272672
rect 457312 272632 460020 272660
rect 457312 272620 457318 272632
rect 460014 272620 460020 272632
rect 460072 272620 460078 272672
rect 460198 272620 460204 272672
rect 460256 272660 460262 272672
rect 460256 272632 465764 272660
rect 460256 272620 460262 272632
rect 319070 272552 319076 272604
rect 319128 272592 319134 272604
rect 319622 272592 319628 272604
rect 319128 272564 319628 272592
rect 319128 272552 319134 272564
rect 319622 272552 319628 272564
rect 319680 272552 319686 272604
rect 65886 272484 65892 272536
rect 65944 272524 65950 272536
rect 136818 272524 136824 272536
rect 65944 272496 136824 272524
rect 65944 272484 65950 272496
rect 136818 272484 136824 272496
rect 136876 272484 136882 272536
rect 137922 272484 137928 272536
rect 137980 272524 137986 272536
rect 137980 272496 180794 272524
rect 137980 272484 137986 272496
rect 116670 272348 116676 272400
rect 116728 272388 116734 272400
rect 172514 272388 172520 272400
rect 116728 272360 172520 272388
rect 116728 272348 116734 272360
rect 172514 272348 172520 272360
rect 172572 272348 172578 272400
rect 180766 272388 180794 272496
rect 181714 272484 181720 272536
rect 181772 272524 181778 272536
rect 186958 272524 186964 272536
rect 181772 272496 186964 272524
rect 181772 272484 181778 272496
rect 186958 272484 186964 272496
rect 187016 272484 187022 272536
rect 195882 272484 195888 272536
rect 195940 272524 195946 272536
rect 227898 272524 227904 272536
rect 195940 272496 227904 272524
rect 195940 272484 195946 272496
rect 227898 272484 227904 272496
rect 227956 272484 227962 272536
rect 228082 272484 228088 272536
rect 228140 272524 228146 272536
rect 249058 272524 249064 272536
rect 228140 272496 249064 272524
rect 228140 272484 228146 272496
rect 249058 272484 249064 272496
rect 249116 272484 249122 272536
rect 254946 272484 254952 272536
rect 255004 272524 255010 272536
rect 269298 272524 269304 272536
rect 255004 272496 269304 272524
rect 255004 272484 255010 272496
rect 269298 272484 269304 272496
rect 269356 272484 269362 272536
rect 270310 272484 270316 272536
rect 270368 272524 270374 272536
rect 280522 272524 280528 272536
rect 270368 272496 280528 272524
rect 270368 272484 270374 272496
rect 280522 272484 280528 272496
rect 280580 272484 280586 272536
rect 329742 272484 329748 272536
rect 329800 272524 329806 272536
rect 338850 272524 338856 272536
rect 329800 272496 338856 272524
rect 329800 272484 329806 272496
rect 338850 272484 338856 272496
rect 338908 272484 338914 272536
rect 339218 272484 339224 272536
rect 339276 272524 339282 272536
rect 354214 272524 354220 272536
rect 339276 272496 354220 272524
rect 339276 272484 339282 272496
rect 354214 272484 354220 272496
rect 354272 272484 354278 272536
rect 354490 272484 354496 272536
rect 354548 272524 354554 272536
rect 375558 272524 375564 272536
rect 354548 272496 375564 272524
rect 354548 272484 354554 272496
rect 375558 272484 375564 272496
rect 375616 272484 375622 272536
rect 379422 272484 379428 272536
rect 379480 272524 379486 272536
rect 410978 272524 410984 272536
rect 379480 272496 410984 272524
rect 379480 272484 379486 272496
rect 410978 272484 410984 272496
rect 411036 272484 411042 272536
rect 416590 272484 416596 272536
rect 416648 272524 416654 272536
rect 460842 272524 460848 272536
rect 416648 272496 460848 272524
rect 416648 272484 416654 272496
rect 460842 272484 460848 272496
rect 460900 272484 460906 272536
rect 461394 272484 461400 272536
rect 461452 272524 461458 272536
rect 465534 272524 465540 272536
rect 461452 272496 465540 272524
rect 461452 272484 461458 272496
rect 465534 272484 465540 272496
rect 465592 272484 465598 272536
rect 465736 272524 465764 272632
rect 465902 272620 465908 272672
rect 465960 272660 465966 272672
rect 522114 272660 522120 272672
rect 465960 272632 522120 272660
rect 465960 272620 465966 272632
rect 522114 272620 522120 272632
rect 522172 272620 522178 272672
rect 526806 272620 526812 272672
rect 526864 272660 526870 272672
rect 621382 272660 621388 272672
rect 526864 272632 621388 272660
rect 526864 272620 526870 272632
rect 621382 272620 621388 272632
rect 621440 272620 621446 272672
rect 470548 272524 470554 272536
rect 465736 272496 470554 272524
rect 470548 272484 470554 272496
rect 470606 272484 470612 272536
rect 470686 272484 470692 272536
rect 470744 272524 470750 272536
rect 532694 272524 532700 272536
rect 470744 272496 532700 272524
rect 470744 272484 470750 272496
rect 532694 272484 532700 272496
rect 532752 272484 532758 272536
rect 532878 272484 532884 272536
rect 532936 272524 532942 272536
rect 538490 272524 538496 272536
rect 532936 272496 538496 272524
rect 532936 272484 532942 272496
rect 538490 272484 538496 272496
rect 538548 272484 538554 272536
rect 538674 272484 538680 272536
rect 538732 272524 538738 272536
rect 628668 272524 628696 272904
rect 632054 272892 632060 272904
rect 632112 272892 632118 272944
rect 635550 272796 635556 272808
rect 538732 272496 628696 272524
rect 629956 272768 635556 272796
rect 538732 272484 538738 272496
rect 318702 272416 318708 272468
rect 318760 272456 318766 272468
rect 324682 272456 324688 272468
rect 318760 272428 324688 272456
rect 318760 272416 318766 272428
rect 324682 272416 324688 272428
rect 324740 272416 324746 272468
rect 187694 272388 187700 272400
rect 180766 272360 187700 272388
rect 187694 272348 187700 272360
rect 187752 272348 187758 272400
rect 194962 272348 194968 272400
rect 195020 272388 195026 272400
rect 227162 272388 227168 272400
rect 195020 272360 227168 272388
rect 195020 272348 195026 272360
rect 227162 272348 227168 272360
rect 227220 272348 227226 272400
rect 395982 272348 395988 272400
rect 396040 272388 396046 272400
rect 434622 272388 434628 272400
rect 396040 272360 434628 272388
rect 396040 272348 396046 272360
rect 434622 272348 434628 272360
rect 434680 272348 434686 272400
rect 449710 272348 449716 272400
rect 449768 272388 449774 272400
rect 504174 272388 504180 272400
rect 449768 272360 504180 272388
rect 449768 272348 449774 272360
rect 504174 272348 504180 272360
rect 504232 272348 504238 272400
rect 504358 272348 504364 272400
rect 504416 272388 504422 272400
rect 513742 272388 513748 272400
rect 504416 272360 513748 272388
rect 504416 272348 504422 272360
rect 513742 272348 513748 272360
rect 513800 272348 513806 272400
rect 517422 272348 517428 272400
rect 517480 272388 517486 272400
rect 600774 272388 600780 272400
rect 517480 272360 600780 272388
rect 517480 272348 517486 272360
rect 600774 272348 600780 272360
rect 600832 272348 600838 272400
rect 600958 272348 600964 272400
rect 601016 272388 601022 272400
rect 629956 272388 629984 272768
rect 635550 272756 635556 272768
rect 635608 272756 635614 272808
rect 634078 272620 634084 272672
rect 634136 272660 634142 272672
rect 640334 272660 640340 272672
rect 634136 272632 640340 272660
rect 634136 272620 634142 272632
rect 640334 272620 640340 272632
rect 640392 272620 640398 272672
rect 601016 272360 629984 272388
rect 601016 272348 601022 272360
rect 127342 272212 127348 272264
rect 127400 272252 127406 272264
rect 179874 272252 179880 272264
rect 127400 272224 179880 272252
rect 127400 272212 127406 272224
rect 179874 272212 179880 272224
rect 179932 272212 179938 272264
rect 189074 272212 189080 272264
rect 189132 272252 189138 272264
rect 196434 272252 196440 272264
rect 189132 272224 196440 272252
rect 189132 272212 189138 272224
rect 196434 272212 196440 272224
rect 196492 272212 196498 272264
rect 391842 272212 391848 272264
rect 391900 272252 391906 272264
rect 428734 272252 428740 272264
rect 391900 272224 428740 272252
rect 391900 272212 391906 272224
rect 428734 272212 428740 272224
rect 428792 272212 428798 272264
rect 450538 272212 450544 272264
rect 450596 272252 450602 272264
rect 510246 272252 510252 272264
rect 450596 272224 510252 272252
rect 450596 272212 450602 272224
rect 510246 272212 510252 272224
rect 510304 272212 510310 272264
rect 510430 272212 510436 272264
rect 510488 272252 510494 272264
rect 518710 272252 518716 272264
rect 510488 272224 518716 272252
rect 510488 272212 510494 272224
rect 518710 272212 518716 272224
rect 518768 272212 518774 272264
rect 520090 272212 520096 272264
rect 520148 272252 520154 272264
rect 610710 272252 610716 272264
rect 520148 272224 610716 272252
rect 520148 272212 520154 272224
rect 610710 272212 610716 272224
rect 610768 272212 610774 272264
rect 145098 272076 145104 272128
rect 145156 272116 145162 272128
rect 192386 272116 192392 272128
rect 145156 272088 192392 272116
rect 145156 272076 145162 272088
rect 192386 272076 192392 272088
rect 192444 272076 192450 272128
rect 384942 272076 384948 272128
rect 385000 272116 385006 272128
rect 418062 272116 418068 272128
rect 385000 272088 418068 272116
rect 385000 272076 385006 272088
rect 418062 272076 418068 272088
rect 418120 272076 418126 272128
rect 428458 272076 428464 272128
rect 428516 272116 428522 272128
rect 470548 272116 470554 272128
rect 428516 272088 470554 272116
rect 428516 272076 428522 272088
rect 470548 272076 470554 272088
rect 470606 272076 470612 272128
rect 470778 272076 470784 272128
rect 470836 272116 470842 272128
rect 470836 272088 485268 272116
rect 470836 272076 470842 272088
rect 124950 271940 124956 271992
rect 125008 271980 125014 271992
rect 151078 271980 151084 271992
rect 125008 271952 151084 271980
rect 125008 271940 125014 271952
rect 151078 271940 151084 271952
rect 151136 271940 151142 271992
rect 431678 271940 431684 271992
rect 431736 271980 431742 271992
rect 431736 271952 480392 271980
rect 431736 271940 431742 271952
rect 105998 271804 106004 271856
rect 106056 271844 106062 271856
rect 164970 271844 164976 271856
rect 106056 271816 164976 271844
rect 106056 271804 106062 271816
rect 164970 271804 164976 271816
rect 165028 271804 165034 271856
rect 174262 271804 174268 271856
rect 174320 271844 174326 271856
rect 189166 271844 189172 271856
rect 174320 271816 189172 271844
rect 174320 271804 174326 271816
rect 189166 271804 189172 271816
rect 189224 271804 189230 271856
rect 202966 271804 202972 271856
rect 203024 271844 203030 271856
rect 233234 271844 233240 271856
rect 203024 271816 233240 271844
rect 203024 271804 203030 271816
rect 233234 271804 233240 271816
rect 233292 271804 233298 271856
rect 274634 271804 274640 271856
rect 274692 271844 274698 271856
rect 279234 271844 279240 271856
rect 274692 271816 279240 271844
rect 274692 271804 274698 271816
rect 279234 271804 279240 271816
rect 279292 271804 279298 271856
rect 355318 271804 355324 271856
rect 355376 271844 355382 271856
rect 356606 271844 356612 271856
rect 355376 271816 356612 271844
rect 355376 271804 355382 271816
rect 356606 271804 356612 271816
rect 356664 271804 356670 271856
rect 375282 271804 375288 271856
rect 375340 271844 375346 271856
rect 403894 271844 403900 271856
rect 375340 271816 403900 271844
rect 375340 271804 375346 271816
rect 403894 271804 403900 271816
rect 403952 271804 403958 271856
rect 433150 271804 433156 271856
rect 433208 271844 433214 271856
rect 480162 271844 480168 271856
rect 433208 271816 480168 271844
rect 433208 271804 433214 271816
rect 480162 271804 480168 271816
rect 480220 271804 480226 271856
rect 480364 271844 480392 271952
rect 480530 271940 480536 271992
rect 480588 271980 480594 271992
rect 485038 271980 485044 271992
rect 480588 271952 485044 271980
rect 480588 271940 480594 271952
rect 485038 271940 485044 271952
rect 485096 271940 485102 271992
rect 485240 271980 485268 272088
rect 485406 272076 485412 272128
rect 485464 272116 485470 272128
rect 547506 272116 547512 272128
rect 485464 272088 547512 272116
rect 485464 272076 485470 272088
rect 547506 272076 547512 272088
rect 547564 272076 547570 272128
rect 547690 272076 547696 272128
rect 547748 272116 547754 272128
rect 547748 272088 586514 272116
rect 547748 272076 547754 272088
rect 504358 271980 504364 271992
rect 485240 271952 504364 271980
rect 504358 271940 504364 271952
rect 504416 271940 504422 271992
rect 504542 271940 504548 271992
rect 504600 271980 504606 271992
rect 562318 271980 562324 271992
rect 504600 271952 562324 271980
rect 504600 271940 504606 271952
rect 562318 271940 562324 271952
rect 562376 271940 562382 271992
rect 586486 271980 586514 272088
rect 600774 272076 600780 272128
rect 600832 272116 600838 272128
rect 607214 272116 607220 272128
rect 600832 272088 607220 272116
rect 600832 272076 600838 272088
rect 607214 272076 607220 272088
rect 607272 272076 607278 272128
rect 600958 271980 600964 271992
rect 586486 271952 600964 271980
rect 600958 271940 600964 271952
rect 601016 271940 601022 271992
rect 484670 271844 484676 271856
rect 480364 271816 484676 271844
rect 484670 271804 484676 271816
rect 484728 271804 484734 271856
rect 494698 271804 494704 271856
rect 494756 271844 494762 271856
rect 501414 271844 501420 271856
rect 494756 271816 501420 271844
rect 494756 271804 494762 271816
rect 501414 271804 501420 271816
rect 501472 271804 501478 271856
rect 504358 271804 504364 271856
rect 504416 271844 504422 271856
rect 578510 271844 578516 271856
rect 504416 271816 578516 271844
rect 504416 271804 504422 271816
rect 578510 271804 578516 271816
rect 578568 271804 578574 271856
rect 578878 271804 578884 271856
rect 578936 271844 578942 271856
rect 604822 271844 604828 271856
rect 578936 271816 604828 271844
rect 578936 271804 578942 271816
rect 604822 271804 604828 271816
rect 604880 271804 604886 271856
rect 97810 271668 97816 271720
rect 97868 271708 97874 271720
rect 158806 271708 158812 271720
rect 97868 271680 158812 271708
rect 97868 271668 97874 271680
rect 158806 271668 158812 271680
rect 158864 271668 158870 271720
rect 169846 271668 169852 271720
rect 169904 271708 169910 271720
rect 209958 271708 209964 271720
rect 169904 271680 209964 271708
rect 169904 271668 169910 271680
rect 209958 271668 209964 271680
rect 210016 271668 210022 271720
rect 225414 271668 225420 271720
rect 225472 271708 225478 271720
rect 228358 271708 228364 271720
rect 225472 271680 228364 271708
rect 225472 271668 225478 271680
rect 228358 271668 228364 271680
rect 228416 271668 228422 271720
rect 351178 271668 351184 271720
rect 351236 271708 351242 271720
rect 366082 271708 366088 271720
rect 351236 271680 366088 271708
rect 351236 271668 351242 271680
rect 366082 271668 366088 271680
rect 366140 271668 366146 271720
rect 381998 271668 382004 271720
rect 382056 271708 382062 271720
rect 414566 271708 414572 271720
rect 382056 271680 414572 271708
rect 382056 271668 382062 271680
rect 414566 271668 414572 271680
rect 414624 271668 414630 271720
rect 421650 271708 421656 271720
rect 417160 271680 421656 271708
rect 87138 271532 87144 271584
rect 87196 271572 87202 271584
rect 151998 271572 152004 271584
rect 87196 271544 152004 271572
rect 87196 271532 87202 271544
rect 151998 271532 152004 271544
rect 152056 271532 152062 271584
rect 165154 271532 165160 271584
rect 165212 271572 165218 271584
rect 205634 271572 205640 271584
rect 165212 271544 205640 271572
rect 165212 271532 165218 271544
rect 205634 271532 205640 271544
rect 205692 271532 205698 271584
rect 215938 271532 215944 271584
rect 215996 271572 216002 271584
rect 242066 271572 242072 271584
rect 215996 271544 242072 271572
rect 215996 271532 216002 271544
rect 242066 271532 242072 271544
rect 242124 271532 242130 271584
rect 337930 271532 337936 271584
rect 337988 271572 337994 271584
rect 350718 271572 350724 271584
rect 337988 271544 350724 271572
rect 337988 271532 337994 271544
rect 350718 271532 350724 271544
rect 350776 271532 350782 271584
rect 360838 271532 360844 271584
rect 360896 271572 360902 271584
rect 377858 271572 377864 271584
rect 360896 271544 377864 271572
rect 360896 271532 360902 271544
rect 377858 271532 377864 271544
rect 377916 271532 377922 271584
rect 387702 271532 387708 271584
rect 387760 271572 387766 271584
rect 417160 271572 417188 271680
rect 421650 271668 421656 271680
rect 421708 271668 421714 271720
rect 430390 271668 430396 271720
rect 430448 271708 430454 271720
rect 483198 271708 483204 271720
rect 430448 271680 483204 271708
rect 430448 271668 430454 271680
rect 483198 271668 483204 271680
rect 483256 271668 483262 271720
rect 499298 271668 499304 271720
rect 499356 271708 499362 271720
rect 582374 271708 582380 271720
rect 499356 271680 582380 271708
rect 499356 271668 499362 271680
rect 582374 271668 582380 271680
rect 582432 271668 582438 271720
rect 583018 271668 583024 271720
rect 583076 271708 583082 271720
rect 611906 271708 611912 271720
rect 583076 271680 611912 271708
rect 583076 271668 583082 271680
rect 611906 271668 611912 271680
rect 611964 271668 611970 271720
rect 387760 271544 417188 271572
rect 387760 271532 387766 271544
rect 420178 271532 420184 271584
rect 420236 271572 420242 271584
rect 431126 271572 431132 271584
rect 420236 271544 431132 271572
rect 420236 271532 420242 271544
rect 431126 271532 431132 271544
rect 431184 271532 431190 271584
rect 437198 271532 437204 271584
rect 437256 271572 437262 271584
rect 493686 271572 493692 271584
rect 437256 271544 493692 271572
rect 437256 271532 437262 271544
rect 493686 271532 493692 271544
rect 493744 271532 493750 271584
rect 497274 271572 497280 271584
rect 493888 271544 497280 271572
rect 75362 271396 75368 271448
rect 75420 271436 75426 271448
rect 142706 271436 142712 271448
rect 75420 271408 142712 271436
rect 75420 271396 75426 271408
rect 142706 271396 142712 271408
rect 142764 271396 142770 271448
rect 162670 271396 162676 271448
rect 162728 271436 162734 271448
rect 204714 271436 204720 271448
rect 162728 271408 204720 271436
rect 162728 271396 162734 271408
rect 204714 271396 204720 271408
rect 204772 271396 204778 271448
rect 213638 271396 213644 271448
rect 213696 271436 213702 271448
rect 240410 271436 240416 271448
rect 213696 271408 240416 271436
rect 213696 271396 213702 271408
rect 240410 271396 240416 271408
rect 240468 271396 240474 271448
rect 240778 271396 240784 271448
rect 240836 271436 240842 271448
rect 259638 271436 259644 271448
rect 240836 271408 259644 271436
rect 240836 271396 240842 271408
rect 259638 271396 259644 271408
rect 259696 271396 259702 271448
rect 259822 271396 259828 271448
rect 259880 271436 259886 271448
rect 272610 271436 272616 271448
rect 259880 271408 272616 271436
rect 259880 271396 259886 271408
rect 272610 271396 272616 271408
rect 272668 271396 272674 271448
rect 325510 271396 325516 271448
rect 325568 271436 325574 271448
rect 334158 271436 334164 271448
rect 325568 271408 334164 271436
rect 325568 271396 325574 271408
rect 334158 271396 334164 271408
rect 334216 271396 334222 271448
rect 347682 271396 347688 271448
rect 347740 271436 347746 271448
rect 364886 271436 364892 271448
rect 347740 271408 364892 271436
rect 347740 271396 347746 271408
rect 364886 271396 364892 271408
rect 364944 271396 364950 271448
rect 366358 271396 366364 271448
rect 366416 271436 366422 271448
rect 383838 271436 383844 271448
rect 366416 271408 383844 271436
rect 366416 271396 366422 271408
rect 383838 271396 383844 271408
rect 383896 271396 383902 271448
rect 384758 271396 384764 271448
rect 384816 271436 384822 271448
rect 419258 271436 419264 271448
rect 384816 271408 419264 271436
rect 384816 271396 384822 271408
rect 419258 271396 419264 271408
rect 419316 271396 419322 271448
rect 426342 271436 426348 271448
rect 424336 271408 426348 271436
rect 76834 271260 76840 271312
rect 76892 271300 76898 271312
rect 143534 271300 143540 271312
rect 76892 271272 143540 271300
rect 76892 271260 76898 271272
rect 143534 271260 143540 271272
rect 143592 271260 143598 271312
rect 152182 271260 152188 271312
rect 152240 271300 152246 271312
rect 197354 271300 197360 271312
rect 152240 271272 197360 271300
rect 152240 271260 152246 271272
rect 197354 271260 197360 271272
rect 197412 271260 197418 271312
rect 198274 271260 198280 271312
rect 198332 271300 198338 271312
rect 229554 271300 229560 271312
rect 198332 271272 229560 271300
rect 198332 271260 198338 271272
rect 229554 271260 229560 271272
rect 229612 271260 229618 271312
rect 235258 271260 235264 271312
rect 235316 271300 235322 271312
rect 255314 271300 255320 271312
rect 235316 271272 255320 271300
rect 235316 271260 235322 271272
rect 255314 271260 255320 271272
rect 255372 271260 255378 271312
rect 256694 271260 256700 271312
rect 256752 271300 256758 271312
rect 261018 271300 261024 271312
rect 256752 271272 261024 271300
rect 256752 271260 256758 271272
rect 261018 271260 261024 271272
rect 261076 271260 261082 271312
rect 262030 271260 262036 271312
rect 262088 271300 262094 271312
rect 274634 271300 274640 271312
rect 262088 271272 274640 271300
rect 262088 271260 262094 271272
rect 274634 271260 274640 271272
rect 274692 271260 274698 271312
rect 329558 271260 329564 271312
rect 329616 271300 329622 271312
rect 340046 271300 340052 271312
rect 329616 271272 340052 271300
rect 329616 271260 329622 271272
rect 340046 271260 340052 271272
rect 340104 271260 340110 271312
rect 340598 271260 340604 271312
rect 340656 271300 340662 271312
rect 355134 271300 355140 271312
rect 340656 271272 355140 271300
rect 340656 271260 340662 271272
rect 355134 271260 355140 271272
rect 355192 271260 355198 271312
rect 357158 271260 357164 271312
rect 357216 271300 357222 271312
rect 379054 271300 379060 271312
rect 357216 271272 379060 271300
rect 357216 271260 357222 271272
rect 379054 271260 379060 271272
rect 379112 271260 379118 271312
rect 390278 271260 390284 271312
rect 390336 271300 390342 271312
rect 424336 271300 424364 271408
rect 426342 271396 426348 271408
rect 426400 271396 426406 271448
rect 439958 271396 439964 271448
rect 440016 271436 440022 271448
rect 493888 271436 493916 271544
rect 497274 271532 497280 271544
rect 497332 271532 497338 271584
rect 501966 271532 501972 271584
rect 502024 271572 502030 271584
rect 585962 271572 585968 271584
rect 502024 271544 585968 271572
rect 502024 271532 502030 271544
rect 585962 271532 585968 271544
rect 586020 271532 586026 271584
rect 611998 271532 612004 271584
rect 612056 271572 612062 271584
rect 618990 271572 618996 271584
rect 612056 271544 618996 271572
rect 612056 271532 612062 271544
rect 618990 271532 618996 271544
rect 619048 271532 619054 271584
rect 440016 271408 493916 271436
rect 440016 271396 440022 271408
rect 496538 271396 496544 271448
rect 496596 271436 496602 271448
rect 504358 271436 504364 271448
rect 496596 271408 504364 271436
rect 496596 271396 496602 271408
rect 504358 271396 504364 271408
rect 504416 271396 504422 271448
rect 505002 271396 505008 271448
rect 505060 271436 505066 271448
rect 589458 271436 589464 271448
rect 505060 271408 589464 271436
rect 505060 271396 505066 271408
rect 589458 271396 589464 271408
rect 589516 271396 589522 271448
rect 589918 271396 589924 271448
rect 589976 271436 589982 271448
rect 633250 271436 633256 271448
rect 589976 271408 633256 271436
rect 589976 271396 589982 271408
rect 633250 271396 633256 271408
rect 633308 271396 633314 271448
rect 432230 271300 432236 271312
rect 390336 271272 424364 271300
rect 425992 271272 432236 271300
rect 390336 271260 390342 271272
rect 68186 271124 68192 271176
rect 68244 271164 68250 271176
rect 138474 271164 138480 271176
rect 68244 271136 138480 271164
rect 68244 271124 68250 271136
rect 138474 271124 138480 271136
rect 138532 271124 138538 271176
rect 141510 271124 141516 271176
rect 141568 271164 141574 271176
rect 189810 271164 189816 271176
rect 141568 271136 189816 271164
rect 141568 271124 141574 271136
rect 189810 271124 189816 271136
rect 189868 271124 189874 271176
rect 191190 271124 191196 271176
rect 191248 271164 191254 271176
rect 225138 271164 225144 271176
rect 191248 271136 225144 271164
rect 191248 271124 191254 271136
rect 225138 271124 225144 271136
rect 225196 271124 225202 271176
rect 230198 271124 230204 271176
rect 230256 271164 230262 271176
rect 252002 271164 252008 271176
rect 230256 271136 252008 271164
rect 230256 271124 230262 271136
rect 252002 271124 252008 271136
rect 252060 271124 252066 271176
rect 268010 271124 268016 271176
rect 268068 271164 268074 271176
rect 278774 271164 278780 271176
rect 268068 271136 278780 271164
rect 268068 271124 268074 271136
rect 278774 271124 278780 271136
rect 278832 271124 278838 271176
rect 279786 271124 279792 271176
rect 279844 271164 279850 271176
rect 287054 271164 287060 271176
rect 279844 271136 287060 271164
rect 279844 271124 279850 271136
rect 287054 271124 287060 271136
rect 287112 271124 287118 271176
rect 331122 271124 331128 271176
rect 331180 271164 331186 271176
rect 342438 271164 342444 271176
rect 331180 271136 342444 271164
rect 331180 271124 331186 271136
rect 342438 271124 342444 271136
rect 342496 271124 342502 271176
rect 343542 271124 343548 271176
rect 343600 271164 343606 271176
rect 360194 271164 360200 271176
rect 343600 271136 360200 271164
rect 343600 271124 343606 271136
rect 360194 271124 360200 271136
rect 360252 271124 360258 271176
rect 364150 271124 364156 271176
rect 364208 271164 364214 271176
rect 389726 271164 389732 271176
rect 364208 271136 389732 271164
rect 364208 271124 364214 271136
rect 389726 271124 389732 271136
rect 389784 271124 389790 271176
rect 394326 271124 394332 271176
rect 394384 271164 394390 271176
rect 425992 271164 426020 271272
rect 432230 271260 432236 271272
rect 432288 271260 432294 271312
rect 442902 271260 442908 271312
rect 442960 271300 442966 271312
rect 500862 271300 500868 271312
rect 442960 271272 500868 271300
rect 442960 271260 442966 271272
rect 500862 271260 500868 271272
rect 500920 271260 500926 271312
rect 507670 271260 507676 271312
rect 507728 271300 507734 271312
rect 593046 271300 593052 271312
rect 507728 271272 593052 271300
rect 507728 271260 507734 271272
rect 593046 271260 593052 271272
rect 593104 271260 593110 271312
rect 598198 271260 598204 271312
rect 598256 271300 598262 271312
rect 645026 271300 645032 271312
rect 598256 271272 645032 271300
rect 598256 271260 598262 271272
rect 645026 271260 645032 271272
rect 645084 271260 645090 271312
rect 437934 271164 437940 271176
rect 394384 271136 426020 271164
rect 427096 271136 437940 271164
rect 394384 271124 394390 271136
rect 113450 270988 113456 271040
rect 113508 271028 113514 271040
rect 169938 271028 169944 271040
rect 113508 271000 169944 271028
rect 113508 270988 113514 271000
rect 169938 270988 169944 271000
rect 169996 270988 170002 271040
rect 187418 270988 187424 271040
rect 187476 271028 187482 271040
rect 215938 271028 215944 271040
rect 187476 271000 215944 271028
rect 187476 270988 187482 271000
rect 215938 270988 215944 271000
rect 215996 270988 216002 271040
rect 251450 270988 251456 271040
rect 251508 271028 251514 271040
rect 266906 271028 266912 271040
rect 251508 271000 266912 271028
rect 251508 270988 251514 271000
rect 266906 270988 266912 271000
rect 266964 270988 266970 271040
rect 417418 270988 417424 271040
rect 417476 271028 417482 271040
rect 427096 271028 427124 271136
rect 437934 271124 437940 271136
rect 437992 271124 437998 271176
rect 441338 271124 441344 271176
rect 441396 271164 441402 271176
rect 445018 271164 445024 271176
rect 441396 271136 445024 271164
rect 441396 271124 441402 271136
rect 445018 271124 445024 271136
rect 445076 271124 445082 271176
rect 445662 271124 445668 271176
rect 445720 271164 445726 271176
rect 503990 271164 503996 271176
rect 445720 271136 503996 271164
rect 445720 271124 445726 271136
rect 503990 271124 503996 271136
rect 504048 271124 504054 271176
rect 524046 271124 524052 271176
rect 524104 271164 524110 271176
rect 617334 271164 617340 271176
rect 524104 271136 617340 271164
rect 524104 271124 524110 271136
rect 617334 271124 617340 271136
rect 617392 271124 617398 271176
rect 617518 271124 617524 271176
rect 617576 271164 617582 271176
rect 626074 271164 626080 271176
rect 617576 271136 626080 271164
rect 617576 271124 617582 271136
rect 626074 271124 626080 271136
rect 626132 271124 626138 271176
rect 417476 271000 427124 271028
rect 417476 270988 417482 271000
rect 427446 270988 427452 271040
rect 427504 271028 427510 271040
rect 479150 271028 479156 271040
rect 427504 271000 479156 271028
rect 427504 270988 427510 271000
rect 479150 270988 479156 271000
rect 479208 270988 479214 271040
rect 485038 270988 485044 271040
rect 485096 271028 485102 271040
rect 494698 271028 494704 271040
rect 485096 271000 494704 271028
rect 485096 270988 485102 271000
rect 494698 270988 494704 271000
rect 494756 270988 494762 271040
rect 495066 270988 495072 271040
rect 495124 271028 495130 271040
rect 575290 271028 575296 271040
rect 495124 271000 575296 271028
rect 495124 270988 495130 271000
rect 575290 270988 575296 271000
rect 575348 270988 575354 271040
rect 123754 270852 123760 270904
rect 123812 270892 123818 270904
rect 177482 270892 177488 270904
rect 123812 270864 177488 270892
rect 123812 270852 123818 270864
rect 177482 270852 177488 270864
rect 177540 270852 177546 270904
rect 407758 270852 407764 270904
rect 407816 270892 407822 270904
rect 440510 270892 440516 270904
rect 407816 270864 440516 270892
rect 407816 270852 407822 270864
rect 440510 270852 440516 270864
rect 440568 270852 440574 270904
rect 449158 270852 449164 270904
rect 449216 270892 449222 270904
rect 490190 270892 490196 270904
rect 449216 270864 490196 270892
rect 449216 270852 449222 270864
rect 490190 270852 490196 270864
rect 490248 270852 490254 270904
rect 492582 270852 492588 270904
rect 492640 270892 492646 270904
rect 571702 270892 571708 270904
rect 492640 270864 571708 270892
rect 492640 270852 492646 270864
rect 571702 270852 571708 270864
rect 571760 270852 571766 270904
rect 134426 270716 134432 270768
rect 134484 270756 134490 270768
rect 185118 270756 185124 270768
rect 134484 270728 185124 270756
rect 134484 270716 134490 270728
rect 185118 270716 185124 270728
rect 185176 270716 185182 270768
rect 321370 270716 321376 270768
rect 321428 270756 321434 270768
rect 327074 270756 327080 270768
rect 321428 270728 327080 270756
rect 321428 270716 321434 270728
rect 327074 270716 327080 270728
rect 327132 270716 327138 270768
rect 414658 270716 414664 270768
rect 414716 270756 414722 270768
rect 450814 270756 450820 270768
rect 414716 270728 450820 270756
rect 414716 270716 414722 270728
rect 450814 270716 450820 270728
rect 450872 270716 450878 270768
rect 480254 270716 480260 270768
rect 480312 270756 480318 270768
rect 486602 270756 486608 270768
rect 480312 270728 486608 270756
rect 480312 270716 480318 270728
rect 486602 270716 486608 270728
rect 486660 270716 486666 270768
rect 486970 270716 486976 270768
rect 487028 270756 487034 270768
rect 564618 270756 564624 270768
rect 487028 270728 564624 270756
rect 487028 270716 487034 270728
rect 564618 270716 564624 270728
rect 564676 270716 564682 270768
rect 567838 270716 567844 270768
rect 567896 270756 567902 270768
rect 597738 270756 597744 270768
rect 567896 270728 597744 270756
rect 567896 270716 567902 270728
rect 597738 270716 597744 270728
rect 597796 270716 597802 270768
rect 121454 270580 121460 270632
rect 121512 270620 121518 270632
rect 168098 270620 168104 270632
rect 121512 270592 168104 270620
rect 121512 270580 121518 270592
rect 168098 270580 168104 270592
rect 168156 270580 168162 270632
rect 403618 270580 403624 270632
rect 403676 270620 403682 270632
rect 433426 270620 433432 270632
rect 403676 270592 433432 270620
rect 403676 270580 403682 270592
rect 433426 270580 433432 270592
rect 433484 270580 433490 270632
rect 453298 270580 453304 270632
rect 453356 270620 453362 270632
rect 487798 270620 487804 270632
rect 453356 270592 487804 270620
rect 453356 270580 453362 270592
rect 487798 270580 487804 270592
rect 487856 270580 487862 270632
rect 489638 270580 489644 270632
rect 489696 270620 489702 270632
rect 568206 270620 568212 270632
rect 489696 270592 568212 270620
rect 489696 270580 489702 270592
rect 568206 270580 568212 270592
rect 568264 270580 568270 270632
rect 84102 270444 84108 270496
rect 84160 270484 84166 270496
rect 137462 270484 137468 270496
rect 84160 270456 137468 270484
rect 84160 270444 84166 270456
rect 137462 270444 137468 270456
rect 137520 270444 137526 270496
rect 137646 270444 137652 270496
rect 137704 270484 137710 270496
rect 186130 270484 186136 270496
rect 137704 270456 186136 270484
rect 137704 270444 137710 270456
rect 186130 270444 186136 270456
rect 186188 270444 186194 270496
rect 201034 270444 201040 270496
rect 201092 270484 201098 270496
rect 201862 270484 201868 270496
rect 201092 270456 201868 270484
rect 201092 270444 201098 270456
rect 201862 270444 201868 270456
rect 201920 270444 201926 270496
rect 206830 270444 206836 270496
rect 206888 270484 206894 270496
rect 235810 270484 235816 270496
rect 206888 270456 235816 270484
rect 206888 270444 206894 270456
rect 235810 270444 235816 270456
rect 235868 270444 235874 270496
rect 278038 270444 278044 270496
rect 278096 270484 278102 270496
rect 283834 270484 283840 270496
rect 278096 270456 283840 270484
rect 278096 270444 278102 270456
rect 283834 270444 283840 270456
rect 283892 270444 283898 270496
rect 400858 270444 400864 270496
rect 400916 270484 400922 270496
rect 441614 270484 441620 270496
rect 400916 270456 441620 270484
rect 400916 270444 400922 270456
rect 441614 270444 441620 270456
rect 441672 270444 441678 270496
rect 456426 270444 456432 270496
rect 456484 270484 456490 270496
rect 520274 270484 520280 270496
rect 456484 270456 520280 270484
rect 456484 270444 456490 270456
rect 520274 270444 520280 270456
rect 520332 270444 520338 270496
rect 523126 270444 523132 270496
rect 523184 270484 523190 270496
rect 532786 270484 532792 270496
rect 523184 270456 532792 270484
rect 523184 270444 523190 270456
rect 532786 270444 532792 270456
rect 532844 270444 532850 270496
rect 619634 270484 619640 270496
rect 533356 270456 619640 270484
rect 533356 270416 533384 270456
rect 619634 270444 619640 270456
rect 619692 270444 619698 270496
rect 533172 270388 533384 270416
rect 78858 270308 78864 270360
rect 78916 270348 78922 270360
rect 132494 270348 132500 270360
rect 78916 270320 132500 270348
rect 78916 270308 78922 270320
rect 132494 270308 132500 270320
rect 132552 270308 132558 270360
rect 133782 270308 133788 270360
rect 133840 270348 133846 270360
rect 183646 270348 183652 270360
rect 133840 270320 183652 270348
rect 133840 270308 133846 270320
rect 183646 270308 183652 270320
rect 183704 270308 183710 270360
rect 185302 270308 185308 270360
rect 185360 270348 185366 270360
rect 194410 270348 194416 270360
rect 185360 270320 194416 270348
rect 185360 270308 185366 270320
rect 194410 270308 194416 270320
rect 194468 270308 194474 270360
rect 199930 270308 199936 270360
rect 199988 270348 199994 270360
rect 230842 270348 230848 270360
rect 199988 270320 230848 270348
rect 199988 270308 199994 270320
rect 230842 270308 230848 270320
rect 230900 270308 230906 270360
rect 232682 270308 232688 270360
rect 232740 270348 232746 270360
rect 248230 270348 248236 270360
rect 232740 270320 248236 270348
rect 232740 270308 232746 270320
rect 248230 270308 248236 270320
rect 248288 270308 248294 270360
rect 283098 270308 283104 270360
rect 283156 270348 283162 270360
rect 284662 270348 284668 270360
rect 283156 270320 284668 270348
rect 283156 270308 283162 270320
rect 284662 270308 284668 270320
rect 284720 270308 284726 270360
rect 355042 270308 355048 270360
rect 355100 270348 355106 270360
rect 376754 270348 376760 270360
rect 355100 270320 376760 270348
rect 355100 270308 355106 270320
rect 376754 270308 376760 270320
rect 376812 270308 376818 270360
rect 380526 270308 380532 270360
rect 380584 270348 380590 270360
rect 404354 270348 404360 270360
rect 380584 270320 404360 270348
rect 380584 270308 380590 270320
rect 404354 270308 404360 270320
rect 404412 270308 404418 270360
rect 415026 270308 415032 270360
rect 415084 270348 415090 270360
rect 461210 270348 461216 270360
rect 415084 270320 461216 270348
rect 415084 270308 415090 270320
rect 461210 270308 461216 270320
rect 461268 270308 461274 270360
rect 461394 270308 461400 270360
rect 461452 270348 461458 270360
rect 461452 270320 524644 270348
rect 461452 270308 461458 270320
rect 111978 270172 111984 270224
rect 112036 270212 112042 270224
rect 168742 270212 168748 270224
rect 112036 270184 168748 270212
rect 112036 270172 112042 270184
rect 168742 270172 168748 270184
rect 168800 270172 168806 270224
rect 184842 270172 184848 270224
rect 184900 270212 184906 270224
rect 219342 270212 219348 270224
rect 184900 270184 219348 270212
rect 184900 270172 184906 270184
rect 219342 270172 219348 270184
rect 219400 270172 219406 270224
rect 244366 270172 244372 270224
rect 244424 270212 244430 270224
rect 262306 270212 262312 270224
rect 244424 270184 262312 270212
rect 244424 270172 244430 270184
rect 262306 270172 262312 270184
rect 262364 270172 262370 270224
rect 334342 270172 334348 270224
rect 334400 270212 334406 270224
rect 346394 270212 346400 270224
rect 334400 270184 346400 270212
rect 334400 270172 334406 270184
rect 346394 270172 346400 270184
rect 346452 270172 346458 270224
rect 372246 270172 372252 270224
rect 372304 270212 372310 270224
rect 397454 270212 397460 270224
rect 372304 270184 397460 270212
rect 372304 270172 372310 270184
rect 397454 270172 397460 270184
rect 397512 270172 397518 270224
rect 409598 270172 409604 270224
rect 409656 270212 409662 270224
rect 454034 270212 454040 270224
rect 409656 270184 454040 270212
rect 409656 270172 409662 270184
rect 454034 270172 454040 270184
rect 454092 270172 454098 270224
rect 458818 270172 458824 270224
rect 458876 270212 458882 270224
rect 524414 270212 524420 270224
rect 458876 270184 524420 270212
rect 458876 270172 458882 270184
rect 524414 270172 524420 270184
rect 524472 270172 524478 270224
rect 524616 270212 524644 270320
rect 525610 270308 525616 270360
rect 525668 270348 525674 270360
rect 533172 270348 533200 270388
rect 525668 270320 533200 270348
rect 525668 270308 525674 270320
rect 533522 270308 533528 270360
rect 533580 270348 533586 270360
rect 626534 270348 626540 270360
rect 533580 270320 626540 270348
rect 533580 270308 533586 270320
rect 626534 270308 626540 270320
rect 626592 270308 626598 270360
rect 527174 270212 527180 270224
rect 524616 270184 527180 270212
rect 527174 270172 527180 270184
rect 527232 270172 527238 270224
rect 528370 270172 528376 270224
rect 528428 270212 528434 270224
rect 533246 270212 533252 270224
rect 528428 270184 533252 270212
rect 528428 270172 528434 270184
rect 533246 270172 533252 270184
rect 533304 270172 533310 270224
rect 533522 270172 533528 270224
rect 533580 270212 533586 270224
rect 623958 270212 623964 270224
rect 533580 270184 623964 270212
rect 533580 270172 533586 270184
rect 623958 270172 623964 270184
rect 624016 270172 624022 270224
rect 89622 270036 89628 270088
rect 89680 270076 89686 270088
rect 153010 270076 153016 270088
rect 89680 270048 153016 270076
rect 89680 270036 89686 270048
rect 153010 270036 153016 270048
rect 153068 270036 153074 270088
rect 176562 270036 176568 270088
rect 176620 270076 176626 270088
rect 211154 270076 211160 270088
rect 176620 270048 211160 270076
rect 176620 270036 176626 270048
rect 211154 270036 211160 270048
rect 211212 270036 211218 270088
rect 212442 270036 212448 270088
rect 212500 270076 212506 270088
rect 239950 270076 239956 270088
rect 212500 270048 239956 270076
rect 212500 270036 212506 270048
rect 239950 270036 239956 270048
rect 240008 270036 240014 270088
rect 241882 270036 241888 270088
rect 241940 270076 241946 270088
rect 260650 270076 260656 270088
rect 241940 270048 260656 270076
rect 241940 270036 241946 270048
rect 260650 270036 260656 270048
rect 260708 270036 260714 270088
rect 266170 270036 266176 270088
rect 266228 270076 266234 270088
rect 277210 270076 277216 270088
rect 266228 270048 277216 270076
rect 266228 270036 266234 270048
rect 277210 270036 277216 270048
rect 277268 270036 277274 270088
rect 345290 270036 345296 270088
rect 345348 270076 345354 270088
rect 358814 270076 358820 270088
rect 345348 270048 358820 270076
rect 345348 270036 345354 270048
rect 358814 270036 358820 270048
rect 358872 270036 358878 270088
rect 366634 270036 366640 270088
rect 366692 270076 366698 270088
rect 393314 270076 393320 270088
rect 366692 270048 393320 270076
rect 366692 270036 366698 270048
rect 393314 270036 393320 270048
rect 393372 270036 393378 270088
rect 394694 270036 394700 270088
rect 394752 270076 394758 270088
rect 408770 270076 408776 270088
rect 394752 270048 408776 270076
rect 394752 270036 394758 270048
rect 408770 270036 408776 270048
rect 408828 270036 408834 270088
rect 412450 270036 412456 270088
rect 412508 270076 412514 270088
rect 458174 270076 458180 270088
rect 412508 270048 458180 270076
rect 412508 270036 412514 270048
rect 458174 270036 458180 270048
rect 458232 270036 458238 270088
rect 463510 270036 463516 270088
rect 463568 270076 463574 270088
rect 530762 270076 530768 270088
rect 463568 270048 530768 270076
rect 463568 270036 463574 270048
rect 530762 270036 530768 270048
rect 530820 270036 530826 270088
rect 530946 270036 530952 270088
rect 531004 270076 531010 270088
rect 532970 270076 532976 270088
rect 531004 270048 532976 270076
rect 531004 270036 531010 270048
rect 532970 270036 532976 270048
rect 533028 270036 533034 270088
rect 538306 270076 538312 270088
rect 533356 270048 538312 270076
rect 85482 269900 85488 269952
rect 85540 269940 85546 269952
rect 149422 269940 149428 269952
rect 85540 269912 149428 269940
rect 85540 269900 85546 269912
rect 149422 269900 149428 269912
rect 149480 269900 149486 269952
rect 152826 269900 152832 269952
rect 152884 269940 152890 269952
rect 157150 269940 157156 269952
rect 152884 269912 157156 269940
rect 152884 269900 152890 269912
rect 157150 269900 157156 269912
rect 157208 269900 157214 269952
rect 173802 269900 173808 269952
rect 173860 269940 173866 269952
rect 212626 269940 212632 269952
rect 173860 269912 212632 269940
rect 173860 269900 173866 269912
rect 212626 269900 212632 269912
rect 212684 269900 212690 269952
rect 226610 269900 226616 269952
rect 226668 269940 226674 269952
rect 249886 269940 249892 269952
rect 226668 269912 249892 269940
rect 226668 269900 226674 269912
rect 249886 269900 249892 269912
rect 249944 269900 249950 269952
rect 256878 269900 256884 269952
rect 256936 269940 256942 269952
rect 268930 269940 268936 269952
rect 256936 269912 268936 269940
rect 256936 269900 256942 269912
rect 268930 269900 268936 269912
rect 268988 269900 268994 269952
rect 330202 269900 330208 269952
rect 330260 269940 330266 269952
rect 340874 269940 340880 269952
rect 330260 269912 340880 269940
rect 330260 269900 330266 269912
rect 340874 269900 340880 269912
rect 340932 269900 340938 269952
rect 341794 269900 341800 269952
rect 341852 269940 341858 269952
rect 357434 269940 357440 269952
rect 341852 269912 357440 269940
rect 341852 269900 341858 269912
rect 357434 269900 357440 269912
rect 357492 269900 357498 269952
rect 359182 269900 359188 269952
rect 359240 269940 359246 269952
rect 382274 269940 382280 269952
rect 359240 269912 382280 269940
rect 359240 269900 359246 269912
rect 382274 269900 382280 269912
rect 382332 269900 382338 269952
rect 383010 269900 383016 269952
rect 383068 269940 383074 269952
rect 411254 269940 411260 269952
rect 383068 269912 411260 269940
rect 383068 269900 383074 269912
rect 411254 269900 411260 269912
rect 411312 269900 411318 269952
rect 419626 269900 419632 269952
rect 419684 269940 419690 269952
rect 468018 269940 468024 269952
rect 419684 269912 468024 269940
rect 419684 269900 419690 269912
rect 468018 269900 468024 269912
rect 468076 269900 468082 269952
rect 468478 269900 468484 269952
rect 468536 269940 468542 269952
rect 533356 269940 533384 270048
rect 538306 270036 538312 270048
rect 538364 270036 538370 270088
rect 630674 270076 630680 270088
rect 538876 270048 630680 270076
rect 468536 269912 533384 269940
rect 468536 269900 468542 269912
rect 533982 269900 533988 269952
rect 534040 269940 534046 269952
rect 538876 269940 538904 270048
rect 630674 270036 630680 270048
rect 630732 270036 630738 270088
rect 534040 269912 538904 269940
rect 534040 269900 534046 269912
rect 539042 269900 539048 269952
rect 539100 269940 539106 269952
rect 541526 269940 541532 269952
rect 539100 269912 541532 269940
rect 539100 269900 539106 269912
rect 541526 269900 541532 269912
rect 541584 269900 541590 269952
rect 640518 269940 640524 269952
rect 542188 269912 640524 269940
rect 70578 269764 70584 269816
rect 70636 269804 70642 269816
rect 79318 269804 79324 269816
rect 70636 269776 79324 269804
rect 70636 269764 70642 269776
rect 79318 269764 79324 269776
rect 79376 269764 79382 269816
rect 80054 269764 80060 269816
rect 80112 269804 80118 269816
rect 146386 269804 146392 269816
rect 80112 269776 146392 269804
rect 80112 269764 80118 269776
rect 146386 269764 146392 269776
rect 146444 269764 146450 269816
rect 158622 269764 158628 269816
rect 158680 269804 158686 269816
rect 201034 269804 201040 269816
rect 158680 269776 201040 269804
rect 158680 269764 158686 269776
rect 201034 269764 201040 269776
rect 201092 269764 201098 269816
rect 201678 269764 201684 269816
rect 201736 269804 201742 269816
rect 232498 269804 232504 269816
rect 201736 269776 232504 269804
rect 201736 269764 201742 269776
rect 232498 269764 232504 269776
rect 232556 269764 232562 269816
rect 237282 269764 237288 269816
rect 237340 269804 237346 269816
rect 257338 269804 257344 269816
rect 237340 269776 257344 269804
rect 237340 269764 237346 269776
rect 257338 269764 257344 269776
rect 257396 269764 257402 269816
rect 258534 269764 258540 269816
rect 258592 269804 258598 269816
rect 272242 269804 272248 269816
rect 258592 269776 272248 269804
rect 258592 269764 258598 269776
rect 272242 269764 272248 269776
rect 272300 269764 272306 269816
rect 273070 269764 273076 269816
rect 273128 269804 273134 269816
rect 282178 269804 282184 269816
rect 273128 269776 282184 269804
rect 273128 269764 273134 269776
rect 282178 269764 282184 269776
rect 282236 269764 282242 269816
rect 326890 269764 326896 269816
rect 326948 269804 326954 269816
rect 335538 269804 335544 269816
rect 326948 269776 335544 269804
rect 326948 269764 326954 269776
rect 335538 269764 335544 269776
rect 335596 269764 335602 269816
rect 335998 269764 336004 269816
rect 336056 269804 336062 269816
rect 349154 269804 349160 269816
rect 336056 269776 349160 269804
rect 336056 269764 336062 269776
rect 349154 269764 349160 269776
rect 349212 269764 349218 269816
rect 351730 269764 351736 269816
rect 351788 269804 351794 269816
rect 371234 269804 371240 269816
rect 351788 269776 371240 269804
rect 351788 269764 351794 269776
rect 371234 269764 371240 269776
rect 371292 269764 371298 269816
rect 376570 269764 376576 269816
rect 376628 269804 376634 269816
rect 407114 269804 407120 269816
rect 376628 269776 407120 269804
rect 376628 269764 376634 269776
rect 407114 269764 407120 269776
rect 407172 269764 407178 269816
rect 417142 269764 417148 269816
rect 417200 269804 417206 269816
rect 465074 269804 465080 269816
rect 417200 269776 465080 269804
rect 417200 269764 417206 269776
rect 465074 269764 465080 269776
rect 465132 269764 465138 269816
rect 465994 269764 466000 269816
rect 466052 269804 466058 269816
rect 532234 269804 532240 269816
rect 466052 269776 532240 269804
rect 466052 269764 466058 269776
rect 532234 269764 532240 269776
rect 532292 269764 532298 269816
rect 538858 269804 538864 269816
rect 532436 269776 538864 269804
rect 122742 269628 122748 269680
rect 122800 269668 122806 269680
rect 176194 269668 176200 269680
rect 122800 269640 176200 269668
rect 122800 269628 122806 269640
rect 176194 269628 176200 269640
rect 176252 269628 176258 269680
rect 183462 269628 183468 269680
rect 183520 269668 183526 269680
rect 205450 269668 205456 269680
rect 183520 269640 205456 269668
rect 183520 269628 183526 269640
rect 205450 269628 205456 269640
rect 205508 269628 205514 269680
rect 392026 269628 392032 269680
rect 392084 269668 392090 269680
rect 401686 269668 401692 269680
rect 392084 269640 401692 269668
rect 392084 269628 392090 269640
rect 401686 269628 401692 269640
rect 401744 269628 401750 269680
rect 404354 269628 404360 269680
rect 404412 269668 404418 269680
rect 423674 269668 423680 269680
rect 404412 269640 423680 269668
rect 404412 269628 404418 269640
rect 423674 269628 423680 269640
rect 423732 269628 423738 269680
rect 423950 269628 423956 269680
rect 424008 269668 424014 269680
rect 451366 269668 451372 269680
rect 424008 269640 451372 269668
rect 424008 269628 424014 269640
rect 451366 269628 451372 269640
rect 451424 269628 451430 269680
rect 453574 269628 453580 269680
rect 453632 269668 453638 269680
rect 509234 269668 509240 269680
rect 453632 269640 509240 269668
rect 453632 269628 453638 269640
rect 509234 269628 509240 269640
rect 509292 269628 509298 269680
rect 532436 269668 532464 269776
rect 538858 269764 538864 269776
rect 538916 269764 538922 269816
rect 540514 269764 540520 269816
rect 540572 269804 540578 269816
rect 542188 269804 542216 269912
rect 640518 269900 640524 269912
rect 640576 269900 640582 269952
rect 540572 269776 542216 269804
rect 540572 269764 540578 269776
rect 542446 269764 542452 269816
rect 542504 269804 542510 269816
rect 637666 269804 637672 269816
rect 542504 269776 637672 269804
rect 542504 269764 542510 269776
rect 637666 269764 637672 269776
rect 637724 269764 637730 269816
rect 509712 269640 532464 269668
rect 129642 269492 129648 269544
rect 129700 269532 129706 269544
rect 181162 269532 181168 269544
rect 129700 269504 181168 269532
rect 129700 269492 129706 269504
rect 181162 269492 181168 269504
rect 181220 269492 181226 269544
rect 204162 269492 204168 269544
rect 204220 269532 204226 269544
rect 223482 269532 223488 269544
rect 204220 269504 223488 269532
rect 204220 269492 204226 269504
rect 223482 269492 223488 269504
rect 223540 269492 223546 269544
rect 398742 269492 398748 269544
rect 398800 269532 398806 269544
rect 412634 269532 412640 269544
rect 398800 269504 412640 269532
rect 398800 269492 398806 269504
rect 412634 269492 412640 269504
rect 412692 269492 412698 269544
rect 424594 269492 424600 269544
rect 424652 269532 424658 269544
rect 475010 269532 475016 269544
rect 424652 269504 475016 269532
rect 424652 269492 424658 269504
rect 475010 269492 475016 269504
rect 475068 269492 475074 269544
rect 495250 269492 495256 269544
rect 495308 269532 495314 269544
rect 509712 269532 509740 269640
rect 532786 269628 532792 269680
rect 532844 269668 532850 269680
rect 616414 269668 616420 269680
rect 532844 269640 616420 269668
rect 532844 269628 532850 269640
rect 616414 269628 616420 269640
rect 616472 269628 616478 269680
rect 495308 269504 509740 269532
rect 495308 269492 495314 269504
rect 509878 269492 509884 269544
rect 509936 269532 509942 269544
rect 596174 269532 596180 269544
rect 509936 269504 596180 269532
rect 509936 269492 509942 269504
rect 596174 269492 596180 269504
rect 596232 269492 596238 269544
rect 126882 269356 126888 269408
rect 126940 269396 126946 269408
rect 178310 269396 178316 269408
rect 126940 269368 178316 269396
rect 126940 269356 126946 269368
rect 178310 269356 178316 269368
rect 178368 269356 178374 269408
rect 408310 269356 408316 269408
rect 408368 269396 408374 269408
rect 426526 269396 426532 269408
rect 408368 269368 426532 269396
rect 408368 269356 408374 269368
rect 426526 269356 426532 269368
rect 426584 269356 426590 269408
rect 441614 269356 441620 269408
rect 441672 269396 441678 269408
rect 458450 269396 458456 269408
rect 441672 269368 458456 269396
rect 441672 269356 441678 269368
rect 458450 269356 458456 269368
rect 458508 269356 458514 269408
rect 470962 269356 470968 269408
rect 471020 269396 471026 269408
rect 538674 269396 538680 269408
rect 471020 269368 538680 269396
rect 471020 269356 471026 269368
rect 538674 269356 538680 269368
rect 538732 269356 538738 269408
rect 538858 269356 538864 269408
rect 538916 269396 538922 269408
rect 575474 269396 575480 269408
rect 538916 269368 575480 269396
rect 538916 269356 538922 269368
rect 575474 269356 575480 269368
rect 575532 269356 575538 269408
rect 143902 269220 143908 269272
rect 143960 269260 143966 269272
rect 191098 269260 191104 269272
rect 143960 269232 191104 269260
rect 143960 269220 143966 269232
rect 191098 269220 191104 269232
rect 191156 269220 191162 269272
rect 282730 269220 282736 269272
rect 282788 269260 282794 269272
rect 288802 269260 288808 269272
rect 282788 269232 288808 269260
rect 282788 269220 282794 269232
rect 288802 269220 288808 269232
rect 288860 269220 288866 269272
rect 401686 269220 401692 269272
rect 401744 269260 401750 269272
rect 416774 269260 416780 269272
rect 401744 269232 416780 269260
rect 401744 269220 401750 269232
rect 416774 269220 416780 269232
rect 416832 269220 416838 269272
rect 474274 269220 474280 269272
rect 474332 269260 474338 269272
rect 546494 269260 546500 269272
rect 474332 269232 546500 269260
rect 474332 269220 474338 269232
rect 546494 269220 546500 269232
rect 546552 269220 546558 269272
rect 319438 269084 319444 269136
rect 319496 269124 319502 269136
rect 325694 269124 325700 269136
rect 319496 269096 325700 269124
rect 319496 269084 319502 269096
rect 325694 269084 325700 269096
rect 325752 269084 325758 269136
rect 118602 269016 118608 269068
rect 118660 269056 118666 269068
rect 174538 269056 174544 269068
rect 118660 269028 174544 269056
rect 118660 269016 118666 269028
rect 174538 269016 174544 269028
rect 174596 269016 174602 269068
rect 175090 269016 175096 269068
rect 175148 269056 175154 269068
rect 177666 269056 177672 269068
rect 175148 269028 177672 269056
rect 175148 269016 175154 269028
rect 177666 269016 177672 269028
rect 177724 269016 177730 269068
rect 273254 269016 273260 269068
rect 273312 269056 273318 269068
rect 275554 269056 275560 269068
rect 273312 269028 275560 269056
rect 273312 269016 273318 269028
rect 275554 269016 275560 269028
rect 275612 269016 275618 269068
rect 436554 269016 436560 269068
rect 436612 269056 436618 269068
rect 491662 269056 491668 269068
rect 436612 269028 491668 269056
rect 436612 269016 436618 269028
rect 491662 269016 491668 269028
rect 491720 269016 491726 269068
rect 495802 269016 495808 269068
rect 495860 269056 495866 269068
rect 576854 269056 576860 269068
rect 495860 269028 576860 269056
rect 495860 269016 495866 269028
rect 576854 269016 576860 269028
rect 576912 269016 576918 269068
rect 115842 268880 115848 268932
rect 115900 268920 115906 268932
rect 171226 268920 171232 268932
rect 115900 268892 171232 268920
rect 115900 268880 115906 268892
rect 171226 268880 171232 268892
rect 171284 268880 171290 268932
rect 382366 268880 382372 268932
rect 382424 268920 382430 268932
rect 415394 268920 415400 268932
rect 382424 268892 415400 268920
rect 382424 268880 382430 268892
rect 415394 268880 415400 268892
rect 415452 268880 415458 268932
rect 433702 268880 433708 268932
rect 433760 268920 433766 268932
rect 488534 268920 488540 268932
rect 433760 268892 488540 268920
rect 433760 268880 433766 268892
rect 488534 268880 488540 268892
rect 488592 268880 488598 268932
rect 498286 268880 498292 268932
rect 498344 268920 498350 268932
rect 580994 268920 581000 268932
rect 498344 268892 581000 268920
rect 498344 268880 498350 268892
rect 580994 268880 581000 268892
rect 581052 268880 581058 268932
rect 110322 268744 110328 268796
rect 110380 268784 110386 268796
rect 167914 268784 167920 268796
rect 110380 268756 167920 268784
rect 110380 268744 110386 268756
rect 167914 268744 167920 268756
rect 167972 268744 167978 268796
rect 168282 268744 168288 268796
rect 168340 268784 168346 268796
rect 181990 268784 181996 268796
rect 168340 268756 181996 268784
rect 168340 268744 168346 268756
rect 181990 268744 181996 268756
rect 182048 268744 182054 268796
rect 188890 268744 188896 268796
rect 188948 268784 188954 268796
rect 190454 268784 190460 268796
rect 188948 268756 190460 268784
rect 188948 268744 188954 268756
rect 190454 268744 190460 268756
rect 190512 268744 190518 268796
rect 200574 268744 200580 268796
rect 200632 268784 200638 268796
rect 231302 268784 231308 268796
rect 200632 268756 231308 268784
rect 200632 268744 200638 268756
rect 231302 268744 231308 268756
rect 231360 268744 231366 268796
rect 387334 268744 387340 268796
rect 387392 268784 387398 268796
rect 422294 268784 422300 268796
rect 387392 268756 422300 268784
rect 387392 268744 387398 268756
rect 422294 268744 422300 268756
rect 422352 268744 422358 268796
rect 438670 268744 438676 268796
rect 438728 268784 438734 268796
rect 495434 268784 495440 268796
rect 438728 268756 495440 268784
rect 438728 268744 438734 268756
rect 495434 268744 495440 268756
rect 495492 268744 495498 268796
rect 500770 268744 500776 268796
rect 500828 268784 500834 268796
rect 583754 268784 583760 268796
rect 500828 268756 583760 268784
rect 500828 268744 500834 268756
rect 583754 268744 583760 268756
rect 583812 268744 583818 268796
rect 104986 268608 104992 268660
rect 105044 268648 105050 268660
rect 163774 268648 163780 268660
rect 105044 268620 163780 268648
rect 105044 268608 105050 268620
rect 163774 268608 163780 268620
rect 163832 268608 163838 268660
rect 176930 268608 176936 268660
rect 176988 268648 176994 268660
rect 215110 268648 215116 268660
rect 176988 268620 215116 268648
rect 176988 268608 176994 268620
rect 215110 268608 215116 268620
rect 215168 268608 215174 268660
rect 224218 268608 224224 268660
rect 224276 268648 224282 268660
rect 243262 268648 243268 268660
rect 224276 268620 243268 268648
rect 224276 268608 224282 268620
rect 243262 268608 243268 268620
rect 243320 268608 243326 268660
rect 352558 268608 352564 268660
rect 352616 268648 352622 268660
rect 372614 268648 372620 268660
rect 352616 268620 372620 268648
rect 352616 268608 352622 268620
rect 372614 268608 372620 268620
rect 372672 268608 372678 268660
rect 393682 268608 393688 268660
rect 393740 268648 393746 268660
rect 429194 268648 429200 268660
rect 393740 268620 429200 268648
rect 393740 268608 393746 268620
rect 429194 268608 429200 268620
rect 429252 268608 429258 268660
rect 441154 268608 441160 268660
rect 441212 268648 441218 268660
rect 499574 268648 499580 268660
rect 441212 268620 499580 268648
rect 441212 268608 441218 268620
rect 499574 268608 499580 268620
rect 499632 268608 499638 268660
rect 503254 268608 503260 268660
rect 503312 268648 503318 268660
rect 587894 268648 587900 268660
rect 503312 268620 587900 268648
rect 503312 268608 503318 268620
rect 587894 268608 587900 268620
rect 587952 268608 587958 268660
rect 99282 268472 99288 268524
rect 99340 268512 99346 268524
rect 160462 268512 160468 268524
rect 99340 268484 160468 268512
rect 99340 268472 99346 268484
rect 160462 268472 160468 268484
rect 160520 268472 160526 268524
rect 180702 268472 180708 268524
rect 180760 268512 180766 268524
rect 217594 268512 217600 268524
rect 180760 268484 217600 268512
rect 180760 268472 180766 268484
rect 217594 268472 217600 268484
rect 217652 268472 217658 268524
rect 231670 268472 231676 268524
rect 231728 268512 231734 268524
rect 253198 268512 253204 268524
rect 231728 268484 253204 268512
rect 231728 268472 231734 268484
rect 253198 268472 253204 268484
rect 253256 268472 253262 268524
rect 338482 268472 338488 268524
rect 338540 268512 338546 268524
rect 352098 268512 352104 268524
rect 338540 268484 352104 268512
rect 338540 268472 338546 268484
rect 352098 268472 352104 268484
rect 352156 268472 352162 268524
rect 367462 268472 367468 268524
rect 367520 268512 367526 268524
rect 393498 268512 393504 268524
rect 367520 268484 393504 268512
rect 367520 268472 367526 268484
rect 393498 268472 393504 268484
rect 393556 268472 393562 268524
rect 397270 268472 397276 268524
rect 397328 268512 397334 268524
rect 436094 268512 436100 268524
rect 397328 268484 436100 268512
rect 397328 268472 397334 268484
rect 436094 268472 436100 268484
rect 436152 268472 436158 268524
rect 446122 268472 446128 268524
rect 446180 268512 446186 268524
rect 506474 268512 506480 268524
rect 446180 268484 506480 268512
rect 446180 268472 446186 268484
rect 506474 268472 506480 268484
rect 506532 268472 506538 268524
rect 508222 268472 508228 268524
rect 508280 268512 508286 268524
rect 594794 268512 594800 268524
rect 508280 268484 594800 268512
rect 508280 268472 508286 268484
rect 594794 268472 594800 268484
rect 594852 268472 594858 268524
rect 92382 268336 92388 268388
rect 92440 268376 92446 268388
rect 155494 268376 155500 268388
rect 92440 268348 155500 268376
rect 92440 268336 92446 268348
rect 155494 268336 155500 268348
rect 155552 268336 155558 268388
rect 161566 268336 161572 268388
rect 161624 268376 161630 268388
rect 203518 268376 203524 268388
rect 161624 268348 203524 268376
rect 161624 268336 161630 268348
rect 203518 268336 203524 268348
rect 203576 268336 203582 268388
rect 210694 268336 210700 268388
rect 210752 268376 210758 268388
rect 236638 268376 236644 268388
rect 210752 268348 236644 268376
rect 210752 268336 210758 268348
rect 236638 268336 236644 268348
rect 236696 268336 236702 268388
rect 252646 268336 252652 268388
rect 252704 268376 252710 268388
rect 268102 268376 268108 268388
rect 252704 268348 268108 268376
rect 252704 268336 252710 268348
rect 268102 268336 268108 268348
rect 268160 268336 268166 268388
rect 348786 268336 348792 268388
rect 348844 268376 348850 268388
rect 367094 268376 367100 268388
rect 348844 268348 367100 268376
rect 348844 268336 348850 268348
rect 367094 268336 367100 268348
rect 367152 268336 367158 268388
rect 372430 268336 372436 268388
rect 372488 268376 372494 268388
rect 400490 268376 400496 268388
rect 372488 268348 400496 268376
rect 372488 268336 372494 268348
rect 400490 268336 400496 268348
rect 400548 268336 400554 268388
rect 402238 268336 402244 268388
rect 402296 268376 402302 268388
rect 443086 268376 443092 268388
rect 402296 268348 443092 268376
rect 402296 268336 402302 268348
rect 443086 268336 443092 268348
rect 443144 268336 443150 268388
rect 461854 268336 461860 268388
rect 461912 268376 461918 268388
rect 528554 268376 528560 268388
rect 461912 268348 528560 268376
rect 461912 268336 461918 268348
rect 528554 268336 528560 268348
rect 528612 268336 528618 268388
rect 541342 268336 541348 268388
rect 541400 268376 541406 268388
rect 641714 268376 641720 268388
rect 541400 268348 641720 268376
rect 541400 268336 541406 268348
rect 641714 268336 641720 268348
rect 641772 268336 641778 268388
rect 135622 268200 135628 268252
rect 135680 268240 135686 268252
rect 140682 268240 140688 268252
rect 135680 268212 140688 268240
rect 135680 268200 135686 268212
rect 140682 268200 140688 268212
rect 140740 268200 140746 268252
rect 140866 268200 140872 268252
rect 140924 268240 140930 268252
rect 188614 268240 188620 268252
rect 140924 268212 188620 268240
rect 140924 268200 140930 268212
rect 188614 268200 188620 268212
rect 188672 268200 188678 268252
rect 416222 268200 416228 268252
rect 416280 268240 416286 268252
rect 447134 268240 447140 268252
rect 416280 268212 447140 268240
rect 416280 268200 416286 268212
rect 447134 268200 447140 268212
rect 447192 268200 447198 268252
rect 493318 268200 493324 268252
rect 493376 268240 493382 268252
rect 574094 268240 574100 268252
rect 493376 268212 574100 268240
rect 493376 268200 493382 268212
rect 574094 268200 574100 268212
rect 574152 268200 574158 268252
rect 151722 268064 151728 268116
rect 151780 268104 151786 268116
rect 196066 268104 196072 268116
rect 151780 268076 196072 268104
rect 151780 268064 151786 268076
rect 196066 268064 196072 268076
rect 196124 268064 196130 268116
rect 422294 268064 422300 268116
rect 422352 268104 422358 268116
rect 444374 268104 444380 268116
rect 422352 268076 444380 268104
rect 422352 268064 422358 268076
rect 444374 268064 444380 268076
rect 444432 268064 444438 268116
rect 448422 268064 448428 268116
rect 448480 268104 448486 268116
rect 494054 268104 494060 268116
rect 448480 268076 494060 268104
rect 448480 268064 448486 268076
rect 494054 268064 494060 268076
rect 494112 268064 494118 268116
rect 527174 268064 527180 268116
rect 527232 268104 527238 268116
rect 607398 268104 607404 268116
rect 527232 268076 607404 268104
rect 527232 268064 527238 268076
rect 607398 268064 607404 268076
rect 607456 268064 607462 268116
rect 490834 267928 490840 267980
rect 490892 267968 490898 267980
rect 569954 267968 569960 267980
rect 490892 267940 569960 267968
rect 490892 267928 490898 267940
rect 569954 267928 569960 267940
rect 570012 267928 570018 267980
rect 276474 267724 276480 267776
rect 276532 267764 276538 267776
rect 278038 267764 278044 267776
rect 276532 267736 278044 267764
rect 276532 267724 276538 267736
rect 278038 267724 278044 267736
rect 278096 267724 278102 267776
rect 119338 267656 119344 267708
rect 119396 267696 119402 267708
rect 153470 267696 153476 267708
rect 119396 267668 153476 267696
rect 119396 267656 119402 267668
rect 153470 267656 153476 267668
rect 153528 267656 153534 267708
rect 169570 267696 169576 267708
rect 161446 267668 169576 267696
rect 111702 267520 111708 267572
rect 111760 267560 111766 267572
rect 161446 267560 161474 267668
rect 169570 267656 169576 267668
rect 169628 267656 169634 267708
rect 178678 267656 178684 267708
rect 178736 267696 178742 267708
rect 209314 267696 209320 267708
rect 178736 267668 209320 267696
rect 178736 267656 178742 267668
rect 209314 267656 209320 267668
rect 209372 267656 209378 267708
rect 390646 267656 390652 267708
rect 390704 267696 390710 267708
rect 408310 267696 408316 267708
rect 390704 267668 408316 267696
rect 390704 267656 390710 267668
rect 408310 267656 408316 267668
rect 408368 267656 408374 267708
rect 422938 267656 422944 267708
rect 422996 267696 423002 267708
rect 438118 267696 438124 267708
rect 422996 267668 438124 267696
rect 422996 267656 423002 267668
rect 438118 267656 438124 267668
rect 438176 267656 438182 267708
rect 445294 267656 445300 267708
rect 445352 267696 445358 267708
rect 490558 267696 490564 267708
rect 445352 267668 490564 267696
rect 445352 267656 445358 267668
rect 490558 267656 490564 267668
rect 490616 267656 490622 267708
rect 509878 267656 509884 267708
rect 509936 267696 509942 267708
rect 567838 267696 567844 267708
rect 509936 267668 567844 267696
rect 509936 267656 509942 267668
rect 567838 267656 567844 267668
rect 567896 267656 567902 267708
rect 111760 267532 161474 267560
rect 111760 267520 111766 267532
rect 169018 267520 169024 267572
rect 169076 267560 169082 267572
rect 199378 267560 199384 267572
rect 169076 267532 199384 267560
rect 169076 267520 169082 267532
rect 199378 267520 199384 267532
rect 199436 267520 199442 267572
rect 215938 267520 215944 267572
rect 215996 267560 216002 267572
rect 222562 267560 222568 267572
rect 215996 267532 222568 267560
rect 215996 267520 216002 267532
rect 222562 267520 222568 267532
rect 222620 267520 222626 267572
rect 362494 267520 362500 267572
rect 362552 267560 362558 267572
rect 369118 267560 369124 267572
rect 362552 267532 369124 267560
rect 362552 267520 362558 267532
rect 369118 267520 369124 267532
rect 369176 267520 369182 267572
rect 380710 267520 380716 267572
rect 380768 267560 380774 267572
rect 398742 267560 398748 267572
rect 380768 267532 398748 267560
rect 380768 267520 380774 267532
rect 398742 267520 398748 267532
rect 398800 267520 398806 267572
rect 404722 267520 404728 267572
rect 404780 267560 404786 267572
rect 416222 267560 416228 267572
rect 404780 267532 416228 267560
rect 404780 267520 404786 267532
rect 416222 267520 416228 267532
rect 416280 267520 416286 267572
rect 421282 267520 421288 267572
rect 421340 267560 421346 267572
rect 440878 267560 440884 267572
rect 421340 267532 440884 267560
rect 421340 267520 421346 267532
rect 440878 267520 440884 267532
rect 440936 267520 440942 267572
rect 450262 267520 450268 267572
rect 450320 267560 450326 267572
rect 498838 267560 498844 267572
rect 450320 267532 498844 267560
rect 450320 267520 450326 267532
rect 498838 267520 498844 267532
rect 498896 267520 498902 267572
rect 514846 267520 514852 267572
rect 514904 267560 514910 267572
rect 578878 267560 578884 267572
rect 514904 267532 578884 267560
rect 514904 267520 514910 267532
rect 578878 267520 578884 267532
rect 578936 267520 578942 267572
rect 86218 267384 86224 267436
rect 86276 267424 86282 267436
rect 144730 267424 144736 267436
rect 86276 267396 144736 267424
rect 86276 267384 86282 267396
rect 144730 267384 144736 267396
rect 144788 267384 144794 267436
rect 145558 267384 145564 267436
rect 145616 267424 145622 267436
rect 191926 267424 191932 267436
rect 145616 267396 191932 267424
rect 145616 267384 145622 267396
rect 191926 267384 191932 267396
rect 191984 267384 191990 267436
rect 199562 267384 199568 267436
rect 199620 267424 199626 267436
rect 204346 267424 204352 267436
rect 199620 267396 204352 267424
rect 199620 267384 199626 267396
rect 204346 267384 204352 267396
rect 204404 267384 204410 267436
rect 205450 267384 205456 267436
rect 205508 267424 205514 267436
rect 218422 267424 218428 267436
rect 205508 267396 218428 267424
rect 205508 267384 205514 267396
rect 218422 267384 218428 267396
rect 218480 267384 218486 267436
rect 233878 267384 233884 267436
rect 233936 267424 233942 267436
rect 233936 267396 238754 267424
rect 233936 267384 233942 267396
rect 104802 267248 104808 267300
rect 104860 267288 104866 267300
rect 164602 267288 164608 267300
rect 104860 267260 164608 267288
rect 104860 267248 104866 267260
rect 164602 267248 164608 267260
rect 164660 267248 164666 267300
rect 186958 267248 186964 267300
rect 187016 267288 187022 267300
rect 219250 267288 219256 267300
rect 187016 267260 219256 267288
rect 187016 267248 187022 267260
rect 219250 267248 219256 267260
rect 219308 267248 219314 267300
rect 223482 267248 223488 267300
rect 223540 267288 223546 267300
rect 234154 267288 234160 267300
rect 223540 267260 234160 267288
rect 223540 267248 223546 267260
rect 234154 267248 234160 267260
rect 234212 267248 234218 267300
rect 238726 267288 238754 267396
rect 243722 267384 243728 267436
rect 243780 267424 243786 267436
rect 251542 267424 251548 267436
rect 243780 267396 251548 267424
rect 243780 267384 243786 267396
rect 251542 267384 251548 267396
rect 251600 267384 251606 267436
rect 315298 267384 315304 267436
rect 315356 267424 315362 267436
rect 319070 267424 319076 267436
rect 315356 267396 319076 267424
rect 315356 267384 315362 267396
rect 319070 267384 319076 267396
rect 319128 267384 319134 267436
rect 340966 267384 340972 267436
rect 341024 267424 341030 267436
rect 355318 267424 355324 267436
rect 341024 267396 355324 267424
rect 341024 267384 341030 267396
rect 355318 267384 355324 267396
rect 355376 267384 355382 267436
rect 365806 267384 365812 267436
rect 365864 267424 365870 267436
rect 381538 267424 381544 267436
rect 365864 267396 381544 267424
rect 365864 267384 365870 267396
rect 381538 267384 381544 267396
rect 381596 267384 381602 267436
rect 383194 267384 383200 267436
rect 383252 267424 383258 267436
rect 401686 267424 401692 267436
rect 383252 267396 401692 267424
rect 383252 267384 383258 267396
rect 401686 267384 401692 267396
rect 401744 267384 401750 267436
rect 403066 267384 403072 267436
rect 403124 267424 403130 267436
rect 422294 267424 422300 267436
rect 403124 267396 422300 267424
rect 403124 267384 403130 267396
rect 422294 267384 422300 267396
rect 422352 267384 422358 267436
rect 428734 267384 428740 267436
rect 428792 267424 428798 267436
rect 447778 267424 447784 267436
rect 428792 267396 447784 267424
rect 428792 267384 428798 267396
rect 447778 267384 447784 267396
rect 447836 267384 447842 267436
rect 460474 267384 460480 267436
rect 460532 267424 460538 267436
rect 516778 267424 516784 267436
rect 460532 267396 516784 267424
rect 460532 267384 460538 267396
rect 516778 267384 516784 267396
rect 516836 267384 516842 267436
rect 519814 267384 519820 267436
rect 519872 267424 519878 267436
rect 583018 267424 583024 267436
rect 519872 267396 583024 267424
rect 519872 267384 519878 267396
rect 583018 267384 583024 267396
rect 583076 267384 583082 267436
rect 244090 267288 244096 267300
rect 238726 267260 244096 267288
rect 244090 267248 244096 267260
rect 244148 267248 244154 267300
rect 321922 267248 321928 267300
rect 321980 267288 321986 267300
rect 327718 267288 327724 267300
rect 321980 267260 327724 267288
rect 321980 267248 321986 267260
rect 327718 267248 327724 267260
rect 327776 267248 327782 267300
rect 350902 267248 350908 267300
rect 350960 267288 350966 267300
rect 362218 267288 362224 267300
rect 350960 267260 362224 267288
rect 350960 267248 350966 267260
rect 362218 267248 362224 267260
rect 362276 267248 362282 267300
rect 374454 267288 374460 267300
rect 369136 267260 374460 267288
rect 90358 267112 90364 267164
rect 90416 267152 90422 267164
rect 151354 267152 151360 267164
rect 90416 267124 151360 267152
rect 90416 267112 90422 267124
rect 151354 267112 151360 267124
rect 151412 267112 151418 267164
rect 159450 267112 159456 267164
rect 159508 267152 159514 267164
rect 162118 267152 162124 267164
rect 159508 267124 162124 267152
rect 159508 267112 159514 267124
rect 162118 267112 162124 267124
rect 162176 267112 162182 267164
rect 168098 267112 168104 267164
rect 168156 267152 168162 267164
rect 177022 267152 177028 267164
rect 168156 267124 177028 267152
rect 168156 267112 168162 267124
rect 177022 267112 177028 267124
rect 177080 267112 177086 267164
rect 177666 267112 177672 267164
rect 177724 267152 177730 267164
rect 214282 267152 214288 267164
rect 177724 267124 214288 267152
rect 177724 267112 177730 267124
rect 214282 267112 214288 267124
rect 214340 267112 214346 267164
rect 220078 267112 220084 267164
rect 220136 267152 220142 267164
rect 239122 267152 239128 267164
rect 220136 267124 239128 267152
rect 220136 267112 220142 267124
rect 239122 267112 239128 267124
rect 239180 267112 239186 267164
rect 246942 267112 246948 267164
rect 247000 267152 247006 267164
rect 263962 267152 263968 267164
rect 247000 267124 263968 267152
rect 247000 267112 247006 267124
rect 263962 267112 263968 267124
rect 264020 267112 264026 267164
rect 314470 267112 314476 267164
rect 314528 267152 314534 267164
rect 319254 267152 319260 267164
rect 314528 267124 319260 267152
rect 314528 267112 314534 267124
rect 319254 267112 319260 267124
rect 319312 267112 319318 267164
rect 360010 267112 360016 267164
rect 360068 267152 360074 267164
rect 366358 267152 366364 267164
rect 360068 267124 366364 267152
rect 360068 267112 360074 267124
rect 366358 267112 366364 267124
rect 366416 267112 366422 267164
rect 79318 266976 79324 267028
rect 79376 267016 79382 267028
rect 140222 267016 140228 267028
rect 79376 266988 140228 267016
rect 79376 266976 79382 266988
rect 140222 266976 140228 266988
rect 140280 266976 140286 267028
rect 140682 266976 140688 267028
rect 140740 267016 140746 267028
rect 186958 267016 186964 267028
rect 140740 266988 186964 267016
rect 140740 266976 140746 266988
rect 186958 266976 186964 266988
rect 187016 266976 187022 267028
rect 190454 266976 190460 267028
rect 190512 267016 190518 267028
rect 224218 267016 224224 267028
rect 190512 266988 224224 267016
rect 190512 266976 190518 266988
rect 224218 266976 224224 266988
rect 224276 266976 224282 267028
rect 228358 266976 228364 267028
rect 228416 267016 228422 267028
rect 248782 267016 248788 267028
rect 228416 266988 248788 267016
rect 228416 266976 228422 266988
rect 248782 266976 248788 266988
rect 248840 266976 248846 267028
rect 255958 266976 255964 267028
rect 256016 267016 256022 267028
rect 258994 267016 259000 267028
rect 256016 266988 259000 267016
rect 256016 266976 256022 266988
rect 258994 266976 259000 266988
rect 259052 266976 259058 267028
rect 286318 266976 286324 267028
rect 286376 267016 286382 267028
rect 287974 267016 287980 267028
rect 286376 266988 287980 267016
rect 286376 266976 286382 266988
rect 287974 266976 287980 266988
rect 288032 266976 288038 267028
rect 313642 266976 313648 267028
rect 313700 267016 313706 267028
rect 317414 267016 317420 267028
rect 313700 266988 317420 267016
rect 313700 266976 313706 266988
rect 317414 266976 317420 266988
rect 317472 266976 317478 267028
rect 353386 266976 353392 267028
rect 353444 267016 353450 267028
rect 369136 267016 369164 267260
rect 374454 267248 374460 267260
rect 374512 267248 374518 267300
rect 378778 267248 378784 267300
rect 378836 267288 378842 267300
rect 385678 267288 385684 267300
rect 378836 267260 385684 267288
rect 378836 267248 378842 267260
rect 385678 267248 385684 267260
rect 385736 267248 385742 267300
rect 398098 267248 398104 267300
rect 398156 267288 398162 267300
rect 417418 267288 417424 267300
rect 398156 267260 417424 267288
rect 398156 267248 398162 267260
rect 417418 267248 417424 267260
rect 417476 267248 417482 267300
rect 432874 267248 432880 267300
rect 432932 267288 432938 267300
rect 453298 267288 453304 267300
rect 432932 267260 453304 267288
rect 432932 267248 432938 267260
rect 453298 267248 453304 267260
rect 453356 267248 453362 267300
rect 462958 267288 462964 267300
rect 454972 267260 462964 267288
rect 373626 267112 373632 267164
rect 373684 267152 373690 267164
rect 392026 267152 392032 267164
rect 373684 267124 392032 267152
rect 373684 267112 373690 267124
rect 392026 267112 392032 267124
rect 392084 267112 392090 267164
rect 399754 267112 399760 267164
rect 399812 267152 399818 267164
rect 407758 267152 407764 267164
rect 399812 267124 407764 267152
rect 399812 267112 399818 267124
rect 407758 267112 407764 267124
rect 407816 267112 407822 267164
rect 413002 267112 413008 267164
rect 413060 267152 413066 267164
rect 441614 267152 441620 267164
rect 413060 267124 441620 267152
rect 413060 267112 413066 267124
rect 441614 267112 441620 267124
rect 441672 267112 441678 267164
rect 447134 267112 447140 267164
rect 447192 267152 447198 267164
rect 448422 267152 448428 267164
rect 447192 267124 448428 267152
rect 447192 267112 447198 267124
rect 448422 267112 448428 267124
rect 448480 267112 448486 267164
rect 452746 267112 452752 267164
rect 452804 267152 452810 267164
rect 454972 267152 455000 267260
rect 462958 267248 462964 267260
rect 463016 267248 463022 267300
rect 465166 267248 465172 267300
rect 465224 267288 465230 267300
rect 523678 267288 523684 267300
rect 465224 267260 523684 267288
rect 465224 267248 465230 267260
rect 523678 267248 523684 267260
rect 523736 267248 523742 267300
rect 524782 267248 524788 267300
rect 524840 267288 524846 267300
rect 611998 267288 612004 267300
rect 524840 267260 612004 267288
rect 524840 267248 524846 267260
rect 611998 267248 612004 267260
rect 612056 267248 612062 267300
rect 452804 267124 455000 267152
rect 452804 267112 452810 267124
rect 455138 267112 455144 267164
rect 455196 267152 455202 267164
rect 515398 267152 515404 267164
rect 455196 267124 515404 267152
rect 455196 267112 455202 267124
rect 515398 267112 515404 267124
rect 515456 267112 515462 267164
rect 517238 267112 517244 267164
rect 517296 267152 517302 267164
rect 527174 267152 527180 267164
rect 517296 267124 527180 267152
rect 517296 267112 517302 267124
rect 527174 267112 527180 267124
rect 527232 267112 527238 267164
rect 529658 267112 529664 267164
rect 529716 267152 529722 267164
rect 617518 267152 617524 267164
rect 529716 267124 617524 267152
rect 529716 267112 529722 267124
rect 617518 267112 617524 267124
rect 617576 267112 617582 267164
rect 353444 266988 369164 267016
rect 353444 266976 353450 266988
rect 393130 266976 393136 267028
rect 393188 267016 393194 267028
rect 420178 267016 420184 267028
rect 393188 266988 420184 267016
rect 393188 266976 393194 266988
rect 420178 266976 420184 266988
rect 420236 266976 420242 267028
rect 457438 267016 457444 267028
rect 431926 266988 457444 267016
rect 132494 266840 132500 266892
rect 132552 266880 132558 266892
rect 147214 266880 147220 266892
rect 132552 266852 147220 266880
rect 132552 266840 132558 266852
rect 147214 266840 147220 266852
rect 147272 266840 147278 266892
rect 153838 266840 153844 266892
rect 153896 266880 153902 266892
rect 184474 266880 184480 266892
rect 153896 266852 184480 266880
rect 153896 266840 153902 266852
rect 184474 266840 184480 266852
rect 184532 266840 184538 266892
rect 218698 266840 218704 266892
rect 218756 266880 218762 266892
rect 220906 266880 220912 266892
rect 218756 266852 220912 266880
rect 218756 266840 218762 266852
rect 220906 266840 220912 266852
rect 220964 266840 220970 266892
rect 312814 266840 312820 266892
rect 312872 266880 312878 266892
rect 316034 266880 316040 266892
rect 312872 266852 316040 266880
rect 312872 266840 312878 266852
rect 316034 266840 316040 266852
rect 316092 266840 316098 266892
rect 332686 266840 332692 266892
rect 332744 266880 332750 266892
rect 343818 266880 343824 266892
rect 332744 266852 343824 266880
rect 332744 266840 332750 266852
rect 343818 266840 343824 266852
rect 343876 266840 343882 266892
rect 374914 266840 374920 266892
rect 374972 266880 374978 266892
rect 380526 266880 380532 266892
rect 374972 266852 380532 266880
rect 374972 266840 374978 266852
rect 380526 266840 380532 266852
rect 380584 266840 380590 266892
rect 388162 266840 388168 266892
rect 388220 266880 388226 266892
rect 388220 266852 402974 266880
rect 388220 266840 388226 266852
rect 317782 266772 317788 266824
rect 317840 266812 317846 266824
rect 322934 266812 322940 266824
rect 317840 266784 322940 266812
rect 317840 266772 317846 266784
rect 322934 266772 322940 266784
rect 322992 266772 322998 266824
rect 137462 266704 137468 266756
rect 137520 266744 137526 266756
rect 150526 266744 150532 266756
rect 137520 266716 150532 266744
rect 137520 266704 137526 266716
rect 150526 266704 150532 266716
rect 150584 266704 150590 266756
rect 151078 266704 151084 266756
rect 151136 266744 151142 266756
rect 179506 266744 179512 266756
rect 151136 266716 179512 266744
rect 151136 266704 151142 266716
rect 179506 266704 179512 266716
rect 179564 266704 179570 266756
rect 368290 266704 368296 266756
rect 368348 266744 368354 266756
rect 378778 266744 378784 266756
rect 368348 266716 378784 266744
rect 368348 266704 368354 266716
rect 378778 266704 378784 266716
rect 378836 266704 378842 266756
rect 394694 266744 394700 266756
rect 383626 266716 394700 266744
rect 308674 266636 308680 266688
rect 308732 266676 308738 266688
rect 310606 266676 310612 266688
rect 308732 266648 310612 266676
rect 308732 266636 308738 266648
rect 310606 266636 310612 266648
rect 310664 266636 310670 266688
rect 316954 266636 316960 266688
rect 317012 266676 317018 266688
rect 321554 266676 321560 266688
rect 317012 266648 321560 266676
rect 317012 266636 317018 266648
rect 321554 266636 321560 266648
rect 321612 266636 321618 266688
rect 347498 266636 347504 266688
rect 347556 266676 347562 266688
rect 351178 266676 351184 266688
rect 347556 266648 351184 266676
rect 347556 266636 347562 266648
rect 351178 266636 351184 266648
rect 351236 266636 351242 266688
rect 130378 266568 130384 266620
rect 130436 266608 130442 266620
rect 138106 266608 138112 266620
rect 130436 266580 138112 266608
rect 130436 266568 130442 266580
rect 138106 266568 138112 266580
rect 138164 266568 138170 266620
rect 149606 266568 149612 266620
rect 149664 266608 149670 266620
rect 159634 266608 159640 266620
rect 149664 266580 159640 266608
rect 149664 266568 149670 266580
rect 159634 266568 159640 266580
rect 159692 266568 159698 266620
rect 378226 266568 378232 266620
rect 378284 266608 378290 266620
rect 383626 266608 383654 266716
rect 394694 266704 394700 266716
rect 394752 266704 394758 266756
rect 402946 266744 402974 266852
rect 427906 266840 427912 266892
rect 427964 266880 427970 266892
rect 431926 266880 431954 266988
rect 457438 266976 457444 266988
rect 457496 266976 457502 267028
rect 470134 266976 470140 267028
rect 470192 267016 470198 267028
rect 534718 267016 534724 267028
rect 470192 266988 534724 267016
rect 470192 266976 470198 266988
rect 534718 266976 534724 266988
rect 534776 266976 534782 267028
rect 535546 266976 535552 267028
rect 535604 267016 535610 267028
rect 536742 267016 536748 267028
rect 535604 266988 536748 267016
rect 535604 266976 535610 266988
rect 536742 266976 536748 266988
rect 536800 266976 536806 267028
rect 539686 266976 539692 267028
rect 539744 267016 539750 267028
rect 634078 267016 634084 267028
rect 539744 266988 634084 267016
rect 539744 266976 539750 266988
rect 634078 266976 634084 266988
rect 634136 266976 634142 267028
rect 427964 266852 431954 266880
rect 427964 266840 427970 266852
rect 442718 266840 442724 266892
rect 442776 266880 442782 266892
rect 485038 266880 485044 266892
rect 442776 266852 485044 266880
rect 442776 266840 442782 266852
rect 485038 266840 485044 266852
rect 485096 266840 485102 266892
rect 499942 266840 499948 266892
rect 500000 266880 500006 266892
rect 507854 266880 507860 266892
rect 500000 266852 507860 266880
rect 500000 266840 500006 266852
rect 507854 266840 507860 266852
rect 507912 266840 507918 266892
rect 534718 266840 534724 266892
rect 534776 266880 534782 266892
rect 589918 266880 589924 266892
rect 534776 266852 589924 266880
rect 534776 266840 534782 266852
rect 589918 266840 589924 266852
rect 589976 266840 589982 266892
rect 404354 266744 404360 266756
rect 402946 266716 404360 266744
rect 404354 266704 404360 266716
rect 404412 266704 404418 266756
rect 408034 266704 408040 266756
rect 408092 266744 408098 266756
rect 423950 266744 423956 266756
rect 408092 266716 423956 266744
rect 408092 266704 408098 266716
rect 423950 266704 423956 266716
rect 424008 266704 424014 266756
rect 434530 266704 434536 266756
rect 434588 266744 434594 266756
rect 449158 266744 449164 266756
rect 434588 266716 449164 266744
rect 434588 266704 434594 266716
rect 449158 266704 449164 266716
rect 449216 266704 449222 266756
rect 457714 266704 457720 266756
rect 457772 266744 457778 266756
rect 476758 266744 476764 266756
rect 457772 266716 476764 266744
rect 457772 266704 457778 266716
rect 476758 266704 476764 266716
rect 476816 266704 476822 266756
rect 485038 266704 485044 266756
rect 485096 266744 485102 266756
rect 485096 266716 489914 266744
rect 485096 266704 485102 266716
rect 378284 266580 383654 266608
rect 378284 266568 378290 266580
rect 394786 266568 394792 266620
rect 394844 266608 394850 266620
rect 403618 266608 403624 266620
rect 394844 266580 403624 266608
rect 394844 266568 394850 266580
rect 403618 266568 403624 266580
rect 403676 266568 403682 266620
rect 407206 266568 407212 266620
rect 407264 266608 407270 266620
rect 414658 266608 414664 266620
rect 407264 266580 414664 266608
rect 407264 266568 407270 266580
rect 414658 266568 414664 266580
rect 414716 266568 414722 266620
rect 437842 266568 437848 266620
rect 437900 266608 437906 266620
rect 447134 266608 447140 266620
rect 437900 266580 447140 266608
rect 437900 266568 437906 266580
rect 447134 266568 447140 266580
rect 447192 266568 447198 266620
rect 489886 266608 489914 266716
rect 490006 266704 490012 266756
rect 490064 266744 490070 266756
rect 509694 266744 509700 266756
rect 490064 266716 509700 266744
rect 490064 266704 490070 266716
rect 509694 266704 509700 266716
rect 509752 266704 509758 266756
rect 510706 266704 510712 266756
rect 510764 266744 510770 266756
rect 511810 266744 511816 266756
rect 510764 266716 511816 266744
rect 510764 266704 510770 266716
rect 511810 266704 511816 266716
rect 511868 266704 511874 266756
rect 512362 266704 512368 266756
rect 512420 266744 512426 266756
rect 513190 266744 513196 266756
rect 512420 266716 513196 266744
rect 512420 266704 512426 266716
rect 513190 266704 513196 266716
rect 513248 266704 513254 266756
rect 516502 266704 516508 266756
rect 516560 266744 516566 266756
rect 517422 266744 517428 266756
rect 516560 266716 517428 266744
rect 516560 266704 516566 266716
rect 517422 266704 517428 266716
rect 517480 266704 517486 266756
rect 518986 266704 518992 266756
rect 519044 266744 519050 266756
rect 520090 266744 520096 266756
rect 519044 266716 520096 266744
rect 519044 266704 519050 266716
rect 520090 266704 520096 266716
rect 520148 266704 520154 266756
rect 527266 266704 527272 266756
rect 527324 266744 527330 266756
rect 528186 266744 528192 266756
rect 527324 266716 528192 266744
rect 527324 266704 527330 266716
rect 528186 266704 528192 266716
rect 528244 266704 528250 266756
rect 528922 266704 528928 266756
rect 528980 266744 528986 266756
rect 529842 266744 529848 266756
rect 528980 266716 529848 266744
rect 528980 266704 528986 266716
rect 529842 266704 529848 266716
rect 529900 266704 529906 266756
rect 531406 266704 531412 266756
rect 531464 266744 531470 266756
rect 532602 266744 532608 266756
rect 531464 266716 532608 266744
rect 531464 266704 531470 266716
rect 532602 266704 532608 266716
rect 532660 266704 532666 266756
rect 533062 266704 533068 266756
rect 533120 266744 533126 266756
rect 533982 266744 533988 266756
rect 533120 266716 533988 266744
rect 533120 266704 533126 266716
rect 533982 266704 533988 266716
rect 534040 266704 534046 266756
rect 542998 266704 543004 266756
rect 543056 266744 543062 266756
rect 598198 266744 598204 266756
rect 543056 266716 598204 266744
rect 543056 266704 543062 266716
rect 598198 266704 598204 266716
rect 598256 266704 598262 266756
rect 501598 266608 501604 266620
rect 489886 266580 501604 266608
rect 501598 266568 501604 266580
rect 501656 266568 501662 266620
rect 504818 266568 504824 266620
rect 504876 266608 504882 266620
rect 556798 266608 556804 266620
rect 504876 266580 556804 266608
rect 504876 266568 504882 266580
rect 556798 266568 556804 266580
rect 556856 266568 556862 266620
rect 250438 266500 250444 266552
rect 250496 266540 250502 266552
rect 256510 266540 256516 266552
rect 250496 266512 256516 266540
rect 250496 266500 250502 266512
rect 256510 266500 256516 266512
rect 256568 266500 256574 266552
rect 310330 266500 310336 266552
rect 310388 266540 310394 266552
rect 311894 266540 311900 266552
rect 310388 266512 311900 266540
rect 310388 266500 310394 266512
rect 311894 266500 311900 266512
rect 311952 266500 311958 266552
rect 312354 266500 312360 266552
rect 312412 266540 312418 266552
rect 314654 266540 314660 266552
rect 312412 266512 314660 266540
rect 312412 266500 312418 266512
rect 314654 266500 314660 266512
rect 314712 266500 314718 266552
rect 316126 266500 316132 266552
rect 316184 266540 316190 266552
rect 320174 266540 320180 266552
rect 316184 266512 320180 266540
rect 316184 266500 316190 266512
rect 320174 266500 320180 266512
rect 320232 266500 320238 266552
rect 327718 266500 327724 266552
rect 327776 266540 327782 266552
rect 331950 266540 331956 266552
rect 327776 266512 331956 266540
rect 327776 266500 327782 266512
rect 331950 266500 331956 266512
rect 332008 266500 332014 266552
rect 345106 266500 345112 266552
rect 345164 266540 345170 266552
rect 348418 266540 348424 266552
rect 345164 266512 348424 266540
rect 345164 266500 345170 266512
rect 348418 266500 348424 266512
rect 348476 266500 348482 266552
rect 350074 266500 350080 266552
rect 350132 266540 350138 266552
rect 353938 266540 353944 266552
rect 350132 266512 353944 266540
rect 350132 266500 350138 266512
rect 353938 266500 353944 266512
rect 353996 266500 354002 266552
rect 355870 266500 355876 266552
rect 355928 266540 355934 266552
rect 360838 266540 360844 266552
rect 355928 266512 360844 266540
rect 355928 266500 355934 266512
rect 360838 266500 360844 266512
rect 360896 266500 360902 266552
rect 369946 266500 369952 266552
rect 370004 266540 370010 266552
rect 372246 266540 372252 266552
rect 370004 266512 372252 266540
rect 370004 266500 370010 266512
rect 372246 266500 372252 266512
rect 372304 266500 372310 266552
rect 423766 266500 423772 266552
rect 423824 266540 423830 266552
rect 425698 266540 425704 266552
rect 423824 266512 425704 266540
rect 423824 266500 423830 266512
rect 425698 266500 425704 266512
rect 425756 266500 425762 266552
rect 426250 266500 426256 266552
rect 426308 266540 426314 266552
rect 428458 266540 428464 266552
rect 426308 266512 428464 266540
rect 426308 266500 426314 266512
rect 428458 266500 428464 266512
rect 428516 266500 428522 266552
rect 447778 266500 447784 266552
rect 447836 266540 447842 266552
rect 456058 266540 456064 266552
rect 447836 266512 456064 266540
rect 447836 266500 447842 266512
rect 456058 266500 456064 266512
rect 456116 266500 456122 266552
rect 491662 266432 491668 266484
rect 491720 266472 491726 266484
rect 492582 266472 492588 266484
rect 491720 266444 492588 266472
rect 491720 266432 491726 266444
rect 492582 266432 492588 266444
rect 492640 266432 492646 266484
rect 494146 266432 494152 266484
rect 494204 266472 494210 266484
rect 495066 266472 495072 266484
rect 494204 266444 495072 266472
rect 494204 266432 494210 266444
rect 495066 266432 495072 266444
rect 495124 266432 495130 266484
rect 502426 266432 502432 266484
rect 502484 266472 502490 266484
rect 503438 266472 503444 266484
rect 502484 266444 503444 266472
rect 502484 266432 502490 266444
rect 503438 266432 503444 266444
rect 503496 266432 503502 266484
rect 504082 266432 504088 266484
rect 504140 266472 504146 266484
rect 505002 266472 505008 266484
rect 504140 266444 505008 266472
rect 504140 266432 504146 266444
rect 505002 266432 505008 266444
rect 505060 266432 505066 266484
rect 506566 266432 506572 266484
rect 506624 266472 506630 266484
rect 507670 266472 507676 266484
rect 506624 266444 507676 266472
rect 506624 266432 506630 266444
rect 507670 266432 507676 266444
rect 507728 266432 507734 266484
rect 507854 266432 507860 266484
rect 507912 266472 507918 266484
rect 549898 266472 549904 266484
rect 507912 266444 549904 266472
rect 507912 266432 507918 266444
rect 549898 266432 549904 266444
rect 549956 266432 549962 266484
rect 163498 266364 163504 266416
rect 163556 266404 163562 266416
rect 167086 266404 167092 266416
rect 163556 266376 167092 266404
rect 163556 266364 163562 266376
rect 167086 266364 167092 266376
rect 167144 266364 167150 266416
rect 211154 266364 211160 266416
rect 211212 266404 211218 266416
rect 213454 266404 213460 266416
rect 211212 266376 213460 266404
rect 211212 266364 211218 266376
rect 213454 266364 213460 266376
rect 213512 266364 213518 266416
rect 214558 266364 214564 266416
rect 214616 266404 214622 266416
rect 215938 266404 215944 266416
rect 214616 266376 215944 266404
rect 214616 266364 214622 266376
rect 215938 266364 215944 266376
rect 215996 266364 216002 266416
rect 239398 266364 239404 266416
rect 239456 266404 239462 266416
rect 241606 266404 241612 266416
rect 239456 266376 241612 266404
rect 239456 266364 239462 266376
rect 241606 266364 241612 266376
rect 241664 266364 241670 266416
rect 243538 266364 243544 266416
rect 243596 266404 243602 266416
rect 246574 266404 246580 266416
rect 243596 266376 246580 266404
rect 243596 266364 243602 266376
rect 246574 266364 246580 266376
rect 246632 266364 246638 266416
rect 249058 266364 249064 266416
rect 249116 266404 249122 266416
rect 250714 266404 250720 266416
rect 249116 266376 250720 266404
rect 249116 266364 249122 266376
rect 250714 266364 250720 266376
rect 250772 266364 250778 266416
rect 300946 266364 300952 266416
rect 301004 266404 301010 266416
rect 302050 266404 302056 266416
rect 301004 266376 302056 266404
rect 301004 266364 301010 266376
rect 302050 266364 302056 266376
rect 302108 266364 302114 266416
rect 303706 266364 303712 266416
rect 303764 266404 303770 266416
rect 304534 266404 304540 266416
rect 303764 266376 304540 266404
rect 303764 266364 303770 266376
rect 304534 266364 304540 266376
rect 304592 266364 304598 266416
rect 307846 266364 307852 266416
rect 307904 266404 307910 266416
rect 309134 266404 309140 266416
rect 307904 266376 309140 266404
rect 307904 266364 307910 266376
rect 309134 266364 309140 266376
rect 309192 266364 309198 266416
rect 309502 266364 309508 266416
rect 309560 266404 309566 266416
rect 310790 266404 310796 266416
rect 309560 266376 310796 266404
rect 309560 266364 309566 266376
rect 310790 266364 310796 266376
rect 310848 266364 310854 266416
rect 311158 266364 311164 266416
rect 311216 266404 311222 266416
rect 313274 266404 313280 266416
rect 311216 266376 313280 266404
rect 311216 266364 311222 266376
rect 313274 266364 313280 266376
rect 313332 266364 313338 266416
rect 320266 266364 320272 266416
rect 320324 266404 320330 266416
rect 321370 266404 321376 266416
rect 320324 266376 321376 266404
rect 320324 266364 320330 266376
rect 321370 266364 321376 266376
rect 321428 266364 321434 266416
rect 324406 266364 324412 266416
rect 324464 266404 324470 266416
rect 325326 266404 325332 266416
rect 324464 266376 325332 266404
rect 324464 266364 324470 266376
rect 325326 266364 325332 266376
rect 325384 266364 325390 266416
rect 328546 266364 328552 266416
rect 328604 266404 328610 266416
rect 329742 266404 329748 266416
rect 328604 266376 329748 266404
rect 328604 266364 328610 266376
rect 329742 266364 329748 266376
rect 329800 266364 329806 266416
rect 336826 266364 336832 266416
rect 336884 266404 336890 266416
rect 337930 266404 337936 266416
rect 336884 266376 337936 266404
rect 336884 266364 336890 266376
rect 337930 266364 337936 266376
rect 337988 266364 337994 266416
rect 342622 266364 342628 266416
rect 342680 266404 342686 266416
rect 345290 266404 345296 266416
rect 342680 266376 345296 266404
rect 342680 266364 342686 266376
rect 345290 266364 345296 266376
rect 345348 266364 345354 266416
rect 346762 266364 346768 266416
rect 346820 266404 346826 266416
rect 347682 266404 347688 266416
rect 346820 266376 347688 266404
rect 346820 266364 346826 266376
rect 347682 266364 347688 266376
rect 347740 266364 347746 266416
rect 349246 266364 349252 266416
rect 349304 266404 349310 266416
rect 350350 266404 350356 266416
rect 349304 266376 350356 266404
rect 349304 266364 349310 266376
rect 350350 266364 350356 266376
rect 350408 266364 350414 266416
rect 357526 266364 357532 266416
rect 357584 266404 357590 266416
rect 359458 266404 359464 266416
rect 357584 266376 359464 266404
rect 357584 266364 357590 266376
rect 359458 266364 359464 266376
rect 359516 266364 359522 266416
rect 361666 266364 361672 266416
rect 361724 266404 361730 266416
rect 362770 266404 362776 266416
rect 361724 266376 362776 266404
rect 361724 266364 361730 266376
rect 362770 266364 362776 266376
rect 362828 266364 362834 266416
rect 369118 266364 369124 266416
rect 369176 266404 369182 266416
rect 370498 266404 370504 266416
rect 369176 266376 370504 266404
rect 369176 266364 369182 266376
rect 370498 266364 370504 266376
rect 370556 266364 370562 266416
rect 371602 266364 371608 266416
rect 371660 266404 371666 266416
rect 373258 266404 373264 266416
rect 371660 266376 373264 266404
rect 371660 266364 371666 266376
rect 373258 266364 373264 266376
rect 373316 266364 373322 266416
rect 374086 266364 374092 266416
rect 374144 266404 374150 266416
rect 375282 266404 375288 266416
rect 374144 266376 375288 266404
rect 374144 266364 374150 266376
rect 375282 266364 375288 266376
rect 375340 266364 375346 266416
rect 379882 266364 379888 266416
rect 379940 266404 379946 266416
rect 383010 266404 383016 266416
rect 379940 266376 383016 266404
rect 379940 266364 379946 266376
rect 383010 266364 383016 266376
rect 383068 266364 383074 266416
rect 384022 266364 384028 266416
rect 384080 266404 384086 266416
rect 384942 266404 384948 266416
rect 384080 266376 384948 266404
rect 384080 266364 384086 266376
rect 384942 266364 384948 266376
rect 385000 266364 385006 266416
rect 386506 266364 386512 266416
rect 386564 266404 386570 266416
rect 387702 266404 387708 266416
rect 386564 266376 387708 266404
rect 386564 266364 386570 266376
rect 387702 266364 387708 266376
rect 387760 266364 387766 266416
rect 392302 266364 392308 266416
rect 392360 266404 392366 266416
rect 393682 266404 393688 266416
rect 392360 266376 393688 266404
rect 392360 266364 392366 266376
rect 393682 266364 393688 266376
rect 393740 266364 393746 266416
rect 398926 266364 398932 266416
rect 398984 266404 398990 266416
rect 400030 266404 400036 266416
rect 398984 266376 400036 266404
rect 398984 266364 398990 266376
rect 400030 266364 400036 266376
rect 400088 266364 400094 266416
rect 408862 266364 408868 266416
rect 408920 266404 408926 266416
rect 409782 266404 409788 266416
rect 408920 266376 409788 266404
rect 408920 266364 408926 266376
rect 409782 266364 409788 266376
rect 409840 266364 409846 266416
rect 411346 266364 411352 266416
rect 411404 266404 411410 266416
rect 412266 266404 412272 266416
rect 411404 266376 412272 266404
rect 411404 266364 411410 266376
rect 412266 266364 412272 266376
rect 412324 266364 412330 266416
rect 415486 266364 415492 266416
rect 415544 266404 415550 266416
rect 416406 266404 416412 266416
rect 415544 266376 416412 266404
rect 415544 266364 415550 266376
rect 416406 266364 416412 266376
rect 416464 266364 416470 266416
rect 417970 266364 417976 266416
rect 418028 266404 418034 266416
rect 418798 266404 418804 266416
rect 418028 266376 418804 266404
rect 418028 266364 418034 266376
rect 418798 266364 418804 266376
rect 418856 266364 418862 266416
rect 425422 266364 425428 266416
rect 425480 266404 425486 266416
rect 427078 266404 427084 266416
rect 425480 266376 427084 266404
rect 425480 266364 425486 266376
rect 427078 266364 427084 266376
rect 427136 266364 427142 266416
rect 429562 266364 429568 266416
rect 429620 266404 429626 266416
rect 430390 266404 430396 266416
rect 429620 266376 430396 266404
rect 429620 266364 429626 266376
rect 430390 266364 430396 266376
rect 430448 266364 430454 266416
rect 432046 266364 432052 266416
rect 432104 266404 432110 266416
rect 433150 266404 433156 266416
rect 432104 266376 433156 266404
rect 432104 266364 432110 266376
rect 433150 266364 433156 266376
rect 433208 266364 433214 266416
rect 440326 266364 440332 266416
rect 440384 266404 440390 266416
rect 441338 266404 441344 266416
rect 440384 266376 441344 266404
rect 440384 266364 440390 266376
rect 441338 266364 441344 266376
rect 441396 266364 441402 266416
rect 441982 266364 441988 266416
rect 442040 266404 442046 266416
rect 442902 266404 442908 266416
rect 442040 266376 442908 266404
rect 442040 266364 442046 266376
rect 442902 266364 442908 266376
rect 442960 266364 442966 266416
rect 444466 266364 444472 266416
rect 444524 266404 444530 266416
rect 445662 266404 445668 266416
rect 444524 266376 445668 266404
rect 444524 266364 444530 266376
rect 445662 266364 445668 266376
rect 445720 266364 445726 266416
rect 448606 266364 448612 266416
rect 448664 266404 448670 266416
rect 450538 266404 450544 266416
rect 448664 266376 450544 266404
rect 448664 266364 448670 266376
rect 450538 266364 450544 266376
rect 450596 266364 450602 266416
rect 454402 266364 454408 266416
rect 454460 266404 454466 266416
rect 455322 266404 455328 266416
rect 454460 266376 455328 266404
rect 454460 266364 454466 266376
rect 455322 266364 455328 266376
rect 455380 266364 455386 266416
rect 456886 266364 456892 266416
rect 456944 266404 456950 266416
rect 457990 266404 457996 266416
rect 456944 266376 457996 266404
rect 456944 266364 456950 266376
rect 457990 266364 457996 266376
rect 458048 266364 458054 266416
rect 459370 266364 459376 266416
rect 459428 266404 459434 266416
rect 460198 266404 460204 266416
rect 459428 266376 460204 266404
rect 459428 266364 459434 266376
rect 460198 266364 460204 266376
rect 460256 266364 460262 266416
rect 473446 266364 473452 266416
rect 473504 266404 473510 266416
rect 474642 266404 474648 266416
rect 473504 266376 474648 266404
rect 473504 266364 473510 266376
rect 474642 266364 474648 266376
rect 474700 266364 474706 266416
rect 475102 266364 475108 266416
rect 475160 266404 475166 266416
rect 479518 266404 479524 266416
rect 475160 266376 479524 266404
rect 475160 266364 475166 266376
rect 479518 266364 479524 266376
rect 479576 266364 479582 266416
rect 481726 266364 481732 266416
rect 481784 266404 481790 266416
rect 482830 266404 482836 266416
rect 481784 266376 482836 266404
rect 481784 266364 481790 266376
rect 482830 266364 482836 266376
rect 482888 266364 482894 266416
rect 483382 266364 483388 266416
rect 483440 266404 483446 266416
rect 484210 266404 484216 266416
rect 483440 266376 484216 266404
rect 483440 266364 483446 266376
rect 484210 266364 484216 266376
rect 484268 266364 484274 266416
rect 485866 266364 485872 266416
rect 485924 266404 485930 266416
rect 486786 266404 486792 266416
rect 485924 266376 486792 266404
rect 485924 266364 485930 266376
rect 486786 266364 486792 266376
rect 486844 266364 486850 266416
rect 487154 266296 487160 266348
rect 487212 266336 487218 266348
rect 557718 266336 557724 266348
rect 487212 266308 557724 266336
rect 487212 266296 487218 266308
rect 557718 266296 557724 266308
rect 557776 266296 557782 266348
rect 484210 266160 484216 266212
rect 484268 266200 484274 266212
rect 560294 266200 560300 266212
rect 484268 266172 560300 266200
rect 484268 266160 484274 266172
rect 560294 266160 560300 266172
rect 560352 266160 560358 266212
rect 482554 266024 482560 266076
rect 482612 266064 482618 266076
rect 487154 266064 487160 266076
rect 482612 266036 487160 266064
rect 482612 266024 482618 266036
rect 487154 266024 487160 266036
rect 487212 266024 487218 266076
rect 492490 266024 492496 266076
rect 492548 266064 492554 266076
rect 572714 266064 572720 266076
rect 492548 266036 572720 266064
rect 492548 266024 492554 266036
rect 572714 266024 572720 266036
rect 572772 266024 572778 266076
rect 513190 265888 513196 265940
rect 513248 265928 513254 265940
rect 601694 265928 601700 265940
rect 513248 265900 601700 265928
rect 513248 265888 513254 265900
rect 601694 265888 601700 265900
rect 601752 265888 601758 265940
rect 515674 265752 515680 265804
rect 515732 265792 515738 265804
rect 605834 265792 605840 265804
rect 515732 265764 605840 265792
rect 515732 265752 515738 265764
rect 605834 265752 605840 265764
rect 605892 265752 605898 265804
rect 209774 265616 209780 265668
rect 209832 265656 209838 265668
rect 210694 265656 210700 265668
rect 209832 265628 210700 265656
rect 209832 265616 209838 265628
rect 210694 265616 210700 265628
rect 210752 265616 210758 265668
rect 224954 265616 224960 265668
rect 225012 265656 225018 265668
rect 225598 265656 225604 265668
rect 225012 265628 225604 265656
rect 225012 265616 225018 265628
rect 225598 265616 225604 265628
rect 225656 265616 225662 265668
rect 280338 265616 280344 265668
rect 280396 265656 280402 265668
rect 280982 265656 280988 265668
rect 280396 265628 280988 265656
rect 280396 265616 280402 265628
rect 280982 265616 280988 265628
rect 281040 265616 281046 265668
rect 292666 265616 292672 265668
rect 292724 265656 292730 265668
rect 293494 265656 293500 265668
rect 292724 265628 293500 265656
rect 292724 265616 292730 265628
rect 293494 265616 293500 265628
rect 293552 265616 293558 265668
rect 520642 265616 520648 265668
rect 520700 265656 520706 265668
rect 612734 265656 612740 265668
rect 520700 265628 612740 265656
rect 520700 265616 520706 265628
rect 612734 265616 612740 265628
rect 612792 265616 612798 265668
rect 479242 265480 479248 265532
rect 479300 265520 479306 265532
rect 553394 265520 553400 265532
rect 479300 265492 553400 265520
rect 479300 265480 479306 265492
rect 553394 265480 553400 265492
rect 553452 265480 553458 265532
rect 477586 265344 477592 265396
rect 477644 265384 477650 265396
rect 550634 265384 550640 265396
rect 477644 265356 550640 265384
rect 477644 265344 477650 265356
rect 550634 265344 550640 265356
rect 550692 265344 550698 265396
rect 469306 265208 469312 265260
rect 469364 265248 469370 265260
rect 539962 265248 539968 265260
rect 469364 265220 539968 265248
rect 469364 265208 469370 265220
rect 539962 265208 539968 265220
rect 540020 265208 540026 265260
rect 466822 265072 466828 265124
rect 466880 265112 466886 265124
rect 535730 265112 535736 265124
rect 466880 265084 535736 265112
rect 466880 265072 466886 265084
rect 535730 265072 535736 265084
rect 535788 265072 535794 265124
rect 58618 264460 58624 264512
rect 58676 264500 58682 264512
rect 669130 264500 669136 264512
rect 58676 264472 669136 264500
rect 58676 264460 58682 264472
rect 669130 264460 669136 264472
rect 669188 264460 669194 264512
rect 53098 264324 53104 264376
rect 53156 264364 53162 264376
rect 668210 264364 668216 264376
rect 53156 264336 668216 264364
rect 53156 264324 53162 264336
rect 668210 264324 668216 264336
rect 668268 264324 668274 264376
rect 46198 264188 46204 264240
rect 46256 264228 46262 264240
rect 668946 264228 668952 264240
rect 46256 264200 668952 264228
rect 46256 264188 46262 264200
rect 668946 264188 668952 264200
rect 669004 264188 669010 264240
rect 570598 261468 570604 261520
rect 570656 261508 570662 261520
rect 645854 261508 645860 261520
rect 570656 261480 645860 261508
rect 570656 261468 570662 261480
rect 645854 261468 645860 261480
rect 645912 261468 645918 261520
rect 554406 260856 554412 260908
rect 554464 260896 554470 260908
rect 568574 260896 568580 260908
rect 554464 260868 568580 260896
rect 554464 260856 554470 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 554314 259428 554320 259480
rect 554372 259468 554378 259480
rect 563698 259468 563704 259480
rect 554372 259440 563704 259468
rect 554372 259428 554378 259440
rect 563698 259428 563704 259440
rect 563756 259428 563762 259480
rect 675846 259428 675852 259480
rect 675904 259468 675910 259480
rect 676398 259468 676404 259480
rect 675904 259440 676404 259468
rect 675904 259428 675910 259440
rect 676398 259428 676404 259440
rect 676456 259428 676462 259480
rect 35802 256776 35808 256828
rect 35860 256816 35866 256828
rect 39574 256816 39580 256828
rect 35860 256788 39580 256816
rect 35860 256776 35866 256788
rect 39574 256776 39580 256788
rect 39632 256776 39638 256828
rect 553946 256708 553952 256760
rect 554004 256748 554010 256760
rect 560938 256748 560944 256760
rect 554004 256720 560944 256748
rect 554004 256708 554010 256720
rect 560938 256708 560944 256720
rect 560996 256708 561002 256760
rect 554498 255552 554504 255604
rect 554556 255592 554562 255604
rect 558178 255592 558184 255604
rect 554556 255564 558184 255592
rect 554556 255552 554562 255564
rect 558178 255552 558184 255564
rect 558236 255552 558242 255604
rect 35802 255416 35808 255468
rect 35860 255456 35866 255468
rect 40494 255456 40500 255468
rect 35860 255428 40500 255456
rect 35860 255416 35866 255428
rect 40494 255416 40500 255428
rect 40552 255416 40558 255468
rect 35618 255280 35624 255332
rect 35676 255320 35682 255332
rect 41690 255320 41696 255332
rect 35676 255292 41696 255320
rect 35676 255280 35682 255292
rect 41690 255280 41696 255292
rect 41748 255280 41754 255332
rect 42058 255280 42064 255332
rect 42116 255320 42122 255332
rect 42794 255320 42800 255332
rect 42116 255292 42800 255320
rect 42116 255280 42122 255292
rect 42794 255280 42800 255292
rect 42852 255280 42858 255332
rect 35802 254328 35808 254380
rect 35860 254368 35866 254380
rect 40678 254368 40684 254380
rect 35860 254340 40684 254368
rect 35860 254328 35866 254340
rect 40678 254328 40684 254340
rect 40736 254328 40742 254380
rect 35802 254056 35808 254108
rect 35860 254096 35866 254108
rect 41506 254096 41512 254108
rect 35860 254068 41512 254096
rect 35860 254056 35866 254068
rect 41506 254056 41512 254068
rect 41564 254056 41570 254108
rect 35618 253920 35624 253972
rect 35676 253960 35682 253972
rect 39942 253960 39948 253972
rect 35676 253932 39948 253960
rect 35676 253920 35682 253932
rect 39942 253920 39948 253932
rect 40000 253920 40006 253972
rect 675846 253104 675852 253156
rect 675904 253144 675910 253156
rect 679618 253144 679624 253156
rect 675904 253116 679624 253144
rect 675904 253104 675910 253116
rect 679618 253104 679624 253116
rect 679676 253104 679682 253156
rect 35802 252696 35808 252748
rect 35860 252736 35866 252748
rect 41322 252736 41328 252748
rect 35860 252708 41328 252736
rect 35860 252696 35866 252708
rect 41322 252696 41328 252708
rect 41380 252696 41386 252748
rect 35618 252560 35624 252612
rect 35676 252600 35682 252612
rect 41690 252600 41696 252612
rect 35676 252572 41696 252600
rect 35676 252560 35682 252572
rect 41690 252560 41696 252572
rect 41748 252560 41754 252612
rect 42058 252560 42064 252612
rect 42116 252600 42122 252612
rect 42702 252600 42708 252612
rect 42116 252572 42708 252600
rect 42116 252560 42122 252572
rect 42702 252560 42708 252572
rect 42760 252560 42766 252612
rect 554406 252560 554412 252612
rect 554464 252600 554470 252612
rect 562318 252600 562324 252612
rect 554464 252572 562324 252600
rect 554464 252560 554470 252572
rect 562318 252560 562324 252572
rect 562376 252560 562382 252612
rect 35802 251200 35808 251252
rect 35860 251240 35866 251252
rect 37918 251240 37924 251252
rect 35860 251212 37924 251240
rect 35860 251200 35866 251212
rect 37918 251200 37924 251212
rect 37976 251200 37982 251252
rect 554130 251200 554136 251252
rect 554188 251240 554194 251252
rect 556798 251240 556804 251252
rect 554188 251212 556804 251240
rect 554188 251200 554194 251212
rect 556798 251200 556804 251212
rect 556856 251200 556862 251252
rect 35802 249908 35808 249960
rect 35860 249948 35866 249960
rect 40310 249948 40316 249960
rect 35860 249920 40316 249948
rect 35860 249908 35866 249920
rect 40310 249908 40316 249920
rect 40368 249908 40374 249960
rect 675386 249568 675392 249620
rect 675444 249568 675450 249620
rect 675404 248532 675432 249568
rect 675386 248480 675392 248532
rect 675444 248480 675450 248532
rect 559558 246304 559564 246356
rect 559616 246344 559622 246356
rect 647234 246344 647240 246356
rect 559616 246316 647240 246344
rect 559616 246304 559622 246316
rect 647234 246304 647240 246316
rect 647292 246304 647298 246356
rect 553854 245624 553860 245676
rect 553912 245664 553918 245676
rect 596818 245664 596824 245676
rect 553912 245636 596824 245664
rect 553912 245624 553918 245636
rect 596818 245624 596824 245636
rect 596876 245624 596882 245676
rect 553486 244264 553492 244316
rect 553544 244304 553550 244316
rect 555418 244304 555424 244316
rect 553544 244276 555424 244304
rect 553544 244264 553550 244276
rect 555418 244264 555424 244276
rect 555476 244264 555482 244316
rect 674650 243652 674656 243704
rect 674708 243692 674714 243704
rect 675202 243692 675208 243704
rect 674708 243664 675208 243692
rect 674708 243652 674714 243664
rect 675202 243652 675208 243664
rect 675260 243652 675266 243704
rect 674834 243176 674840 243228
rect 674892 243216 674898 243228
rect 674892 243188 675248 243216
rect 674892 243176 674898 243188
rect 675220 242956 675248 243188
rect 675202 242904 675208 242956
rect 675260 242904 675266 242956
rect 37918 242836 37924 242888
rect 37976 242876 37982 242888
rect 41690 242876 41696 242888
rect 37976 242848 41696 242876
rect 37976 242836 37982 242848
rect 41690 242836 41696 242848
rect 41748 242836 41754 242888
rect 576118 242156 576124 242208
rect 576176 242196 576182 242208
rect 648614 242196 648620 242208
rect 576176 242168 648620 242196
rect 576176 242156 576182 242168
rect 648614 242156 648620 242168
rect 648672 242156 648678 242208
rect 553670 241476 553676 241528
rect 553728 241516 553734 241528
rect 629938 241516 629944 241528
rect 553728 241488 629944 241516
rect 553728 241476 553734 241488
rect 629938 241476 629944 241488
rect 629996 241476 630002 241528
rect 554498 240116 554504 240168
rect 554556 240156 554562 240168
rect 577498 240156 577504 240168
rect 554556 240128 577504 240156
rect 554556 240116 554562 240128
rect 577498 240116 577504 240128
rect 577556 240116 577562 240168
rect 554314 238688 554320 238740
rect 554372 238728 554378 238740
rect 576118 238728 576124 238740
rect 554372 238700 576124 238728
rect 554372 238688 554378 238700
rect 576118 238688 576124 238700
rect 576176 238688 576182 238740
rect 672166 237056 672172 237108
rect 672224 237096 672230 237108
rect 672224 237068 672770 237096
rect 672224 237056 672230 237068
rect 553762 236784 553768 236836
rect 553820 236824 553826 236836
rect 559558 236824 559564 236836
rect 553820 236796 559564 236824
rect 553820 236784 553826 236796
rect 559558 236784 559564 236796
rect 559616 236784 559622 236836
rect 672874 236756 672902 236878
rect 672828 236728 672902 236756
rect 671154 236580 671160 236632
rect 671212 236620 671218 236632
rect 672828 236620 672856 236728
rect 672954 236700 673006 236706
rect 672954 236642 673006 236648
rect 671212 236592 672856 236620
rect 671212 236580 671218 236592
rect 671982 236444 671988 236496
rect 672040 236484 672046 236496
rect 672040 236456 673118 236484
rect 672040 236444 672046 236456
rect 673184 236292 673236 236298
rect 673184 236234 673236 236240
rect 672276 236116 673330 236144
rect 670970 235900 670976 235952
rect 671028 235940 671034 235952
rect 672276 235940 672304 236116
rect 671028 235912 672304 235940
rect 671028 235900 671034 235912
rect 672902 235900 672908 235952
rect 672960 235940 672966 235952
rect 672960 235912 673440 235940
rect 672960 235900 672966 235912
rect 672994 235696 673000 235748
rect 673052 235736 673058 235748
rect 673052 235708 673554 235736
rect 673052 235696 673058 235708
rect 673178 235492 673184 235544
rect 673236 235532 673242 235544
rect 673236 235504 673670 235532
rect 673236 235492 673242 235504
rect 671982 235288 671988 235340
rect 672040 235328 672046 235340
rect 672040 235300 673778 235328
rect 672040 235288 672046 235300
rect 673874 235136 673926 235142
rect 673874 235078 673926 235084
rect 669682 234812 669688 234864
rect 669740 234852 669746 234864
rect 673978 234852 674006 234906
rect 669740 234824 674006 234852
rect 669740 234812 669746 234824
rect 674100 234648 674128 234702
rect 673886 234620 674128 234648
rect 554406 234540 554412 234592
rect 554464 234580 554470 234592
rect 570598 234580 570604 234592
rect 554464 234552 570604 234580
rect 554464 234540 554470 234552
rect 570598 234540 570604 234552
rect 570656 234540 570662 234592
rect 672166 234472 672172 234524
rect 672224 234512 672230 234524
rect 673546 234512 673552 234524
rect 672224 234484 673552 234512
rect 672224 234472 672230 234484
rect 673546 234472 673552 234484
rect 673604 234472 673610 234524
rect 671338 234336 671344 234388
rect 671396 234376 671402 234388
rect 673886 234376 673914 234620
rect 671396 234348 673914 234376
rect 671396 234336 671402 234348
rect 670326 234132 670332 234184
rect 670384 234172 670390 234184
rect 674208 234172 674236 234498
rect 670384 234144 674236 234172
rect 670384 234132 670390 234144
rect 652202 233860 652208 233912
rect 652260 233900 652266 233912
rect 675478 233900 675484 233912
rect 652260 233872 675484 233900
rect 652260 233860 652266 233872
rect 675478 233860 675484 233872
rect 675536 233860 675542 233912
rect 675846 233860 675852 233912
rect 675904 233900 675910 233912
rect 678238 233900 678244 233912
rect 675904 233872 678244 233900
rect 675904 233860 675910 233872
rect 678238 233860 678244 233872
rect 678296 233860 678302 233912
rect 672994 233384 673000 233436
rect 673052 233384 673058 233436
rect 42334 233248 42340 233300
rect 42392 233288 42398 233300
rect 42702 233288 42708 233300
rect 42392 233260 42708 233288
rect 42392 233248 42398 233260
rect 42702 233248 42708 233260
rect 42760 233248 42766 233300
rect 670878 233180 670884 233232
rect 670936 233220 670942 233232
rect 673012 233220 673040 233384
rect 670936 233192 673040 233220
rect 670936 233180 670942 233192
rect 670050 232840 670056 232892
rect 670108 232880 670114 232892
rect 671982 232880 671988 232892
rect 670108 232852 671988 232880
rect 670108 232840 670114 232852
rect 671982 232840 671988 232852
rect 672040 232840 672046 232892
rect 663058 232636 663064 232688
rect 663116 232676 663122 232688
rect 675478 232676 675484 232688
rect 663116 232648 675484 232676
rect 663116 232636 663122 232648
rect 675478 232636 675484 232648
rect 675536 232636 675542 232688
rect 675846 232636 675852 232688
rect 675904 232676 675910 232688
rect 683114 232676 683120 232688
rect 675904 232648 683120 232676
rect 675904 232636 675910 232648
rect 683114 232636 683120 232648
rect 683172 232636 683178 232688
rect 660298 232500 660304 232552
rect 660356 232540 660362 232552
rect 675478 232540 675484 232552
rect 660356 232512 675484 232540
rect 660356 232500 660362 232512
rect 675478 232500 675484 232512
rect 675536 232500 675542 232552
rect 675846 232500 675852 232552
rect 675904 232540 675910 232552
rect 683298 232540 683304 232552
rect 675904 232512 683304 232540
rect 675904 232500 675910 232512
rect 683298 232500 683304 232512
rect 683356 232500 683362 232552
rect 155126 231752 155132 231804
rect 155184 231792 155190 231804
rect 156966 231792 156972 231804
rect 155184 231764 156972 231792
rect 155184 231752 155190 231764
rect 156966 231752 156972 231764
rect 157024 231752 157030 231804
rect 134886 231616 134892 231668
rect 134944 231656 134950 231668
rect 142062 231656 142068 231668
rect 134944 231628 142068 231656
rect 134944 231616 134950 231628
rect 142062 231616 142068 231628
rect 142120 231616 142126 231668
rect 155494 231616 155500 231668
rect 155552 231656 155558 231668
rect 162670 231656 162676 231668
rect 155552 231628 162676 231656
rect 155552 231616 155558 231628
rect 162670 231616 162676 231628
rect 162728 231616 162734 231668
rect 92382 231480 92388 231532
rect 92440 231520 92446 231532
rect 170766 231520 170772 231532
rect 92440 231492 170772 231520
rect 92440 231480 92446 231492
rect 170766 231480 170772 231492
rect 170824 231480 170830 231532
rect 662506 231480 662512 231532
rect 662564 231520 662570 231532
rect 668578 231520 668584 231532
rect 662564 231492 668584 231520
rect 662564 231480 662570 231492
rect 668578 231480 668584 231492
rect 668636 231480 668642 231532
rect 128262 231344 128268 231396
rect 128320 231384 128326 231396
rect 195882 231384 195888 231396
rect 128320 231356 195888 231384
rect 128320 231344 128326 231356
rect 195882 231344 195888 231356
rect 195940 231344 195946 231396
rect 674834 231316 674840 231328
rect 668596 231288 674840 231316
rect 64322 231208 64328 231260
rect 64380 231248 64386 231260
rect 668026 231248 668032 231260
rect 64380 231220 668032 231248
rect 64380 231208 64386 231220
rect 668026 231208 668032 231220
rect 668084 231208 668090 231260
rect 57238 231072 57244 231124
rect 57296 231112 57302 231124
rect 668596 231112 668624 231288
rect 674834 231276 674840 231288
rect 674892 231276 674898 231328
rect 57296 231084 668624 231112
rect 668688 231152 675326 231180
rect 57296 231072 57302 231084
rect 665082 230936 665088 230988
rect 665140 230976 665146 230988
rect 668688 230976 668716 231152
rect 665140 230948 668716 230976
rect 665140 230936 665146 230948
rect 672166 230936 672172 230988
rect 672224 230976 672230 230988
rect 672224 230948 675142 230976
rect 672224 230936 672230 230948
rect 94498 230868 94504 230920
rect 94556 230908 94562 230920
rect 171410 230908 171416 230920
rect 94556 230880 171416 230908
rect 94556 230868 94562 230880
rect 171410 230868 171416 230880
rect 171468 230868 171474 230920
rect 668578 230800 668584 230852
rect 668636 230840 668642 230852
rect 668636 230812 674880 230840
rect 668636 230800 668642 230812
rect 104802 230732 104808 230784
rect 104860 230772 104866 230784
rect 179138 230772 179144 230784
rect 104860 230744 179144 230772
rect 104860 230732 104866 230744
rect 179138 230732 179144 230744
rect 179196 230732 179202 230784
rect 674852 230772 674880 230812
rect 674852 230744 674982 230772
rect 118602 230596 118608 230648
rect 118660 230636 118666 230648
rect 188154 230636 188160 230648
rect 118660 230608 188160 230636
rect 118660 230596 118666 230608
rect 188154 230596 188160 230608
rect 188212 230596 188218 230648
rect 665266 230596 665272 230648
rect 665324 230636 665330 230648
rect 665324 230608 674820 230636
rect 665324 230596 665330 230608
rect 439314 230528 439320 230580
rect 439372 230568 439378 230580
rect 439372 230540 439544 230568
rect 439372 230528 439378 230540
rect 142154 230460 142160 230512
rect 142212 230500 142218 230512
rect 201034 230500 201040 230512
rect 142212 230472 201040 230500
rect 142212 230460 142218 230472
rect 201034 230460 201040 230472
rect 201092 230460 201098 230512
rect 42334 230392 42340 230444
rect 42392 230432 42398 230444
rect 43070 230432 43076 230444
rect 42392 230404 43076 230432
rect 42392 230392 42398 230404
rect 43070 230392 43076 230404
rect 43128 230392 43134 230444
rect 126882 230392 126888 230444
rect 126940 230432 126946 230444
rect 141970 230432 141976 230444
rect 126940 230404 141976 230432
rect 126940 230392 126946 230404
rect 141970 230392 141976 230404
rect 142028 230392 142034 230444
rect 213086 230392 213092 230444
rect 213144 230432 213150 230444
rect 261570 230432 261576 230444
rect 213144 230404 261576 230432
rect 213144 230392 213150 230404
rect 261570 230392 261576 230404
rect 261628 230392 261634 230444
rect 311986 230392 311992 230444
rect 312044 230432 312050 230444
rect 313090 230432 313096 230444
rect 312044 230404 313096 230432
rect 312044 230392 312050 230404
rect 313090 230392 313096 230404
rect 313148 230392 313154 230444
rect 374638 230392 374644 230444
rect 374696 230432 374702 230444
rect 376202 230432 376208 230444
rect 374696 230404 376208 230432
rect 374696 230392 374702 230404
rect 376202 230392 376208 230404
rect 376260 230392 376266 230444
rect 439516 230432 439544 230540
rect 674676 230444 674728 230450
rect 440694 230432 440700 230444
rect 439516 230404 440700 230432
rect 440694 230392 440700 230404
rect 440752 230392 440758 230444
rect 441890 230392 441896 230444
rect 441948 230432 441954 230444
rect 443454 230432 443460 230444
rect 441948 230404 443460 230432
rect 441948 230392 441954 230404
rect 443454 230392 443460 230404
rect 443512 230392 443518 230444
rect 444466 230392 444472 230444
rect 444524 230432 444530 230444
rect 447594 230432 447600 230444
rect 444524 230404 447600 230432
rect 444524 230392 444530 230404
rect 447594 230392 447600 230404
rect 447652 230392 447658 230444
rect 451550 230392 451556 230444
rect 451608 230432 451614 230444
rect 453298 230432 453304 230444
rect 451608 230404 453304 230432
rect 451608 230392 451614 230404
rect 453298 230392 453304 230404
rect 453356 230392 453362 230444
rect 476114 230392 476120 230444
rect 476172 230432 476178 230444
rect 478598 230432 478604 230444
rect 476172 230404 478604 230432
rect 476172 230392 476178 230404
rect 478598 230392 478604 230404
rect 478656 230392 478662 230444
rect 539594 230432 539600 230444
rect 532528 230404 539600 230432
rect 387426 230324 387432 230376
rect 387484 230364 387490 230376
rect 388438 230364 388444 230376
rect 387484 230336 388444 230364
rect 387484 230324 387490 230336
rect 388438 230324 388444 230336
rect 388496 230324 388502 230376
rect 398098 230324 398104 230376
rect 398156 230364 398162 230376
rect 399386 230364 399392 230376
rect 398156 230336 399392 230364
rect 398156 230324 398162 230336
rect 399386 230324 399392 230336
rect 399444 230324 399450 230376
rect 438670 230324 438676 230376
rect 438728 230364 438734 230376
rect 439314 230364 439320 230376
rect 438728 230336 439320 230364
rect 438728 230324 438734 230336
rect 439314 230324 439320 230336
rect 439372 230324 439378 230376
rect 455414 230324 455420 230376
rect 455472 230364 455478 230376
rect 457162 230364 457168 230376
rect 455472 230336 457168 230364
rect 455472 230324 455478 230336
rect 457162 230324 457168 230336
rect 457220 230324 457226 230376
rect 470870 230324 470876 230376
rect 470928 230364 470934 230376
rect 471882 230364 471888 230376
rect 470928 230336 471888 230364
rect 470928 230324 470934 230336
rect 471882 230324 471888 230336
rect 471940 230324 471946 230376
rect 493410 230324 493416 230376
rect 493468 230364 493474 230376
rect 496354 230364 496360 230376
rect 493468 230336 496360 230364
rect 493468 230324 493474 230336
rect 496354 230324 496360 230336
rect 496412 230324 496418 230376
rect 497274 230324 497280 230376
rect 497332 230364 497338 230376
rect 498102 230364 498108 230376
rect 497332 230336 498108 230364
rect 497332 230324 497338 230336
rect 498102 230324 498108 230336
rect 498160 230324 498166 230376
rect 510798 230324 510804 230376
rect 510856 230364 510862 230376
rect 511902 230364 511908 230376
rect 510856 230336 511908 230364
rect 510856 230324 510862 230336
rect 511902 230324 511908 230336
rect 511960 230324 511966 230376
rect 521102 230324 521108 230376
rect 521160 230364 521166 230376
rect 526438 230364 526444 230376
rect 521160 230336 526444 230364
rect 521160 230324 521166 230336
rect 526438 230324 526444 230336
rect 526496 230324 526502 230376
rect 530118 230324 530124 230376
rect 530176 230364 530182 230376
rect 531130 230364 531136 230376
rect 530176 230336 531136 230364
rect 530176 230324 530182 230336
rect 531130 230324 531136 230336
rect 531188 230324 531194 230376
rect 133782 230256 133788 230308
rect 133840 230296 133846 230308
rect 202322 230296 202328 230308
rect 133840 230268 202328 230296
rect 133840 230256 133846 230268
rect 202322 230256 202328 230268
rect 202380 230256 202386 230308
rect 206278 230256 206284 230308
rect 206336 230296 206342 230308
rect 256418 230296 256424 230308
rect 206336 230268 256424 230296
rect 206336 230256 206342 230268
rect 256418 230256 256424 230268
rect 256476 230256 256482 230308
rect 256602 230256 256608 230308
rect 256660 230296 256666 230308
rect 297634 230296 297640 230308
rect 256660 230268 297640 230296
rect 256660 230256 256666 230268
rect 297634 230256 297640 230268
rect 297692 230256 297698 230308
rect 297818 230256 297824 230308
rect 297876 230296 297882 230308
rect 323394 230296 323400 230308
rect 297876 230268 323400 230296
rect 297876 230256 297882 230268
rect 323394 230256 323400 230268
rect 323452 230256 323458 230308
rect 443822 230188 443828 230240
rect 443880 230228 443886 230240
rect 444650 230228 444656 230240
rect 443880 230200 444656 230228
rect 443880 230188 443886 230200
rect 444650 230188 444656 230200
rect 444708 230188 444714 230240
rect 452838 230188 452844 230240
rect 452896 230228 452902 230240
rect 454310 230228 454316 230240
rect 452896 230200 454316 230228
rect 452896 230188 452902 230200
rect 454310 230188 454316 230200
rect 454368 230188 454374 230240
rect 468294 230188 468300 230240
rect 468352 230228 468358 230240
rect 469122 230228 469128 230240
rect 468352 230200 469128 230228
rect 468352 230188 468358 230200
rect 469122 230188 469128 230200
rect 469180 230188 469186 230240
rect 487614 230188 487620 230240
rect 487672 230228 487678 230240
rect 488442 230228 488448 230240
rect 487672 230200 488448 230228
rect 487672 230188 487678 230200
rect 488442 230188 488448 230200
rect 488500 230188 488506 230240
rect 495158 230228 495164 230240
rect 489886 230200 495164 230228
rect 95234 230120 95240 230172
rect 95292 230160 95298 230172
rect 95292 230132 157334 230160
rect 95292 230120 95298 230132
rect 86218 229984 86224 230036
rect 86276 230024 86282 230036
rect 157150 230024 157156 230036
rect 86276 229996 157156 230024
rect 86276 229984 86282 229996
rect 157150 229984 157156 229996
rect 157208 229984 157214 230036
rect 157306 230024 157334 230132
rect 157426 230120 157432 230172
rect 157484 230160 157490 230172
rect 161106 230160 161112 230172
rect 157484 230132 161112 230160
rect 157484 230120 157490 230132
rect 161106 230120 161112 230132
rect 161164 230120 161170 230172
rect 161290 230120 161296 230172
rect 161348 230160 161354 230172
rect 166258 230160 166264 230172
rect 161348 230132 166264 230160
rect 161348 230120 161354 230132
rect 166258 230120 166264 230132
rect 166316 230120 166322 230172
rect 176470 230120 176476 230172
rect 176528 230160 176534 230172
rect 235810 230160 235816 230172
rect 176528 230132 235816 230160
rect 176528 230120 176534 230132
rect 235810 230120 235816 230132
rect 235868 230120 235874 230172
rect 240318 230120 240324 230172
rect 240376 230160 240382 230172
rect 282178 230160 282184 230172
rect 240376 230132 282184 230160
rect 240376 230120 240382 230132
rect 282178 230120 282184 230132
rect 282236 230120 282242 230172
rect 282638 230120 282644 230172
rect 282696 230160 282702 230172
rect 307938 230160 307944 230172
rect 282696 230132 307944 230160
rect 282696 230120 282702 230132
rect 307938 230120 307944 230132
rect 307996 230120 308002 230172
rect 308122 230120 308128 230172
rect 308180 230160 308186 230172
rect 334986 230160 334992 230172
rect 308180 230132 334992 230160
rect 308180 230120 308186 230132
rect 334986 230120 334992 230132
rect 335044 230120 335050 230172
rect 335170 230120 335176 230172
rect 335228 230160 335234 230172
rect 350442 230160 350448 230172
rect 335228 230132 350448 230160
rect 335228 230120 335234 230132
rect 350442 230120 350448 230132
rect 350500 230120 350506 230172
rect 454126 230052 454132 230104
rect 454184 230092 454190 230104
rect 455322 230092 455328 230104
rect 454184 230064 455328 230092
rect 454184 230052 454190 230064
rect 455322 230052 455328 230064
rect 455380 230052 455386 230104
rect 157794 230024 157800 230036
rect 157306 229996 157800 230024
rect 157794 229984 157800 229996
rect 157852 229984 157858 230036
rect 157978 229984 157984 230036
rect 158036 230024 158042 230036
rect 163682 230024 163688 230036
rect 158036 229996 163688 230024
rect 158036 229984 158042 229996
rect 163682 229984 163688 229996
rect 163740 229984 163746 230036
rect 170950 229984 170956 230036
rect 171008 230024 171014 230036
rect 230658 230024 230664 230036
rect 171008 229996 230664 230024
rect 171008 229984 171014 229996
rect 230658 229984 230664 229996
rect 230716 229984 230722 230036
rect 277026 230024 277032 230036
rect 230860 229996 277032 230024
rect 130378 229848 130384 229900
rect 130436 229888 130442 229900
rect 130436 229860 142384 229888
rect 130436 229848 130442 229860
rect 68278 229712 68284 229764
rect 68336 229752 68342 229764
rect 142154 229752 142160 229764
rect 68336 229724 142160 229752
rect 68336 229712 68342 229724
rect 142154 229712 142160 229724
rect 142212 229712 142218 229764
rect 142356 229752 142384 229860
rect 142614 229848 142620 229900
rect 142672 229888 142678 229900
rect 195054 229888 195060 229900
rect 142672 229860 195060 229888
rect 142672 229848 142678 229860
rect 195054 229848 195060 229860
rect 195112 229848 195118 229900
rect 195422 229848 195428 229900
rect 195480 229888 195486 229900
rect 195480 229860 229094 229888
rect 195480 229848 195486 229860
rect 145006 229752 145012 229764
rect 142356 229724 145012 229752
rect 145006 229712 145012 229724
rect 145064 229712 145070 229764
rect 146938 229712 146944 229764
rect 146996 229752 147002 229764
rect 146996 229724 147996 229752
rect 146996 229712 147002 229724
rect 82078 229576 82084 229628
rect 82136 229616 82142 229628
rect 147766 229616 147772 229628
rect 82136 229588 147772 229616
rect 82136 229576 82142 229588
rect 147766 229576 147772 229588
rect 147824 229576 147830 229628
rect 147968 229616 147996 229724
rect 148134 229712 148140 229764
rect 148192 229752 148198 229764
rect 155954 229752 155960 229764
rect 148192 229724 155960 229752
rect 148192 229712 148198 229724
rect 155954 229712 155960 229724
rect 156012 229712 156018 229764
rect 156322 229712 156328 229764
rect 156380 229752 156386 229764
rect 157288 229752 157294 229764
rect 156380 229724 157294 229752
rect 156380 229712 156386 229724
rect 157288 229712 157294 229724
rect 157346 229712 157352 229764
rect 157426 229712 157432 229764
rect 157484 229752 157490 229764
rect 162578 229752 162584 229764
rect 157484 229724 162584 229752
rect 157484 229712 157490 229724
rect 162578 229712 162584 229724
rect 162636 229712 162642 229764
rect 164050 229712 164056 229764
rect 164108 229752 164114 229764
rect 225506 229752 225512 229764
rect 164108 229724 225512 229752
rect 164108 229712 164114 229724
rect 225506 229712 225512 229724
rect 225564 229712 225570 229764
rect 229066 229752 229094 229860
rect 230474 229848 230480 229900
rect 230532 229888 230538 229900
rect 230860 229888 230888 229996
rect 277026 229984 277032 229996
rect 277084 229984 277090 230036
rect 277210 229984 277216 230036
rect 277268 230024 277274 230036
rect 302786 230024 302792 230036
rect 277268 229996 302792 230024
rect 277268 229984 277274 229996
rect 302786 229984 302792 229996
rect 302844 229984 302850 230036
rect 303246 229984 303252 230036
rect 303304 230024 303310 230036
rect 329834 230024 329840 230036
rect 303304 229996 329840 230024
rect 303304 229984 303310 229996
rect 329834 229984 329840 229996
rect 329892 229984 329898 230036
rect 330938 229984 330944 230036
rect 330996 230024 331002 230036
rect 355594 230024 355600 230036
rect 330996 229996 355600 230024
rect 330996 229984 331002 229996
rect 355594 229984 355600 229996
rect 355652 229984 355658 230036
rect 476666 229984 476672 230036
rect 476724 230024 476730 230036
rect 481634 230024 481640 230036
rect 476724 229996 481640 230024
rect 476724 229984 476730 229996
rect 481634 229984 481640 229996
rect 481692 229984 481698 230036
rect 484394 229984 484400 230036
rect 484452 230024 484458 230036
rect 489886 230024 489914 230200
rect 495158 230188 495164 230200
rect 495216 230188 495222 230240
rect 511442 230188 511448 230240
rect 511500 230228 511506 230240
rect 517514 230228 517520 230240
rect 511500 230200 517520 230228
rect 511500 230188 511506 230200
rect 517514 230188 517520 230200
rect 517572 230188 517578 230240
rect 530762 230188 530768 230240
rect 530820 230228 530826 230240
rect 532528 230228 532556 230404
rect 539594 230392 539600 230404
rect 539652 230392 539658 230444
rect 674676 230386 674728 230392
rect 533522 230256 533528 230308
rect 533580 230296 533586 230308
rect 538306 230296 538312 230308
rect 533580 230268 538312 230296
rect 533580 230256 533586 230268
rect 538306 230256 538312 230268
rect 538364 230256 538370 230308
rect 530820 230200 532556 230228
rect 530820 230188 530826 230200
rect 673086 230188 673092 230240
rect 673144 230228 673150 230240
rect 673144 230200 674590 230228
rect 673144 230188 673150 230200
rect 532694 230120 532700 230172
rect 532752 230160 532758 230172
rect 547138 230160 547144 230172
rect 532752 230132 547144 230160
rect 532752 230120 532758 230132
rect 547138 230120 547144 230132
rect 547196 230120 547202 230172
rect 491478 230052 491484 230104
rect 491536 230092 491542 230104
rect 492490 230092 492496 230104
rect 491536 230064 492496 230092
rect 491536 230052 491542 230064
rect 492490 230052 492496 230064
rect 492548 230052 492554 230104
rect 560938 230052 560944 230104
rect 560996 230092 561002 230104
rect 568114 230092 568120 230104
rect 560996 230064 568120 230092
rect 560996 230052 561002 230064
rect 568114 230052 568120 230064
rect 568172 230052 568178 230104
rect 484452 229996 489914 230024
rect 484452 229984 484458 229996
rect 517238 229984 517244 230036
rect 517296 230024 517302 230036
rect 524598 230024 524604 230036
rect 517296 229996 524604 230024
rect 517296 229984 517302 229996
rect 524598 229984 524604 229996
rect 524656 229984 524662 230036
rect 528830 229984 528836 230036
rect 528888 230024 528894 230036
rect 533522 230024 533528 230036
rect 528888 229996 533528 230024
rect 528888 229984 528894 229996
rect 533522 229984 533528 229996
rect 533580 229984 533586 230036
rect 534626 229984 534632 230036
rect 534684 230024 534690 230036
rect 549254 230024 549260 230036
rect 534684 229996 549260 230024
rect 534684 229984 534690 229996
rect 549254 229984 549260 229996
rect 549312 229984 549318 230036
rect 673270 229984 673276 230036
rect 673328 230024 673334 230036
rect 673328 229996 674478 230024
rect 673328 229984 673334 229996
rect 453482 229916 453488 229968
rect 453540 229956 453546 229968
rect 455782 229956 455788 229968
rect 453540 229928 455788 229956
rect 453540 229916 453546 229928
rect 455782 229916 455788 229928
rect 455840 229916 455846 229968
rect 230532 229860 230888 229888
rect 230532 229848 230538 229860
rect 233694 229848 233700 229900
rect 233752 229888 233758 229900
rect 271874 229888 271880 229900
rect 233752 229860 271880 229888
rect 233752 229848 233758 229860
rect 271874 229848 271880 229860
rect 271932 229848 271938 229900
rect 275646 229848 275652 229900
rect 275704 229888 275710 229900
rect 311986 229888 311992 229900
rect 275704 229860 311992 229888
rect 275704 229848 275710 229860
rect 311986 229848 311992 229860
rect 312044 229848 312050 229900
rect 312630 229848 312636 229900
rect 312688 229888 312694 229900
rect 340138 229888 340144 229900
rect 312688 229860 340144 229888
rect 312688 229848 312694 229860
rect 340138 229848 340144 229860
rect 340196 229848 340202 229900
rect 345658 229848 345664 229900
rect 345716 229888 345722 229900
rect 360746 229888 360752 229900
rect 345716 229860 360752 229888
rect 345716 229848 345722 229860
rect 360746 229848 360752 229860
rect 360804 229848 360810 229900
rect 361206 229848 361212 229900
rect 361264 229888 361270 229900
rect 378778 229888 378784 229900
rect 361264 229860 378784 229888
rect 361264 229848 361270 229860
rect 378778 229848 378784 229860
rect 378836 229848 378842 229900
rect 410886 229848 410892 229900
rect 410944 229888 410950 229900
rect 417418 229888 417424 229900
rect 410944 229860 417424 229888
rect 410944 229848 410950 229860
rect 417418 229848 417424 229860
rect 417476 229848 417482 229900
rect 449618 229848 449624 229900
rect 449676 229888 449682 229900
rect 450538 229888 450544 229900
rect 449676 229860 450544 229888
rect 449676 229848 449682 229860
rect 450538 229848 450544 229860
rect 450596 229848 450602 229900
rect 457346 229848 457352 229900
rect 457404 229888 457410 229900
rect 464062 229888 464068 229900
rect 457404 229860 464068 229888
rect 457404 229848 457410 229860
rect 464062 229848 464068 229860
rect 464120 229848 464126 229900
rect 469582 229848 469588 229900
rect 469640 229888 469646 229900
rect 476758 229888 476764 229900
rect 469640 229860 476764 229888
rect 469640 229848 469646 229860
rect 476758 229848 476764 229860
rect 476816 229848 476822 229900
rect 481818 229848 481824 229900
rect 481876 229888 481882 229900
rect 493686 229888 493692 229900
rect 481876 229860 493692 229888
rect 481876 229848 481882 229860
rect 493686 229848 493692 229860
rect 493744 229848 493750 229900
rect 495986 229848 495992 229900
rect 496044 229888 496050 229900
rect 506382 229888 506388 229900
rect 496044 229860 506388 229888
rect 496044 229848 496050 229860
rect 506382 229848 506388 229860
rect 506440 229848 506446 229900
rect 507578 229848 507584 229900
rect 507636 229888 507642 229900
rect 516778 229888 516784 229900
rect 507636 229860 516784 229888
rect 507636 229848 507642 229860
rect 516778 229848 516784 229860
rect 516836 229848 516842 229900
rect 519170 229848 519176 229900
rect 519228 229888 519234 229900
rect 528554 229888 528560 229900
rect 519228 229860 528560 229888
rect 519228 229848 519234 229860
rect 528554 229848 528560 229860
rect 528612 229848 528618 229900
rect 536558 229848 536564 229900
rect 536616 229888 536622 229900
rect 559558 229888 559564 229900
rect 536616 229860 559564 229888
rect 536616 229848 536622 229860
rect 559558 229848 559564 229860
rect 559616 229848 559622 229900
rect 433518 229780 433524 229832
rect 433576 229820 433582 229832
rect 434162 229820 434168 229832
rect 433576 229792 434168 229820
rect 433576 229780 433582 229792
rect 434162 229780 434168 229792
rect 434220 229780 434226 229832
rect 673868 229780 673874 229832
rect 673926 229820 673932 229832
rect 673926 229792 674360 229820
rect 673926 229780 673932 229792
rect 246114 229752 246120 229764
rect 229066 229724 246120 229752
rect 246114 229712 246120 229724
rect 246172 229712 246178 229764
rect 246482 229712 246488 229764
rect 246540 229752 246546 229764
rect 287330 229752 287336 229764
rect 246540 229724 287336 229752
rect 246540 229712 246546 229724
rect 287330 229712 287336 229724
rect 287388 229712 287394 229764
rect 287698 229712 287704 229764
rect 287756 229752 287762 229764
rect 318242 229752 318248 229764
rect 287756 229724 318248 229752
rect 287756 229712 287762 229724
rect 318242 229712 318248 229724
rect 318300 229712 318306 229764
rect 345290 229752 345296 229764
rect 325666 229724 345296 229752
rect 153378 229616 153384 229628
rect 147968 229588 153384 229616
rect 153378 229576 153384 229588
rect 153436 229576 153442 229628
rect 153838 229576 153844 229628
rect 153896 229616 153902 229628
rect 158530 229616 158536 229628
rect 153896 229588 158536 229616
rect 153896 229576 153902 229588
rect 158530 229576 158536 229588
rect 158588 229576 158594 229628
rect 158714 229576 158720 229628
rect 158772 229616 158778 229628
rect 161750 229616 161756 229628
rect 158772 229588 161756 229616
rect 158772 229576 158778 229588
rect 161750 229576 161756 229588
rect 161808 229576 161814 229628
rect 161934 229576 161940 229628
rect 161992 229616 161998 229628
rect 220354 229616 220360 229628
rect 161992 229588 220360 229616
rect 161992 229576 161998 229588
rect 220354 229576 220360 229588
rect 220412 229576 220418 229628
rect 251266 229616 251272 229628
rect 224926 229588 251272 229616
rect 102134 229440 102140 229492
rect 102192 229480 102198 229492
rect 145650 229480 145656 229492
rect 102192 229452 145656 229480
rect 102192 229440 102198 229452
rect 145650 229440 145656 229452
rect 145708 229440 145714 229492
rect 145834 229440 145840 229492
rect 145892 229480 145898 229492
rect 210050 229480 210056 229492
rect 145892 229452 210056 229480
rect 145892 229440 145898 229452
rect 210050 229440 210056 229452
rect 210108 229440 210114 229492
rect 220262 229440 220268 229492
rect 220320 229480 220326 229492
rect 224926 229480 224954 229588
rect 251266 229576 251272 229588
rect 251324 229576 251330 229628
rect 251726 229576 251732 229628
rect 251784 229616 251790 229628
rect 292482 229616 292488 229628
rect 251784 229588 292488 229616
rect 251784 229576 251790 229588
rect 292482 229576 292488 229588
rect 292540 229576 292546 229628
rect 318058 229576 318064 229628
rect 318116 229616 318122 229628
rect 325666 229616 325694 229724
rect 345290 229712 345296 229724
rect 345348 229712 345354 229764
rect 351730 229712 351736 229764
rect 351788 229752 351794 229764
rect 371050 229752 371056 229764
rect 351788 229724 371056 229752
rect 351788 229712 351794 229724
rect 371050 229712 371056 229724
rect 371108 229712 371114 229764
rect 377674 229712 377680 229764
rect 377732 229752 377738 229764
rect 389082 229752 389088 229764
rect 377732 229724 389088 229752
rect 377732 229712 377738 229724
rect 389082 229712 389088 229724
rect 389140 229712 389146 229764
rect 399846 229712 399852 229764
rect 399904 229752 399910 229764
rect 409690 229752 409696 229764
rect 399904 229724 409696 229752
rect 399904 229712 399910 229724
rect 409690 229712 409696 229724
rect 409748 229712 409754 229764
rect 467006 229712 467012 229764
rect 467064 229752 467070 229764
rect 473998 229752 474004 229764
rect 467064 229724 474004 229752
rect 467064 229712 467070 229724
rect 473998 229712 474004 229724
rect 474056 229712 474062 229764
rect 479242 229712 479248 229764
rect 479300 229752 479306 229764
rect 489914 229752 489920 229764
rect 479300 229724 489920 229752
rect 479300 229712 479306 229724
rect 489914 229712 489920 229724
rect 489972 229712 489978 229764
rect 492122 229712 492128 229764
rect 492180 229752 492186 229764
rect 507118 229752 507124 229764
rect 492180 229724 507124 229752
rect 492180 229712 492186 229724
rect 507118 229712 507124 229724
rect 507176 229712 507182 229764
rect 523034 229712 523040 229764
rect 523092 229752 523098 229764
rect 534718 229752 534724 229764
rect 523092 229724 534724 229752
rect 523092 229712 523098 229724
rect 534718 229712 534724 229724
rect 534776 229712 534782 229764
rect 538490 229712 538496 229764
rect 538548 229752 538554 229764
rect 566826 229752 566832 229764
rect 538548 229724 566832 229752
rect 538548 229712 538554 229724
rect 566826 229712 566832 229724
rect 566884 229712 566890 229764
rect 662322 229712 662328 229764
rect 662380 229752 662386 229764
rect 672166 229752 672172 229764
rect 662380 229724 672172 229752
rect 662380 229712 662386 229724
rect 672166 229712 672172 229724
rect 672224 229712 672230 229764
rect 509510 229644 509516 229696
rect 509568 229684 509574 229696
rect 515490 229684 515496 229696
rect 509568 229656 515496 229684
rect 509568 229644 509574 229656
rect 515490 229644 515496 229656
rect 515548 229644 515554 229696
rect 318116 229588 325694 229616
rect 318116 229576 318122 229588
rect 388622 229576 388628 229628
rect 388680 229616 388686 229628
rect 398742 229616 398748 229628
rect 388680 229588 398748 229616
rect 388680 229576 388686 229588
rect 398742 229576 398748 229588
rect 398800 229576 398806 229628
rect 463786 229576 463792 229628
rect 463844 229616 463850 229628
rect 465718 229616 465724 229628
rect 463844 229588 465724 229616
rect 463844 229576 463850 229588
rect 465718 229576 465724 229588
rect 465776 229576 465782 229628
rect 526898 229576 526904 229628
rect 526956 229616 526962 229628
rect 536098 229616 536104 229628
rect 526956 229588 536104 229616
rect 526956 229576 526962 229588
rect 536098 229576 536104 229588
rect 536156 229576 536162 229628
rect 660942 229576 660948 229628
rect 661000 229616 661006 229628
rect 662506 229616 662512 229628
rect 661000 229588 662512 229616
rect 661000 229576 661006 229588
rect 662506 229576 662512 229588
rect 662564 229576 662570 229628
rect 672902 229576 672908 229628
rect 672960 229616 672966 229628
rect 672960 229588 674268 229616
rect 672960 229576 672966 229588
rect 448974 229508 448980 229560
rect 449032 229548 449038 229560
rect 451366 229548 451372 229560
rect 449032 229520 451372 229548
rect 449032 229508 449038 229520
rect 451366 229508 451372 229520
rect 451424 229508 451430 229560
rect 220320 229452 224954 229480
rect 220320 229440 220326 229452
rect 225598 229440 225604 229492
rect 225656 229480 225662 229492
rect 233694 229480 233700 229492
rect 225656 229452 233700 229480
rect 225656 229440 225662 229452
rect 233694 229440 233700 229452
rect 233752 229440 233758 229492
rect 465442 229440 465448 229492
rect 465500 229480 465506 229492
rect 467466 229480 467472 229492
rect 465500 229452 467472 229480
rect 465500 229440 465506 229452
rect 467466 229440 467472 229452
rect 467524 229440 467530 229492
rect 446398 229372 446404 229424
rect 446456 229412 446462 229424
rect 448974 229412 448980 229424
rect 446456 229384 448980 229412
rect 446456 229372 446462 229384
rect 448974 229372 448980 229384
rect 449032 229372 449038 229424
rect 450906 229372 450912 229424
rect 450964 229412 450970 229424
rect 452654 229412 452660 229424
rect 450964 229384 452660 229412
rect 450964 229372 450970 229384
rect 452654 229372 452660 229384
rect 452712 229372 452718 229424
rect 673454 229372 673460 229424
rect 673512 229412 673518 229424
rect 673512 229384 674130 229412
rect 673512 229372 673518 229384
rect 110138 229304 110144 229356
rect 110196 229344 110202 229356
rect 144638 229344 144644 229356
rect 110196 229316 144644 229344
rect 110196 229304 110202 229316
rect 144638 229304 144644 229316
rect 144696 229304 144702 229356
rect 144822 229304 144828 229356
rect 144880 229344 144886 229356
rect 151446 229344 151452 229356
rect 144880 229316 151452 229344
rect 144880 229304 144886 229316
rect 151446 229304 151452 229316
rect 151504 229304 151510 229356
rect 151630 229304 151636 229356
rect 151688 229344 151694 229356
rect 151688 229316 154252 229344
rect 151688 229304 151694 229316
rect 123478 229168 123484 229220
rect 123536 229208 123542 229220
rect 146938 229208 146944 229220
rect 123536 229180 146944 229208
rect 123536 229168 123542 229180
rect 146938 229168 146944 229180
rect 146996 229168 147002 229220
rect 148318 229168 148324 229220
rect 148376 229208 148382 229220
rect 154022 229208 154028 229220
rect 148376 229180 154028 229208
rect 148376 229168 148382 229180
rect 154022 229168 154028 229180
rect 154080 229168 154086 229220
rect 154224 229208 154252 229316
rect 154390 229304 154396 229356
rect 154448 229344 154454 229356
rect 157150 229344 157156 229356
rect 154448 229316 157156 229344
rect 154448 229304 154454 229316
rect 157150 229304 157156 229316
rect 157208 229304 157214 229356
rect 157334 229304 157340 229356
rect 157392 229344 157398 229356
rect 215202 229344 215208 229356
rect 157392 229316 215208 229344
rect 157392 229304 157398 229316
rect 215202 229304 215208 229316
rect 215260 229304 215266 229356
rect 413830 229304 413836 229356
rect 413888 229344 413894 229356
rect 419994 229344 420000 229356
rect 413888 229316 420000 229344
rect 413888 229304 413894 229316
rect 419994 229304 420000 229316
rect 420052 229304 420058 229356
rect 472158 229304 472164 229356
rect 472216 229344 472222 229356
rect 472986 229344 472992 229356
rect 472216 229316 472992 229344
rect 472216 229304 472222 229316
rect 472986 229304 472992 229316
rect 473044 229304 473050 229356
rect 450262 229236 450268 229288
rect 450320 229276 450326 229288
rect 451734 229276 451740 229288
rect 450320 229248 451740 229276
rect 450320 229236 450326 229248
rect 451734 229236 451740 229248
rect 451792 229236 451798 229288
rect 495342 229236 495348 229288
rect 495400 229276 495406 229288
rect 500218 229276 500224 229288
rect 495400 229248 500224 229276
rect 495400 229236 495406 229248
rect 500218 229236 500224 229248
rect 500276 229236 500282 229288
rect 505646 229236 505652 229288
rect 505704 229276 505710 229288
rect 510614 229276 510620 229288
rect 505704 229248 510620 229276
rect 505704 229236 505710 229248
rect 510614 229236 510620 229248
rect 510672 229236 510678 229288
rect 513374 229236 513380 229288
rect 513432 229276 513438 229288
rect 519078 229276 519084 229288
rect 513432 229248 519084 229276
rect 513432 229236 513438 229248
rect 519078 229236 519084 229248
rect 519136 229236 519142 229288
rect 156322 229208 156328 229220
rect 154224 229180 156328 229208
rect 156322 229168 156328 229180
rect 156380 229168 156386 229220
rect 162578 229168 162584 229220
rect 162636 229208 162642 229220
rect 180426 229208 180432 229220
rect 162636 229180 180432 229208
rect 162636 229168 162642 229180
rect 180426 229168 180432 229180
rect 180484 229168 180490 229220
rect 183370 229168 183376 229220
rect 183428 229208 183434 229220
rect 240962 229208 240968 229220
rect 183428 229180 240968 229208
rect 183428 229168 183434 229180
rect 240962 229168 240968 229180
rect 241020 229168 241026 229220
rect 423490 229100 423496 229152
rect 423548 229140 423554 229152
rect 427722 229140 427728 229152
rect 423548 229112 427728 229140
rect 423548 229100 423554 229112
rect 427722 229100 427728 229112
rect 427780 229100 427786 229152
rect 441246 229100 441252 229152
rect 441304 229140 441310 229152
rect 442074 229140 442080 229152
rect 441304 229112 442080 229140
rect 441304 229100 441310 229112
rect 442074 229100 442080 229112
rect 442132 229100 442138 229152
rect 503714 229100 503720 229152
rect 503772 229140 503778 229152
rect 509878 229140 509884 229152
rect 503772 229112 509884 229140
rect 503772 229100 503778 229112
rect 509878 229100 509884 229112
rect 509936 229100 509942 229152
rect 515306 229100 515312 229152
rect 515364 229140 515370 229152
rect 520918 229140 520924 229152
rect 515364 229112 520924 229140
rect 515364 229100 515370 229112
rect 520918 229100 520924 229112
rect 520976 229100 520982 229152
rect 524966 229100 524972 229152
rect 525024 229140 525030 229152
rect 529934 229140 529940 229152
rect 525024 229112 529940 229140
rect 525024 229100 525030 229112
rect 529934 229100 529940 229112
rect 529992 229100 529998 229152
rect 673868 229100 673874 229152
rect 673926 229140 673932 229152
rect 673926 229112 674038 229140
rect 673926 229100 673932 229112
rect 100662 229032 100668 229084
rect 100720 229072 100726 229084
rect 167362 229072 167368 229084
rect 100720 229044 167368 229072
rect 100720 229032 100726 229044
rect 167362 229032 167368 229044
rect 167420 229032 167426 229084
rect 167546 229032 167552 229084
rect 167604 229072 167610 229084
rect 169478 229072 169484 229084
rect 167604 229044 169484 229072
rect 167604 229032 167610 229044
rect 169478 229032 169484 229044
rect 169536 229032 169542 229084
rect 179782 229072 179788 229084
rect 171796 229044 179788 229072
rect 106182 228896 106188 228948
rect 106240 228936 106246 228948
rect 171796 228936 171824 229044
rect 179782 229032 179788 229044
rect 179840 229032 179846 229084
rect 180058 229032 180064 229084
rect 180116 229072 180122 229084
rect 185578 229072 185584 229084
rect 180116 229044 185584 229072
rect 180116 229032 180122 229044
rect 185578 229032 185584 229044
rect 185636 229032 185642 229084
rect 189718 229032 189724 229084
rect 189776 229072 189782 229084
rect 189776 229044 190454 229072
rect 189776 229032 189782 229044
rect 184934 228936 184940 228948
rect 106240 228908 171824 228936
rect 171888 228908 184940 228936
rect 106240 228896 106246 228908
rect 93762 228760 93768 228812
rect 93820 228800 93826 228812
rect 166350 228800 166356 228812
rect 93820 228772 166356 228800
rect 93820 228760 93826 228772
rect 166350 228760 166356 228772
rect 166408 228760 166414 228812
rect 171888 228800 171916 228908
rect 184934 228896 184940 228908
rect 184992 228896 184998 228948
rect 185394 228896 185400 228948
rect 185452 228936 185458 228948
rect 190086 228936 190092 228948
rect 185452 228908 190092 228936
rect 185452 228896 185458 228908
rect 190086 228896 190092 228908
rect 190144 228896 190150 228948
rect 190426 228936 190454 229044
rect 192478 229032 192484 229084
rect 192536 229072 192542 229084
rect 200390 229072 200396 229084
rect 192536 229044 200396 229072
rect 192536 229032 192542 229044
rect 200390 229032 200396 229044
rect 200448 229032 200454 229084
rect 201402 229032 201408 229084
rect 201460 229072 201466 229084
rect 252554 229072 252560 229084
rect 201460 229044 252560 229072
rect 201460 229032 201466 229044
rect 252554 229032 252560 229044
rect 252612 229032 252618 229084
rect 255222 229032 255228 229084
rect 255280 229072 255286 229084
rect 295702 229072 295708 229084
rect 255280 229044 295708 229072
rect 255280 229032 255286 229044
rect 295702 229032 295708 229044
rect 295760 229032 295766 229084
rect 305546 229032 305552 229084
rect 305604 229072 305610 229084
rect 315666 229072 315672 229084
rect 305604 229044 315672 229072
rect 305604 229032 305610 229044
rect 315666 229032 315672 229044
rect 315724 229032 315730 229084
rect 326890 229032 326896 229084
rect 326948 229072 326954 229084
rect 351086 229072 351092 229084
rect 326948 229044 351092 229072
rect 326948 229032 326954 229044
rect 351086 229032 351092 229044
rect 351144 229032 351150 229084
rect 195238 228936 195244 228948
rect 190426 228908 195244 228936
rect 195238 228896 195244 228908
rect 195296 228896 195302 228948
rect 195606 228896 195612 228948
rect 195664 228936 195670 228948
rect 246758 228936 246764 228948
rect 195664 228908 246764 228936
rect 195664 228896 195670 228908
rect 246758 228896 246764 228908
rect 246816 228896 246822 228948
rect 248230 228896 248236 228948
rect 248288 228936 248294 228948
rect 291838 228936 291844 228948
rect 248288 228908 291844 228936
rect 248288 228896 248294 228908
rect 291838 228896 291844 228908
rect 291896 228896 291902 228948
rect 302142 228896 302148 228948
rect 302200 228936 302206 228948
rect 331214 228936 331220 228948
rect 302200 228908 331220 228936
rect 302200 228896 302206 228908
rect 331214 228896 331220 228908
rect 331272 228896 331278 228948
rect 506382 228896 506388 228948
rect 506440 228936 506446 228948
rect 512730 228936 512736 228948
rect 506440 228908 512736 228936
rect 506440 228896 506446 228908
rect 512730 228896 512736 228908
rect 512788 228896 512794 228948
rect 526438 228896 526444 228948
rect 526496 228936 526502 228948
rect 544010 228936 544016 228948
rect 526496 228908 544016 228936
rect 526496 228896 526502 228908
rect 544010 228896 544016 228908
rect 544068 228896 544074 228948
rect 166552 228772 171916 228800
rect 67542 228624 67548 228676
rect 67600 228664 67606 228676
rect 146018 228664 146024 228676
rect 67600 228636 146024 228664
rect 67600 228624 67606 228636
rect 146018 228624 146024 228636
rect 146076 228624 146082 228676
rect 166552 228664 166580 228772
rect 173158 228760 173164 228812
rect 173216 228800 173222 228812
rect 231302 228800 231308 228812
rect 173216 228772 231308 228800
rect 173216 228760 173222 228772
rect 231302 228760 231308 228772
rect 231360 228760 231366 228812
rect 238570 228760 238576 228812
rect 238628 228800 238634 228812
rect 282822 228800 282828 228812
rect 238628 228772 282828 228800
rect 238628 228760 238634 228772
rect 282822 228760 282828 228772
rect 282880 228760 282886 228812
rect 291838 228760 291844 228812
rect 291896 228800 291902 228812
rect 300210 228800 300216 228812
rect 291896 228772 300216 228800
rect 291896 228760 291902 228772
rect 300210 228760 300216 228772
rect 300268 228760 300274 228812
rect 300670 228760 300676 228812
rect 300728 228800 300734 228812
rect 330478 228800 330484 228812
rect 300728 228772 330484 228800
rect 300728 228760 300734 228772
rect 330478 228760 330484 228772
rect 330536 228760 330542 228812
rect 376018 228760 376024 228812
rect 376076 228800 376082 228812
rect 387794 228800 387800 228812
rect 376076 228772 387800 228800
rect 376076 228760 376082 228772
rect 387794 228760 387800 228772
rect 387852 228760 387858 228812
rect 478874 228760 478880 228812
rect 478932 228800 478938 228812
rect 490374 228800 490380 228812
rect 478932 228772 490380 228800
rect 478932 228760 478938 228772
rect 490374 228760 490380 228772
rect 490432 228760 490438 228812
rect 499850 228760 499856 228812
rect 499908 228800 499914 228812
rect 518158 228800 518164 228812
rect 499908 228772 518164 228800
rect 499908 228760 499914 228772
rect 518158 228760 518164 228772
rect 518216 228760 518222 228812
rect 518526 228760 518532 228812
rect 518584 228800 518590 228812
rect 541618 228800 541624 228812
rect 518584 228772 541624 228800
rect 518584 228760 518590 228772
rect 541618 228760 541624 228772
rect 541676 228760 541682 228812
rect 146956 228636 166580 228664
rect 61378 228488 61384 228540
rect 61436 228528 61442 228540
rect 61436 228500 137232 228528
rect 61436 228488 61442 228500
rect 57238 228352 57244 228404
rect 57296 228392 57302 228404
rect 136818 228392 136824 228404
rect 57296 228364 136824 228392
rect 57296 228352 57302 228364
rect 136818 228352 136824 228364
rect 136876 228352 136882 228404
rect 137204 228392 137232 228500
rect 137370 228488 137376 228540
rect 137428 228528 137434 228540
rect 146956 228528 146984 228636
rect 166948 228624 166954 228676
rect 167006 228664 167012 228676
rect 181438 228664 181444 228676
rect 167006 228636 181444 228664
rect 167006 228624 167012 228636
rect 181438 228624 181444 228636
rect 181496 228624 181502 228676
rect 181622 228624 181628 228676
rect 181680 228664 181686 228676
rect 185394 228664 185400 228676
rect 181680 228636 185400 228664
rect 181680 228624 181686 228636
rect 185394 228624 185400 228636
rect 185452 228624 185458 228676
rect 185578 228624 185584 228676
rect 185636 228664 185642 228676
rect 226150 228664 226156 228676
rect 185636 228636 226156 228664
rect 185636 228624 185642 228636
rect 226150 228624 226156 228636
rect 226208 228624 226214 228676
rect 226334 228624 226340 228676
rect 226392 228664 226398 228676
rect 272518 228664 272524 228676
rect 226392 228636 272524 228664
rect 226392 228624 226398 228636
rect 272518 228624 272524 228636
rect 272576 228624 272582 228676
rect 296622 228624 296628 228676
rect 296680 228664 296686 228676
rect 329190 228664 329196 228676
rect 296680 228636 329196 228664
rect 296680 228624 296686 228636
rect 329190 228624 329196 228636
rect 329248 228624 329254 228676
rect 336458 228624 336464 228676
rect 336516 228664 336522 228676
rect 358814 228664 358820 228676
rect 336516 228636 358820 228664
rect 336516 228624 336522 228636
rect 358814 228624 358820 228636
rect 358872 228624 358878 228676
rect 359918 228624 359924 228676
rect 359976 228664 359982 228676
rect 376846 228664 376852 228676
rect 359976 228636 376852 228664
rect 359976 228624 359982 228636
rect 376846 228624 376852 228636
rect 376904 228624 376910 228676
rect 485682 228624 485688 228676
rect 485740 228664 485746 228676
rect 498286 228664 498292 228676
rect 485740 228636 498292 228664
rect 485740 228624 485746 228636
rect 498286 228624 498292 228636
rect 498344 228624 498350 228676
rect 498562 228624 498568 228676
rect 498620 228664 498626 228676
rect 515766 228664 515772 228676
rect 498620 228636 515772 228664
rect 498620 228624 498626 228636
rect 515766 228624 515772 228636
rect 515824 228624 515830 228676
rect 517882 228624 517888 228676
rect 517940 228664 517946 228676
rect 539410 228664 539416 228676
rect 517940 228636 539416 228664
rect 517940 228624 517946 228636
rect 539410 228624 539416 228636
rect 539468 228624 539474 228676
rect 539594 228624 539600 228676
rect 539652 228664 539658 228676
rect 557166 228664 557172 228676
rect 539652 228636 557172 228664
rect 539652 228624 539658 228636
rect 557166 228624 557172 228636
rect 557224 228624 557230 228676
rect 137428 228500 146984 228528
rect 137428 228488 137434 228500
rect 147122 228488 147128 228540
rect 147180 228528 147186 228540
rect 200114 228528 200120 228540
rect 147180 228500 200120 228528
rect 147180 228488 147186 228500
rect 200114 228488 200120 228500
rect 200172 228488 200178 228540
rect 200298 228488 200304 228540
rect 200356 228528 200362 228540
rect 220998 228528 221004 228540
rect 200356 228500 221004 228528
rect 200356 228488 200362 228500
rect 220998 228488 221004 228500
rect 221056 228488 221062 228540
rect 264790 228528 264796 228540
rect 221200 228500 264796 228528
rect 137204 228364 137416 228392
rect 112990 228216 112996 228268
rect 113048 228256 113054 228268
rect 137186 228256 137192 228268
rect 113048 228228 137192 228256
rect 113048 228216 113054 228228
rect 137186 228216 137192 228228
rect 137244 228216 137250 228268
rect 137388 228256 137416 228364
rect 139302 228352 139308 228404
rect 139360 228392 139366 228404
rect 139360 228364 152504 228392
rect 139360 228352 139366 228364
rect 143074 228256 143080 228268
rect 137388 228228 143080 228256
rect 143074 228216 143080 228228
rect 143132 228216 143138 228268
rect 143442 228216 143448 228268
rect 143500 228256 143506 228268
rect 145834 228256 145840 228268
rect 143500 228228 145840 228256
rect 143500 228216 143506 228228
rect 145834 228216 145840 228228
rect 145892 228216 145898 228268
rect 146018 228216 146024 228268
rect 146076 228256 146082 228268
rect 148870 228256 148876 228268
rect 146076 228228 148876 228256
rect 146076 228216 146082 228228
rect 148870 228216 148876 228228
rect 148928 228216 148934 228268
rect 152476 228256 152504 228364
rect 153102 228352 153108 228404
rect 153160 228392 153166 228404
rect 215846 228392 215852 228404
rect 153160 228364 215852 228392
rect 153160 228352 153166 228364
rect 215846 228352 215852 228364
rect 215904 228352 215910 228404
rect 216490 228352 216496 228404
rect 216548 228392 216554 228404
rect 221200 228392 221228 228500
rect 264790 228488 264796 228500
rect 264848 228488 264854 228540
rect 272518 228488 272524 228540
rect 272576 228528 272582 228540
rect 309870 228528 309876 228540
rect 272576 228500 309876 228528
rect 272576 228488 272582 228500
rect 309870 228488 309876 228500
rect 309928 228488 309934 228540
rect 313918 228488 313924 228540
rect 313976 228528 313982 228540
rect 320818 228528 320824 228540
rect 313976 228500 320824 228528
rect 313976 228488 313982 228500
rect 320818 228488 320824 228500
rect 320876 228488 320882 228540
rect 325418 228488 325424 228540
rect 325476 228528 325482 228540
rect 349154 228528 349160 228540
rect 325476 228500 349160 228528
rect 325476 228488 325482 228500
rect 349154 228488 349160 228500
rect 349212 228488 349218 228540
rect 350442 228488 350448 228540
rect 350500 228528 350506 228540
rect 369118 228528 369124 228540
rect 350500 228500 369124 228528
rect 350500 228488 350506 228500
rect 369118 228488 369124 228500
rect 369176 228488 369182 228540
rect 371050 228488 371056 228540
rect 371108 228528 371114 228540
rect 385218 228528 385224 228540
rect 371108 228500 385224 228528
rect 371108 228488 371114 228500
rect 385218 228488 385224 228500
rect 385276 228488 385282 228540
rect 386046 228488 386052 228540
rect 386104 228528 386110 228540
rect 397454 228528 397460 228540
rect 386104 228500 397460 228528
rect 386104 228488 386110 228500
rect 397454 228488 397460 228500
rect 397512 228488 397518 228540
rect 407758 228528 407764 228540
rect 400232 228500 407764 228528
rect 216548 228364 221228 228392
rect 216548 228352 216554 228364
rect 224770 228352 224776 228404
rect 224828 228392 224834 228404
rect 273806 228392 273812 228404
rect 224828 228364 273812 228392
rect 224828 228352 224834 228364
rect 273806 228352 273812 228364
rect 273864 228352 273870 228404
rect 285490 228352 285496 228404
rect 285548 228392 285554 228404
rect 318886 228392 318892 228404
rect 285548 228364 318892 228392
rect 285548 228352 285554 228364
rect 318886 228352 318892 228364
rect 318944 228352 318950 228404
rect 330478 228352 330484 228404
rect 330536 228392 330542 228404
rect 354950 228392 354956 228404
rect 330536 228364 354956 228392
rect 330536 228352 330542 228364
rect 354950 228352 354956 228364
rect 355008 228352 355014 228404
rect 355318 228352 355324 228404
rect 355376 228392 355382 228404
rect 372982 228392 372988 228404
rect 355376 228364 372988 228392
rect 355376 228352 355382 228364
rect 372982 228352 372988 228364
rect 373040 228352 373046 228404
rect 373442 228352 373448 228404
rect 373500 228392 373506 228404
rect 387150 228392 387156 228404
rect 373500 228364 387156 228392
rect 373500 228352 373506 228364
rect 387150 228352 387156 228364
rect 387208 228352 387214 228404
rect 390002 228352 390008 228404
rect 390060 228392 390066 228404
rect 400030 228392 400036 228404
rect 390060 228364 400036 228392
rect 390060 228352 390066 228364
rect 400030 228352 400036 228364
rect 400088 228352 400094 228404
rect 205542 228256 205548 228268
rect 152476 228228 205548 228256
rect 205542 228216 205548 228228
rect 205600 228216 205606 228268
rect 205726 228216 205732 228268
rect 205784 228256 205790 228268
rect 257062 228256 257068 228268
rect 205784 228228 257068 228256
rect 205784 228216 205790 228228
rect 257062 228216 257068 228228
rect 257120 228216 257126 228268
rect 257614 228216 257620 228268
rect 257672 228256 257678 228268
rect 296346 228256 296352 228268
rect 257672 228228 296352 228256
rect 257672 228216 257678 228228
rect 296346 228216 296352 228228
rect 296404 228216 296410 228268
rect 400232 228256 400260 228500
rect 407758 228488 407764 228500
rect 407816 228488 407822 228540
rect 409782 228488 409788 228540
rect 409840 228528 409846 228540
rect 415486 228528 415492 228540
rect 409840 228500 415492 228528
rect 409840 228488 409846 228500
rect 415486 228488 415492 228500
rect 415544 228488 415550 228540
rect 485038 228488 485044 228540
rect 485096 228528 485102 228540
rect 498654 228528 498660 228540
rect 485096 228500 498660 228528
rect 485096 228488 485102 228500
rect 498654 228488 498660 228500
rect 498712 228488 498718 228540
rect 502426 228488 502432 228540
rect 502484 228528 502490 228540
rect 521102 228528 521108 228540
rect 502484 228500 521108 228528
rect 502484 228488 502490 228500
rect 521102 228488 521108 228500
rect 521160 228488 521166 228540
rect 527542 228488 527548 228540
rect 527600 228528 527606 228540
rect 553302 228528 553308 228540
rect 527600 228500 553308 228528
rect 527600 228488 527606 228500
rect 553302 228488 553308 228500
rect 553360 228488 553366 228540
rect 556798 228488 556804 228540
rect 556856 228528 556862 228540
rect 570598 228528 570604 228540
rect 556856 228500 570604 228528
rect 556856 228488 556862 228500
rect 570598 228488 570604 228500
rect 570656 228488 570662 228540
rect 402790 228352 402796 228404
rect 402848 228392 402854 228404
rect 411622 228392 411628 228404
rect 402848 228364 411628 228392
rect 402848 228352 402854 228364
rect 411622 228352 411628 228364
rect 411680 228352 411686 228404
rect 474458 228352 474464 228404
rect 474516 228392 474522 228404
rect 484486 228392 484492 228404
rect 474516 228364 484492 228392
rect 474516 228352 474522 228364
rect 484486 228352 484492 228364
rect 484544 228352 484550 228404
rect 490190 228352 490196 228404
rect 490248 228392 490254 228404
rect 505186 228392 505192 228404
rect 490248 228364 505192 228392
rect 490248 228352 490254 228364
rect 505186 228352 505192 228364
rect 505244 228352 505250 228404
rect 512086 228352 512092 228404
rect 512144 228392 512150 228404
rect 533522 228392 533528 228404
rect 512144 228364 533528 228392
rect 512144 228352 512150 228364
rect 533522 228352 533528 228364
rect 533580 228352 533586 228404
rect 537202 228352 537208 228404
rect 537260 228392 537266 228404
rect 565630 228392 565636 228404
rect 537260 228364 565636 228392
rect 537260 228352 537266 228364
rect 565630 228352 565636 228364
rect 565688 228352 565694 228404
rect 672488 228352 672494 228404
rect 672546 228392 672552 228404
rect 673086 228392 673092 228404
rect 672546 228364 673092 228392
rect 672546 228352 672552 228364
rect 673086 228352 673092 228364
rect 673144 228352 673150 228404
rect 400140 228228 400260 228256
rect 400140 228132 400168 228228
rect 539410 228216 539416 228268
rect 539468 228256 539474 228268
rect 540790 228256 540796 228268
rect 539468 228228 540796 228256
rect 539468 228216 539474 228228
rect 540790 228216 540796 228228
rect 540848 228216 540854 228268
rect 119982 228080 119988 228132
rect 120040 228120 120046 228132
rect 181254 228120 181260 228132
rect 120040 228092 181260 228120
rect 120040 228080 120046 228092
rect 181254 228080 181260 228092
rect 181312 228080 181318 228132
rect 181438 228080 181444 228132
rect 181496 228120 181502 228132
rect 181496 228092 194180 228120
rect 181496 228080 181502 228092
rect 126698 227944 126704 227996
rect 126756 227984 126762 227996
rect 194152 227984 194180 228092
rect 195238 228080 195244 228132
rect 195296 228120 195302 228132
rect 239030 228120 239036 228132
rect 195296 228092 239036 228120
rect 195296 228080 195302 228092
rect 239030 228080 239036 228092
rect 239088 228080 239094 228132
rect 246298 228080 246304 228132
rect 246356 228120 246362 228132
rect 253842 228120 253848 228132
rect 246356 228092 253848 228120
rect 246356 228080 246362 228092
rect 253842 228080 253848 228092
rect 253900 228080 253906 228132
rect 268930 228080 268936 228132
rect 268988 228120 268994 228132
rect 306006 228120 306012 228132
rect 268988 228092 306012 228120
rect 268988 228080 268994 228092
rect 306006 228080 306012 228092
rect 306064 228080 306070 228132
rect 400122 228080 400128 228132
rect 400180 228080 400186 228132
rect 415026 228012 415032 228064
rect 415084 228052 415090 228064
rect 421926 228052 421932 228064
rect 415084 228024 421932 228052
rect 415084 228012 415090 228024
rect 421926 228012 421932 228024
rect 421984 228012 421990 228064
rect 200298 227984 200304 227996
rect 126756 227956 192892 227984
rect 194152 227956 200304 227984
rect 126756 227944 126762 227956
rect 88242 227808 88248 227860
rect 88300 227848 88306 227860
rect 95234 227848 95240 227860
rect 88300 227820 95240 227848
rect 88300 227808 88306 227820
rect 95234 227808 95240 227820
rect 95292 227808 95298 227860
rect 133506 227808 133512 227860
rect 133564 227848 133570 227860
rect 136634 227848 136640 227860
rect 133564 227820 136640 227848
rect 133564 227808 133570 227820
rect 136634 227808 136640 227820
rect 136692 227808 136698 227860
rect 136818 227808 136824 227860
rect 136876 227848 136882 227860
rect 141142 227848 141148 227860
rect 136876 227820 141148 227848
rect 136876 227808 136882 227820
rect 141142 227808 141148 227820
rect 141200 227808 141206 227860
rect 141510 227808 141516 227860
rect 141568 227848 141574 227860
rect 192478 227848 192484 227860
rect 141568 227820 192484 227848
rect 141568 227808 141574 227820
rect 192478 227808 192484 227820
rect 192536 227808 192542 227860
rect 192864 227848 192892 227956
rect 200298 227944 200304 227956
rect 200356 227944 200362 227996
rect 210418 227944 210424 227996
rect 210476 227984 210482 227996
rect 238386 227984 238392 227996
rect 210476 227956 238392 227984
rect 210476 227944 210482 227956
rect 238386 227944 238392 227956
rect 238444 227944 238450 227996
rect 416682 227876 416688 227928
rect 416740 227916 416746 227928
rect 420638 227916 420644 227928
rect 416740 227888 420644 227916
rect 416740 227876 416746 227888
rect 420638 227876 420644 227888
rect 420696 227876 420702 227928
rect 447042 227876 447048 227928
rect 447100 227916 447106 227928
rect 450538 227916 450544 227928
rect 447100 227888 450544 227916
rect 447100 227876 447106 227888
rect 450538 227876 450544 227888
rect 450596 227876 450602 227928
rect 195054 227848 195060 227860
rect 192864 227820 195060 227848
rect 195054 227808 195060 227820
rect 195112 227808 195118 227860
rect 200114 227808 200120 227860
rect 200172 227848 200178 227860
rect 210234 227848 210240 227860
rect 200172 227820 210240 227848
rect 200172 227808 200178 227820
rect 210234 227808 210240 227820
rect 210292 227808 210298 227860
rect 409046 227740 409052 227792
rect 409104 227780 409110 227792
rect 410334 227780 410340 227792
rect 409104 227752 410340 227780
rect 409104 227740 409110 227752
rect 410334 227740 410340 227752
rect 410392 227740 410398 227792
rect 411898 227740 411904 227792
rect 411956 227780 411962 227792
rect 413554 227780 413560 227792
rect 411956 227752 413560 227780
rect 411956 227740 411962 227752
rect 413554 227740 413560 227752
rect 413612 227740 413618 227792
rect 420638 227740 420644 227792
rect 420696 227780 420702 227792
rect 423858 227780 423864 227792
rect 420696 227752 423864 227780
rect 420696 227740 420702 227752
rect 423858 227740 423864 227752
rect 423916 227740 423922 227792
rect 471514 227740 471520 227792
rect 471572 227780 471578 227792
rect 479518 227780 479524 227792
rect 471572 227752 479524 227780
rect 471572 227740 471578 227752
rect 479518 227740 479524 227752
rect 479576 227740 479582 227792
rect 75178 227672 75184 227724
rect 75236 227712 75242 227724
rect 146294 227712 146300 227724
rect 75236 227684 146300 227712
rect 75236 227672 75242 227684
rect 146294 227672 146300 227684
rect 146352 227672 146358 227724
rect 150066 227672 150072 227724
rect 150124 227712 150130 227724
rect 213362 227712 213368 227724
rect 150124 227684 213368 227712
rect 150124 227672 150130 227684
rect 213362 227672 213368 227684
rect 213420 227672 213426 227724
rect 213822 227672 213828 227724
rect 213880 227712 213886 227724
rect 262858 227712 262864 227724
rect 213880 227684 262864 227712
rect 213880 227672 213886 227684
rect 262858 227672 262864 227684
rect 262916 227672 262922 227724
rect 263502 227672 263508 227724
rect 263560 227712 263566 227724
rect 277210 227712 277216 227724
rect 263560 227684 277216 227712
rect 263560 227672 263566 227684
rect 277210 227672 277216 227684
rect 277268 227672 277274 227724
rect 311802 227712 311808 227724
rect 277366 227684 311808 227712
rect 64782 227536 64788 227588
rect 64840 227576 64846 227588
rect 110138 227576 110144 227588
rect 64840 227548 110144 227576
rect 64840 227536 64846 227548
rect 110138 227536 110144 227548
rect 110196 227536 110202 227588
rect 110322 227536 110328 227588
rect 110380 227576 110386 227588
rect 182358 227576 182364 227588
rect 110380 227548 182364 227576
rect 110380 227536 110386 227548
rect 182358 227536 182364 227548
rect 182416 227536 182422 227588
rect 185394 227536 185400 227588
rect 185452 227576 185458 227588
rect 192662 227576 192668 227588
rect 185452 227548 192668 227576
rect 185452 227536 185458 227548
rect 192662 227536 192668 227548
rect 192720 227536 192726 227588
rect 200022 227536 200028 227588
rect 200080 227576 200086 227588
rect 200080 227548 205036 227576
rect 200080 227536 200086 227548
rect 205008 227508 205036 227548
rect 205634 227536 205640 227588
rect 205692 227576 205698 227588
rect 214558 227576 214564 227588
rect 205692 227548 214564 227576
rect 205692 227536 205698 227548
rect 214558 227536 214564 227548
rect 214616 227536 214622 227588
rect 214742 227536 214748 227588
rect 214800 227576 214806 227588
rect 262214 227576 262220 227588
rect 214800 227548 262220 227576
rect 214800 227536 214806 227548
rect 262214 227536 262220 227548
rect 262272 227536 262278 227588
rect 277210 227536 277216 227588
rect 277268 227576 277274 227588
rect 277366 227576 277394 227684
rect 311802 227672 311808 227684
rect 311860 227672 311866 227724
rect 465902 227604 465908 227656
rect 465960 227644 465966 227656
rect 469858 227644 469864 227656
rect 465960 227616 469864 227644
rect 465960 227604 465966 227616
rect 469858 227604 469864 227616
rect 469916 227604 469922 227656
rect 277268 227548 277394 227576
rect 277268 227536 277274 227548
rect 282178 227536 282184 227588
rect 282236 227576 282242 227588
rect 308582 227576 308588 227588
rect 282236 227548 308588 227576
rect 282236 227536 282242 227548
rect 308582 227536 308588 227548
rect 308640 227536 308646 227588
rect 524598 227536 524604 227588
rect 524656 227576 524662 227588
rect 539962 227576 539968 227588
rect 524656 227548 539968 227576
rect 524656 227536 524662 227548
rect 539962 227536 539968 227548
rect 540020 227536 540026 227588
rect 205008 227480 205220 227508
rect 60642 227400 60648 227452
rect 60700 227440 60706 227452
rect 102134 227440 102140 227452
rect 60700 227412 102140 227440
rect 60700 227400 60706 227412
rect 102134 227400 102140 227412
rect 102192 227400 102198 227452
rect 103422 227400 103428 227452
rect 103480 227440 103486 227452
rect 177206 227440 177212 227452
rect 103480 227412 177212 227440
rect 103480 227400 103486 227412
rect 177206 227400 177212 227412
rect 177264 227400 177270 227452
rect 181254 227400 181260 227452
rect 181312 227440 181318 227452
rect 181312 227412 185808 227440
rect 181312 227400 181318 227412
rect 96522 227264 96528 227316
rect 96580 227304 96586 227316
rect 169386 227304 169392 227316
rect 96580 227276 169392 227304
rect 96580 227264 96586 227276
rect 169386 227264 169392 227276
rect 169444 227264 169450 227316
rect 169570 227264 169576 227316
rect 169628 227304 169634 227316
rect 169628 227276 171732 227304
rect 169628 227264 169634 227276
rect 171704 227236 171732 227276
rect 172054 227264 172060 227316
rect 172112 227304 172118 227316
rect 185578 227304 185584 227316
rect 172112 227276 185584 227304
rect 172112 227264 172118 227276
rect 185578 227264 185584 227276
rect 185636 227264 185642 227316
rect 185780 227304 185808 227412
rect 186130 227400 186136 227452
rect 186188 227440 186194 227452
rect 204806 227440 204812 227452
rect 186188 227412 204812 227440
rect 186188 227400 186194 227412
rect 204806 227400 204812 227412
rect 204864 227400 204870 227452
rect 205192 227440 205220 227480
rect 251910 227440 251916 227452
rect 205192 227412 251916 227440
rect 251910 227400 251916 227412
rect 251968 227400 251974 227452
rect 259270 227400 259276 227452
rect 259328 227440 259334 227452
rect 298278 227440 298284 227452
rect 259328 227412 298284 227440
rect 259328 227400 259334 227412
rect 298278 227400 298284 227412
rect 298336 227400 298342 227452
rect 304902 227400 304908 227452
rect 304960 227440 304966 227452
rect 333698 227440 333704 227452
rect 304960 227412 333704 227440
rect 304960 227400 304966 227412
rect 333698 227400 333704 227412
rect 333756 227400 333762 227452
rect 333882 227400 333888 227452
rect 333940 227440 333946 227452
rect 356238 227440 356244 227452
rect 333940 227412 356244 227440
rect 333940 227400 333946 227412
rect 356238 227400 356244 227412
rect 356296 227400 356302 227452
rect 357066 227400 357072 227452
rect 357124 227440 357130 227452
rect 374270 227440 374276 227452
rect 357124 227412 374276 227440
rect 357124 227400 357130 227412
rect 374270 227400 374276 227412
rect 374328 227400 374334 227452
rect 514018 227400 514024 227452
rect 514076 227440 514082 227452
rect 535730 227440 535736 227452
rect 514076 227412 535736 227440
rect 514076 227400 514082 227412
rect 535730 227400 535736 227412
rect 535788 227400 535794 227452
rect 538306 227400 538312 227452
rect 538364 227440 538370 227452
rect 556062 227440 556068 227452
rect 538364 227412 556068 227440
rect 538364 227400 538370 227412
rect 556062 227400 556068 227412
rect 556120 227400 556126 227452
rect 219158 227304 219164 227316
rect 185780 227276 219164 227304
rect 219158 227264 219164 227276
rect 219216 227264 219222 227316
rect 220078 227264 220084 227316
rect 220136 227304 220142 227316
rect 241606 227304 241612 227316
rect 220136 227276 241612 227304
rect 220136 227264 220142 227276
rect 241606 227264 241612 227276
rect 241664 227264 241670 227316
rect 257798 227264 257804 227316
rect 257856 227304 257862 227316
rect 299566 227304 299572 227316
rect 257856 227276 299572 227304
rect 257856 227264 257862 227276
rect 299566 227264 299572 227276
rect 299624 227264 299630 227316
rect 310422 227264 310428 227316
rect 310480 227304 310486 227316
rect 338206 227304 338212 227316
rect 310480 227276 338212 227304
rect 310480 227264 310486 227276
rect 338206 227264 338212 227276
rect 338264 227264 338270 227316
rect 340690 227264 340696 227316
rect 340748 227304 340754 227316
rect 361390 227304 361396 227316
rect 340748 227276 361396 227304
rect 340748 227264 340754 227276
rect 361390 227264 361396 227276
rect 361448 227264 361454 227316
rect 402606 227304 402612 227316
rect 393286 227276 402612 227304
rect 171704 227208 171916 227236
rect 89622 227128 89628 227180
rect 89680 227168 89686 227180
rect 157288 227168 157294 227180
rect 89680 227140 157294 227168
rect 89680 227128 89686 227140
rect 157288 227128 157294 227140
rect 157346 227128 157352 227180
rect 157426 227128 157432 227180
rect 157484 227168 157490 227180
rect 171502 227168 171508 227180
rect 157484 227140 171508 227168
rect 157484 227128 157490 227140
rect 171502 227128 171508 227140
rect 171560 227128 171566 227180
rect 171888 227168 171916 227208
rect 171888 227140 224954 227168
rect 56502 226992 56508 227044
rect 56560 227032 56566 227044
rect 142430 227032 142436 227044
rect 56560 227004 142436 227032
rect 56560 226992 56566 227004
rect 142430 226992 142436 227004
rect 142488 226992 142494 227044
rect 143258 226992 143264 227044
rect 143316 227032 143322 227044
rect 208118 227032 208124 227044
rect 143316 227004 208124 227032
rect 143316 226992 143322 227004
rect 208118 226992 208124 227004
rect 208176 226992 208182 227044
rect 214558 226992 214564 227044
rect 214616 227032 214622 227044
rect 220078 227032 220084 227044
rect 214616 227004 220084 227032
rect 214616 226992 214622 227004
rect 220078 226992 220084 227004
rect 220136 226992 220142 227044
rect 220446 226992 220452 227044
rect 220504 227032 220510 227044
rect 222930 227032 222936 227044
rect 220504 227004 222936 227032
rect 220504 226992 220510 227004
rect 222930 226992 222936 227004
rect 222988 226992 222994 227044
rect 224926 227032 224954 227140
rect 235810 227128 235816 227180
rect 235868 227168 235874 227180
rect 280246 227168 280252 227180
rect 235868 227140 280252 227168
rect 235868 227128 235874 227140
rect 280246 227128 280252 227140
rect 280304 227128 280310 227180
rect 306190 227128 306196 227180
rect 306248 227168 306254 227180
rect 336918 227168 336924 227180
rect 306248 227140 336924 227168
rect 306248 227128 306254 227140
rect 336918 227128 336924 227140
rect 336976 227128 336982 227180
rect 338666 227128 338672 227180
rect 338724 227168 338730 227180
rect 360102 227168 360108 227180
rect 338724 227140 360108 227168
rect 338724 227128 338730 227140
rect 360102 227128 360108 227140
rect 360160 227128 360166 227180
rect 362770 227128 362776 227180
rect 362828 227168 362834 227180
rect 379422 227168 379428 227180
rect 362828 227140 379428 227168
rect 362828 227128 362834 227140
rect 379422 227128 379428 227140
rect 379480 227128 379486 227180
rect 382090 227128 382096 227180
rect 382148 227168 382154 227180
rect 392946 227168 392952 227180
rect 382148 227140 392952 227168
rect 382148 227128 382154 227140
rect 392946 227128 392952 227140
rect 393004 227128 393010 227180
rect 393130 227128 393136 227180
rect 393188 227168 393194 227180
rect 393286 227168 393314 227276
rect 402606 227264 402612 227276
rect 402664 227264 402670 227316
rect 494698 227264 494704 227316
rect 494756 227304 494762 227316
rect 494756 227276 504404 227304
rect 494756 227264 494762 227276
rect 393188 227140 393314 227168
rect 393188 227128 393194 227140
rect 402238 227128 402244 227180
rect 402296 227168 402302 227180
rect 408402 227168 408408 227180
rect 402296 227140 408408 227168
rect 402296 227128 402302 227140
rect 408402 227128 408408 227140
rect 408460 227128 408466 227180
rect 478598 227128 478604 227180
rect 478656 227168 478662 227180
rect 486786 227168 486792 227180
rect 478656 227140 486792 227168
rect 478656 227128 478662 227140
rect 486786 227128 486792 227140
rect 486844 227128 486850 227180
rect 489546 227128 489552 227180
rect 489604 227168 489610 227180
rect 504174 227168 504180 227180
rect 489604 227140 504180 227168
rect 489604 227128 489610 227140
rect 504174 227128 504180 227140
rect 504232 227128 504238 227180
rect 228726 227032 228732 227044
rect 224926 227004 228732 227032
rect 228726 226992 228732 227004
rect 228784 226992 228790 227044
rect 228910 226992 228916 227044
rect 228968 227032 228974 227044
rect 271230 227032 271236 227044
rect 228968 227004 271236 227032
rect 228968 226992 228974 227004
rect 271230 226992 271236 227004
rect 271288 226992 271294 227044
rect 271782 226992 271788 227044
rect 271840 227032 271846 227044
rect 282178 227032 282184 227044
rect 271840 227004 282184 227032
rect 271840 226992 271846 227004
rect 282178 226992 282184 227004
rect 282236 226992 282242 227044
rect 317598 227032 317604 227044
rect 287026 227004 317604 227032
rect 122742 226856 122748 226908
rect 122800 226896 122806 226908
rect 185394 226896 185400 226908
rect 122800 226868 185400 226896
rect 122800 226856 122806 226868
rect 185394 226856 185400 226868
rect 185452 226856 185458 226908
rect 185578 226856 185584 226908
rect 185636 226896 185642 226908
rect 218422 226896 218428 226908
rect 185636 226868 218428 226896
rect 185636 226856 185642 226868
rect 218422 226856 218428 226868
rect 218480 226856 218486 226908
rect 219342 226856 219348 226908
rect 219400 226896 219406 226908
rect 267366 226896 267372 226908
rect 219400 226868 267372 226896
rect 219400 226856 219406 226868
rect 267366 226856 267372 226868
rect 267424 226856 267430 226908
rect 281350 226856 281356 226908
rect 281408 226896 281414 226908
rect 287026 226896 287054 227004
rect 317598 226992 317604 227004
rect 317656 226992 317662 227044
rect 322842 226992 322848 227044
rect 322900 227032 322906 227044
rect 349798 227032 349804 227044
rect 322900 227004 349804 227032
rect 322900 226992 322906 227004
rect 349798 226992 349804 227004
rect 349856 226992 349862 227044
rect 355870 226992 355876 227044
rect 355928 227032 355934 227044
rect 375558 227032 375564 227044
rect 355928 227004 375564 227032
rect 355928 226992 355934 227004
rect 375558 226992 375564 227004
rect 375616 226992 375622 227044
rect 376662 226992 376668 227044
rect 376720 227032 376726 227044
rect 389726 227032 389732 227044
rect 376720 227004 389732 227032
rect 376720 226992 376726 227004
rect 389726 226992 389732 227004
rect 389784 226992 389790 227044
rect 391842 226992 391848 227044
rect 391900 227032 391906 227044
rect 403526 227032 403532 227044
rect 391900 227004 403532 227032
rect 391900 226992 391906 227004
rect 403526 226992 403532 227004
rect 403584 226992 403590 227044
rect 412542 226992 412548 227044
rect 412600 227032 412606 227044
rect 419350 227032 419356 227044
rect 412600 227004 419356 227032
rect 412600 226992 412606 227004
rect 419350 226992 419356 227004
rect 419408 226992 419414 227044
rect 486970 226992 486976 227044
rect 487028 227032 487034 227044
rect 500954 227032 500960 227044
rect 487028 227004 500960 227032
rect 487028 226992 487034 227004
rect 500954 226992 500960 227004
rect 501012 226992 501018 227044
rect 281408 226868 287054 226896
rect 281408 226856 281414 226868
rect 293770 226856 293776 226908
rect 293828 226896 293834 226908
rect 324958 226896 324964 226908
rect 293828 226868 324964 226896
rect 293828 226856 293834 226868
rect 324958 226856 324964 226868
rect 325016 226856 325022 226908
rect 504376 226896 504404 227276
rect 510614 227264 510620 227316
rect 510672 227304 510678 227316
rect 524414 227304 524420 227316
rect 510672 227276 524420 227304
rect 510672 227264 510678 227276
rect 524414 227264 524420 227276
rect 524472 227264 524478 227316
rect 526254 227264 526260 227316
rect 526312 227304 526318 227316
rect 551554 227304 551560 227316
rect 526312 227276 551560 227304
rect 526312 227264 526318 227276
rect 551554 227264 551560 227276
rect 551612 227264 551618 227316
rect 506198 227128 506204 227180
rect 506256 227168 506262 227180
rect 525978 227168 525984 227180
rect 506256 227140 525984 227168
rect 506256 227128 506262 227140
rect 525978 227128 525984 227140
rect 526036 227128 526042 227180
rect 533338 227128 533344 227180
rect 533396 227168 533402 227180
rect 560938 227168 560944 227180
rect 533396 227140 560944 227168
rect 533396 227128 533402 227140
rect 560938 227128 560944 227140
rect 560996 227128 561002 227180
rect 669222 227128 669228 227180
rect 669280 227168 669286 227180
rect 669866 227168 669872 227180
rect 669280 227140 669872 227168
rect 669280 227128 669286 227140
rect 669866 227128 669872 227140
rect 669924 227128 669930 227180
rect 505002 226992 505008 227044
rect 505060 227032 505066 227044
rect 523034 227032 523040 227044
rect 505060 227004 523040 227032
rect 505060 226992 505066 227004
rect 523034 226992 523040 227004
rect 523092 226992 523098 227044
rect 523678 226992 523684 227044
rect 523736 227032 523742 227044
rect 548334 227032 548340 227044
rect 523736 227004 548340 227032
rect 523736 226992 523742 227004
rect 548334 226992 548340 227004
rect 548392 226992 548398 227044
rect 555418 226992 555424 227044
rect 555476 227032 555482 227044
rect 633710 227032 633716 227044
rect 555476 227004 633716 227032
rect 555476 226992 555482 227004
rect 633710 226992 633716 227004
rect 633768 226992 633774 227044
rect 672534 227032 672540 227044
rect 669286 227004 672540 227032
rect 510982 226896 510988 226908
rect 504376 226868 510988 226896
rect 510982 226856 510988 226868
rect 511040 226856 511046 226908
rect 117222 226720 117228 226772
rect 117280 226760 117286 226772
rect 187510 226760 187516 226772
rect 117280 226732 187516 226760
rect 117280 226720 117286 226732
rect 187510 226720 187516 226732
rect 187568 226720 187574 226772
rect 189994 226720 190000 226772
rect 190052 226760 190058 226772
rect 233878 226760 233884 226772
rect 190052 226732 233884 226760
rect 190052 226720 190058 226732
rect 233878 226720 233884 226732
rect 233936 226720 233942 226772
rect 249610 226720 249616 226772
rect 249668 226760 249674 226772
rect 290550 226760 290556 226772
rect 249668 226732 290556 226760
rect 249668 226720 249674 226732
rect 290550 226720 290556 226732
rect 290608 226720 290614 226772
rect 668394 226720 668400 226772
rect 668452 226760 668458 226772
rect 669286 226760 669314 227004
rect 672534 226992 672540 227004
rect 672592 226992 672598 227044
rect 668452 226732 669314 226760
rect 668452 226720 668458 226732
rect 243446 226652 243452 226704
rect 243504 226692 243510 226704
rect 248690 226692 248696 226704
rect 243504 226664 248696 226692
rect 243504 226652 243510 226664
rect 248690 226652 248696 226664
rect 248748 226652 248754 226704
rect 129550 226584 129556 226636
rect 129608 226624 129614 226636
rect 197354 226624 197360 226636
rect 129608 226596 197360 226624
rect 129608 226584 129614 226596
rect 197354 226584 197360 226596
rect 197412 226584 197418 226636
rect 203518 226584 203524 226636
rect 203576 226624 203582 226636
rect 203576 226596 215294 226624
rect 203576 226584 203582 226596
rect 136542 226448 136548 226500
rect 136600 226488 136606 226500
rect 141786 226488 141792 226500
rect 136600 226460 141792 226488
rect 136600 226448 136606 226460
rect 141786 226448 141792 226460
rect 141844 226448 141850 226500
rect 142246 226448 142252 226500
rect 142304 226488 142310 226500
rect 202966 226488 202972 226500
rect 142304 226460 202972 226488
rect 142304 226448 142310 226460
rect 202966 226448 202972 226460
rect 203024 226448 203030 226500
rect 212166 226448 212172 226500
rect 212224 226488 212230 226500
rect 214742 226488 214748 226500
rect 212224 226460 214748 226488
rect 212224 226448 212230 226460
rect 214742 226448 214748 226460
rect 214800 226448 214806 226500
rect 215266 226488 215294 226596
rect 219158 226584 219164 226636
rect 219216 226624 219222 226636
rect 223574 226624 223580 226636
rect 219216 226596 223580 226624
rect 219216 226584 219222 226596
rect 223574 226584 223580 226596
rect 223632 226584 223638 226636
rect 231026 226584 231032 226636
rect 231084 226624 231090 226636
rect 243262 226624 243268 226636
rect 231084 226596 243268 226624
rect 231084 226584 231090 226596
rect 243262 226584 243268 226596
rect 243320 226584 243326 226636
rect 264146 226584 264152 226636
rect 264204 226624 264210 226636
rect 269298 226624 269304 226636
rect 264204 226596 269304 226624
rect 264204 226584 264210 226596
rect 269298 226584 269304 226596
rect 269356 226584 269362 226636
rect 669866 226584 669872 226636
rect 669924 226624 669930 226636
rect 670510 226624 670516 226636
rect 669924 226596 670516 226624
rect 669924 226584 669930 226596
rect 670510 226584 670516 226596
rect 670568 226584 670574 226636
rect 673270 226556 673276 226568
rect 672842 226528 673276 226556
rect 673270 226516 673276 226528
rect 673328 226516 673334 226568
rect 220446 226488 220452 226500
rect 215266 226460 220452 226488
rect 220446 226448 220452 226460
rect 220504 226448 220510 226500
rect 221826 226448 221832 226500
rect 221884 226488 221890 226500
rect 228910 226488 228916 226500
rect 221884 226460 228916 226488
rect 221884 226448 221890 226460
rect 228910 226448 228916 226460
rect 228968 226448 228974 226500
rect 351086 226448 351092 226500
rect 351144 226488 351150 226500
rect 353018 226488 353024 226500
rect 351144 226460 353024 226488
rect 351144 226448 351150 226460
rect 353018 226448 353024 226460
rect 353076 226448 353082 226500
rect 403986 226448 403992 226500
rect 404044 226488 404050 226500
rect 412266 226488 412272 226500
rect 404044 226460 412272 226488
rect 404044 226448 404050 226460
rect 412266 226448 412272 226460
rect 412324 226448 412330 226500
rect 474734 226448 474740 226500
rect 474792 226488 474798 226500
rect 482738 226488 482744 226500
rect 474792 226460 482744 226488
rect 474792 226448 474798 226460
rect 482738 226448 482744 226460
rect 482796 226448 482802 226500
rect 672724 226432 672776 226438
rect 141970 226380 141976 226432
rect 142028 226420 142034 226432
rect 142108 226420 142114 226432
rect 142028 226392 142114 226420
rect 142028 226380 142034 226392
rect 142108 226380 142114 226392
rect 142166 226380 142172 226432
rect 271138 226380 271144 226432
rect 271196 226420 271202 226432
rect 279602 226420 279608 226432
rect 271196 226392 279608 226420
rect 271196 226380 271202 226392
rect 279602 226380 279608 226392
rect 279660 226380 279666 226432
rect 672724 226374 672776 226380
rect 350258 226312 350264 226364
rect 350316 226352 350322 226364
rect 351730 226352 351736 226364
rect 350316 226324 351736 226352
rect 350316 226312 350322 226324
rect 351730 226312 351736 226324
rect 351788 226312 351794 226364
rect 388530 226312 388536 226364
rect 388588 226352 388594 226364
rect 391658 226352 391664 226364
rect 388588 226324 391664 226352
rect 388588 226312 388594 226324
rect 391658 226312 391664 226324
rect 391716 226312 391722 226364
rect 407758 226312 407764 226364
rect 407816 226352 407822 226364
rect 408678 226352 408684 226364
rect 407816 226324 408684 226352
rect 407816 226312 407822 226324
rect 408678 226312 408684 226324
rect 408736 226312 408742 226364
rect 481634 226312 481640 226364
rect 481692 226352 481698 226364
rect 487798 226352 487804 226364
rect 481692 226324 487804 226352
rect 481692 226312 481698 226324
rect 487798 226312 487804 226324
rect 487856 226312 487862 226364
rect 663426 226312 663432 226364
rect 663484 226352 663490 226364
rect 665266 226352 665272 226364
rect 663484 226324 665272 226352
rect 663484 226312 663490 226324
rect 665266 226312 665272 226324
rect 665324 226312 665330 226364
rect 58986 226244 58992 226296
rect 59044 226284 59050 226296
rect 130378 226284 130384 226296
rect 59044 226256 130384 226284
rect 59044 226244 59050 226256
rect 130378 226244 130384 226256
rect 130436 226244 130442 226296
rect 135070 226244 135076 226296
rect 135128 226284 135134 226296
rect 204254 226284 204260 226296
rect 135128 226256 204260 226284
rect 135128 226244 135134 226256
rect 204254 226244 204260 226256
rect 204312 226244 204318 226296
rect 208118 226244 208124 226296
rect 208176 226284 208182 226296
rect 257430 226284 257436 226296
rect 208176 226256 257436 226284
rect 208176 226244 208182 226256
rect 257430 226244 257436 226256
rect 257488 226244 257494 226296
rect 266998 226244 267004 226296
rect 267056 226284 267062 226296
rect 274450 226284 274456 226296
rect 267056 226256 274456 226284
rect 267056 226244 267062 226256
rect 274450 226244 274456 226256
rect 274508 226244 274514 226296
rect 286318 226244 286324 226296
rect 286376 226284 286382 226296
rect 289906 226284 289912 226296
rect 286376 226256 289912 226284
rect 286376 226244 286382 226256
rect 289906 226244 289912 226256
rect 289964 226244 289970 226296
rect 291010 226244 291016 226296
rect 291068 226284 291074 226296
rect 322106 226284 322112 226296
rect 291068 226256 322112 226284
rect 291068 226244 291074 226256
rect 322106 226244 322112 226256
rect 322164 226244 322170 226296
rect 458634 226244 458640 226296
rect 458692 226284 458698 226296
rect 462958 226284 462964 226296
rect 458692 226256 462964 226284
rect 458692 226244 458698 226256
rect 462958 226244 462964 226256
rect 463016 226244 463022 226296
rect 672604 226160 672656 226166
rect 127434 226108 127440 226160
rect 127492 226148 127498 226160
rect 142108 226148 142114 226160
rect 127492 226120 142114 226148
rect 127492 226108 127498 226120
rect 142108 226108 142114 226120
rect 142166 226108 142172 226160
rect 142246 226108 142252 226160
rect 142304 226148 142310 226160
rect 209406 226148 209412 226160
rect 142304 226120 209412 226148
rect 142304 226108 142310 226120
rect 209406 226108 209412 226120
rect 209464 226108 209470 226160
rect 209682 226108 209688 226160
rect 209740 226148 209746 226160
rect 259638 226148 259644 226160
rect 209740 226120 259644 226148
rect 209740 226108 209746 226120
rect 259638 226108 259644 226120
rect 259696 226108 259702 226160
rect 261846 226108 261852 226160
rect 261904 226148 261910 226160
rect 300854 226148 300860 226160
rect 261904 226120 300860 226148
rect 261904 226108 261910 226120
rect 300854 226108 300860 226120
rect 300912 226108 300918 226160
rect 309042 226108 309048 226160
rect 309100 226148 309106 226160
rect 336274 226148 336280 226160
rect 309100 226120 336280 226148
rect 309100 226108 309106 226120
rect 336274 226108 336280 226120
rect 336332 226108 336338 226160
rect 528554 226108 528560 226160
rect 528612 226148 528618 226160
rect 542630 226148 542636 226160
rect 528612 226120 542636 226148
rect 528612 226108 528618 226120
rect 542630 226108 542636 226120
rect 542688 226108 542694 226160
rect 672604 226102 672656 226108
rect 66162 225972 66168 226024
rect 66220 226012 66226 226024
rect 142614 226012 142620 226024
rect 66220 225984 142620 226012
rect 66220 225972 66226 225984
rect 142614 225972 142620 225984
rect 142672 225972 142678 226024
rect 142798 225972 142804 226024
rect 142856 226012 142862 226024
rect 147582 226012 147588 226024
rect 142856 225984 147588 226012
rect 142856 225972 142862 225984
rect 147582 225972 147588 225984
rect 147640 225972 147646 226024
rect 147766 225972 147772 226024
rect 147824 226012 147830 226024
rect 147824 225984 157104 226012
rect 147824 225972 147830 225984
rect 83458 225836 83464 225888
rect 83516 225876 83522 225888
rect 155494 225876 155500 225888
rect 83516 225848 155500 225876
rect 83516 225836 83522 225848
rect 155494 225836 155500 225848
rect 155552 225836 155558 225888
rect 157076 225808 157104 225984
rect 157334 225972 157340 226024
rect 157392 226012 157398 226024
rect 217134 226012 217140 226024
rect 157392 225984 217140 226012
rect 157392 225972 157398 225984
rect 217134 225972 217140 225984
rect 217192 225972 217198 226024
rect 222010 225972 222016 226024
rect 222068 226012 222074 226024
rect 269942 226012 269948 226024
rect 222068 225984 269948 226012
rect 222068 225972 222074 225984
rect 269942 225972 269948 225984
rect 270000 225972 270006 226024
rect 278406 225972 278412 226024
rect 278464 226012 278470 226024
rect 313274 226012 313280 226024
rect 278464 225984 313280 226012
rect 278464 225972 278470 225984
rect 313274 225972 313280 225984
rect 313332 225972 313338 226024
rect 329742 225972 329748 226024
rect 329800 226012 329806 226024
rect 353662 226012 353668 226024
rect 329800 225984 353668 226012
rect 329800 225972 329806 225984
rect 353662 225972 353668 225984
rect 353720 225972 353726 226024
rect 354582 225972 354588 226024
rect 354640 226012 354646 226024
rect 372338 226012 372344 226024
rect 354640 225984 372344 226012
rect 354640 225972 354646 225984
rect 372338 225972 372344 225984
rect 372396 225972 372402 226024
rect 498102 225972 498108 226024
rect 498160 226012 498166 226024
rect 514294 226012 514300 226024
rect 498160 225984 514300 226012
rect 498160 225972 498166 225984
rect 514294 225972 514300 225984
rect 514352 225972 514358 226024
rect 516594 225972 516600 226024
rect 516652 226012 516658 226024
rect 538674 226012 538680 226024
rect 516652 225984 538680 226012
rect 516652 225972 516658 225984
rect 538674 225972 538680 225984
rect 538732 225972 538738 226024
rect 672494 225956 672546 225962
rect 672494 225898 672546 225904
rect 197998 225836 198004 225888
rect 198056 225876 198062 225888
rect 249334 225876 249340 225888
rect 198056 225848 249340 225876
rect 198056 225836 198062 225848
rect 249334 225836 249340 225848
rect 249392 225836 249398 225888
rect 252462 225836 252468 225888
rect 252520 225876 252526 225888
rect 293126 225876 293132 225888
rect 252520 225848 293132 225876
rect 252520 225836 252526 225848
rect 293126 225836 293132 225848
rect 293184 225836 293190 225888
rect 296438 225836 296444 225888
rect 296496 225876 296502 225888
rect 327534 225876 327540 225888
rect 296496 225848 327540 225876
rect 296496 225836 296502 225848
rect 327534 225836 327540 225848
rect 327592 225836 327598 225888
rect 332226 225836 332232 225888
rect 332284 225876 332290 225888
rect 357526 225876 357532 225888
rect 332284 225848 357532 225876
rect 332284 225836 332290 225848
rect 357526 225836 357532 225848
rect 357584 225836 357590 225888
rect 373810 225836 373816 225888
rect 373868 225876 373874 225888
rect 377674 225876 377680 225888
rect 373868 225848 377680 225876
rect 373868 225836 373874 225848
rect 377674 225836 377680 225848
rect 377732 225836 377738 225888
rect 377858 225836 377864 225888
rect 377916 225876 377922 225888
rect 390370 225876 390376 225888
rect 377916 225848 390376 225876
rect 377916 225836 377922 225848
rect 390370 225836 390376 225848
rect 390428 225836 390434 225888
rect 394326 225836 394332 225888
rect 394384 225876 394390 225888
rect 403250 225876 403256 225888
rect 394384 225848 403256 225876
rect 394384 225836 394390 225848
rect 403250 225836 403256 225848
rect 403308 225836 403314 225888
rect 483750 225836 483756 225888
rect 483808 225876 483814 225888
rect 497274 225876 497280 225888
rect 483808 225848 497280 225876
rect 483808 225836 483814 225848
rect 497274 225836 497280 225848
rect 497332 225836 497338 225888
rect 501138 225836 501144 225888
rect 501196 225876 501202 225888
rect 519262 225876 519268 225888
rect 501196 225848 519268 225876
rect 501196 225836 501202 225848
rect 519262 225836 519268 225848
rect 519320 225836 519326 225888
rect 521746 225836 521752 225888
rect 521804 225876 521810 225888
rect 545758 225876 545764 225888
rect 521804 225848 545764 225876
rect 521804 225836 521810 225848
rect 545758 225836 545764 225848
rect 545816 225836 545822 225888
rect 558178 225836 558184 225888
rect 558236 225876 558242 225888
rect 572254 225876 572260 225888
rect 558236 225848 572260 225876
rect 558236 225836 558242 225848
rect 572254 225836 572260 225848
rect 572312 225836 572318 225888
rect 672166 225836 672172 225888
rect 672224 225876 672230 225888
rect 672224 225848 672406 225876
rect 672224 225836 672230 225848
rect 157076 225780 164234 225808
rect 76558 225700 76564 225752
rect 76616 225740 76622 225752
rect 164206 225740 164234 225780
rect 184014 225740 184020 225752
rect 76616 225712 147904 225740
rect 164206 225712 184020 225740
rect 76616 225700 76622 225712
rect 147876 225672 147904 225712
rect 184014 225700 184020 225712
rect 184072 225700 184078 225752
rect 184198 225700 184204 225752
rect 184256 225740 184262 225752
rect 212626 225740 212632 225752
rect 184256 225712 212632 225740
rect 184256 225700 184262 225712
rect 212626 225700 212632 225712
rect 212684 225700 212690 225752
rect 237282 225700 237288 225752
rect 237340 225740 237346 225752
rect 240318 225740 240324 225752
rect 237340 225712 240324 225740
rect 237340 225700 237346 225712
rect 240318 225700 240324 225712
rect 240376 225700 240382 225752
rect 255038 225700 255044 225752
rect 255096 225740 255102 225752
rect 296990 225740 296996 225752
rect 255096 225712 296996 225740
rect 255096 225700 255102 225712
rect 296990 225700 296996 225712
rect 297048 225700 297054 225752
rect 315666 225700 315672 225752
rect 315724 225740 315730 225752
rect 344646 225740 344652 225752
rect 315724 225712 344652 225740
rect 315724 225700 315730 225712
rect 344646 225700 344652 225712
rect 344704 225700 344710 225752
rect 352926 225700 352932 225752
rect 352984 225740 352990 225752
rect 371602 225740 371608 225752
rect 352984 225712 371608 225740
rect 352984 225700 352990 225712
rect 371602 225700 371608 225712
rect 371660 225700 371666 225752
rect 371786 225700 371792 225752
rect 371844 225740 371850 225752
rect 382734 225740 382740 225752
rect 371844 225712 382740 225740
rect 371844 225700 371850 225712
rect 382734 225700 382740 225712
rect 382792 225700 382798 225752
rect 382918 225700 382924 225752
rect 382976 225740 382982 225752
rect 396166 225740 396172 225752
rect 382976 225712 396172 225740
rect 382976 225700 382982 225712
rect 396166 225700 396172 225712
rect 396224 225700 396230 225752
rect 488902 225700 488908 225752
rect 488960 225740 488966 225752
rect 503622 225740 503628 225752
rect 488960 225712 503628 225740
rect 488960 225700 488966 225712
rect 503622 225700 503628 225712
rect 503680 225700 503686 225752
rect 508866 225700 508872 225752
rect 508924 225740 508930 225752
rect 529198 225740 529204 225752
rect 508924 225712 529204 225740
rect 508924 225700 508930 225712
rect 529198 225700 529204 225712
rect 529256 225700 529262 225752
rect 535914 225700 535920 225752
rect 535972 225740 535978 225752
rect 563974 225740 563980 225752
rect 535972 225712 563980 225740
rect 535972 225700 535978 225712
rect 563974 225700 563980 225712
rect 564032 225700 564038 225752
rect 156598 225672 156604 225684
rect 147876 225644 156604 225672
rect 156598 225632 156604 225644
rect 156656 225632 156662 225684
rect 72418 225564 72424 225616
rect 72476 225604 72482 225616
rect 142108 225604 142114 225616
rect 72476 225576 142114 225604
rect 72476 225564 72482 225576
rect 142108 225564 142114 225576
rect 142166 225564 142172 225616
rect 142246 225564 142252 225616
rect 142304 225604 142310 225616
rect 147674 225604 147680 225616
rect 142304 225576 147680 225604
rect 142304 225564 142310 225576
rect 147674 225564 147680 225576
rect 147732 225564 147738 225616
rect 157334 225564 157340 225616
rect 157392 225604 157398 225616
rect 214374 225604 214380 225616
rect 157392 225576 214380 225604
rect 157392 225564 157398 225576
rect 214374 225564 214380 225576
rect 214432 225564 214438 225616
rect 215202 225564 215208 225616
rect 215260 225604 215266 225616
rect 266078 225604 266084 225616
rect 215260 225576 266084 225604
rect 215260 225564 215266 225576
rect 266078 225564 266084 225576
rect 266136 225564 266142 225616
rect 270034 225564 270040 225616
rect 270092 225604 270098 225616
rect 282638 225604 282644 225616
rect 270092 225576 282644 225604
rect 270092 225564 270098 225576
rect 282638 225564 282644 225576
rect 282696 225564 282702 225616
rect 284110 225564 284116 225616
rect 284168 225604 284174 225616
rect 320174 225604 320180 225616
rect 284168 225576 320180 225604
rect 284168 225564 284174 225576
rect 320174 225564 320180 225576
rect 320232 225564 320238 225616
rect 321370 225564 321376 225616
rect 321428 225604 321434 225616
rect 346578 225604 346584 225616
rect 321428 225576 346584 225604
rect 321428 225564 321434 225576
rect 346578 225564 346584 225576
rect 346636 225564 346642 225616
rect 347038 225564 347044 225616
rect 347096 225604 347102 225616
rect 367830 225604 367836 225616
rect 347096 225576 367836 225604
rect 347096 225564 347102 225576
rect 367830 225564 367836 225576
rect 367888 225564 367894 225616
rect 372522 225564 372528 225616
rect 372580 225604 372586 225616
rect 387426 225604 387432 225616
rect 372580 225576 387432 225604
rect 372580 225564 372586 225576
rect 387426 225564 387432 225576
rect 387484 225564 387490 225616
rect 390186 225564 390192 225616
rect 390244 225604 390250 225616
rect 401962 225604 401968 225616
rect 390244 225576 401968 225604
rect 390244 225564 390250 225576
rect 401962 225564 401968 225576
rect 402020 225564 402026 225616
rect 410978 225564 410984 225616
rect 411036 225604 411042 225616
rect 416130 225604 416136 225616
rect 411036 225576 416136 225604
rect 411036 225564 411042 225576
rect 416130 225564 416136 225576
rect 416188 225564 416194 225616
rect 467650 225564 467656 225616
rect 467708 225604 467714 225616
rect 476574 225604 476580 225616
rect 467708 225576 476580 225604
rect 467708 225564 467714 225576
rect 476574 225564 476580 225576
rect 476632 225564 476638 225616
rect 477310 225564 477316 225616
rect 477368 225604 477374 225616
rect 488810 225604 488816 225616
rect 477368 225576 488816 225604
rect 477368 225564 477374 225576
rect 488810 225564 488816 225576
rect 488868 225564 488874 225616
rect 494054 225564 494060 225616
rect 494112 225604 494118 225616
rect 509694 225604 509700 225616
rect 494112 225576 509700 225604
rect 494112 225564 494118 225576
rect 509694 225564 509700 225576
rect 509752 225564 509758 225616
rect 510154 225564 510160 225616
rect 510212 225604 510218 225616
rect 530946 225604 530952 225616
rect 510212 225576 530952 225604
rect 510212 225564 510218 225576
rect 530946 225564 530952 225576
rect 531004 225564 531010 225616
rect 531406 225564 531412 225616
rect 531464 225604 531470 225616
rect 558270 225604 558276 225616
rect 531464 225576 558276 225604
rect 531464 225564 531470 225576
rect 558270 225564 558276 225576
rect 558328 225564 558334 225616
rect 672264 225548 672316 225554
rect 672264 225490 672316 225496
rect 110138 225428 110144 225480
rect 110196 225468 110202 225480
rect 127434 225468 127440 225480
rect 110196 225440 127440 225468
rect 110196 225428 110202 225440
rect 127434 225428 127440 225440
rect 127492 225428 127498 225480
rect 193582 225468 193588 225480
rect 127636 225440 193588 225468
rect 122558 225156 122564 225208
rect 122616 225196 122622 225208
rect 127636 225196 127664 225440
rect 193582 225428 193588 225440
rect 193640 225428 193646 225480
rect 193766 225428 193772 225480
rect 193824 225468 193830 225480
rect 244182 225468 244188 225480
rect 193824 225440 244188 225468
rect 193824 225428 193830 225440
rect 244182 225428 244188 225440
rect 244240 225428 244246 225480
rect 672156 225412 672208 225418
rect 463142 225360 463148 225412
rect 463200 225400 463206 225412
rect 467282 225400 467288 225412
rect 463200 225372 467288 225400
rect 463200 225360 463206 225372
rect 467282 225360 467288 225372
rect 467340 225360 467346 225412
rect 672156 225354 672208 225360
rect 196158 225332 196164 225344
rect 122616 225168 127664 225196
rect 127728 225304 196164 225332
rect 122616 225156 122622 225168
rect 125226 225020 125232 225072
rect 125284 225060 125290 225072
rect 127728 225060 127756 225304
rect 196158 225292 196164 225304
rect 196216 225292 196222 225344
rect 196618 225292 196624 225344
rect 196676 225332 196682 225344
rect 236454 225332 236460 225344
rect 196676 225304 236460 225332
rect 196676 225292 196682 225304
rect 236454 225292 236460 225304
rect 236512 225292 236518 225344
rect 241146 225292 241152 225344
rect 241204 225332 241210 225344
rect 286686 225332 286692 225344
rect 241204 225304 286692 225332
rect 241204 225292 241210 225304
rect 286686 225292 286692 225304
rect 286744 225292 286750 225344
rect 563026 225304 572714 225332
rect 129366 225156 129372 225208
rect 129424 225196 129430 225208
rect 199102 225196 199108 225208
rect 129424 225168 199108 225196
rect 129424 225156 129430 225168
rect 199102 225156 199108 225168
rect 199160 225156 199166 225208
rect 242710 225156 242716 225208
rect 242768 225196 242774 225208
rect 285030 225196 285036 225208
rect 242768 225168 285036 225196
rect 242768 225156 242774 225168
rect 285030 225156 285036 225168
rect 285088 225156 285094 225208
rect 125284 225032 127756 225060
rect 125284 225020 125290 225032
rect 132402 225020 132408 225072
rect 132460 225060 132466 225072
rect 201678 225060 201684 225072
rect 132460 225032 201684 225060
rect 132460 225020 132466 225032
rect 201678 225020 201684 225032
rect 201736 225020 201742 225072
rect 202230 225020 202236 225072
rect 202288 225060 202294 225072
rect 254486 225060 254492 225072
rect 202288 225032 254492 225060
rect 202288 225020 202294 225032
rect 254486 225020 254492 225032
rect 254544 225020 254550 225072
rect 297266 224952 297272 225004
rect 297324 224992 297330 225004
rect 305362 224992 305368 225004
rect 297324 224964 305368 224992
rect 297324 224952 297330 224964
rect 305362 224952 305368 224964
rect 305420 224952 305426 225004
rect 327718 224952 327724 225004
rect 327776 224992 327782 225004
rect 332042 224992 332048 225004
rect 327776 224964 332048 224992
rect 327776 224952 327782 224964
rect 332042 224952 332048 224964
rect 332100 224952 332106 225004
rect 369118 224952 369124 225004
rect 369176 224992 369182 225004
rect 373626 224992 373632 225004
rect 369176 224964 373632 224992
rect 369176 224952 369182 224964
rect 373626 224952 373632 224964
rect 373684 224952 373690 225004
rect 404170 224952 404176 225004
rect 404228 224992 404234 225004
rect 410610 224992 410616 225004
rect 404228 224964 410616 224992
rect 404228 224952 404234 224964
rect 410610 224952 410616 224964
rect 410668 224952 410674 225004
rect 416498 224952 416504 225004
rect 416556 224992 416562 225004
rect 422202 224992 422208 225004
rect 416556 224964 422208 224992
rect 416556 224952 416562 224964
rect 422202 224952 422208 224964
rect 422260 224952 422266 225004
rect 493686 224952 493692 225004
rect 493744 224992 493750 225004
rect 494698 224992 494704 225004
rect 493744 224964 494704 224992
rect 493744 224952 493750 224964
rect 494698 224952 494704 224964
rect 494756 224952 494762 225004
rect 495158 224952 495164 225004
rect 495216 224992 495222 225004
rect 563026 224992 563054 225304
rect 567010 225088 567016 225140
rect 567068 225128 567074 225140
rect 571426 225128 571432 225140
rect 567068 225100 571432 225128
rect 567068 225088 567074 225100
rect 571426 225088 571432 225100
rect 571484 225088 571490 225140
rect 495216 224964 563054 224992
rect 495216 224952 495222 224964
rect 563698 224952 563704 225004
rect 563756 224992 563762 225004
rect 572686 224992 572714 225304
rect 672034 225276 672086 225282
rect 672034 225218 672086 225224
rect 666462 225156 666468 225208
rect 666520 225196 666526 225208
rect 666520 225168 669314 225196
rect 666520 225156 666526 225168
rect 669286 225060 669314 225168
rect 669286 225032 671968 225060
rect 630858 224992 630864 225004
rect 563756 224964 567148 224992
rect 572686 224964 630864 224992
rect 563756 224952 563762 224964
rect 96062 224884 96068 224936
rect 96120 224924 96126 224936
rect 172974 224924 172980 224936
rect 96120 224896 172980 224924
rect 96120 224884 96126 224896
rect 172974 224884 172980 224896
rect 173032 224884 173038 224936
rect 174906 224884 174912 224936
rect 174964 224924 174970 224936
rect 185578 224924 185584 224936
rect 174964 224896 185584 224924
rect 174964 224884 174970 224896
rect 185578 224884 185584 224896
rect 185636 224884 185642 224936
rect 185762 224884 185768 224936
rect 185820 224924 185826 224936
rect 195238 224924 195244 224936
rect 185820 224896 195244 224924
rect 185820 224884 185826 224896
rect 195238 224884 195244 224896
rect 195296 224884 195302 224936
rect 195606 224884 195612 224936
rect 195664 224924 195670 224936
rect 242894 224924 242900 224936
rect 195664 224896 242900 224924
rect 195664 224884 195670 224896
rect 242894 224884 242900 224896
rect 242952 224884 242958 224936
rect 266170 224884 266176 224936
rect 266228 224924 266234 224936
rect 567120 224924 567148 224964
rect 630858 224952 630864 224964
rect 630916 224952 630922 225004
rect 568942 224924 568948 224936
rect 266228 224896 296714 224924
rect 567120 224896 568948 224924
rect 266228 224884 266234 224896
rect 296686 224856 296714 224896
rect 568942 224884 568948 224896
rect 569000 224884 569006 224936
rect 303430 224856 303436 224868
rect 296686 224828 303436 224856
rect 303430 224816 303436 224828
rect 303488 224816 303494 224868
rect 549254 224816 549260 224868
rect 549312 224856 549318 224868
rect 554774 224856 554780 224868
rect 549312 224828 554780 224856
rect 549312 224816 549318 224828
rect 554774 224816 554780 224828
rect 554832 224816 554838 224868
rect 610986 224816 610992 224868
rect 611044 224856 611050 224868
rect 614942 224856 614948 224868
rect 611044 224828 614948 224856
rect 611044 224816 611050 224828
rect 614942 224816 614948 224828
rect 615000 224816 615006 224868
rect 670712 224828 671846 224856
rect 102042 224748 102048 224800
rect 102100 224788 102106 224800
rect 178494 224788 178500 224800
rect 102100 224760 178500 224788
rect 102100 224748 102106 224760
rect 178494 224748 178500 224760
rect 178552 224748 178558 224800
rect 178678 224748 178684 224800
rect 178736 224788 178742 224800
rect 204530 224788 204536 224800
rect 178736 224760 204536 224788
rect 178736 224748 178742 224760
rect 204530 224748 204536 224760
rect 204588 224748 204594 224800
rect 204714 224748 204720 224800
rect 204772 224788 204778 224800
rect 204772 224760 224264 224788
rect 204772 224748 204778 224760
rect 79962 224612 79968 224664
rect 80020 224652 80026 224664
rect 160462 224652 160468 224664
rect 80020 224624 160468 224652
rect 80020 224612 80026 224624
rect 160462 224612 160468 224624
rect 160520 224612 160526 224664
rect 162762 224612 162768 224664
rect 162820 224652 162826 224664
rect 224034 224652 224040 224664
rect 162820 224624 224040 224652
rect 162820 224612 162826 224624
rect 224034 224612 224040 224624
rect 224092 224612 224098 224664
rect 224236 224652 224264 224760
rect 224586 224748 224592 224800
rect 224644 224788 224650 224800
rect 224644 224760 238754 224788
rect 224644 224748 224650 224760
rect 237742 224652 237748 224664
rect 224236 224624 237748 224652
rect 237742 224612 237748 224624
rect 237800 224612 237806 224664
rect 238726 224652 238754 224760
rect 245286 224748 245292 224800
rect 245344 224788 245350 224800
rect 287974 224788 287980 224800
rect 245344 224760 287980 224788
rect 245344 224748 245350 224760
rect 287974 224748 287980 224760
rect 288032 224748 288038 224800
rect 311526 224748 311532 224800
rect 311584 224788 311590 224800
rect 338850 224788 338856 224800
rect 311584 224760 338856 224788
rect 311584 224748 311590 224760
rect 338850 224748 338856 224760
rect 338908 224748 338914 224800
rect 462498 224748 462504 224800
rect 462556 224788 462562 224800
rect 469306 224788 469312 224800
rect 462556 224760 469312 224788
rect 462556 224748 462562 224760
rect 469306 224748 469312 224760
rect 469364 224748 469370 224800
rect 506934 224748 506940 224800
rect 506992 224788 506998 224800
rect 526714 224788 526720 224800
rect 506992 224760 526720 224788
rect 506992 224748 506998 224760
rect 526714 224748 526720 224760
rect 526772 224748 526778 224800
rect 529934 224748 529940 224800
rect 529992 224788 529998 224800
rect 549070 224788 549076 224800
rect 529992 224760 549076 224788
rect 529992 224748 529998 224760
rect 549070 224748 549076 224760
rect 549128 224748 549134 224800
rect 554958 224748 554964 224800
rect 555016 224788 555022 224800
rect 555786 224788 555792 224800
rect 555016 224760 555792 224788
rect 555016 224748 555022 224760
rect 555786 224748 555792 224760
rect 555844 224748 555850 224800
rect 555970 224748 555976 224800
rect 556028 224788 556034 224800
rect 562134 224788 562140 224800
rect 556028 224760 562140 224788
rect 556028 224748 556034 224760
rect 562134 224748 562140 224760
rect 562192 224748 562198 224800
rect 562318 224748 562324 224800
rect 562376 224788 562382 224800
rect 567010 224788 567016 224800
rect 562376 224760 567016 224788
rect 562376 224748 562382 224760
rect 567010 224748 567016 224760
rect 567068 224748 567074 224800
rect 567838 224748 567844 224800
rect 567896 224788 567902 224800
rect 610802 224788 610808 224800
rect 567896 224760 610808 224788
rect 567896 224748 567902 224760
rect 610802 224748 610808 224760
rect 610860 224748 610866 224800
rect 670510 224748 670516 224800
rect 670568 224788 670574 224800
rect 670712 224788 670740 224828
rect 670568 224760 670740 224788
rect 670568 224748 670574 224760
rect 270586 224652 270592 224664
rect 238726 224624 270592 224652
rect 270586 224612 270592 224624
rect 270644 224612 270650 224664
rect 274266 224612 274272 224664
rect 274324 224652 274330 224664
rect 312446 224652 312452 224664
rect 274324 224624 312452 224652
rect 274324 224612 274330 224624
rect 312446 224612 312452 224624
rect 312504 224612 312510 224664
rect 319990 224612 319996 224664
rect 320048 224652 320054 224664
rect 345934 224652 345940 224664
rect 320048 224624 345940 224652
rect 320048 224612 320054 224624
rect 345934 224612 345940 224624
rect 345992 224612 345998 224664
rect 346210 224612 346216 224664
rect 346268 224652 346274 224664
rect 366542 224652 366548 224664
rect 346268 224624 366548 224652
rect 346268 224612 346274 224624
rect 366542 224612 366548 224624
rect 366600 224612 366606 224664
rect 505186 224612 505192 224664
rect 505244 224652 505250 224664
rect 610434 224652 610440 224664
rect 505244 224624 610440 224652
rect 505244 224612 505250 224624
rect 610434 224612 610440 224624
rect 610492 224612 610498 224664
rect 610618 224612 610624 224664
rect 610676 224652 610682 224664
rect 616046 224652 616052 224664
rect 610676 224624 616052 224652
rect 610676 224612 610682 224624
rect 616046 224612 616052 224624
rect 616104 224612 616110 224664
rect 668578 224612 668584 224664
rect 668636 224652 668642 224664
rect 668636 224624 671738 224652
rect 668636 224612 668642 224624
rect 85482 224476 85488 224528
rect 85540 224516 85546 224528
rect 165614 224516 165620 224528
rect 85540 224488 165620 224516
rect 85540 224476 85546 224488
rect 165614 224476 165620 224488
rect 165672 224476 165678 224528
rect 179322 224476 179328 224528
rect 179380 224516 179386 224528
rect 185394 224516 185400 224528
rect 179380 224488 185400 224516
rect 179380 224476 179386 224488
rect 185394 224476 185400 224488
rect 185452 224476 185458 224528
rect 185578 224476 185584 224528
rect 185636 224516 185642 224528
rect 235166 224516 235172 224528
rect 185636 224488 235172 224516
rect 185636 224476 185642 224488
rect 235166 224476 235172 224488
rect 235224 224476 235230 224528
rect 251082 224476 251088 224528
rect 251140 224516 251146 224528
rect 294414 224516 294420 224528
rect 251140 224488 294420 224516
rect 251140 224476 251146 224488
rect 294414 224476 294420 224488
rect 294472 224476 294478 224528
rect 299290 224476 299296 224528
rect 299348 224516 299354 224528
rect 331766 224516 331772 224528
rect 299348 224488 331772 224516
rect 299348 224476 299354 224488
rect 331766 224476 331772 224488
rect 331824 224476 331830 224528
rect 335170 224476 335176 224528
rect 335228 224516 335234 224528
rect 356882 224516 356888 224528
rect 335228 224488 356888 224516
rect 335228 224476 335234 224488
rect 356882 224476 356888 224488
rect 356940 224476 356946 224528
rect 366726 224476 366732 224528
rect 366784 224516 366790 224528
rect 381630 224516 381636 224528
rect 366784 224488 381636 224516
rect 366784 224476 366790 224488
rect 381630 224476 381636 224488
rect 381688 224476 381694 224528
rect 456058 224476 456064 224528
rect 456116 224516 456122 224528
rect 459738 224516 459744 224528
rect 456116 224488 459744 224516
rect 456116 224476 456122 224488
rect 459738 224476 459744 224488
rect 459796 224476 459802 224528
rect 491294 224476 491300 224528
rect 491352 224516 491358 224528
rect 506014 224516 506020 224528
rect 491352 224488 506020 224516
rect 491352 224476 491358 224488
rect 506014 224476 506020 224488
rect 506072 224476 506078 224528
rect 515950 224476 515956 224528
rect 516008 224516 516014 224528
rect 538306 224516 538312 224528
rect 516008 224488 538312 224516
rect 516008 224476 516014 224488
rect 538306 224476 538312 224488
rect 538364 224476 538370 224528
rect 538858 224476 538864 224528
rect 538916 224516 538922 224528
rect 538916 224488 552704 224516
rect 538916 224476 538922 224488
rect 73706 224340 73712 224392
rect 73764 224380 73770 224392
rect 155310 224380 155316 224392
rect 73764 224352 155316 224380
rect 73764 224340 73770 224352
rect 155310 224340 155316 224352
rect 155368 224340 155374 224392
rect 157242 224340 157248 224392
rect 157300 224380 157306 224392
rect 161934 224380 161940 224392
rect 157300 224352 161940 224380
rect 157300 224340 157306 224352
rect 161934 224340 161940 224352
rect 161992 224340 161998 224392
rect 165522 224340 165528 224392
rect 165580 224380 165586 224392
rect 227438 224380 227444 224392
rect 165580 224352 227444 224380
rect 165580 224340 165586 224352
rect 227438 224340 227444 224352
rect 227496 224340 227502 224392
rect 228726 224340 228732 224392
rect 228784 224380 228790 224392
rect 274910 224380 274916 224392
rect 228784 224352 274916 224380
rect 228784 224340 228790 224352
rect 274910 224340 274916 224352
rect 274968 224340 274974 224392
rect 275094 224340 275100 224392
rect 275152 224380 275158 224392
rect 311158 224380 311164 224392
rect 275152 224352 311164 224380
rect 275152 224340 275158 224352
rect 311158 224340 311164 224352
rect 311216 224340 311222 224392
rect 319806 224340 319812 224392
rect 319864 224380 319870 224392
rect 347222 224380 347228 224392
rect 319864 224352 347228 224380
rect 319864 224340 319870 224352
rect 347222 224340 347228 224352
rect 347280 224340 347286 224392
rect 361206 224340 361212 224392
rect 361264 224380 361270 224392
rect 377490 224380 377496 224392
rect 361264 224352 377496 224380
rect 361264 224340 361270 224352
rect 377490 224340 377496 224352
rect 377548 224340 377554 224392
rect 387702 224340 387708 224392
rect 387760 224380 387766 224392
rect 397822 224380 397828 224392
rect 387760 224352 397828 224380
rect 387760 224340 387766 224352
rect 397822 224340 397828 224352
rect 397880 224340 397886 224392
rect 480530 224340 480536 224392
rect 480588 224380 480594 224392
rect 492766 224380 492772 224392
rect 480588 224352 492772 224380
rect 480588 224340 480594 224352
rect 492766 224340 492772 224352
rect 492824 224340 492830 224392
rect 499206 224340 499212 224392
rect 499264 224380 499270 224392
rect 516778 224380 516784 224392
rect 499264 224352 516784 224380
rect 499264 224340 499270 224352
rect 516778 224340 516784 224352
rect 516836 224340 516842 224392
rect 525610 224340 525616 224392
rect 525668 224380 525674 224392
rect 550818 224380 550824 224392
rect 525668 224352 550824 224380
rect 525668 224340 525674 224352
rect 550818 224340 550824 224352
rect 550876 224340 550882 224392
rect 552676 224380 552704 224488
rect 552842 224476 552848 224528
rect 552900 224516 552906 224528
rect 625430 224516 625436 224528
rect 552900 224488 625436 224516
rect 552900 224476 552906 224488
rect 625430 224476 625436 224488
rect 625488 224476 625494 224528
rect 671596 224392 671648 224398
rect 552676 224352 556200 224380
rect 68922 224204 68928 224256
rect 68980 224244 68986 224256
rect 96246 224244 96252 224256
rect 68980 224216 96252 224244
rect 68980 224204 68986 224216
rect 96246 224204 96252 224216
rect 96304 224204 96310 224256
rect 167822 224244 167828 224256
rect 96448 224216 167828 224244
rect 89438 224068 89444 224120
rect 89496 224108 89502 224120
rect 96448 224108 96476 224216
rect 167822 224204 167828 224216
rect 167880 224204 167886 224256
rect 168282 224204 168288 224256
rect 168340 224244 168346 224256
rect 230014 224244 230020 224256
rect 168340 224216 230020 224244
rect 168340 224204 168346 224216
rect 230014 224204 230020 224216
rect 230072 224204 230078 224256
rect 231670 224204 231676 224256
rect 231728 224244 231734 224256
rect 278958 224244 278964 224256
rect 231728 224216 278964 224244
rect 231728 224204 231734 224216
rect 278958 224204 278964 224216
rect 279016 224204 279022 224256
rect 290826 224204 290832 224256
rect 290884 224244 290890 224256
rect 323670 224244 323676 224256
rect 290884 224216 323676 224244
rect 290884 224204 290890 224216
rect 323670 224204 323676 224216
rect 323728 224204 323734 224256
rect 323946 224204 323952 224256
rect 324004 224244 324010 224256
rect 334986 224244 334992 224256
rect 324004 224216 334992 224244
rect 324004 224204 324010 224216
rect 334986 224204 334992 224216
rect 335044 224204 335050 224256
rect 339402 224204 339408 224256
rect 339460 224244 339466 224256
rect 362310 224244 362316 224256
rect 339460 224216 362316 224244
rect 339460 224204 339466 224216
rect 362310 224204 362316 224216
rect 362368 224204 362374 224256
rect 363598 224204 363604 224256
rect 363656 224244 363662 224256
rect 368474 224244 368480 224256
rect 363656 224216 368480 224244
rect 363656 224204 363662 224216
rect 368474 224204 368480 224216
rect 368532 224204 368538 224256
rect 379238 224204 379244 224256
rect 379296 224244 379302 224256
rect 393590 224244 393596 224256
rect 379296 224216 393596 224244
rect 379296 224204 379302 224216
rect 393590 224204 393596 224216
rect 393648 224204 393654 224256
rect 394510 224204 394516 224256
rect 394568 224244 394574 224256
rect 404538 224244 404544 224256
rect 394568 224216 404544 224244
rect 394568 224204 394574 224216
rect 404538 224204 404544 224216
rect 404596 224204 404602 224256
rect 405550 224204 405556 224256
rect 405608 224244 405614 224256
rect 414198 224244 414204 224256
rect 405608 224216 414204 224244
rect 405608 224204 405614 224216
rect 414198 224204 414204 224216
rect 414256 224204 414262 224256
rect 470226 224204 470232 224256
rect 470284 224244 470290 224256
rect 480438 224244 480444 224256
rect 470284 224216 480444 224244
rect 470284 224204 470290 224216
rect 480438 224204 480444 224216
rect 480496 224204 480502 224256
rect 486602 224204 486608 224256
rect 486660 224244 486666 224256
rect 500402 224244 500408 224256
rect 486660 224216 500408 224244
rect 486660 224204 486666 224216
rect 500402 224204 500408 224216
rect 500460 224204 500466 224256
rect 504358 224204 504364 224256
rect 504416 224244 504422 224256
rect 523494 224244 523500 224256
rect 504416 224216 523500 224244
rect 504416 224204 504422 224216
rect 523494 224204 523500 224216
rect 523552 224204 523558 224256
rect 524414 224204 524420 224256
rect 524472 224244 524478 224256
rect 525058 224244 525064 224256
rect 524472 224216 525064 224244
rect 524472 224204 524478 224216
rect 525058 224204 525064 224216
rect 525116 224244 525122 224256
rect 538858 224244 538864 224256
rect 525116 224216 538864 224244
rect 525116 224204 525122 224216
rect 538858 224204 538864 224216
rect 538916 224204 538922 224256
rect 539318 224204 539324 224256
rect 539376 224244 539382 224256
rect 555970 224244 555976 224256
rect 539376 224216 555976 224244
rect 539376 224204 539382 224216
rect 555970 224204 555976 224216
rect 556028 224204 556034 224256
rect 556172 224244 556200 224352
rect 556338 224340 556344 224392
rect 556396 224380 556402 224392
rect 625246 224380 625252 224392
rect 556396 224352 625252 224380
rect 556396 224340 556402 224352
rect 625246 224340 625252 224352
rect 625304 224340 625310 224392
rect 671596 224334 671648 224340
rect 671482 224324 671534 224330
rect 671482 224266 671534 224272
rect 619634 224244 619640 224256
rect 556172 224216 619640 224244
rect 619634 224204 619640 224216
rect 619692 224204 619698 224256
rect 137968 224108 137974 224120
rect 89496 224080 96476 224108
rect 103486 224080 137974 224108
rect 89496 224068 89502 224080
rect 96246 223932 96252 223984
rect 96304 223972 96310 223984
rect 103486 223972 103514 224080
rect 137968 224068 137974 224080
rect 138026 224068 138032 224120
rect 138106 224068 138112 224120
rect 138164 224108 138170 224120
rect 194594 224108 194600 224120
rect 138164 224080 194600 224108
rect 138164 224068 138170 224080
rect 194594 224068 194600 224080
rect 194652 224068 194658 224120
rect 195238 224068 195244 224120
rect 195296 224108 195302 224120
rect 204714 224108 204720 224120
rect 195296 224080 204720 224108
rect 195296 224068 195302 224080
rect 204714 224068 204720 224080
rect 204772 224068 204778 224120
rect 204898 224068 204904 224120
rect 204956 224108 204962 224120
rect 250622 224108 250628 224120
rect 204956 224080 250628 224108
rect 204956 224068 204962 224080
rect 250622 224068 250628 224080
rect 250680 224068 250686 224120
rect 286686 224068 286692 224120
rect 286744 224108 286750 224120
rect 319530 224108 319536 224120
rect 286744 224080 319536 224108
rect 286744 224068 286750 224080
rect 319530 224068 319536 224080
rect 319588 224068 319594 224120
rect 358078 224068 358084 224120
rect 358136 224108 358142 224120
rect 363230 224108 363236 224120
rect 358136 224080 363236 224108
rect 358136 224068 358142 224080
rect 363230 224068 363236 224080
rect 363288 224068 363294 224120
rect 509694 224068 509700 224120
rect 509752 224108 509758 224120
rect 510154 224108 510160 224120
rect 509752 224080 510160 224108
rect 509752 224068 509758 224080
rect 510154 224068 510160 224080
rect 510212 224108 510218 224120
rect 610618 224108 610624 224120
rect 510212 224080 610624 224108
rect 510212 224068 510218 224080
rect 610618 224068 610624 224080
rect 610676 224068 610682 224120
rect 377398 224000 377404 224052
rect 377456 224040 377462 224052
rect 385862 224040 385868 224052
rect 377456 224012 385868 224040
rect 377456 224000 377462 224012
rect 385862 224000 385868 224012
rect 385920 224000 385926 224052
rect 610802 224000 610808 224052
rect 610860 224040 610866 224052
rect 623774 224040 623780 224052
rect 610860 224012 623780 224040
rect 610860 224000 610866 224012
rect 623774 224000 623780 224012
rect 623832 224000 623838 224052
rect 669222 224040 669228 224052
rect 669056 224012 669228 224040
rect 96304 223944 103514 223972
rect 96304 223932 96310 223944
rect 105998 223932 106004 223984
rect 106056 223972 106062 223984
rect 181070 223972 181076 223984
rect 106056 223944 181076 223972
rect 106056 223932 106062 223944
rect 181070 223932 181076 223944
rect 181128 223932 181134 223984
rect 201218 223932 201224 223984
rect 201276 223972 201282 223984
rect 255774 223972 255780 223984
rect 201276 223944 255780 223972
rect 201276 223932 201282 223944
rect 255774 223932 255780 223944
rect 255832 223932 255838 223984
rect 279418 223932 279424 223984
rect 279476 223972 279482 223984
rect 284754 223972 284760 223984
rect 279476 223944 284760 223972
rect 279476 223932 279482 223944
rect 284754 223932 284760 223944
rect 284812 223932 284818 223984
rect 519078 223932 519084 223984
rect 519136 223972 519142 223984
rect 519136 223944 528554 223972
rect 519136 223932 519142 223944
rect 108666 223796 108672 223848
rect 108724 223836 108730 223848
rect 183830 223836 183836 223848
rect 108724 223808 183836 223836
rect 108724 223796 108730 223808
rect 183830 223796 183836 223808
rect 183888 223796 183894 223848
rect 185946 223836 185952 223848
rect 184032 223808 185952 223836
rect 112806 223660 112812 223712
rect 112864 223700 112870 223712
rect 184032 223700 184060 223808
rect 185946 223796 185952 223808
rect 186004 223796 186010 223848
rect 186958 223796 186964 223848
rect 187016 223836 187022 223848
rect 217778 223836 217784 223848
rect 187016 223808 217784 223836
rect 187016 223796 187022 223808
rect 217778 223796 217784 223808
rect 217836 223796 217842 223848
rect 233142 223796 233148 223848
rect 233200 223836 233206 223848
rect 277670 223836 277676 223848
rect 233200 223808 277676 223836
rect 233200 223796 233206 223808
rect 277670 223796 277676 223808
rect 277728 223796 277734 223848
rect 528526 223768 528554 223944
rect 535270 223932 535276 223984
rect 535328 223972 535334 223984
rect 539318 223972 539324 223984
rect 535328 223944 539324 223972
rect 535328 223932 535334 223944
rect 539318 223932 539324 223944
rect 539376 223932 539382 223984
rect 539962 223864 539968 223916
rect 540020 223904 540026 223916
rect 622670 223904 622676 223916
rect 540020 223876 622676 223904
rect 540020 223864 540026 223876
rect 622670 223864 622676 223876
rect 622728 223864 622734 223916
rect 535086 223768 535092 223780
rect 528526 223740 535092 223768
rect 535086 223728 535092 223740
rect 535144 223768 535150 223780
rect 621566 223768 621572 223780
rect 535144 223740 621572 223768
rect 535144 223728 535150 223740
rect 621566 223728 621572 223740
rect 621624 223728 621630 223780
rect 112864 223672 184060 223700
rect 112864 223660 112870 223672
rect 184842 223660 184848 223712
rect 184900 223700 184906 223712
rect 195606 223700 195612 223712
rect 184900 223672 195612 223700
rect 184900 223660 184906 223672
rect 195606 223660 195612 223672
rect 195664 223660 195670 223712
rect 195882 223660 195888 223712
rect 195940 223700 195946 223712
rect 204898 223700 204904 223712
rect 195940 223672 204904 223700
rect 195940 223660 195946 223672
rect 204898 223660 204904 223672
rect 204956 223660 204962 223712
rect 238018 223660 238024 223712
rect 238076 223700 238082 223712
rect 266722 223700 266728 223712
rect 238076 223672 266728 223700
rect 238076 223660 238082 223672
rect 266722 223660 266728 223672
rect 266780 223660 266786 223712
rect 460566 223660 460572 223712
rect 460624 223700 460630 223712
rect 463142 223700 463148 223712
rect 460624 223672 463148 223700
rect 460624 223660 460630 223672
rect 463142 223660 463148 223672
rect 463200 223660 463206 223712
rect 520458 223592 520464 223644
rect 520516 223632 520522 223644
rect 543826 223632 543832 223644
rect 520516 223604 543832 223632
rect 520516 223592 520522 223604
rect 543826 223592 543832 223604
rect 543884 223592 543890 223644
rect 544010 223592 544016 223644
rect 544068 223632 544074 223644
rect 544930 223632 544936 223644
rect 544068 223604 544936 223632
rect 544068 223592 544074 223604
rect 544930 223592 544936 223604
rect 544988 223632 544994 223644
rect 567838 223632 567844 223644
rect 544988 223604 567844 223632
rect 544988 223592 544994 223604
rect 567838 223592 567844 223604
rect 567896 223592 567902 223644
rect 628742 223632 628748 223644
rect 568040 223604 628748 223632
rect 81342 223524 81348 223576
rect 81400 223564 81406 223576
rect 159818 223564 159824 223576
rect 81400 223536 159824 223564
rect 81400 223524 81406 223536
rect 159818 223524 159824 223536
rect 159876 223524 159882 223576
rect 162118 223524 162124 223576
rect 162176 223564 162182 223576
rect 186590 223564 186596 223576
rect 162176 223536 186596 223564
rect 162176 223524 162182 223536
rect 186590 223524 186596 223536
rect 186648 223524 186654 223576
rect 187326 223524 187332 223576
rect 187384 223564 187390 223576
rect 242250 223564 242256 223576
rect 187384 223536 242256 223564
rect 187384 223524 187390 223536
rect 242250 223524 242256 223536
rect 242308 223524 242314 223576
rect 250898 223524 250904 223576
rect 250956 223564 250962 223576
rect 291194 223564 291200 223576
rect 250956 223536 291200 223564
rect 250956 223524 250962 223536
rect 291194 223524 291200 223536
rect 291252 223524 291258 223576
rect 297910 223524 297916 223576
rect 297968 223564 297974 223576
rect 303246 223564 303252 223576
rect 297968 223536 303252 223564
rect 297968 223524 297974 223536
rect 303246 223524 303252 223536
rect 303304 223524 303310 223576
rect 307662 223524 307668 223576
rect 307720 223564 307726 223576
rect 335630 223564 335636 223576
rect 307720 223536 335636 223564
rect 307720 223524 307726 223536
rect 335630 223524 335636 223536
rect 335688 223524 335694 223576
rect 406746 223524 406752 223576
rect 406804 223564 406810 223576
rect 414842 223564 414848 223576
rect 406804 223536 414848 223564
rect 406804 223524 406810 223536
rect 414842 223524 414848 223536
rect 414900 223524 414906 223576
rect 454862 223524 454868 223576
rect 454920 223564 454926 223576
rect 460474 223564 460480 223576
rect 454920 223536 460480 223564
rect 454920 223524 454926 223536
rect 460474 223524 460480 223536
rect 460532 223524 460538 223576
rect 473446 223524 473452 223576
rect 473504 223564 473510 223576
rect 475562 223564 475568 223576
rect 473504 223536 475568 223564
rect 473504 223524 473510 223536
rect 475562 223524 475568 223536
rect 475620 223524 475626 223576
rect 342070 223496 342076 223508
rect 335832 223468 342076 223496
rect 75822 223388 75828 223440
rect 75880 223428 75886 223440
rect 154666 223428 154672 223440
rect 75880 223400 154672 223428
rect 75880 223388 75886 223400
rect 154666 223388 154672 223400
rect 154724 223388 154730 223440
rect 159358 223388 159364 223440
rect 159416 223428 159422 223440
rect 175918 223428 175924 223440
rect 159416 223400 175924 223428
rect 159416 223388 159422 223400
rect 175918 223388 175924 223400
rect 175976 223388 175982 223440
rect 184658 223388 184664 223440
rect 184716 223428 184722 223440
rect 239674 223428 239680 223440
rect 184716 223400 239680 223428
rect 184716 223388 184722 223400
rect 239674 223388 239680 223400
rect 239732 223388 239738 223440
rect 244090 223388 244096 223440
rect 244148 223428 244154 223440
rect 286042 223428 286048 223440
rect 244148 223400 286048 223428
rect 244148 223388 244154 223400
rect 286042 223388 286048 223400
rect 286100 223388 286106 223440
rect 312906 223388 312912 223440
rect 312964 223428 312970 223440
rect 312964 223400 335354 223428
rect 312964 223388 312970 223400
rect 335326 223360 335354 223400
rect 335832 223360 335860 223468
rect 342070 223456 342076 223468
rect 342128 223456 342134 223508
rect 566826 223456 566832 223508
rect 566884 223496 566890 223508
rect 568040 223496 568068 223604
rect 628742 223592 628748 223604
rect 628800 223592 628806 223644
rect 566884 223468 568068 223496
rect 566884 223456 566890 223468
rect 342806 223388 342812 223440
rect 342864 223428 342870 223440
rect 347866 223428 347872 223440
rect 342864 223400 347872 223428
rect 342864 223388 342870 223400
rect 347866 223388 347872 223400
rect 347924 223388 347930 223440
rect 493042 223388 493048 223440
rect 493100 223428 493106 223440
rect 508590 223428 508596 223440
rect 493100 223400 508596 223428
rect 493100 223388 493106 223400
rect 508590 223388 508596 223400
rect 508648 223388 508654 223440
rect 517514 223388 517520 223440
rect 517572 223428 517578 223440
rect 531498 223428 531504 223440
rect 517572 223400 531504 223428
rect 517572 223388 517578 223400
rect 531498 223388 531504 223400
rect 531556 223388 531562 223440
rect 534718 223388 534724 223440
rect 534776 223428 534782 223440
rect 547414 223428 547420 223440
rect 534776 223400 547420 223428
rect 534776 223388 534782 223400
rect 547414 223388 547420 223400
rect 547472 223388 547478 223440
rect 335326 223332 335860 223360
rect 335998 223320 336004 223372
rect 336056 223360 336062 223372
rect 342254 223360 342260 223372
rect 336056 223332 342260 223360
rect 336056 223320 336062 223332
rect 342254 223320 342260 223332
rect 342312 223320 342318 223372
rect 69566 223252 69572 223304
rect 69624 223292 69630 223304
rect 69624 223264 143028 223292
rect 69624 223252 69630 223264
rect 66898 223116 66904 223168
rect 66956 223156 66962 223168
rect 142522 223156 142528 223168
rect 66956 223128 142528 223156
rect 66956 223116 66962 223128
rect 142522 223116 142528 223128
rect 142580 223116 142586 223168
rect 143000 223156 143028 223264
rect 143810 223252 143816 223304
rect 143868 223292 143874 223304
rect 152090 223292 152096 223304
rect 143868 223264 152096 223292
rect 143868 223252 143874 223264
rect 152090 223252 152096 223264
rect 152148 223252 152154 223304
rect 156414 223252 156420 223304
rect 156472 223292 156478 223304
rect 162394 223292 162400 223304
rect 156472 223264 162400 223292
rect 156472 223252 156478 223264
rect 162394 223252 162400 223264
rect 162452 223252 162458 223304
rect 171778 223252 171784 223304
rect 171836 223292 171842 223304
rect 199746 223292 199752 223304
rect 171836 223264 199752 223292
rect 171836 223252 171842 223264
rect 199746 223252 199752 223264
rect 199804 223252 199810 223304
rect 204714 223252 204720 223304
rect 204772 223292 204778 223304
rect 204772 223264 209774 223292
rect 204772 223252 204778 223264
rect 143000 223128 143212 223156
rect 51902 222980 51908 223032
rect 51960 223020 51966 223032
rect 63126 223020 63132 223032
rect 51960 222992 63132 223020
rect 51960 222980 51966 222992
rect 63126 222980 63132 222992
rect 63184 222980 63190 223032
rect 71406 222980 71412 223032
rect 71464 223020 71470 223032
rect 139854 223020 139860 223032
rect 71464 222992 139860 223020
rect 71464 222980 71470 222992
rect 139854 222980 139860 222992
rect 139912 222980 139918 223032
rect 143184 223020 143212 223128
rect 143626 223116 143632 223168
rect 143684 223156 143690 223168
rect 146570 223156 146576 223168
rect 143684 223128 146576 223156
rect 143684 223116 143690 223128
rect 146570 223116 146576 223128
rect 146628 223116 146634 223168
rect 146754 223116 146760 223168
rect 146812 223156 146818 223168
rect 173342 223156 173348 223168
rect 146812 223128 173348 223156
rect 146812 223116 146818 223128
rect 173342 223116 173348 223128
rect 173400 223116 173406 223168
rect 173526 223116 173532 223168
rect 173584 223156 173590 223168
rect 185762 223156 185768 223168
rect 173584 223128 185768 223156
rect 173584 223116 173590 223128
rect 185762 223116 185768 223128
rect 185820 223116 185826 223168
rect 194502 223116 194508 223168
rect 194560 223156 194566 223168
rect 204898 223156 204904 223168
rect 194560 223128 204904 223156
rect 194560 223116 194566 223128
rect 204898 223116 204904 223128
rect 204956 223116 204962 223168
rect 209746 223156 209774 223264
rect 211430 223252 211436 223304
rect 211488 223292 211494 223304
rect 214374 223292 214380 223304
rect 211488 223264 214380 223292
rect 211488 223252 211494 223264
rect 214374 223252 214380 223264
rect 214432 223252 214438 223304
rect 219526 223292 219532 223304
rect 214576 223264 219532 223292
rect 211614 223156 211620 223168
rect 209746 223128 211620 223156
rect 211614 223116 211620 223128
rect 211672 223116 211678 223168
rect 149514 223020 149520 223032
rect 143184 222992 149520 223020
rect 149514 222980 149520 222992
rect 149572 222980 149578 223032
rect 166258 223020 166264 223032
rect 151786 222992 166264 223020
rect 62758 222844 62764 222896
rect 62816 222884 62822 222896
rect 143994 222884 144000 222896
rect 62816 222856 144000 222884
rect 62816 222844 62822 222856
rect 143994 222844 144000 222856
rect 144052 222844 144058 222896
rect 145098 222844 145104 222896
rect 145156 222884 145162 222896
rect 151786 222884 151814 222992
rect 166258 222980 166264 222992
rect 166316 222980 166322 223032
rect 166442 222980 166448 223032
rect 166500 223020 166506 223032
rect 214576 223020 214604 223264
rect 219526 223252 219532 223264
rect 219584 223252 219590 223304
rect 246850 223252 246856 223304
rect 246908 223292 246914 223304
rect 288618 223292 288624 223304
rect 246908 223264 288624 223292
rect 246908 223252 246914 223264
rect 288618 223252 288624 223264
rect 288676 223252 288682 223304
rect 289722 223252 289728 223304
rect 289780 223292 289786 223304
rect 297726 223292 297732 223304
rect 289780 223264 297732 223292
rect 289780 223252 289786 223264
rect 297726 223252 297732 223264
rect 297784 223252 297790 223304
rect 299106 223252 299112 223304
rect 299164 223292 299170 223304
rect 328546 223292 328552 223304
rect 299164 223264 328552 223292
rect 299164 223252 299170 223264
rect 328546 223252 328552 223264
rect 328604 223252 328610 223304
rect 347222 223252 347228 223304
rect 347280 223292 347286 223304
rect 357894 223292 357900 223304
rect 347280 223264 357900 223292
rect 347280 223252 347286 223264
rect 357894 223252 357900 223264
rect 357952 223252 357958 223304
rect 483106 223252 483112 223304
rect 483164 223292 483170 223304
rect 496078 223292 496084 223304
rect 483164 223264 496084 223292
rect 483164 223252 483170 223264
rect 496078 223252 496084 223264
rect 496136 223252 496142 223304
rect 514662 223252 514668 223304
rect 514720 223292 514726 223304
rect 536650 223292 536656 223304
rect 514720 223264 536656 223292
rect 514720 223252 514726 223264
rect 536650 223252 536656 223264
rect 536708 223252 536714 223304
rect 564618 223252 564624 223304
rect 564676 223292 564682 223304
rect 564676 223264 576854 223292
rect 564676 223252 564682 223264
rect 228082 223156 228088 223168
rect 166500 222992 214604 223020
rect 214668 223128 228088 223156
rect 166500 222980 166506 222992
rect 145156 222856 151814 222884
rect 145156 222844 145162 222856
rect 154206 222844 154212 222896
rect 154264 222884 154270 222896
rect 211430 222884 211436 222896
rect 154264 222856 211436 222884
rect 154264 222844 154270 222856
rect 211430 222844 211436 222856
rect 211488 222844 211494 222896
rect 211798 222844 211804 222896
rect 211856 222884 211862 222896
rect 214668 222884 214696 223128
rect 228082 223116 228088 223128
rect 228140 223116 228146 223168
rect 241330 223116 241336 223168
rect 241388 223156 241394 223168
rect 283466 223156 283472 223168
rect 241388 223128 283472 223156
rect 241388 223116 241394 223128
rect 283466 223116 283472 223128
rect 283524 223116 283530 223168
rect 288250 223116 288256 223168
rect 288308 223156 288314 223168
rect 321094 223156 321100 223168
rect 288308 223128 321100 223156
rect 288308 223116 288314 223128
rect 321094 223116 321100 223128
rect 321152 223116 321158 223168
rect 344646 223116 344652 223168
rect 344704 223156 344710 223168
rect 364610 223156 364616 223168
rect 344704 223128 364616 223156
rect 344704 223116 344710 223128
rect 364610 223116 364616 223128
rect 364668 223116 364674 223168
rect 365530 223116 365536 223168
rect 365588 223156 365594 223168
rect 379606 223156 379612 223168
rect 365588 223128 379612 223156
rect 365588 223116 365594 223128
rect 379606 223116 379612 223128
rect 379664 223116 379670 223168
rect 380066 223116 380072 223168
rect 380124 223156 380130 223168
rect 386506 223156 386512 223168
rect 380124 223128 386512 223156
rect 380124 223116 380130 223128
rect 386506 223116 386512 223128
rect 386564 223116 386570 223168
rect 488626 223116 488632 223168
rect 488684 223156 488690 223168
rect 503162 223156 503168 223168
rect 488684 223128 503168 223156
rect 488684 223116 488690 223128
rect 503162 223116 503168 223128
rect 503220 223116 503226 223168
rect 503346 223116 503352 223168
rect 503404 223156 503410 223168
rect 521746 223156 521752 223168
rect 503404 223128 521752 223156
rect 503404 223116 503410 223128
rect 521746 223116 521752 223128
rect 521804 223116 521810 223168
rect 532050 223116 532056 223168
rect 532108 223156 532114 223168
rect 559006 223156 559012 223168
rect 532108 223128 559012 223156
rect 532108 223116 532114 223128
rect 559006 223116 559012 223128
rect 559064 223116 559070 223168
rect 561674 223116 561680 223168
rect 561732 223156 561738 223168
rect 562410 223156 562416 223168
rect 561732 223128 562416 223156
rect 561732 223116 561738 223128
rect 562410 223116 562416 223128
rect 562468 223156 562474 223168
rect 564802 223156 564808 223168
rect 562468 223128 564808 223156
rect 562468 223116 562474 223128
rect 564802 223116 564808 223128
rect 564860 223116 564866 223168
rect 576826 223156 576854 223264
rect 620646 223156 620652 223168
rect 576826 223128 596174 223156
rect 214834 222980 214840 223032
rect 214892 223020 214898 223032
rect 216214 223020 216220 223032
rect 214892 222992 216220 223020
rect 214892 222980 214898 222992
rect 216214 222980 216220 222992
rect 216272 222980 216278 223032
rect 230198 222980 230204 223032
rect 230256 223020 230262 223032
rect 275462 223020 275468 223032
rect 230256 222992 275468 223020
rect 230256 222980 230262 222992
rect 275462 222980 275468 222992
rect 275520 222980 275526 223032
rect 278590 222980 278596 223032
rect 278648 223020 278654 223032
rect 315022 223020 315028 223032
rect 278648 222992 315028 223020
rect 278648 222980 278654 222992
rect 315022 222980 315028 222992
rect 315080 222980 315086 223032
rect 316678 222980 316684 223032
rect 316736 223020 316742 223032
rect 327258 223020 327264 223032
rect 316736 222992 327264 223020
rect 316736 222980 316742 222992
rect 327258 222980 327264 222992
rect 327316 222980 327322 223032
rect 328086 222980 328092 223032
rect 328144 223020 328150 223032
rect 351454 223020 351460 223032
rect 328144 222992 351460 223020
rect 328144 222980 328150 222992
rect 351454 222980 351460 222992
rect 351512 222980 351518 223032
rect 353938 222980 353944 223032
rect 353996 223020 354002 223032
rect 365898 223020 365904 223032
rect 353996 222992 365904 223020
rect 353996 222980 354002 222992
rect 365898 222980 365904 222992
rect 365956 222980 365962 223032
rect 366910 222980 366916 223032
rect 366968 223020 366974 223032
rect 383930 223020 383936 223032
rect 366968 222992 383936 223020
rect 366968 222980 366974 222992
rect 383930 222980 383936 222992
rect 383988 222980 383994 223032
rect 384298 222980 384304 223032
rect 384356 223020 384362 223032
rect 393958 223020 393964 223032
rect 384356 222992 393964 223020
rect 384356 222980 384362 222992
rect 393958 222980 393964 222992
rect 394016 222980 394022 223032
rect 482738 222980 482744 223032
rect 482796 223020 482802 223032
rect 593966 223020 593972 223032
rect 482796 222992 593972 223020
rect 482796 222980 482802 222992
rect 593966 222980 593972 222992
rect 594024 222980 594030 223032
rect 596146 223020 596174 223128
rect 605806 223128 620652 223156
rect 605806 223020 605834 223128
rect 620646 223116 620652 223128
rect 620704 223116 620710 223168
rect 669056 223088 669084 224012
rect 669222 224000 669228 224012
rect 669280 224000 669286 224052
rect 670510 224000 670516 224052
rect 670568 224040 670574 224052
rect 670568 224012 671398 224040
rect 670568 224000 670574 224012
rect 669240 223876 671278 223904
rect 669240 223780 669268 223876
rect 669222 223728 669228 223780
rect 669280 223728 669286 223780
rect 670050 223768 670056 223780
rect 669884 223740 670056 223768
rect 669884 223644 669912 223740
rect 670050 223728 670056 223740
rect 670108 223728 670114 223780
rect 669866 223592 669872 223644
rect 669924 223592 669930 223644
rect 670160 223604 671186 223632
rect 669682 223564 669688 223576
rect 669424 223536 669688 223564
rect 669424 223224 669452 223536
rect 669682 223524 669688 223536
rect 669740 223524 669746 223576
rect 669590 223388 669596 223440
rect 669648 223428 669654 223440
rect 670160 223428 670188 223604
rect 669648 223400 670188 223428
rect 670804 223468 671048 223496
rect 669648 223388 669654 223400
rect 670804 223360 670832 223468
rect 670344 223332 670832 223360
rect 669424 223196 669728 223224
rect 669700 223100 669728 223196
rect 669866 223116 669872 223168
rect 669924 223156 669930 223168
rect 669924 223128 670096 223156
rect 669924 223116 669930 223128
rect 669056 223060 669544 223088
rect 596146 222992 605834 223020
rect 620278 222980 620284 223032
rect 620336 223020 620342 223032
rect 625614 223020 625620 223032
rect 620336 222992 625620 223020
rect 620336 222980 620342 222992
rect 625614 222980 625620 222992
rect 625672 222980 625678 223032
rect 669516 222952 669544 223060
rect 669682 223048 669688 223100
rect 669740 223048 669746 223100
rect 669866 222952 669872 222964
rect 669516 222924 669872 222952
rect 669866 222912 669872 222924
rect 669924 222912 669930 222964
rect 670068 222896 670096 223128
rect 211856 222856 214696 222884
rect 211856 222844 211862 222856
rect 215938 222844 215944 222896
rect 215996 222884 216002 222896
rect 233326 222884 233332 222896
rect 215996 222856 233332 222884
rect 215996 222844 216002 222856
rect 233326 222844 233332 222856
rect 233384 222844 233390 222896
rect 234522 222844 234528 222896
rect 234580 222884 234586 222896
rect 281534 222884 281540 222896
rect 234580 222856 281540 222884
rect 234580 222844 234586 222856
rect 281534 222844 281540 222856
rect 281592 222844 281598 222896
rect 282454 222844 282460 222896
rect 282512 222884 282518 222896
rect 316310 222884 316316 222896
rect 282512 222856 316316 222884
rect 282512 222844 282518 222856
rect 316310 222844 316316 222856
rect 316368 222844 316374 222896
rect 324130 222844 324136 222896
rect 324188 222884 324194 222896
rect 348510 222884 348516 222896
rect 324188 222856 348516 222884
rect 324188 222844 324194 222856
rect 348510 222844 348516 222856
rect 348568 222844 348574 222896
rect 349062 222844 349068 222896
rect 349120 222884 349126 222896
rect 367186 222884 367192 222896
rect 349120 222856 367192 222884
rect 349120 222844 349126 222856
rect 367186 222844 367192 222856
rect 367244 222844 367250 222896
rect 368382 222844 368388 222896
rect 368440 222884 368446 222896
rect 382366 222884 382372 222896
rect 368440 222856 382372 222884
rect 368440 222844 368446 222856
rect 382366 222844 382372 222856
rect 382424 222844 382430 222896
rect 383470 222844 383476 222896
rect 383528 222884 383534 222896
rect 394878 222884 394884 222896
rect 383528 222856 394884 222884
rect 383528 222844 383534 222856
rect 394878 222844 394884 222856
rect 394936 222844 394942 222896
rect 395798 222844 395804 222896
rect 395856 222884 395862 222896
rect 406470 222884 406476 222896
rect 395856 222856 406476 222884
rect 395856 222844 395862 222856
rect 406470 222844 406476 222856
rect 406528 222844 406534 222896
rect 420822 222844 420828 222896
rect 420880 222884 420886 222896
rect 425146 222884 425152 222896
rect 420880 222856 425152 222884
rect 420880 222844 420886 222856
rect 425146 222844 425152 222856
rect 425204 222844 425210 222896
rect 459922 222844 459928 222896
rect 459980 222884 459986 222896
rect 467098 222884 467104 222896
rect 459980 222856 467104 222884
rect 459980 222844 459986 222856
rect 467098 222844 467104 222856
rect 467156 222844 467162 222896
rect 467466 222844 467472 222896
rect 467524 222884 467530 222896
rect 473722 222884 473728 222896
rect 467524 222856 473728 222884
rect 467524 222844 467530 222856
rect 473722 222844 473728 222856
rect 473780 222844 473786 222896
rect 479886 222844 479892 222896
rect 479944 222884 479950 222896
rect 491938 222884 491944 222896
rect 479944 222856 491944 222884
rect 479944 222844 479950 222856
rect 491938 222844 491944 222856
rect 491996 222844 492002 222896
rect 500770 222844 500776 222896
rect 500828 222884 500834 222896
rect 517514 222884 517520 222896
rect 500828 222856 517520 222884
rect 500828 222844 500834 222856
rect 517514 222844 517520 222856
rect 517572 222844 517578 222896
rect 519814 222844 519820 222896
rect 519872 222884 519878 222896
rect 542354 222884 542360 222896
rect 519872 222856 542360 222884
rect 519872 222844 519878 222856
rect 542354 222844 542360 222856
rect 542412 222844 542418 222896
rect 554038 222844 554044 222896
rect 554096 222884 554102 222896
rect 632698 222884 632704 222896
rect 554096 222856 632704 222884
rect 554096 222844 554102 222856
rect 632698 222844 632704 222856
rect 632756 222844 632762 222896
rect 651282 222844 651288 222896
rect 651340 222884 651346 222896
rect 666462 222884 666468 222896
rect 651340 222856 666468 222884
rect 651340 222844 651346 222856
rect 666462 222844 666468 222856
rect 666520 222844 666526 222896
rect 670050 222844 670056 222896
rect 670108 222844 670114 222896
rect 78582 222708 78588 222760
rect 78640 222748 78646 222760
rect 155126 222748 155132 222760
rect 78640 222720 155132 222748
rect 78640 222708 78646 222720
rect 155126 222708 155132 222720
rect 155184 222708 155190 222760
rect 155678 222708 155684 222760
rect 155736 222748 155742 222760
rect 155736 222720 166120 222748
rect 155736 222708 155742 222720
rect 87966 222572 87972 222624
rect 88024 222612 88030 222624
rect 164970 222612 164976 222624
rect 88024 222584 164976 222612
rect 88024 222572 88030 222584
rect 164970 222572 164976 222584
rect 165028 222572 165034 222624
rect 166092 222612 166120 222720
rect 166258 222708 166264 222760
rect 166316 222748 166322 222760
rect 173526 222748 173532 222760
rect 166316 222720 173532 222748
rect 166316 222708 166322 222720
rect 173526 222708 173532 222720
rect 173584 222708 173590 222760
rect 173728 222720 185624 222748
rect 166442 222612 166448 222624
rect 166092 222584 166448 222612
rect 166442 222572 166448 222584
rect 166500 222572 166506 222624
rect 166626 222572 166632 222624
rect 166684 222612 166690 222624
rect 173728 222612 173756 222720
rect 166684 222584 173756 222612
rect 166684 222572 166690 222584
rect 173894 222572 173900 222624
rect 173952 222612 173958 222624
rect 175550 222612 175556 222624
rect 173952 222584 175556 222612
rect 173952 222572 173958 222584
rect 175550 222572 175556 222584
rect 175608 222572 175614 222624
rect 175918 222572 175924 222624
rect 175976 222612 175982 222624
rect 181806 222612 181812 222624
rect 175976 222584 181812 222612
rect 175976 222572 175982 222584
rect 181806 222572 181812 222584
rect 181864 222572 181870 222624
rect 185596 222612 185624 222720
rect 185762 222708 185768 222760
rect 185820 222748 185826 222760
rect 204714 222748 204720 222760
rect 185820 222720 204720 222748
rect 185820 222708 185826 222720
rect 204714 222708 204720 222720
rect 204772 222708 204778 222760
rect 204898 222708 204904 222760
rect 204956 222748 204962 222760
rect 247402 222748 247408 222760
rect 204956 222720 247408 222748
rect 204956 222708 204962 222720
rect 247402 222708 247408 222720
rect 247460 222708 247466 222760
rect 264790 222708 264796 222760
rect 264848 222748 264854 222760
rect 304350 222748 304356 222760
rect 264848 222720 304356 222748
rect 264848 222708 264854 222720
rect 304350 222708 304356 222720
rect 304408 222708 304414 222760
rect 508222 222708 508228 222760
rect 508280 222748 508286 222760
rect 527818 222748 527824 222760
rect 508280 222720 527824 222748
rect 508280 222708 508286 222720
rect 527818 222708 527824 222720
rect 527876 222708 527882 222760
rect 552474 222708 552480 222760
rect 552532 222748 552538 222760
rect 555694 222748 555700 222760
rect 552532 222720 555700 222748
rect 552532 222708 552538 222720
rect 555694 222708 555700 222720
rect 555752 222708 555758 222760
rect 558178 222708 558184 222760
rect 558236 222748 558242 222760
rect 620278 222748 620284 222760
rect 558236 222720 620284 222748
rect 558236 222708 558242 222720
rect 620278 222708 620284 222720
rect 620336 222708 620342 222760
rect 620462 222708 620468 222760
rect 620520 222748 620526 222760
rect 627086 222748 627092 222760
rect 620520 222720 627092 222748
rect 620520 222708 620526 222720
rect 627086 222708 627092 222720
rect 627144 222708 627150 222760
rect 304718 222640 304724 222692
rect 304776 222680 304782 222692
rect 308122 222680 308128 222692
rect 304776 222652 308128 222680
rect 304776 222640 304782 222652
rect 308122 222640 308128 222652
rect 308180 222640 308186 222692
rect 670344 222680 670372 223332
rect 670510 223116 670516 223168
rect 670568 223156 670574 223168
rect 670568 223128 670956 223156
rect 670568 223116 670574 223128
rect 670510 222680 670516 222692
rect 670344 222652 670516 222680
rect 670510 222640 670516 222652
rect 670568 222640 670574 222692
rect 192018 222612 192024 222624
rect 185596 222584 192024 222612
rect 192018 222572 192024 222584
rect 192076 222572 192082 222624
rect 197170 222572 197176 222624
rect 197228 222612 197234 222624
rect 249978 222612 249984 222624
rect 197228 222584 249984 222612
rect 197228 222572 197234 222584
rect 249978 222572 249984 222584
rect 250036 222572 250042 222624
rect 529842 222572 529848 222624
rect 529900 222612 529906 222624
rect 619910 222612 619916 222624
rect 529900 222584 619916 222612
rect 529900 222572 529906 222584
rect 619910 222572 619916 222584
rect 619968 222572 619974 222624
rect 426434 222504 426440 222556
rect 426492 222544 426498 222556
rect 426986 222544 426992 222556
rect 426492 222516 426992 222544
rect 426492 222504 426498 222516
rect 426986 222504 426992 222516
rect 427044 222504 427050 222556
rect 85298 222436 85304 222488
rect 85356 222476 85362 222488
rect 156414 222476 156420 222488
rect 85356 222448 156420 222476
rect 85356 222436 85362 222448
rect 156414 222436 156420 222448
rect 156472 222436 156478 222488
rect 156598 222436 156604 222488
rect 156656 222476 156662 222488
rect 156656 222448 175964 222476
rect 156656 222436 156662 222448
rect 99282 222300 99288 222352
rect 99340 222340 99346 222352
rect 99340 222312 173204 222340
rect 99340 222300 99346 222312
rect 118418 222164 118424 222216
rect 118476 222204 118482 222216
rect 156598 222204 156604 222216
rect 118476 222176 156604 222204
rect 118476 222164 118482 222176
rect 156598 222164 156604 222176
rect 156656 222164 156662 222216
rect 173176 222204 173204 222312
rect 173342 222300 173348 222352
rect 173400 222340 173406 222352
rect 175734 222340 175740 222352
rect 173400 222312 175740 222340
rect 173400 222300 173406 222312
rect 175734 222300 175740 222312
rect 175792 222300 175798 222352
rect 175936 222340 175964 222448
rect 176102 222436 176108 222488
rect 176160 222476 176166 222488
rect 207474 222476 207480 222488
rect 176160 222448 207480 222476
rect 176160 222436 176166 222448
rect 207474 222436 207480 222448
rect 207532 222436 207538 222488
rect 207658 222436 207664 222488
rect 207716 222476 207722 222488
rect 258350 222476 258356 222488
rect 207716 222448 258356 222476
rect 207716 222436 207722 222448
rect 258350 222436 258356 222448
rect 258408 222436 258414 222488
rect 489914 222436 489920 222488
rect 489972 222476 489978 222488
rect 491110 222476 491116 222488
rect 489972 222448 491116 222476
rect 489972 222436 489978 222448
rect 491110 222436 491116 222448
rect 491168 222476 491174 222488
rect 491168 222448 499574 222476
rect 491168 222436 491174 222448
rect 175936 222312 185624 222340
rect 173894 222204 173900 222216
rect 173176 222176 173900 222204
rect 173894 222164 173900 222176
rect 173952 222164 173958 222216
rect 185596 222204 185624 222312
rect 188890 222300 188896 222352
rect 188948 222340 188954 222352
rect 245102 222340 245108 222352
rect 188948 222312 245108 222340
rect 188948 222300 188954 222312
rect 245102 222300 245108 222312
rect 245160 222300 245166 222352
rect 287882 222300 287888 222352
rect 287940 222340 287946 222352
rect 295058 222340 295064 222352
rect 287940 222312 295064 222340
rect 287940 222300 287946 222312
rect 295058 222300 295064 222312
rect 295116 222300 295122 222352
rect 484486 222300 484492 222352
rect 484544 222340 484550 222352
rect 499546 222340 499574 222448
rect 504358 222436 504364 222488
rect 504416 222476 504422 222488
rect 523678 222476 523684 222488
rect 504416 222448 523684 222476
rect 504416 222436 504422 222448
rect 523678 222436 523684 222448
rect 523736 222436 523742 222488
rect 529474 222436 529480 222488
rect 529532 222476 529538 222488
rect 552474 222476 552480 222488
rect 529532 222448 552480 222476
rect 529532 222436 529538 222448
rect 552474 222436 552480 222448
rect 552532 222436 552538 222488
rect 552658 222436 552664 222488
rect 552716 222476 552722 222488
rect 564618 222476 564624 222488
rect 552716 222448 564624 222476
rect 552716 222436 552722 222448
rect 564618 222436 564624 222448
rect 564676 222436 564682 222488
rect 564802 222436 564808 222488
rect 564860 222476 564866 222488
rect 627914 222476 627920 222488
rect 564860 222448 627920 222476
rect 564860 222436 564866 222448
rect 627914 222436 627920 222448
rect 627972 222436 627978 222488
rect 629846 222340 629852 222352
rect 484544 222312 485774 222340
rect 499546 222312 629852 222340
rect 484544 222300 484550 222312
rect 191006 222204 191012 222216
rect 185596 222176 191012 222204
rect 191006 222164 191012 222176
rect 191064 222164 191070 222216
rect 485746 222204 485774 222312
rect 629846 222300 629852 222312
rect 629904 222300 629910 222352
rect 504358 222204 504364 222216
rect 485746 222176 504364 222204
rect 504358 222164 504364 222176
rect 504416 222164 504422 222216
rect 523678 222164 523684 222216
rect 523736 222204 523742 222216
rect 552658 222204 552664 222216
rect 523736 222176 552664 222204
rect 523736 222164 523742 222176
rect 552658 222164 552664 222176
rect 552716 222164 552722 222216
rect 552842 222164 552848 222216
rect 552900 222204 552906 222216
rect 558178 222204 558184 222216
rect 552900 222176 558184 222204
rect 552900 222164 552906 222176
rect 558178 222164 558184 222176
rect 558236 222164 558242 222216
rect 558546 222164 558552 222216
rect 558604 222204 558610 222216
rect 559926 222204 559932 222216
rect 558604 222176 559932 222204
rect 558604 222164 558610 222176
rect 559926 222164 559932 222176
rect 559984 222204 559990 222216
rect 620462 222204 620468 222216
rect 559984 222176 620468 222204
rect 559984 222164 559990 222176
rect 620462 222164 620468 222176
rect 620520 222164 620526 222216
rect 620646 222164 620652 222216
rect 620704 222204 620710 222216
rect 631502 222204 631508 222216
rect 620704 222176 631508 222204
rect 620704 222164 620710 222176
rect 631502 222164 631508 222176
rect 631560 222164 631566 222216
rect 160830 222096 160836 222148
rect 160888 222136 160894 222148
rect 166074 222136 166080 222148
rect 160888 222108 166080 222136
rect 160888 222096 160894 222108
rect 166074 222096 166080 222108
rect 166132 222096 166138 222148
rect 172698 222136 172704 222148
rect 166276 222108 172704 222136
rect 97902 221960 97908 222012
rect 97960 222000 97966 222012
rect 166276 222000 166304 222108
rect 172698 222096 172704 222108
rect 172756 222096 172762 222148
rect 174354 222096 174360 222148
rect 174412 222136 174418 222148
rect 174412 222108 180794 222136
rect 174412 222096 174418 222108
rect 97960 221972 166304 222000
rect 97960 221960 97966 221972
rect 167454 221960 167460 222012
rect 167512 222000 167518 222012
rect 175918 222000 175924 222012
rect 167512 221972 175924 222000
rect 167512 221960 167518 221972
rect 175918 221960 175924 221972
rect 175976 221960 175982 222012
rect 180766 222000 180794 222108
rect 181438 222096 181444 222148
rect 181496 222136 181502 222148
rect 182634 222136 182640 222148
rect 181496 222108 182640 222136
rect 181496 222096 181502 222108
rect 182634 222096 182640 222108
rect 182692 222096 182698 222148
rect 191466 222096 191472 222148
rect 191524 222136 191530 222148
rect 247586 222136 247592 222148
rect 191524 222108 247592 222136
rect 191524 222096 191530 222108
rect 247586 222096 247592 222108
rect 247644 222096 247650 222148
rect 258074 222096 258080 222148
rect 258132 222136 258138 222148
rect 263686 222136 263692 222148
rect 258132 222108 263692 222136
rect 258132 222096 258138 222108
rect 263686 222096 263692 222108
rect 263744 222096 263750 222148
rect 270218 222096 270224 222148
rect 270276 222136 270282 222148
rect 306558 222136 306564 222148
rect 270276 222108 306564 222136
rect 270276 222096 270282 222108
rect 306558 222096 306564 222108
rect 306616 222096 306622 222148
rect 310698 222096 310704 222148
rect 310756 222136 310762 222148
rect 312630 222136 312636 222148
rect 310756 222108 312636 222136
rect 310756 222096 310762 222108
rect 312630 222096 312636 222108
rect 312688 222096 312694 222148
rect 331398 222096 331404 222148
rect 331456 222136 331462 222148
rect 353754 222136 353760 222148
rect 331456 222108 353760 222136
rect 331456 222096 331462 222108
rect 353754 222096 353760 222108
rect 353812 222096 353818 222148
rect 452470 222096 452476 222148
rect 452528 222136 452534 222148
rect 455598 222136 455604 222148
rect 452528 222108 455604 222136
rect 452528 222096 452534 222108
rect 455598 222096 455604 222108
rect 455656 222096 455662 222148
rect 462130 222096 462136 222148
rect 462188 222136 462194 222148
rect 468754 222136 468760 222148
rect 462188 222108 468760 222136
rect 462188 222096 462194 222108
rect 468754 222096 468760 222108
rect 468812 222096 468818 222148
rect 471882 222096 471888 222148
rect 471940 222136 471946 222148
rect 477862 222136 477868 222148
rect 471940 222108 477868 222136
rect 471940 222096 471946 222108
rect 477862 222096 477868 222108
rect 477920 222096 477926 222148
rect 495158 222028 495164 222080
rect 495216 222068 495222 222080
rect 497734 222068 497740 222080
rect 495216 222040 497740 222068
rect 495216 222028 495222 222040
rect 497734 222028 497740 222040
rect 497792 222028 497798 222080
rect 515490 222028 515496 222080
rect 515548 222068 515554 222080
rect 529842 222068 529848 222080
rect 515548 222040 529848 222068
rect 515548 222028 515554 222040
rect 529842 222028 529848 222040
rect 529900 222028 529906 222080
rect 533982 222028 533988 222080
rect 534040 222068 534046 222080
rect 534040 222028 534074 222068
rect 536098 222028 536104 222080
rect 536156 222068 536162 222080
rect 539594 222068 539600 222080
rect 536156 222040 539600 222068
rect 536156 222028 536162 222040
rect 539594 222028 539600 222040
rect 539652 222028 539658 222080
rect 539778 222028 539784 222080
rect 539836 222068 539842 222080
rect 539836 222040 586514 222068
rect 539836 222028 539842 222040
rect 232130 222000 232136 222012
rect 180766 221972 232136 222000
rect 232130 221960 232136 221972
rect 232188 221960 232194 222012
rect 233694 221960 233700 222012
rect 233752 222000 233758 222012
rect 277946 222000 277952 222012
rect 233752 221972 277952 222000
rect 233752 221960 233758 221972
rect 277946 221960 277952 221972
rect 278004 221960 278010 222012
rect 280062 221960 280068 222012
rect 280120 222000 280126 222012
rect 313734 222000 313740 222012
rect 280120 221972 313740 222000
rect 280120 221960 280126 221972
rect 313734 221960 313740 221972
rect 313792 221960 313798 222012
rect 318242 221960 318248 222012
rect 318300 222000 318306 222012
rect 343818 222000 343824 222012
rect 318300 221972 343824 222000
rect 318300 221960 318306 221972
rect 343818 221960 343824 221972
rect 343876 221960 343882 222012
rect 367646 221960 367652 222012
rect 367704 222000 367710 222012
rect 380250 222000 380256 222012
rect 367704 221972 380256 222000
rect 367704 221960 367710 221972
rect 380250 221960 380256 221972
rect 380308 221960 380314 222012
rect 424962 221892 424968 221944
rect 425020 221932 425026 221944
rect 429194 221932 429200 221944
rect 425020 221904 429200 221932
rect 425020 221892 425026 221904
rect 429194 221892 429200 221904
rect 429252 221892 429258 221944
rect 534046 221932 534074 222028
rect 559374 221932 559380 221944
rect 534046 221904 559380 221932
rect 559374 221892 559380 221904
rect 559432 221892 559438 221944
rect 559558 221892 559564 221944
rect 559616 221932 559622 221944
rect 564802 221932 564808 221944
rect 559616 221904 564808 221932
rect 559616 221892 559622 221904
rect 564802 221892 564808 221904
rect 564860 221892 564866 221944
rect 104526 221824 104532 221876
rect 104584 221864 104590 221876
rect 173342 221864 173348 221876
rect 104584 221836 173348 221864
rect 104584 221824 104590 221836
rect 173342 221824 173348 221836
rect 173400 221824 173406 221876
rect 173526 221824 173532 221876
rect 173584 221864 173590 221876
rect 181438 221864 181444 221876
rect 173584 221836 181444 221864
rect 173584 221824 173590 221836
rect 181438 221824 181444 221836
rect 181496 221824 181502 221876
rect 181622 221824 181628 221876
rect 181680 221864 181686 221876
rect 240134 221864 240140 221876
rect 181680 221836 240140 221864
rect 181680 221824 181686 221836
rect 240134 221824 240140 221836
rect 240192 221824 240198 221876
rect 263318 221824 263324 221876
rect 263376 221864 263382 221876
rect 301130 221864 301136 221876
rect 263376 221836 301136 221864
rect 263376 221824 263382 221836
rect 301130 221824 301136 221836
rect 301188 221824 301194 221876
rect 301958 221824 301964 221876
rect 302016 221864 302022 221876
rect 310882 221864 310888 221876
rect 302016 221836 310888 221864
rect 302016 221824 302022 221836
rect 310882 221824 310888 221836
rect 310940 221824 310946 221876
rect 313182 221824 313188 221876
rect 313240 221864 313246 221876
rect 340414 221864 340420 221876
rect 313240 221836 340420 221864
rect 313240 221824 313246 221836
rect 340414 221824 340420 221836
rect 340472 221824 340478 221876
rect 351270 221824 351276 221876
rect 351328 221864 351334 221876
rect 369302 221864 369308 221876
rect 351328 221836 369308 221864
rect 351328 221824 351334 221836
rect 369302 221824 369308 221836
rect 369360 221824 369366 221876
rect 509878 221824 509884 221876
rect 509936 221864 509942 221876
rect 522574 221864 522580 221876
rect 509936 221836 522580 221864
rect 509936 221824 509942 221836
rect 522574 221824 522580 221836
rect 522632 221824 522638 221876
rect 586486 221864 586514 222040
rect 596634 221960 596640 222012
rect 596692 222000 596698 222012
rect 605006 222000 605012 222012
rect 596692 221972 605012 222000
rect 596692 221960 596698 221972
rect 605006 221960 605012 221972
rect 605064 221960 605070 222012
rect 600774 221864 600780 221876
rect 586486 221836 600780 221864
rect 600774 221824 600780 221836
rect 600832 221824 600838 221876
rect 600958 221824 600964 221876
rect 601016 221864 601022 221876
rect 606662 221864 606668 221876
rect 601016 221836 606668 221864
rect 601016 221824 601022 221836
rect 606662 221824 606668 221836
rect 606720 221824 606726 221876
rect 539318 221796 539324 221808
rect 534046 221768 539324 221796
rect 80514 221688 80520 221740
rect 80572 221728 80578 221740
rect 86218 221728 86224 221740
rect 80572 221700 86224 221728
rect 80572 221688 80578 221700
rect 86218 221688 86224 221700
rect 86276 221688 86282 221740
rect 94682 221688 94688 221740
rect 94740 221728 94746 221740
rect 161428 221728 161434 221740
rect 94740 221700 161434 221728
rect 94740 221688 94746 221700
rect 161428 221688 161434 221700
rect 161486 221688 161492 221740
rect 161566 221688 161572 221740
rect 161624 221728 161630 221740
rect 167178 221728 167184 221740
rect 161624 221700 167184 221728
rect 161624 221688 161630 221700
rect 167178 221688 167184 221700
rect 167236 221688 167242 221740
rect 167638 221688 167644 221740
rect 167696 221728 167702 221740
rect 169754 221728 169760 221740
rect 167696 221700 169760 221728
rect 167696 221688 167702 221700
rect 169754 221688 169760 221700
rect 169812 221688 169818 221740
rect 171594 221688 171600 221740
rect 171652 221728 171658 221740
rect 232314 221728 232320 221740
rect 171652 221700 232320 221728
rect 171652 221688 171658 221700
rect 232314 221688 232320 221700
rect 232372 221688 232378 221740
rect 239306 221688 239312 221740
rect 239364 221728 239370 221740
rect 283650 221728 283656 221740
rect 239364 221700 283656 221728
rect 239364 221688 239370 221700
rect 283650 221688 283656 221700
rect 283708 221688 283714 221740
rect 303246 221688 303252 221740
rect 303304 221728 303310 221740
rect 332778 221728 332784 221740
rect 303304 221700 332784 221728
rect 303304 221688 303310 221700
rect 332778 221688 332784 221700
rect 332836 221688 332842 221740
rect 357158 221688 357164 221740
rect 357216 221728 357222 221740
rect 374638 221728 374644 221740
rect 357216 221700 374644 221728
rect 357216 221688 357222 221700
rect 374638 221688 374644 221700
rect 374696 221688 374702 221740
rect 391014 221688 391020 221740
rect 391072 221728 391078 221740
rect 400306 221728 400312 221740
rect 391072 221700 400312 221728
rect 391072 221688 391078 221700
rect 400306 221688 400312 221700
rect 400364 221688 400370 221740
rect 475930 221688 475936 221740
rect 475988 221728 475994 221740
rect 486142 221728 486148 221740
rect 475988 221700 486148 221728
rect 475988 221688 475994 221700
rect 486142 221688 486148 221700
rect 486200 221688 486206 221740
rect 496262 221688 496268 221740
rect 496320 221728 496326 221740
rect 513558 221728 513564 221740
rect 496320 221700 513564 221728
rect 496320 221688 496326 221700
rect 513558 221688 513564 221700
rect 513616 221688 513622 221740
rect 524230 221688 524236 221740
rect 524288 221728 524294 221740
rect 534046 221728 534074 221768
rect 539318 221756 539324 221768
rect 539376 221756 539382 221808
rect 539594 221756 539600 221808
rect 539652 221796 539658 221808
rect 547828 221796 547834 221808
rect 539652 221768 547834 221796
rect 539652 221756 539658 221768
rect 547828 221756 547834 221768
rect 547886 221756 547892 221808
rect 547966 221756 547972 221808
rect 548024 221796 548030 221808
rect 549070 221796 549076 221808
rect 548024 221768 549076 221796
rect 548024 221756 548030 221768
rect 549070 221756 549076 221768
rect 549128 221756 549134 221808
rect 549254 221756 549260 221808
rect 549312 221796 549318 221808
rect 552106 221796 552112 221808
rect 549312 221768 552112 221796
rect 549312 221756 549318 221768
rect 552106 221756 552112 221768
rect 552164 221796 552170 221808
rect 552842 221796 552848 221808
rect 552164 221768 552848 221796
rect 552164 221756 552170 221768
rect 552842 221756 552848 221768
rect 552900 221756 552906 221808
rect 553302 221756 553308 221808
rect 553360 221796 553366 221808
rect 553360 221768 563054 221796
rect 553360 221756 553366 221768
rect 524288 221700 534074 221728
rect 563026 221728 563054 221768
rect 608594 221728 608600 221740
rect 563026 221700 608600 221728
rect 524288 221688 524294 221700
rect 608594 221688 608600 221700
rect 608652 221688 608658 221740
rect 546586 221660 546592 221672
rect 538876 221632 546592 221660
rect 59354 221552 59360 221604
rect 59412 221592 59418 221604
rect 141326 221592 141332 221604
rect 59412 221564 141332 221592
rect 59412 221552 59418 221564
rect 141326 221552 141332 221564
rect 141384 221552 141390 221604
rect 141510 221552 141516 221604
rect 141568 221592 141574 221604
rect 147398 221592 147404 221604
rect 141568 221564 147404 221592
rect 141568 221552 141574 221564
rect 147398 221552 147404 221564
rect 147456 221552 147462 221604
rect 147582 221552 147588 221604
rect 147640 221592 147646 221604
rect 205910 221592 205916 221604
rect 147640 221564 205916 221592
rect 147640 221552 147646 221564
rect 205910 221552 205916 221564
rect 205968 221552 205974 221604
rect 208394 221552 208400 221604
rect 208452 221592 208458 221604
rect 260834 221592 260840 221604
rect 208452 221564 260840 221592
rect 208452 221552 208458 221564
rect 260834 221552 260840 221564
rect 260892 221552 260898 221604
rect 261018 221552 261024 221604
rect 261076 221592 261082 221604
rect 301774 221592 301780 221604
rect 261076 221564 301780 221592
rect 261076 221552 261082 221564
rect 301774 221552 301780 221564
rect 301832 221552 301838 221604
rect 308858 221552 308864 221604
rect 308916 221592 308922 221604
rect 339678 221592 339684 221604
rect 308916 221564 339684 221592
rect 308916 221552 308922 221564
rect 339678 221552 339684 221564
rect 339736 221552 339742 221604
rect 341334 221552 341340 221604
rect 341392 221592 341398 221604
rect 361758 221592 361764 221604
rect 341392 221564 361764 221592
rect 341392 221552 341398 221564
rect 361758 221552 361764 221564
rect 361816 221552 361822 221604
rect 369486 221552 369492 221604
rect 369544 221592 369550 221604
rect 384114 221592 384120 221604
rect 369544 221564 384120 221592
rect 369544 221552 369550 221564
rect 384114 221552 384120 221564
rect 384172 221552 384178 221604
rect 384482 221552 384488 221604
rect 384540 221592 384546 221604
rect 395154 221592 395160 221604
rect 384540 221564 395160 221592
rect 384540 221552 384546 221564
rect 395154 221552 395160 221564
rect 395212 221552 395218 221604
rect 400674 221552 400680 221604
rect 400732 221592 400738 221604
rect 405826 221592 405832 221604
rect 400732 221564 405832 221592
rect 400732 221552 400738 221564
rect 405826 221552 405832 221564
rect 405884 221552 405890 221604
rect 480806 221552 480812 221604
rect 480864 221592 480870 221604
rect 492950 221592 492956 221604
rect 480864 221564 492956 221592
rect 480864 221552 480870 221564
rect 492950 221552 492956 221564
rect 493008 221552 493014 221604
rect 497458 221552 497464 221604
rect 497516 221592 497522 221604
rect 515122 221592 515128 221604
rect 497516 221564 515128 221592
rect 497516 221552 497522 221564
rect 515122 221552 515128 221564
rect 515180 221552 515186 221604
rect 522850 221552 522856 221604
rect 522908 221592 522914 221604
rect 538876 221592 538904 221632
rect 546586 221620 546592 221632
rect 546644 221620 546650 221672
rect 547138 221620 547144 221672
rect 547196 221660 547202 221672
rect 553946 221660 553952 221672
rect 547196 221632 553952 221660
rect 547196 221620 547202 221632
rect 553946 221620 553952 221632
rect 554004 221620 554010 221672
rect 596634 221592 596640 221604
rect 522908 221564 538904 221592
rect 554148 221564 596640 221592
rect 522908 221552 522914 221564
rect 539318 221484 539324 221536
rect 539376 221524 539382 221536
rect 547828 221524 547834 221536
rect 539376 221496 547834 221524
rect 539376 221484 539382 221496
rect 547828 221484 547834 221496
rect 547886 221484 547892 221536
rect 547966 221484 547972 221536
rect 548024 221524 548030 221536
rect 552290 221524 552296 221536
rect 548024 221496 552296 221524
rect 548024 221484 548030 221496
rect 552290 221484 552296 221496
rect 552348 221484 552354 221536
rect 554148 221524 554176 221564
rect 596634 221552 596640 221564
rect 596692 221552 596698 221604
rect 596818 221552 596824 221604
rect 596876 221592 596882 221604
rect 633434 221592 633440 221604
rect 596876 221564 633440 221592
rect 596876 221552 596882 221564
rect 633434 221552 633440 221564
rect 633492 221552 633498 221604
rect 552676 221496 554176 221524
rect 73890 221416 73896 221468
rect 73948 221456 73954 221468
rect 82078 221456 82084 221468
rect 73948 221428 82084 221456
rect 73948 221416 73954 221428
rect 82078 221416 82084 221428
rect 82136 221416 82142 221468
rect 86310 221416 86316 221468
rect 86368 221456 86374 221468
rect 86368 221428 161612 221456
rect 86368 221416 86374 221428
rect 91278 221280 91284 221332
rect 91336 221320 91342 221332
rect 91336 221292 118004 221320
rect 91336 221280 91342 221292
rect 117976 221184 118004 221292
rect 118142 221280 118148 221332
rect 118200 221320 118206 221332
rect 127434 221320 127440 221332
rect 118200 221292 127440 221320
rect 118200 221280 118206 221292
rect 127434 221280 127440 221292
rect 127492 221280 127498 221332
rect 161428 221320 161434 221332
rect 127636 221292 161434 221320
rect 127636 221184 127664 221292
rect 161428 221280 161434 221292
rect 161486 221280 161492 221332
rect 161584 221320 161612 221428
rect 161750 221416 161756 221468
rect 161808 221456 161814 221468
rect 161808 221428 173756 221456
rect 161808 221416 161814 221428
rect 164326 221320 164332 221332
rect 161584 221292 164332 221320
rect 164326 221280 164332 221292
rect 164384 221280 164390 221332
rect 173526 221320 173532 221332
rect 164712 221292 173532 221320
rect 164712 221184 164740 221292
rect 173526 221280 173532 221292
rect 173584 221280 173590 221332
rect 173728 221320 173756 221428
rect 175918 221416 175924 221468
rect 175976 221456 175982 221468
rect 226518 221456 226524 221468
rect 175976 221428 226524 221456
rect 175976 221416 175982 221428
rect 226518 221416 226524 221428
rect 226576 221416 226582 221468
rect 227898 221416 227904 221468
rect 227956 221456 227962 221468
rect 276106 221456 276112 221468
rect 227956 221428 276112 221456
rect 227956 221416 227962 221428
rect 276106 221416 276112 221428
rect 276164 221416 276170 221468
rect 292482 221416 292488 221468
rect 292540 221456 292546 221468
rect 326246 221456 326252 221468
rect 292540 221428 326252 221456
rect 292540 221416 292546 221428
rect 326246 221416 326252 221428
rect 326304 221416 326310 221468
rect 342162 221416 342168 221468
rect 342220 221456 342226 221468
rect 364794 221456 364800 221468
rect 342220 221428 364800 221456
rect 342220 221416 342226 221428
rect 364794 221416 364800 221428
rect 364852 221416 364858 221468
rect 375282 221416 375288 221468
rect 375340 221456 375346 221468
rect 390738 221456 390744 221468
rect 375340 221428 390744 221456
rect 375340 221416 375346 221428
rect 390738 221416 390744 221428
rect 390796 221416 390802 221468
rect 396810 221416 396816 221468
rect 396868 221456 396874 221468
rect 407298 221456 407304 221468
rect 396868 221428 407304 221456
rect 396868 221416 396874 221428
rect 407298 221416 407304 221428
rect 407356 221416 407362 221468
rect 408402 221416 408408 221468
rect 408460 221456 408466 221468
rect 416866 221456 416872 221468
rect 408460 221428 416872 221456
rect 408460 221416 408466 221428
rect 416866 221416 416872 221428
rect 416924 221416 416930 221468
rect 468938 221416 468944 221468
rect 468996 221456 469002 221468
rect 476206 221456 476212 221468
rect 468996 221428 476212 221456
rect 468996 221416 469002 221428
rect 476206 221416 476212 221428
rect 476264 221416 476270 221468
rect 483750 221416 483756 221468
rect 483808 221456 483814 221468
rect 538490 221456 538496 221468
rect 483808 221428 538496 221456
rect 483808 221416 483814 221428
rect 538490 221416 538496 221428
rect 538548 221416 538554 221468
rect 552676 221456 552704 221496
rect 600958 221456 600964 221468
rect 552492 221428 552704 221456
rect 563026 221428 600964 221456
rect 538674 221348 538680 221400
rect 538732 221388 538738 221400
rect 552492 221388 552520 221428
rect 538732 221360 552520 221388
rect 538732 221348 538738 221360
rect 553118 221348 553124 221400
rect 553176 221388 553182 221400
rect 563026 221388 563054 221428
rect 600958 221416 600964 221428
rect 601016 221416 601022 221468
rect 553176 221360 563054 221388
rect 553176 221348 553182 221360
rect 193398 221320 193404 221332
rect 173728 221292 193404 221320
rect 193398 221280 193404 221292
rect 193456 221280 193462 221332
rect 204162 221280 204168 221332
rect 204220 221320 204226 221332
rect 252738 221320 252744 221332
rect 204220 221292 252744 221320
rect 204220 221280 204226 221292
rect 252738 221280 252744 221292
rect 252796 221280 252802 221332
rect 266814 221280 266820 221332
rect 266872 221320 266878 221332
rect 303798 221320 303804 221332
rect 266872 221292 303804 221320
rect 266872 221280 266878 221292
rect 303798 221280 303804 221292
rect 303856 221280 303862 221332
rect 600866 221280 600872 221332
rect 600924 221320 600930 221332
rect 604638 221320 604644 221332
rect 600924 221292 604644 221320
rect 600924 221280 600930 221292
rect 604638 221280 604644 221292
rect 604696 221280 604702 221332
rect 521102 221212 521108 221264
rect 521160 221252 521166 221264
rect 600498 221252 600504 221264
rect 521160 221224 600504 221252
rect 521160 221212 521166 221224
rect 600498 221212 600504 221224
rect 600556 221212 600562 221264
rect 117976 221156 127664 221184
rect 127728 221156 164740 221184
rect 111150 221008 111156 221060
rect 111208 221048 111214 221060
rect 118142 221048 118148 221060
rect 111208 221020 118148 221048
rect 111208 221008 111214 221020
rect 118142 221008 118148 221020
rect 118200 221008 118206 221060
rect 124398 221008 124404 221060
rect 124456 221048 124462 221060
rect 127250 221048 127256 221060
rect 124456 221020 127256 221048
rect 124456 221008 124462 221020
rect 127250 221008 127256 221020
rect 127308 221008 127314 221060
rect 127434 221008 127440 221060
rect 127492 221048 127498 221060
rect 127728 221048 127756 221156
rect 166074 221144 166080 221196
rect 166132 221184 166138 221196
rect 221274 221184 221280 221196
rect 166132 221156 221280 221184
rect 166132 221144 166138 221156
rect 221274 221144 221280 221156
rect 221332 221144 221338 221196
rect 222746 221144 222752 221196
rect 222804 221184 222810 221196
rect 268286 221184 268292 221196
rect 222804 221156 268292 221184
rect 222804 221144 222810 221156
rect 268286 221144 268292 221156
rect 268344 221144 268350 221196
rect 523494 221076 523500 221128
rect 523552 221116 523558 221128
rect 601786 221116 601792 221128
rect 523552 221088 601792 221116
rect 523552 221076 523558 221088
rect 601786 221076 601792 221088
rect 601844 221076 601850 221128
rect 127492 221020 127756 221048
rect 127492 221008 127498 221020
rect 127894 221008 127900 221060
rect 127952 221048 127958 221060
rect 127952 221020 147444 221048
rect 127952 221008 127958 221020
rect 82998 220872 83004 220924
rect 83056 220912 83062 220924
rect 147416 220912 147444 221020
rect 147628 221008 147634 221060
rect 147686 221048 147692 221060
rect 206462 221048 206468 221060
rect 147686 221020 206468 221048
rect 147686 221008 147692 221020
rect 206462 221008 206468 221020
rect 206520 221008 206526 221060
rect 219802 221008 219808 221060
rect 219860 221048 219866 221060
rect 263042 221048 263048 221060
rect 219860 221020 263048 221048
rect 219860 221008 219866 221020
rect 263042 221008 263048 221020
rect 263100 221008 263106 221060
rect 525978 220940 525984 220992
rect 526036 220980 526042 220992
rect 602246 220980 602252 220992
rect 526036 220952 602252 220980
rect 526036 220940 526042 220952
rect 602246 220940 602252 220952
rect 602304 220940 602310 220992
rect 161428 220912 161434 220924
rect 83056 220884 146984 220912
rect 147416 220884 161434 220912
rect 83056 220872 83062 220884
rect 146956 220844 146984 220884
rect 161428 220872 161434 220884
rect 161486 220872 161492 220924
rect 161566 220872 161572 220924
rect 161624 220912 161630 220924
rect 222286 220912 222292 220924
rect 161624 220884 222292 220912
rect 161624 220872 161630 220884
rect 222286 220872 222292 220884
rect 222344 220872 222350 220924
rect 282638 220872 282644 220924
rect 282696 220912 282702 220924
rect 287698 220912 287704 220924
rect 282696 220884 287704 220912
rect 282696 220872 282702 220884
rect 287698 220872 287704 220884
rect 287756 220872 287762 220924
rect 456702 220872 456708 220924
rect 456760 220912 456766 220924
rect 456760 220884 460934 220912
rect 456760 220872 456766 220884
rect 147214 220844 147220 220856
rect 146956 220816 147220 220844
rect 147214 220804 147220 220816
rect 147272 220804 147278 220856
rect 253842 220804 253848 220856
rect 253900 220844 253906 220856
rect 258626 220844 258632 220856
rect 253900 220816 258632 220844
rect 253900 220804 253906 220816
rect 258626 220804 258632 220816
rect 258684 220804 258690 220856
rect 418338 220804 418344 220856
rect 418396 220844 418402 220856
rect 424042 220844 424048 220856
rect 418396 220816 424048 220844
rect 418396 220804 418402 220816
rect 424042 220804 424048 220816
rect 424100 220804 424106 220856
rect 460906 220844 460934 220884
rect 462130 220844 462136 220856
rect 460906 220816 462136 220844
rect 462130 220804 462136 220816
rect 462188 220804 462194 220856
rect 466086 220804 466092 220856
rect 466144 220844 466150 220856
rect 471422 220844 471428 220856
rect 466144 220816 471428 220844
rect 466144 220804 466150 220816
rect 471422 220804 471428 220816
rect 471480 220804 471486 220856
rect 517514 220804 517520 220856
rect 517572 220844 517578 220856
rect 518526 220844 518532 220856
rect 517572 220816 518532 220844
rect 517572 220804 517578 220816
rect 518526 220804 518532 220816
rect 518584 220844 518590 220856
rect 600314 220844 600320 220856
rect 518584 220816 600320 220844
rect 518584 220804 518590 220816
rect 600314 220804 600320 220816
rect 600372 220804 600378 220856
rect 114278 220736 114284 220788
rect 114336 220776 114342 220788
rect 146754 220776 146760 220788
rect 114336 220748 146760 220776
rect 114336 220736 114342 220748
rect 146754 220736 146760 220748
rect 146812 220736 146818 220788
rect 180748 220776 180754 220788
rect 147554 220748 180754 220776
rect 101214 220600 101220 220652
rect 101272 220640 101278 220652
rect 147030 220640 147036 220652
rect 101272 220612 147036 220640
rect 101272 220600 101278 220612
rect 147030 220600 147036 220612
rect 147088 220600 147094 220652
rect 147554 220640 147582 220748
rect 180748 220736 180754 220748
rect 180806 220736 180812 220788
rect 181070 220736 181076 220788
rect 181128 220776 181134 220788
rect 190362 220776 190368 220788
rect 181128 220748 190368 220776
rect 181128 220736 181134 220748
rect 190362 220736 190368 220748
rect 190420 220736 190426 220788
rect 190546 220736 190552 220788
rect 190604 220776 190610 220788
rect 236638 220776 236644 220788
rect 190604 220748 236644 220776
rect 190604 220736 190610 220748
rect 236638 220736 236644 220748
rect 236696 220736 236702 220788
rect 242618 220736 242624 220788
rect 242676 220776 242682 220788
rect 246482 220776 246488 220788
rect 242676 220748 246488 220776
rect 242676 220736 242682 220748
rect 246482 220736 246488 220748
rect 246540 220736 246546 220788
rect 260190 220736 260196 220788
rect 260248 220776 260254 220788
rect 298554 220776 298560 220788
rect 260248 220748 298560 220776
rect 260248 220736 260254 220748
rect 298554 220736 298560 220748
rect 298612 220736 298618 220788
rect 321554 220736 321560 220788
rect 321612 220776 321618 220788
rect 324498 220776 324504 220788
rect 321612 220748 324504 220776
rect 321612 220736 321618 220748
rect 324498 220736 324504 220748
rect 324556 220736 324562 220788
rect 385218 220736 385224 220788
rect 385276 220776 385282 220788
rect 388714 220776 388720 220788
rect 385276 220748 388720 220776
rect 385276 220736 385282 220748
rect 388714 220736 388720 220748
rect 388772 220736 388778 220788
rect 414198 220736 414204 220788
rect 414256 220776 414262 220788
rect 418154 220776 418160 220788
rect 414256 220748 418160 220776
rect 414256 220736 414262 220748
rect 418154 220736 418160 220748
rect 418212 220736 418218 220788
rect 455322 220736 455328 220788
rect 455380 220776 455386 220788
rect 458818 220776 458824 220788
rect 455380 220748 458824 220776
rect 455380 220736 455386 220748
rect 458818 220736 458824 220748
rect 458876 220736 458882 220788
rect 473998 220736 474004 220788
rect 474056 220776 474062 220788
rect 475378 220776 475384 220788
rect 474056 220748 475384 220776
rect 474056 220736 474062 220748
rect 475378 220736 475384 220748
rect 475436 220736 475442 220788
rect 476758 220736 476764 220788
rect 476816 220776 476822 220788
rect 478690 220776 478696 220788
rect 476816 220748 478696 220776
rect 476816 220736 476822 220748
rect 478690 220736 478696 220748
rect 478748 220736 478754 220788
rect 511810 220736 511816 220788
rect 511868 220776 511874 220788
rect 511868 220748 512040 220776
rect 511868 220736 511874 220748
rect 465718 220668 465724 220720
rect 465776 220708 465782 220720
rect 469582 220708 469588 220720
rect 465776 220680 469588 220708
rect 465776 220668 465782 220680
rect 469582 220668 469588 220680
rect 469640 220668 469646 220720
rect 512012 220708 512040 220748
rect 512012 220680 518894 220708
rect 147416 220612 147582 220640
rect 69750 220464 69756 220516
rect 69808 220504 69814 220516
rect 136910 220504 136916 220516
rect 69808 220476 136916 220504
rect 69808 220464 69814 220476
rect 136910 220464 136916 220476
rect 136968 220464 136974 220516
rect 137094 220464 137100 220516
rect 137152 220504 137158 220516
rect 147416 220504 147444 220612
rect 147674 220600 147680 220652
rect 147732 220640 147738 220652
rect 175274 220640 175280 220652
rect 147732 220612 175280 220640
rect 147732 220600 147738 220612
rect 175274 220600 175280 220612
rect 175332 220600 175338 220652
rect 177390 220600 177396 220652
rect 177448 220640 177454 220652
rect 180748 220640 180754 220652
rect 177448 220612 180754 220640
rect 177448 220600 177454 220612
rect 180748 220600 180754 220612
rect 180806 220600 180812 220652
rect 180886 220600 180892 220652
rect 180944 220640 180950 220652
rect 224218 220640 224224 220652
rect 180944 220612 224224 220640
rect 180944 220600 180950 220612
rect 224218 220600 224224 220612
rect 224276 220600 224282 220652
rect 253566 220600 253572 220652
rect 253624 220640 253630 220652
rect 293310 220640 293316 220652
rect 253624 220612 293316 220640
rect 253624 220600 253630 220612
rect 293310 220600 293316 220612
rect 293368 220600 293374 220652
rect 302418 220600 302424 220652
rect 302476 220640 302482 220652
rect 334066 220640 334072 220652
rect 302476 220612 334072 220640
rect 302476 220600 302482 220612
rect 334066 220600 334072 220612
rect 334124 220600 334130 220652
rect 357894 220600 357900 220652
rect 357952 220640 357958 220652
rect 374454 220640 374460 220652
rect 357952 220612 374460 220640
rect 357952 220600 357958 220612
rect 374454 220600 374460 220612
rect 374512 220600 374518 220652
rect 500218 220600 500224 220652
rect 500276 220640 500282 220652
rect 511810 220640 511816 220652
rect 500276 220612 511816 220640
rect 500276 220600 500282 220612
rect 511810 220600 511816 220612
rect 511868 220600 511874 220652
rect 137152 220476 147444 220504
rect 137152 220464 137158 220476
rect 147582 220464 147588 220516
rect 147640 220504 147646 220516
rect 150710 220504 150716 220516
rect 147640 220476 150716 220504
rect 147640 220464 147646 220476
rect 150710 220464 150716 220476
rect 150768 220464 150774 220516
rect 150894 220464 150900 220516
rect 150952 220504 150958 220516
rect 150952 220476 151814 220504
rect 150952 220464 150958 220476
rect 73062 220328 73068 220380
rect 73120 220368 73126 220380
rect 147214 220368 147220 220380
rect 73120 220340 147220 220368
rect 73120 220328 73126 220340
rect 147214 220328 147220 220340
rect 147272 220328 147278 220380
rect 147398 220328 147404 220380
rect 147456 220368 147462 220380
rect 151538 220368 151544 220380
rect 147456 220340 151544 220368
rect 147456 220328 147462 220340
rect 151538 220328 151544 220340
rect 151596 220328 151602 220380
rect 151786 220368 151814 220476
rect 151906 220464 151912 220516
rect 151964 220504 151970 220516
rect 211246 220504 211252 220516
rect 151964 220476 211252 220504
rect 151964 220464 151970 220476
rect 211246 220464 211252 220476
rect 211304 220464 211310 220516
rect 214098 220504 214104 220516
rect 211908 220476 214104 220504
rect 211908 220368 211936 220476
rect 214098 220464 214104 220476
rect 214156 220464 214162 220516
rect 214282 220464 214288 220516
rect 214340 220504 214346 220516
rect 218698 220504 218704 220516
rect 214340 220476 218704 220504
rect 214340 220464 214346 220476
rect 218698 220464 218704 220476
rect 218756 220464 218762 220516
rect 220446 220464 220452 220516
rect 220504 220504 220510 220516
rect 267918 220504 267924 220516
rect 220504 220476 267924 220504
rect 220504 220464 220510 220476
rect 267918 220464 267924 220476
rect 267976 220464 267982 220516
rect 273438 220464 273444 220516
rect 273496 220504 273502 220516
rect 309226 220504 309232 220516
rect 273496 220476 309232 220504
rect 273496 220464 273502 220476
rect 309226 220464 309232 220476
rect 309284 220464 309290 220516
rect 338022 220464 338028 220516
rect 338080 220504 338086 220516
rect 358998 220504 359004 220516
rect 338080 220476 359004 220504
rect 338080 220464 338086 220476
rect 358998 220464 359004 220476
rect 359056 220464 359062 220516
rect 432230 220464 432236 220516
rect 432288 220504 432294 220516
rect 434806 220504 434812 220516
rect 432288 220476 434812 220504
rect 432288 220464 432294 220476
rect 434806 220464 434812 220476
rect 434864 220464 434870 220516
rect 469122 220464 469128 220516
rect 469180 220504 469186 220516
rect 474550 220504 474556 220516
rect 469180 220476 474556 220504
rect 469180 220464 469186 220476
rect 474550 220464 474556 220476
rect 474608 220464 474614 220516
rect 488442 220464 488448 220516
rect 488500 220504 488506 220516
rect 501874 220504 501880 220516
rect 488500 220476 501880 220504
rect 488500 220464 488506 220476
rect 501874 220464 501880 220476
rect 501932 220464 501938 220516
rect 518866 220504 518894 220680
rect 545758 220668 545764 220720
rect 545816 220708 545822 220720
rect 547966 220708 547972 220720
rect 545816 220680 547972 220708
rect 545816 220668 545822 220680
rect 547966 220668 547972 220680
rect 548024 220668 548030 220720
rect 558730 220668 558736 220720
rect 558788 220708 558794 220720
rect 562962 220708 562968 220720
rect 558788 220680 562968 220708
rect 558788 220668 558794 220680
rect 562962 220668 562968 220680
rect 563020 220668 563026 220720
rect 563146 220668 563152 220720
rect 563204 220708 563210 220720
rect 566458 220708 566464 220720
rect 563204 220680 566464 220708
rect 563204 220668 563210 220680
rect 566458 220668 566464 220680
rect 566516 220668 566522 220720
rect 566826 220668 566832 220720
rect 566884 220708 566890 220720
rect 567286 220708 567292 220720
rect 566884 220680 567292 220708
rect 566884 220668 566890 220680
rect 567286 220668 567292 220680
rect 567344 220668 567350 220720
rect 520918 220600 520924 220652
rect 520976 220640 520982 220652
rect 537478 220640 537484 220652
rect 520976 220612 537484 220640
rect 520976 220600 520982 220612
rect 537478 220600 537484 220612
rect 537536 220600 537542 220652
rect 550818 220600 550824 220652
rect 550876 220640 550882 220652
rect 558546 220640 558552 220652
rect 550876 220612 558552 220640
rect 550876 220600 550882 220612
rect 558546 220600 558552 220612
rect 558604 220600 558610 220652
rect 568574 220600 568580 220652
rect 568632 220640 568638 220652
rect 569770 220640 569776 220652
rect 568632 220612 569776 220640
rect 568632 220600 568638 220612
rect 569770 220600 569776 220612
rect 569828 220600 569834 220652
rect 569954 220600 569960 220652
rect 570012 220640 570018 220652
rect 572438 220640 572444 220652
rect 570012 220612 572444 220640
rect 570012 220600 570018 220612
rect 572438 220600 572444 220612
rect 572496 220600 572502 220652
rect 572622 220600 572628 220652
rect 572680 220640 572686 220652
rect 610526 220640 610532 220652
rect 572680 220612 610532 220640
rect 572680 220600 572686 220612
rect 610526 220600 610532 220612
rect 610584 220600 610590 220652
rect 563026 220544 563284 220572
rect 531682 220504 531688 220516
rect 518866 220476 531688 220504
rect 531682 220464 531688 220476
rect 531740 220464 531746 220516
rect 548334 220464 548340 220516
rect 548392 220504 548398 220516
rect 563026 220504 563054 220544
rect 548392 220476 563054 220504
rect 563256 220504 563284 220544
rect 598566 220504 598572 220516
rect 563256 220476 598572 220504
rect 548392 220464 548398 220476
rect 598566 220464 598572 220476
rect 598624 220464 598630 220516
rect 600958 220464 600964 220516
rect 601016 220504 601022 220516
rect 611446 220504 611452 220516
rect 601016 220476 611452 220504
rect 601016 220464 601022 220476
rect 611446 220464 611452 220476
rect 611504 220464 611510 220516
rect 151786 220340 211936 220368
rect 213638 220328 213644 220380
rect 213696 220368 213702 220380
rect 213696 220340 224264 220368
rect 213696 220328 213702 220340
rect 79686 220192 79692 220244
rect 79744 220232 79750 220244
rect 151722 220232 151728 220244
rect 79744 220204 151728 220232
rect 79744 220192 79750 220204
rect 151722 220192 151728 220204
rect 151780 220192 151786 220244
rect 151906 220192 151912 220244
rect 151964 220232 151970 220244
rect 154022 220232 154028 220244
rect 151964 220204 154028 220232
rect 151964 220192 151970 220204
rect 154022 220192 154028 220204
rect 154080 220192 154086 220244
rect 154390 220192 154396 220244
rect 154448 220232 154454 220244
rect 158898 220232 158904 220244
rect 154448 220204 158904 220232
rect 154448 220192 154454 220204
rect 158898 220192 158904 220204
rect 158956 220192 158962 220244
rect 164234 220192 164240 220244
rect 164292 220232 164298 220244
rect 223758 220232 223764 220244
rect 164292 220204 223764 220232
rect 164292 220192 164298 220204
rect 223758 220192 223764 220204
rect 223816 220192 223822 220244
rect 224236 220232 224264 220340
rect 224402 220328 224408 220380
rect 224460 220368 224466 220380
rect 265158 220368 265164 220380
rect 224460 220340 265164 220368
rect 224460 220328 224466 220340
rect 265158 220328 265164 220340
rect 265216 220328 265222 220380
rect 267642 220328 267648 220380
rect 267700 220368 267706 220380
rect 306926 220368 306932 220380
rect 267700 220340 306932 220368
rect 267700 220328 267706 220340
rect 306926 220328 306932 220340
rect 306984 220328 306990 220380
rect 314838 220328 314844 220380
rect 314896 220368 314902 220380
rect 341058 220368 341064 220380
rect 314896 220340 341064 220368
rect 314896 220328 314902 220340
rect 341058 220328 341064 220340
rect 341116 220328 341122 220380
rect 342990 220328 342996 220380
rect 343048 220368 343054 220380
rect 363414 220368 363420 220380
rect 343048 220340 363420 220368
rect 343048 220328 343054 220340
rect 363414 220328 363420 220340
rect 363472 220328 363478 220380
rect 472986 220328 472992 220380
rect 473044 220368 473050 220380
rect 481174 220368 481180 220380
rect 473044 220340 481180 220368
rect 473044 220328 473050 220340
rect 481174 220328 481180 220340
rect 481232 220328 481238 220380
rect 496446 220328 496452 220380
rect 496504 220368 496510 220380
rect 509326 220368 509332 220380
rect 496504 220340 509332 220368
rect 496504 220328 496510 220340
rect 509326 220328 509332 220340
rect 509384 220328 509390 220380
rect 516962 220328 516968 220380
rect 517020 220368 517026 220380
rect 527542 220368 527548 220380
rect 517020 220340 527548 220368
rect 517020 220328 517026 220340
rect 527542 220328 527548 220340
rect 527600 220328 527606 220380
rect 531130 220328 531136 220380
rect 531188 220368 531194 220380
rect 556522 220368 556528 220380
rect 531188 220340 556528 220368
rect 531188 220328 531194 220340
rect 556522 220328 556528 220340
rect 556580 220328 556586 220380
rect 563192 220368 563198 220380
rect 558196 220340 563198 220368
rect 234154 220232 234160 220244
rect 224236 220204 234160 220232
rect 234154 220192 234160 220204
rect 234212 220192 234218 220244
rect 237006 220192 237012 220244
rect 237064 220232 237070 220244
rect 280430 220232 280436 220244
rect 237064 220204 280436 220232
rect 237064 220192 237070 220204
rect 280430 220192 280436 220204
rect 280488 220192 280494 220244
rect 283374 220192 283380 220244
rect 283432 220232 283438 220244
rect 316310 220232 316316 220244
rect 283432 220204 316316 220232
rect 283432 220192 283438 220204
rect 316310 220192 316316 220204
rect 316368 220192 316374 220244
rect 316494 220192 316500 220244
rect 316552 220232 316558 220244
rect 342622 220232 342628 220244
rect 316552 220204 342628 220232
rect 316552 220192 316558 220204
rect 342622 220192 342628 220204
rect 342680 220192 342686 220244
rect 348786 220192 348792 220244
rect 348844 220232 348850 220244
rect 369946 220232 369952 220244
rect 348844 220204 369952 220232
rect 348844 220192 348850 220204
rect 369946 220192 369952 220204
rect 370004 220192 370010 220244
rect 370498 220192 370504 220244
rect 370556 220232 370562 220244
rect 381078 220232 381084 220244
rect 370556 220204 381084 220232
rect 370556 220192 370562 220204
rect 381078 220192 381084 220204
rect 381136 220192 381142 220244
rect 388714 220192 388720 220244
rect 388772 220232 388778 220244
rect 400950 220232 400956 220244
rect 388772 220204 400956 220232
rect 388772 220192 388778 220204
rect 400950 220192 400956 220204
rect 401008 220192 401014 220244
rect 459462 220192 459468 220244
rect 459520 220232 459526 220244
rect 465442 220232 465448 220244
rect 459520 220204 465448 220232
rect 459520 220192 459526 220204
rect 465442 220192 465448 220204
rect 465500 220192 465506 220244
rect 473170 220192 473176 220244
rect 473228 220232 473234 220244
rect 482002 220232 482008 220244
rect 473228 220204 482008 220232
rect 473228 220192 473234 220204
rect 482002 220192 482008 220204
rect 482060 220192 482066 220244
rect 482922 220192 482928 220244
rect 482980 220232 482986 220244
rect 495250 220232 495256 220244
rect 482980 220204 495256 220232
rect 482980 220192 482986 220204
rect 495250 220192 495256 220204
rect 495308 220192 495314 220244
rect 501322 220192 501328 220244
rect 501380 220232 501386 220244
rect 520182 220232 520188 220244
rect 501380 220204 520188 220232
rect 501380 220192 501386 220204
rect 520182 220192 520188 220204
rect 520240 220192 520246 220244
rect 528370 220192 528376 220244
rect 528428 220232 528434 220244
rect 554038 220232 554044 220244
rect 528428 220204 554044 220232
rect 528428 220192 528434 220204
rect 554038 220192 554044 220204
rect 554096 220192 554102 220244
rect 555694 220192 555700 220244
rect 555752 220232 555758 220244
rect 557994 220232 558000 220244
rect 555752 220204 558000 220232
rect 555752 220192 555758 220204
rect 557994 220192 558000 220204
rect 558052 220192 558058 220244
rect 76374 220056 76380 220108
rect 76432 220096 76438 220108
rect 156138 220096 156144 220108
rect 76432 220068 156144 220096
rect 76432 220056 76438 220068
rect 156138 220056 156144 220068
rect 156196 220056 156202 220108
rect 157518 220056 157524 220108
rect 157576 220096 157582 220108
rect 214282 220096 214288 220108
rect 157576 220068 214288 220096
rect 157576 220056 157582 220068
rect 214282 220056 214288 220068
rect 214340 220056 214346 220108
rect 244274 220096 244280 220108
rect 214576 220068 244280 220096
rect 107838 219920 107844 219972
rect 107896 219960 107902 219972
rect 114278 219960 114284 219972
rect 107896 219932 114284 219960
rect 107896 219920 107902 219932
rect 114278 219920 114284 219932
rect 114336 219920 114342 219972
rect 114462 219920 114468 219972
rect 114520 219960 114526 219972
rect 114520 219932 126744 219960
rect 114520 219920 114526 219932
rect 121086 219784 121092 219836
rect 121144 219824 121150 219836
rect 126716 219824 126744 219932
rect 127618 219920 127624 219972
rect 127676 219960 127682 219972
rect 180748 219960 180754 219972
rect 127676 219932 180754 219960
rect 127676 219920 127682 219932
rect 180748 219920 180754 219932
rect 180806 219920 180812 219972
rect 180886 219920 180892 219972
rect 180944 219960 180950 219972
rect 213638 219960 213644 219972
rect 180944 219932 213644 219960
rect 180944 219920 180950 219932
rect 213638 219920 213644 219932
rect 213696 219920 213702 219972
rect 137094 219824 137100 219836
rect 121144 219796 122834 219824
rect 126716 219796 137100 219824
rect 121144 219784 121150 219796
rect 122806 219688 122834 219796
rect 137094 219784 137100 219796
rect 137152 219784 137158 219836
rect 197630 219824 197636 219836
rect 137296 219796 197636 219824
rect 127618 219688 127624 219700
rect 122806 219660 127624 219688
rect 127618 219648 127624 219660
rect 127676 219648 127682 219700
rect 131022 219648 131028 219700
rect 131080 219688 131086 219700
rect 137296 219688 137324 219796
rect 197630 219784 197636 219796
rect 197688 219784 197694 219836
rect 197814 219784 197820 219836
rect 197872 219824 197878 219836
rect 214576 219824 214604 220068
rect 244274 220056 244280 220068
rect 244332 220056 244338 220108
rect 244458 220056 244464 220108
rect 244516 220096 244522 220108
rect 288526 220096 288532 220108
rect 244516 220068 288532 220096
rect 244516 220056 244522 220068
rect 288526 220056 288532 220068
rect 288584 220056 288590 220108
rect 288710 220056 288716 220108
rect 288768 220096 288774 220108
rect 322382 220096 322388 220108
rect 288768 220068 322388 220096
rect 288768 220056 288774 220068
rect 322382 220056 322388 220068
rect 322440 220056 322446 220108
rect 325602 220056 325608 220108
rect 325660 220096 325666 220108
rect 352098 220096 352104 220108
rect 325660 220068 352104 220096
rect 325660 220056 325666 220068
rect 352098 220056 352104 220068
rect 352156 220056 352162 220108
rect 358814 220056 358820 220108
rect 358872 220096 358878 220108
rect 378318 220096 378324 220108
rect 358872 220068 378324 220096
rect 358872 220056 358878 220068
rect 378318 220056 378324 220068
rect 378376 220056 378382 220108
rect 379422 220056 379428 220108
rect 379480 220096 379486 220108
rect 392118 220096 392124 220108
rect 379480 220068 392124 220096
rect 379480 220056 379486 220068
rect 392118 220056 392124 220068
rect 392176 220056 392182 220108
rect 395982 220056 395988 220108
rect 396040 220096 396046 220108
rect 404814 220096 404820 220108
rect 396040 220068 404820 220096
rect 396040 220056 396046 220068
rect 404814 220056 404820 220068
rect 404872 220056 404878 220108
rect 421650 220056 421656 220108
rect 421708 220096 421714 220108
rect 426710 220096 426716 220108
rect 421708 220068 426716 220096
rect 421708 220056 421714 220068
rect 426710 220056 426716 220068
rect 426768 220056 426774 220108
rect 478322 220056 478328 220108
rect 478380 220096 478386 220108
rect 489454 220096 489460 220108
rect 478380 220068 489460 220096
rect 478380 220056 478386 220068
rect 489454 220056 489460 220068
rect 489512 220056 489518 220108
rect 492490 220056 492496 220108
rect 492548 220096 492554 220108
rect 506842 220096 506848 220108
rect 492548 220068 506848 220096
rect 492548 220056 492554 220068
rect 506842 220056 506848 220068
rect 506900 220056 506906 220108
rect 513098 220056 513104 220108
rect 513156 220096 513162 220108
rect 534166 220096 534172 220108
rect 513156 220068 534172 220096
rect 513156 220056 513162 220068
rect 534166 220056 534172 220068
rect 534224 220056 534230 220108
rect 538122 220056 538128 220108
rect 538180 220096 538186 220108
rect 558196 220096 558224 220340
rect 563192 220328 563198 220340
rect 563250 220328 563256 220380
rect 563330 220328 563336 220380
rect 563388 220368 563394 220380
rect 609422 220368 609428 220380
rect 563388 220340 609428 220368
rect 563388 220328 563394 220340
rect 609422 220328 609428 220340
rect 609480 220328 609486 220380
rect 558362 220192 558368 220244
rect 558420 220232 558426 220244
rect 562870 220232 562876 220244
rect 558420 220204 562876 220232
rect 558420 220192 558426 220204
rect 562870 220192 562876 220204
rect 562928 220192 562934 220244
rect 563054 220192 563060 220244
rect 563112 220232 563118 220244
rect 608870 220232 608876 220244
rect 563112 220204 608876 220232
rect 563112 220192 563118 220204
rect 608870 220192 608876 220204
rect 608928 220192 608934 220244
rect 648614 220192 648620 220244
rect 648672 220232 648678 220244
rect 652754 220232 652760 220244
rect 648672 220204 652760 220232
rect 648672 220192 648678 220204
rect 652754 220192 652760 220204
rect 652812 220192 652818 220244
rect 538180 220068 558224 220096
rect 538180 220056 538186 220068
rect 572668 220056 572674 220108
rect 572726 220096 572732 220108
rect 572726 220068 598428 220096
rect 572726 220056 572732 220068
rect 558362 219988 558368 220040
rect 558420 220028 558426 220040
rect 572530 220028 572536 220040
rect 558420 220000 572536 220028
rect 558420 219988 558426 220000
rect 572530 219988 572536 220000
rect 572588 219988 572594 220040
rect 214742 219920 214748 219972
rect 214800 219960 214806 219972
rect 254762 219960 254768 219972
rect 214800 219932 254768 219960
rect 214800 219920 214806 219932
rect 254762 219920 254768 219932
rect 254820 219920 254826 219972
rect 294966 219920 294972 219972
rect 295024 219960 295030 219972
rect 325878 219960 325884 219972
rect 295024 219932 325884 219960
rect 295024 219920 295030 219932
rect 325878 219920 325884 219932
rect 325936 219920 325942 219972
rect 598400 219960 598428 220068
rect 598566 220056 598572 220108
rect 598624 220096 598630 220108
rect 607306 220096 607312 220108
rect 598624 220068 607312 220096
rect 598624 220056 598630 220068
rect 607306 220056 607312 220068
rect 607364 220056 607370 220108
rect 676214 220056 676220 220108
rect 676272 220096 676278 220108
rect 677318 220096 677324 220108
rect 676272 220068 677324 220096
rect 676272 220056 676278 220068
rect 677318 220056 677324 220068
rect 677376 220056 677382 220108
rect 600958 219960 600964 219972
rect 598400 219932 600964 219960
rect 600958 219920 600964 219932
rect 601016 219920 601022 219972
rect 503622 219852 503628 219904
rect 503680 219892 503686 219904
rect 589274 219892 589280 219904
rect 503680 219864 589280 219892
rect 503680 219852 503686 219864
rect 589274 219852 589280 219864
rect 589332 219852 589338 219904
rect 589458 219852 589464 219904
rect 589516 219892 589522 219904
rect 596726 219892 596732 219904
rect 589516 219864 596732 219892
rect 589516 219852 589522 219864
rect 596726 219852 596732 219864
rect 596784 219852 596790 219904
rect 259914 219824 259920 219836
rect 197872 219796 214604 219824
rect 214760 219796 259920 219824
rect 197872 219784 197878 219796
rect 131080 219660 137324 219688
rect 137388 219660 142936 219688
rect 131080 219648 131086 219660
rect 136910 219512 136916 219564
rect 136968 219552 136974 219564
rect 137388 219552 137416 219660
rect 136968 219524 137416 219552
rect 136968 219512 136974 219524
rect 137646 219512 137652 219564
rect 137704 219552 137710 219564
rect 142706 219552 142712 219564
rect 137704 219524 142712 219552
rect 137704 219512 137710 219524
rect 142706 219512 142712 219524
rect 142764 219512 142770 219564
rect 142908 219552 142936 219660
rect 143074 219648 143080 219700
rect 143132 219688 143138 219700
rect 203150 219688 203156 219700
rect 143132 219660 203156 219688
rect 143132 219648 143138 219660
rect 203150 219648 203156 219660
rect 203208 219648 203214 219700
rect 208578 219688 208584 219700
rect 203720 219660 208584 219688
rect 144086 219552 144092 219564
rect 142908 219524 144092 219552
rect 144086 219512 144092 219524
rect 144144 219512 144150 219564
rect 144270 219512 144276 219564
rect 144328 219552 144334 219564
rect 203720 219552 203748 219660
rect 208578 219648 208584 219660
rect 208636 219648 208642 219700
rect 210510 219648 210516 219700
rect 210568 219688 210574 219700
rect 214760 219688 214788 219796
rect 259914 219784 259920 219796
rect 259972 219784 259978 219836
rect 540790 219716 540796 219768
rect 540848 219756 540854 219768
rect 606018 219756 606024 219768
rect 540848 219728 606024 219756
rect 540848 219716 540854 219728
rect 606018 219716 606024 219728
rect 606076 219716 606082 219768
rect 210568 219660 214788 219688
rect 210568 219648 210574 219660
rect 217134 219648 217140 219700
rect 217192 219688 217198 219700
rect 224402 219688 224408 219700
rect 217192 219660 224408 219688
rect 217192 219648 217198 219660
rect 224402 219648 224408 219660
rect 224460 219648 224466 219700
rect 227070 219648 227076 219700
rect 227128 219688 227134 219700
rect 272702 219688 272708 219700
rect 227128 219660 272708 219688
rect 227128 219648 227134 219660
rect 272702 219648 272708 219660
rect 272760 219648 272766 219700
rect 464982 219580 464988 219632
rect 465040 219620 465046 219632
rect 472066 219620 472072 219632
rect 465040 219592 472072 219620
rect 465040 219580 465046 219592
rect 472066 219580 472072 219592
rect 472124 219580 472130 219632
rect 527542 219580 527548 219632
rect 527600 219620 527606 219632
rect 558362 219620 558368 219632
rect 527600 219592 558368 219620
rect 527600 219580 527606 219592
rect 558362 219580 558368 219592
rect 558420 219580 558426 219632
rect 558546 219580 558552 219632
rect 558604 219620 558610 219632
rect 600866 219620 600872 219632
rect 558604 219592 600872 219620
rect 558604 219580 558610 219592
rect 600866 219580 600872 219592
rect 600924 219580 600930 219632
rect 620094 219620 620100 219632
rect 601068 219592 620100 219620
rect 144328 219524 203748 219552
rect 144328 219512 144334 219524
rect 203886 219512 203892 219564
rect 203944 219552 203950 219564
rect 214742 219552 214748 219564
rect 203944 219524 214748 219552
rect 203944 219512 203950 219524
rect 214742 219512 214748 219524
rect 214800 219512 214806 219564
rect 224218 219512 224224 219564
rect 224276 219552 224282 219564
rect 229278 219552 229284 219564
rect 224276 219524 229284 219552
rect 224276 219512 224282 219524
rect 229278 219512 229284 219524
rect 229336 219512 229342 219564
rect 332686 219512 332692 219564
rect 332744 219552 332750 219564
rect 337194 219552 337200 219564
rect 332744 219524 337200 219552
rect 332744 219512 332750 219524
rect 337194 219512 337200 219524
rect 337252 219512 337258 219564
rect 432046 219552 432052 219564
rect 431926 219524 432052 219552
rect 240152 219456 241514 219484
rect 109494 219376 109500 219428
rect 109552 219416 109558 219428
rect 110414 219416 110420 219428
rect 109552 219388 110420 219416
rect 109552 219376 109558 219388
rect 110414 219376 110420 219388
rect 110472 219376 110478 219428
rect 113634 219376 113640 219428
rect 113692 219416 113698 219428
rect 156506 219416 156512 219428
rect 113692 219388 156512 219416
rect 113692 219376 113698 219388
rect 156506 219376 156512 219388
rect 156564 219376 156570 219428
rect 165798 219376 165804 219428
rect 165856 219416 165862 219428
rect 165856 219388 171134 219416
rect 165856 219376 165862 219388
rect 70578 219240 70584 219292
rect 70636 219280 70642 219292
rect 117774 219280 117780 219292
rect 70636 219252 117780 219280
rect 70636 219240 70642 219252
rect 117774 219240 117780 219252
rect 117832 219240 117838 219292
rect 131850 219240 131856 219292
rect 131908 219280 131914 219292
rect 132402 219280 132408 219292
rect 131908 219252 132408 219280
rect 131908 219240 131914 219252
rect 132402 219240 132408 219252
rect 132460 219240 132466 219292
rect 132586 219240 132592 219292
rect 132644 219280 132650 219292
rect 136174 219280 136180 219292
rect 132644 219252 136180 219280
rect 132644 219240 132650 219252
rect 136174 219240 136180 219252
rect 136232 219240 136238 219292
rect 136358 219240 136364 219292
rect 136416 219280 136422 219292
rect 170950 219280 170956 219292
rect 136416 219252 170956 219280
rect 136416 219240 136422 219252
rect 170950 219240 170956 219252
rect 171008 219240 171014 219292
rect 171106 219280 171134 219388
rect 175734 219376 175740 219428
rect 175792 219416 175798 219428
rect 181438 219416 181444 219428
rect 175792 219388 181444 219416
rect 175792 219376 175798 219388
rect 181438 219376 181444 219388
rect 181496 219376 181502 219428
rect 183830 219376 183836 219428
rect 183888 219416 183894 219428
rect 189994 219416 190000 219428
rect 183888 219388 190000 219416
rect 183888 219376 183894 219388
rect 189994 219376 190000 219388
rect 190052 219376 190058 219428
rect 192294 219376 192300 219428
rect 192352 219416 192358 219428
rect 224402 219416 224408 219428
rect 192352 219388 224408 219416
rect 192352 219376 192358 219388
rect 224402 219376 224408 219388
rect 224460 219376 224466 219428
rect 229554 219376 229560 219428
rect 229612 219416 229618 219428
rect 230474 219416 230480 219428
rect 229612 219388 230480 219416
rect 229612 219376 229618 219388
rect 230474 219376 230480 219388
rect 230532 219376 230538 219428
rect 237834 219376 237840 219428
rect 237892 219416 237898 219428
rect 239306 219416 239312 219428
rect 237892 219388 239312 219416
rect 237892 219376 237898 219388
rect 239306 219376 239312 219388
rect 239364 219376 239370 219428
rect 239490 219376 239496 219428
rect 239548 219416 239554 219428
rect 240152 219416 240180 219456
rect 239548 219388 240180 219416
rect 241486 219416 241514 219456
rect 405918 219444 405924 219496
rect 405976 219484 405982 219496
rect 412726 219484 412732 219496
rect 405976 219456 412732 219484
rect 405976 219444 405982 219456
rect 412726 219444 412732 219456
rect 412784 219444 412790 219496
rect 421006 219484 421012 219496
rect 418172 219456 421012 219484
rect 241790 219416 241796 219428
rect 241486 219388 241796 219416
rect 239548 219376 239554 219388
rect 241790 219376 241796 219388
rect 241848 219376 241854 219428
rect 241974 219376 241980 219428
rect 242032 219416 242038 219428
rect 242894 219416 242900 219428
rect 242032 219388 242900 219416
rect 242032 219376 242038 219388
rect 242894 219376 242900 219388
rect 242952 219376 242958 219428
rect 244918 219376 244924 219428
rect 244976 219416 244982 219428
rect 272334 219416 272340 219428
rect 244976 219388 272340 219416
rect 244976 219376 244982 219388
rect 272334 219376 272340 219388
rect 272392 219376 272398 219428
rect 272702 219376 272708 219428
rect 272760 219416 272766 219428
rect 272760 219388 277394 219416
rect 272760 219376 272766 219388
rect 180058 219280 180064 219292
rect 171106 219252 180064 219280
rect 180058 219240 180064 219252
rect 180116 219240 180122 219292
rect 180242 219240 180248 219292
rect 180300 219280 180306 219292
rect 215938 219280 215944 219292
rect 180300 219252 215944 219280
rect 180300 219240 180306 219252
rect 215938 219240 215944 219252
rect 215996 219240 216002 219292
rect 219618 219240 219624 219292
rect 219676 219280 219682 219292
rect 264146 219280 264152 219292
rect 219676 219252 264152 219280
rect 219676 219240 219682 219252
rect 264146 219240 264152 219252
rect 264204 219240 264210 219292
rect 277366 219280 277394 219388
rect 285858 219376 285864 219428
rect 285916 219416 285922 219428
rect 285916 219388 306374 219416
rect 285916 219376 285922 219388
rect 301958 219280 301964 219292
rect 277366 219252 301964 219280
rect 301958 219240 301964 219252
rect 302016 219240 302022 219292
rect 306346 219280 306374 219388
rect 308214 219376 308220 219428
rect 308272 219416 308278 219428
rect 309134 219416 309140 219428
rect 308272 219388 309140 219416
rect 308272 219376 308278 219388
rect 309134 219376 309140 219388
rect 309192 219376 309198 219428
rect 333698 219376 333704 219428
rect 333756 219416 333762 219428
rect 347222 219416 347228 219428
rect 333756 219388 347228 219416
rect 333756 219376 333762 219388
rect 347222 219376 347228 219388
rect 347280 219376 347286 219428
rect 349614 219376 349620 219428
rect 349672 219416 349678 219428
rect 350534 219416 350540 219428
rect 349672 219388 350540 219416
rect 349672 219376 349678 219388
rect 350534 219376 350540 219388
rect 350592 219376 350598 219428
rect 352098 219376 352104 219428
rect 352156 219416 352162 219428
rect 355318 219416 355324 219428
rect 352156 219388 355324 219416
rect 352156 219376 352162 219388
rect 355318 219376 355324 219388
rect 355376 219376 355382 219428
rect 362034 219376 362040 219428
rect 362092 219416 362098 219428
rect 367646 219416 367652 219428
rect 362092 219388 367652 219416
rect 362092 219376 362098 219388
rect 367646 219376 367652 219388
rect 367704 219376 367710 219428
rect 380250 219376 380256 219428
rect 380308 219416 380314 219428
rect 384206 219416 384212 219428
rect 380308 219388 384212 219416
rect 380308 219376 380314 219388
rect 384206 219376 384212 219388
rect 384264 219376 384270 219428
rect 399294 219376 399300 219428
rect 399352 219416 399358 219428
rect 400214 219416 400220 219428
rect 399352 219388 400220 219416
rect 399352 219376 399358 219388
rect 400214 219376 400220 219388
rect 400272 219376 400278 219428
rect 415854 219376 415860 219428
rect 415912 219416 415918 219428
rect 416774 219416 416780 219428
rect 415912 219388 416780 219416
rect 415912 219376 415918 219388
rect 416774 219376 416780 219388
rect 416832 219376 416838 219428
rect 417510 219376 417516 219428
rect 417568 219416 417574 219428
rect 418172 219416 418200 219456
rect 421006 219444 421012 219456
rect 421064 219444 421070 219496
rect 431926 219484 431954 219524
rect 432046 219512 432052 219524
rect 432104 219512 432110 219564
rect 501138 219512 501144 219564
rect 501196 219552 501202 219564
rect 501196 219524 509234 219552
rect 501196 219512 501202 219524
rect 429212 219456 431954 219484
rect 509206 219484 509234 219524
rect 589090 219484 589096 219496
rect 509206 219456 589096 219484
rect 417568 219388 418200 219416
rect 417568 219376 417574 219388
rect 428274 219376 428280 219428
rect 428332 219416 428338 219428
rect 429212 219416 429240 219456
rect 589090 219444 589096 219456
rect 589148 219444 589154 219496
rect 601068 219484 601096 219592
rect 620094 219580 620100 219592
rect 620152 219580 620158 219632
rect 589246 219456 601096 219484
rect 428332 219388 429240 219416
rect 428332 219376 428338 219388
rect 438210 219376 438216 219428
rect 438268 219416 438274 219428
rect 438854 219416 438860 219428
rect 438268 219388 438860 219416
rect 438268 219376 438274 219388
rect 438854 219376 438860 219388
rect 438912 219376 438918 219428
rect 439866 219376 439872 219428
rect 439924 219416 439930 219428
rect 440326 219416 440332 219428
rect 439924 219388 440332 219416
rect 439924 219376 439930 219388
rect 440326 219376 440332 219388
rect 440384 219376 440390 219428
rect 572668 219308 572674 219360
rect 572726 219348 572732 219360
rect 589246 219348 589274 219456
rect 601234 219444 601240 219496
rect 601292 219484 601298 219496
rect 607490 219484 607496 219496
rect 601292 219456 607496 219484
rect 601292 219444 601298 219456
rect 607490 219444 607496 219456
rect 607548 219444 607554 219496
rect 572726 219320 589274 219348
rect 572726 219308 572732 219320
rect 313918 219280 313924 219292
rect 306346 219252 313924 219280
rect 313918 219240 313924 219252
rect 313976 219240 313982 219292
rect 320634 219240 320640 219292
rect 320692 219280 320698 219292
rect 342806 219280 342812 219292
rect 320692 219252 342812 219280
rect 320692 219240 320698 219252
rect 342806 219240 342812 219252
rect 342864 219240 342870 219292
rect 419166 219240 419172 219292
rect 419224 219280 419230 219292
rect 422662 219280 422668 219292
rect 419224 219252 422668 219280
rect 419224 219240 419230 219252
rect 422662 219240 422668 219252
rect 422720 219240 422726 219292
rect 548150 219240 548156 219292
rect 548208 219280 548214 219292
rect 563054 219280 563060 219292
rect 548208 219252 563060 219280
rect 548208 219240 548214 219252
rect 563054 219240 563060 219252
rect 563112 219240 563118 219292
rect 563238 219240 563244 219292
rect 563296 219280 563302 219292
rect 563296 219252 572300 219280
rect 563296 219240 563302 219252
rect 572272 219212 572300 219252
rect 574370 219212 574376 219224
rect 572272 219184 574376 219212
rect 574370 219172 574376 219184
rect 574428 219172 574434 219224
rect 589274 219172 589280 219224
rect 589332 219212 589338 219224
rect 597554 219212 597560 219224
rect 589332 219184 597560 219212
rect 589332 219172 589338 219184
rect 597554 219172 597560 219184
rect 597612 219172 597618 219224
rect 64598 219104 64604 219156
rect 64656 219144 64662 219156
rect 66898 219144 66904 219156
rect 64656 219116 66904 219144
rect 64656 219104 64662 219116
rect 66898 219104 66904 219116
rect 66956 219104 66962 219156
rect 93578 219104 93584 219156
rect 93636 219144 93642 219156
rect 94406 219144 94412 219156
rect 93636 219116 94412 219144
rect 93636 219104 93642 219116
rect 94406 219104 94412 219116
rect 94464 219104 94470 219156
rect 117958 219104 117964 219156
rect 118016 219144 118022 219156
rect 154666 219144 154672 219156
rect 118016 219116 154672 219144
rect 118016 219104 118022 219116
rect 154666 219104 154672 219116
rect 154724 219104 154730 219156
rect 157978 219144 157984 219156
rect 154868 219116 157984 219144
rect 62298 218968 62304 219020
rect 62356 219008 62362 219020
rect 72418 219008 72424 219020
rect 62356 218980 72424 219008
rect 62356 218968 62362 218980
rect 72418 218968 72424 218980
rect 72476 218968 72482 219020
rect 83826 218968 83832 219020
rect 83884 219008 83890 219020
rect 154868 219008 154896 219116
rect 157978 219104 157984 219116
rect 158036 219104 158042 219156
rect 166626 219104 166632 219156
rect 166684 219144 166690 219156
rect 208486 219144 208492 219156
rect 166684 219116 208492 219144
rect 166684 219104 166690 219116
rect 208486 219104 208492 219116
rect 208544 219104 208550 219156
rect 208854 219104 208860 219156
rect 208912 219144 208918 219156
rect 209682 219144 209688 219156
rect 208912 219116 209688 219144
rect 208912 219104 208918 219116
rect 209682 219104 209688 219116
rect 209740 219104 209746 219156
rect 218790 219104 218796 219156
rect 218848 219144 218854 219156
rect 219342 219144 219348 219156
rect 218848 219116 219348 219144
rect 218848 219104 218854 219116
rect 219342 219104 219348 219116
rect 219400 219104 219406 219156
rect 224218 219104 224224 219156
rect 224276 219144 224282 219156
rect 253014 219144 253020 219156
rect 224276 219116 253020 219144
rect 224276 219104 224282 219116
rect 253014 219104 253020 219116
rect 253072 219104 253078 219156
rect 265986 219104 265992 219156
rect 266044 219144 266050 219156
rect 266044 219116 291884 219144
rect 266044 219104 266050 219116
rect 83884 218980 154896 219008
rect 83884 218968 83890 218980
rect 156506 218968 156512 219020
rect 156564 219008 156570 219020
rect 162118 219008 162124 219020
rect 156564 218980 162124 219008
rect 156564 218968 156570 218980
rect 162118 218968 162124 218980
rect 162176 218968 162182 219020
rect 162486 218968 162492 219020
rect 162544 219008 162550 219020
rect 175734 219008 175740 219020
rect 162544 218980 175740 219008
rect 162544 218968 162550 218980
rect 175734 218968 175740 218980
rect 175792 218968 175798 219020
rect 176654 218968 176660 219020
rect 176712 219008 176718 219020
rect 180242 219008 180248 219020
rect 176712 218980 180248 219008
rect 176712 218968 176718 218980
rect 180242 218968 180248 218980
rect 180300 218968 180306 219020
rect 182358 218968 182364 219020
rect 182416 219008 182422 219020
rect 189718 219008 189724 219020
rect 182416 218980 189724 219008
rect 182416 218968 182422 218980
rect 189718 218968 189724 218980
rect 189776 218968 189782 219020
rect 190638 218968 190644 219020
rect 190696 219008 190702 219020
rect 197814 219008 197820 219020
rect 190696 218980 197820 219008
rect 190696 218968 190702 218980
rect 197814 218968 197820 218980
rect 197872 218968 197878 219020
rect 200206 218968 200212 219020
rect 200264 219008 200270 219020
rect 241606 219008 241612 219020
rect 200264 218980 241612 219008
rect 200264 218968 200270 218980
rect 241606 218968 241612 218980
rect 241664 218968 241670 219020
rect 241790 218968 241796 219020
rect 241848 219008 241854 219020
rect 244918 219008 244924 219020
rect 241848 218980 244924 219008
rect 241848 218968 241854 218980
rect 244918 218968 244924 218980
rect 244976 218968 244982 219020
rect 252738 218968 252744 219020
rect 252796 219008 252802 219020
rect 287882 219008 287888 219020
rect 252796 218980 287888 219008
rect 252796 218968 252802 218980
rect 287882 218968 287888 218980
rect 287940 218968 287946 219020
rect 291856 219008 291884 219116
rect 295794 219104 295800 219156
rect 295852 219144 295858 219156
rect 296714 219144 296720 219156
rect 295852 219116 296720 219144
rect 295852 219104 295858 219116
rect 296714 219104 296720 219116
rect 296772 219104 296778 219156
rect 314010 219104 314016 219156
rect 314068 219144 314074 219156
rect 335998 219144 336004 219156
rect 314068 219116 336004 219144
rect 314068 219104 314074 219116
rect 335998 219104 336004 219116
rect 336056 219104 336062 219156
rect 343818 219104 343824 219156
rect 343876 219144 343882 219156
rect 353938 219144 353944 219156
rect 343876 219116 353944 219144
rect 343876 219104 343882 219116
rect 353938 219104 353944 219116
rect 353996 219104 354002 219156
rect 542630 219104 542636 219156
rect 542688 219144 542694 219156
rect 562870 219144 562876 219156
rect 542688 219116 548564 219144
rect 542688 219104 542694 219116
rect 297266 219008 297272 219020
rect 291856 218980 297272 219008
rect 297266 218968 297272 218980
rect 297324 218968 297330 219020
rect 307386 218968 307392 219020
rect 307444 219008 307450 219020
rect 332686 219008 332692 219020
rect 307444 218980 332692 219008
rect 307444 218968 307450 218980
rect 332686 218968 332692 218980
rect 332744 218968 332750 219020
rect 337194 218968 337200 219020
rect 337252 219008 337258 219020
rect 345658 219008 345664 219020
rect 337252 218980 345664 219008
rect 337252 218968 337258 218980
rect 345658 218968 345664 218980
rect 345716 218968 345722 219020
rect 347222 218968 347228 219020
rect 347280 219008 347286 219020
rect 363598 219008 363604 219020
rect 347280 218980 363604 219008
rect 347280 218968 347286 218980
rect 363598 218968 363604 218980
rect 363656 218968 363662 219020
rect 368658 218968 368664 219020
rect 368716 219008 368722 219020
rect 377398 219008 377404 219020
rect 368716 218980 377404 219008
rect 368716 218968 368722 218980
rect 377398 218968 377404 218980
rect 377456 218968 377462 219020
rect 377600 218980 383654 219008
rect 63126 218832 63132 218884
rect 63184 218872 63190 218884
rect 75178 218872 75184 218884
rect 63184 218844 75184 218872
rect 63184 218832 63190 218844
rect 75178 218832 75184 218844
rect 75236 218832 75242 218884
rect 77202 218832 77208 218884
rect 77260 218872 77266 218884
rect 150434 218872 150440 218884
rect 77260 218844 150440 218872
rect 77260 218832 77266 218844
rect 150434 218832 150440 218844
rect 150492 218832 150498 218884
rect 152366 218832 152372 218884
rect 152424 218872 152430 218884
rect 153838 218872 153844 218884
rect 152424 218844 153844 218872
rect 152424 218832 152430 218844
rect 153838 218832 153844 218844
rect 153896 218832 153902 218884
rect 154666 218832 154672 218884
rect 154724 218872 154730 218884
rect 159358 218872 159364 218884
rect 154724 218844 159364 218872
rect 154724 218832 154730 218844
rect 159358 218832 159364 218844
rect 159416 218832 159422 218884
rect 159818 218832 159824 218884
rect 159876 218872 159882 218884
rect 203518 218872 203524 218884
rect 159876 218844 203524 218872
rect 159876 218832 159882 218844
rect 203518 218832 203524 218844
rect 203576 218832 203582 218884
rect 206462 218832 206468 218884
rect 206520 218872 206526 218884
rect 253842 218872 253848 218884
rect 206520 218844 253848 218872
rect 206520 218832 206526 218844
rect 253842 218832 253848 218844
rect 253900 218832 253906 218884
rect 259086 218832 259092 218884
rect 259144 218872 259150 218884
rect 259144 218844 287054 218872
rect 259144 218832 259150 218844
rect 59814 218696 59820 218748
rect 59872 218736 59878 218748
rect 140038 218736 140044 218748
rect 59872 218708 140044 218736
rect 59872 218696 59878 218708
rect 140038 218696 140044 218708
rect 140096 218696 140102 218748
rect 140958 218696 140964 218748
rect 141016 218736 141022 218748
rect 142062 218736 142068 218748
rect 141016 218708 142068 218736
rect 141016 218696 141022 218708
rect 142062 218696 142068 218708
rect 142120 218696 142126 218748
rect 142614 218696 142620 218748
rect 142672 218736 142678 218748
rect 143258 218736 143264 218748
rect 142672 218708 143264 218736
rect 142672 218696 142678 218708
rect 143258 218696 143264 218708
rect 143316 218696 143322 218748
rect 146754 218696 146760 218748
rect 146812 218736 146818 218748
rect 184198 218736 184204 218748
rect 146812 218708 184204 218736
rect 146812 218696 146818 218708
rect 184198 218696 184204 218708
rect 184256 218696 184262 218748
rect 186498 218696 186504 218748
rect 186556 218736 186562 218748
rect 192294 218736 192300 218748
rect 186556 218708 192300 218736
rect 186556 218696 186562 218708
rect 192294 218696 192300 218708
rect 192352 218696 192358 218748
rect 192846 218696 192852 218748
rect 192904 218736 192910 218748
rect 243446 218736 243452 218748
rect 192904 218708 243452 218736
rect 192904 218696 192910 218708
rect 243446 218696 243452 218708
rect 243504 218696 243510 218748
rect 253198 218696 253204 218748
rect 253256 218736 253262 218748
rect 286318 218736 286324 218748
rect 253256 218708 286324 218736
rect 253256 218696 253262 218708
rect 286318 218696 286324 218708
rect 286376 218696 286382 218748
rect 287026 218736 287054 218844
rect 291654 218832 291660 218884
rect 291712 218872 291718 218884
rect 291712 218844 296714 218872
rect 291712 218832 291718 218844
rect 291838 218736 291844 218748
rect 287026 218708 291844 218736
rect 291838 218696 291844 218708
rect 291896 218696 291902 218748
rect 296686 218736 296714 218844
rect 300486 218832 300492 218884
rect 300544 218872 300550 218884
rect 327718 218872 327724 218884
rect 300544 218844 327724 218872
rect 300544 218832 300550 218844
rect 327718 218832 327724 218844
rect 327776 218832 327782 218884
rect 340506 218832 340512 218884
rect 340564 218872 340570 218884
rect 358078 218872 358084 218884
rect 340564 218844 358084 218872
rect 340564 218832 340570 218844
rect 358078 218832 358084 218844
rect 358136 218832 358142 218884
rect 363690 218832 363696 218884
rect 363748 218872 363754 218884
rect 370498 218872 370504 218884
rect 363748 218844 370504 218872
rect 363748 218832 363754 218844
rect 370498 218832 370504 218844
rect 370556 218832 370562 218884
rect 376938 218832 376944 218884
rect 376996 218872 377002 218884
rect 377600 218872 377628 218980
rect 376996 218844 377628 218872
rect 376996 218832 377002 218844
rect 382734 218832 382740 218884
rect 382792 218872 382798 218884
rect 383470 218872 383476 218884
rect 382792 218844 383476 218872
rect 382792 218832 382798 218844
rect 383470 218832 383476 218844
rect 383528 218832 383534 218884
rect 383626 218872 383654 218980
rect 386874 218968 386880 219020
rect 386932 219008 386938 219020
rect 398098 219008 398104 219020
rect 386932 218980 398104 219008
rect 386932 218968 386938 218980
rect 398098 218968 398104 218980
rect 398156 218968 398162 219020
rect 547414 218968 547420 219020
rect 547472 219008 547478 219020
rect 548536 219008 548564 219116
rect 553366 219116 562876 219144
rect 553366 219008 553394 219116
rect 562870 219104 562876 219116
rect 562928 219104 562934 219156
rect 563514 219104 563520 219156
rect 563572 219144 563578 219156
rect 572070 219144 572076 219156
rect 563572 219116 572076 219144
rect 563572 219104 563578 219116
rect 572070 219104 572076 219116
rect 572128 219104 572134 219156
rect 547472 218980 548472 219008
rect 548536 218980 553394 219008
rect 547472 218968 547478 218980
rect 388530 218872 388536 218884
rect 383626 218844 388536 218872
rect 388530 218832 388536 218844
rect 388588 218832 388594 218884
rect 402606 218832 402612 218884
rect 402664 218872 402670 218884
rect 409046 218872 409052 218884
rect 402664 218844 409052 218872
rect 402664 218832 402670 218844
rect 409046 218832 409052 218844
rect 409104 218832 409110 218884
rect 411714 218832 411720 218884
rect 411772 218872 411778 218884
rect 412542 218872 412548 218884
rect 411772 218844 412548 218872
rect 411772 218832 411778 218844
rect 412542 218832 412548 218844
rect 412600 218832 412606 218884
rect 512730 218832 512736 218884
rect 512788 218872 512794 218884
rect 548150 218872 548156 218884
rect 512788 218844 528554 218872
rect 512788 218832 512794 218844
rect 321554 218736 321560 218748
rect 296686 218708 321560 218736
rect 321554 218696 321560 218708
rect 321612 218696 321618 218748
rect 327258 218696 327264 218748
rect 327316 218736 327322 218748
rect 351086 218736 351092 218748
rect 327316 218708 351092 218736
rect 327316 218696 327322 218708
rect 351086 218696 351092 218708
rect 351144 218696 351150 218748
rect 353754 218696 353760 218748
rect 353812 218736 353818 218748
rect 369118 218736 369124 218748
rect 353812 218708 369124 218736
rect 353812 218696 353818 218708
rect 369118 218696 369124 218708
rect 369176 218696 369182 218748
rect 370314 218696 370320 218748
rect 370372 218736 370378 218748
rect 380066 218736 380072 218748
rect 370372 218708 380072 218736
rect 370372 218696 370378 218708
rect 380066 218696 380072 218708
rect 380124 218696 380130 218748
rect 383562 218696 383568 218748
rect 383620 218736 383626 218748
rect 396258 218736 396264 218748
rect 383620 218708 396264 218736
rect 383620 218696 383626 218708
rect 396258 218696 396264 218708
rect 396316 218696 396322 218748
rect 412542 218696 412548 218748
rect 412600 218736 412606 218748
rect 417142 218736 417148 218748
rect 412600 218708 417148 218736
rect 412600 218696 412606 218708
rect 417142 218696 417148 218708
rect 417200 218696 417206 218748
rect 429930 218696 429936 218748
rect 429988 218736 429994 218748
rect 432690 218736 432696 218748
rect 429988 218708 432696 218736
rect 429988 218696 429994 218708
rect 432690 218696 432696 218708
rect 432748 218696 432754 218748
rect 482738 218696 482744 218748
rect 482796 218736 482802 218748
rect 485314 218736 485320 218748
rect 482796 218708 485320 218736
rect 482796 218696 482802 218708
rect 485314 218696 485320 218708
rect 485372 218696 485378 218748
rect 500402 218696 500408 218748
rect 500460 218736 500466 218748
rect 508038 218736 508044 218748
rect 500460 218708 508044 218736
rect 500460 218696 500466 218708
rect 508038 218696 508044 218708
rect 508096 218696 508102 218748
rect 517698 218696 517704 218748
rect 517756 218736 517762 218748
rect 518158 218736 518164 218748
rect 517756 218708 518164 218736
rect 517756 218696 517762 218708
rect 518158 218696 518164 218708
rect 518216 218736 518222 218748
rect 519998 218736 520004 218748
rect 518216 218708 520004 218736
rect 518216 218696 518222 218708
rect 519998 218696 520004 218708
rect 520056 218696 520062 218748
rect 528526 218736 528554 218844
rect 534046 218844 548156 218872
rect 534046 218736 534074 218844
rect 548150 218832 548156 218844
rect 548208 218832 548214 218884
rect 548444 218872 548472 218980
rect 557350 218968 557356 219020
rect 557408 219008 557414 219020
rect 614114 219008 614120 219020
rect 557408 218980 614120 219008
rect 557408 218968 557414 218980
rect 614114 218968 614120 218980
rect 614172 218968 614178 219020
rect 562686 218872 562692 218884
rect 548444 218844 562692 218872
rect 562686 218832 562692 218844
rect 562744 218832 562750 218884
rect 563606 218832 563612 218884
rect 563664 218872 563670 218884
rect 572070 218872 572076 218884
rect 563664 218844 572076 218872
rect 563664 218832 563670 218844
rect 572070 218832 572076 218844
rect 572128 218832 572134 218884
rect 574738 218832 574744 218884
rect 574796 218872 574802 218884
rect 603074 218872 603080 218884
rect 574796 218844 603080 218872
rect 574796 218832 574802 218844
rect 603074 218832 603080 218844
rect 603132 218832 603138 218884
rect 572456 218776 572852 218804
rect 528526 218708 534074 218736
rect 537478 218696 537484 218748
rect 537536 218736 537542 218748
rect 563330 218736 563336 218748
rect 537536 218708 563336 218736
rect 537536 218696 537542 218708
rect 563330 218696 563336 218708
rect 563388 218696 563394 218748
rect 564158 218696 564164 218748
rect 564216 218736 564222 218748
rect 572456 218736 572484 218776
rect 564216 218708 572484 218736
rect 572824 218736 572852 218776
rect 598842 218736 598848 218748
rect 572824 218708 598848 218736
rect 564216 218696 564222 218708
rect 598842 218696 598848 218708
rect 598900 218696 598906 218748
rect 100386 218560 100392 218612
rect 100444 218600 100450 218612
rect 146570 218600 146576 218612
rect 100444 218572 146576 218600
rect 100444 218560 100450 218572
rect 146570 218560 146576 218572
rect 146628 218560 146634 218612
rect 148410 218560 148416 218612
rect 148468 218600 148474 218612
rect 148870 218600 148876 218612
rect 148468 218572 148876 218600
rect 148468 218560 148474 218572
rect 148870 218560 148876 218572
rect 148928 218560 148934 218612
rect 149238 218560 149244 218612
rect 149296 218600 149302 218612
rect 150066 218600 150072 218612
rect 149296 218572 150072 218600
rect 149296 218560 149302 218572
rect 150066 218560 150072 218572
rect 150124 218560 150130 218612
rect 150434 218560 150440 218612
rect 150492 218600 150498 218612
rect 152366 218600 152372 218612
rect 150492 218572 152372 218600
rect 150492 218560 150498 218572
rect 152366 218560 152372 218572
rect 152424 218560 152430 218612
rect 152550 218560 152556 218612
rect 152608 218600 152614 218612
rect 153102 218600 153108 218612
rect 152608 218572 153108 218600
rect 152608 218560 152614 218572
rect 153102 218560 153108 218572
rect 153160 218560 153166 218612
rect 153378 218560 153384 218612
rect 153436 218600 153442 218612
rect 154482 218600 154488 218612
rect 153436 218572 154488 218600
rect 153436 218560 153442 218572
rect 154482 218560 154488 218572
rect 154540 218560 154546 218612
rect 155034 218560 155040 218612
rect 155092 218600 155098 218612
rect 155678 218600 155684 218612
rect 155092 218572 155684 218600
rect 155092 218560 155098 218572
rect 155678 218560 155684 218572
rect 155736 218560 155742 218612
rect 156690 218560 156696 218612
rect 156748 218600 156754 218612
rect 157242 218600 157248 218612
rect 156748 218572 157248 218600
rect 156748 218560 156754 218572
rect 157242 218560 157248 218572
rect 157300 218560 157306 218612
rect 159174 218560 159180 218612
rect 159232 218600 159238 218612
rect 160002 218600 160008 218612
rect 159232 218572 160008 218600
rect 159232 218560 159238 218572
rect 160002 218560 160008 218572
rect 160060 218560 160066 218612
rect 160186 218560 160192 218612
rect 160244 218600 160250 218612
rect 186958 218600 186964 218612
rect 160244 218572 186964 218600
rect 160244 218560 160250 218572
rect 186958 218560 186964 218572
rect 187016 218560 187022 218612
rect 188706 218560 188712 218612
rect 188764 218600 188770 218612
rect 193582 218600 193588 218612
rect 188764 218572 193588 218600
rect 188764 218560 188770 218572
rect 193582 218560 193588 218572
rect 193640 218560 193646 218612
rect 195606 218560 195612 218612
rect 195664 218600 195670 218612
rect 197998 218600 198004 218612
rect 195664 218572 198004 218600
rect 195664 218560 195670 218572
rect 197998 218560 198004 218572
rect 198056 218560 198062 218612
rect 198918 218560 198924 218612
rect 198976 218600 198982 218612
rect 200022 218600 200028 218612
rect 198976 218572 200028 218600
rect 198976 218560 198982 218572
rect 200022 218560 200028 218572
rect 200080 218560 200086 218612
rect 204714 218560 204720 218612
rect 204772 218600 204778 218612
rect 207658 218600 207664 218612
rect 204772 218572 207664 218600
rect 204772 218560 204778 218572
rect 207658 218560 207664 218572
rect 207716 218560 207722 218612
rect 214282 218600 214288 218612
rect 207860 218572 214288 218600
rect 107010 218424 107016 218476
rect 107068 218464 107074 218476
rect 117958 218464 117964 218476
rect 107068 218436 117964 218464
rect 107068 218424 107074 218436
rect 117958 218424 117964 218436
rect 118016 218424 118022 218476
rect 120258 218424 120264 218476
rect 120316 218464 120322 218476
rect 166258 218464 166264 218476
rect 120316 218436 166264 218464
rect 120316 218424 120322 218436
rect 166258 218424 166264 218436
rect 166316 218424 166322 218476
rect 170950 218424 170956 218476
rect 171008 218464 171014 218476
rect 176286 218464 176292 218476
rect 171008 218436 176292 218464
rect 171008 218424 171014 218436
rect 176286 218424 176292 218436
rect 176344 218424 176350 218476
rect 179874 218424 179880 218476
rect 179932 218464 179938 218476
rect 204898 218464 204904 218476
rect 179932 218436 204904 218464
rect 179932 218424 179938 218436
rect 204898 218424 204904 218436
rect 204956 218424 204962 218476
rect 117774 218288 117780 218340
rect 117832 218328 117838 218340
rect 123478 218328 123484 218340
rect 117832 218300 123484 218328
rect 117832 218288 117838 218300
rect 123478 218288 123484 218300
rect 123536 218288 123542 218340
rect 130194 218288 130200 218340
rect 130252 218328 130258 218340
rect 136358 218328 136364 218340
rect 130252 218300 136364 218328
rect 130252 218288 130258 218300
rect 136358 218288 136364 218300
rect 136416 218288 136422 218340
rect 136818 218288 136824 218340
rect 136876 218328 136882 218340
rect 174722 218328 174728 218340
rect 136876 218300 174728 218328
rect 136876 218288 136882 218300
rect 174722 218288 174728 218300
rect 174780 218288 174786 218340
rect 175734 218288 175740 218340
rect 175792 218328 175798 218340
rect 179506 218328 179512 218340
rect 175792 218300 179512 218328
rect 175792 218288 175798 218300
rect 179506 218288 179512 218300
rect 179564 218288 179570 218340
rect 180702 218288 180708 218340
rect 180760 218328 180766 218340
rect 185946 218328 185952 218340
rect 180760 218300 185952 218328
rect 180760 218288 180766 218300
rect 185946 218288 185952 218300
rect 186004 218288 186010 218340
rect 189810 218288 189816 218340
rect 189868 218328 189874 218340
rect 195238 218328 195244 218340
rect 189868 218300 195244 218328
rect 189868 218288 189874 218300
rect 195238 218288 195244 218300
rect 195296 218288 195302 218340
rect 198090 218288 198096 218340
rect 198148 218328 198154 218340
rect 198148 218300 200436 218328
rect 198148 218288 198154 218300
rect 123662 218220 123668 218272
rect 123720 218260 123726 218272
rect 123720 218232 129596 218260
rect 123720 218220 123726 218232
rect 55674 218152 55680 218204
rect 55732 218192 55738 218204
rect 56502 218192 56508 218204
rect 55732 218164 56508 218192
rect 55732 218152 55738 218164
rect 56502 218152 56508 218164
rect 56560 218152 56566 218204
rect 57422 218152 57428 218204
rect 57480 218192 57486 218204
rect 61378 218192 61384 218204
rect 57480 218164 61384 218192
rect 57480 218152 57486 218164
rect 61378 218152 61384 218164
rect 61436 218152 61442 218204
rect 66438 218152 66444 218204
rect 66496 218192 66502 218204
rect 67542 218192 67548 218204
rect 66496 218164 67548 218192
rect 66496 218152 66502 218164
rect 67542 218152 67548 218164
rect 67600 218152 67606 218204
rect 68094 218152 68100 218204
rect 68152 218192 68158 218204
rect 69566 218192 69572 218204
rect 68152 218164 69572 218192
rect 68152 218152 68158 218164
rect 69566 218152 69572 218164
rect 69624 218152 69630 218204
rect 75546 218152 75552 218204
rect 75604 218192 75610 218204
rect 76558 218192 76564 218204
rect 75604 218164 76564 218192
rect 75604 218152 75610 218164
rect 76558 218152 76564 218164
rect 76616 218152 76622 218204
rect 97074 218152 97080 218204
rect 97132 218192 97138 218204
rect 97132 218164 100892 218192
rect 97132 218152 97138 218164
rect 56502 218016 56508 218068
rect 56560 218056 56566 218068
rect 57238 218056 57244 218068
rect 56560 218028 57244 218056
rect 56560 218016 56566 218028
rect 57238 218016 57244 218028
rect 57296 218016 57302 218068
rect 58158 218016 58164 218068
rect 58216 218056 58222 218068
rect 59354 218056 59360 218068
rect 58216 218028 59360 218056
rect 58216 218016 58222 218028
rect 59354 218016 59360 218028
rect 59412 218016 59418 218068
rect 61470 218016 61476 218068
rect 61528 218056 61534 218068
rect 62758 218056 62764 218068
rect 61528 218028 62764 218056
rect 61528 218016 61534 218028
rect 62758 218016 62764 218028
rect 62816 218016 62822 218068
rect 63954 218016 63960 218068
rect 64012 218056 64018 218068
rect 64782 218056 64788 218068
rect 64012 218028 64788 218056
rect 64012 218016 64018 218028
rect 64782 218016 64788 218028
rect 64840 218016 64846 218068
rect 65610 218016 65616 218068
rect 65668 218056 65674 218068
rect 66162 218056 66168 218068
rect 65668 218028 66168 218056
rect 65668 218016 65674 218028
rect 66162 218016 66168 218028
rect 66220 218016 66226 218068
rect 67266 218016 67272 218068
rect 67324 218056 67330 218068
rect 68278 218056 68284 218068
rect 67324 218028 68284 218056
rect 67324 218016 67330 218028
rect 68278 218016 68284 218028
rect 68336 218016 68342 218068
rect 72234 218016 72240 218068
rect 72292 218056 72298 218068
rect 73706 218056 73712 218068
rect 72292 218028 73712 218056
rect 72292 218016 72298 218028
rect 73706 218016 73712 218028
rect 73764 218016 73770 218068
rect 74718 218016 74724 218068
rect 74776 218056 74782 218068
rect 75822 218056 75828 218068
rect 74776 218028 75828 218056
rect 74776 218016 74782 218028
rect 75822 218016 75828 218028
rect 75880 218016 75886 218068
rect 78030 218016 78036 218068
rect 78088 218056 78094 218068
rect 78582 218056 78588 218068
rect 78088 218028 78588 218056
rect 78088 218016 78094 218028
rect 78582 218016 78588 218028
rect 78640 218016 78646 218068
rect 78858 218016 78864 218068
rect 78916 218056 78922 218068
rect 79962 218056 79968 218068
rect 78916 218028 79968 218056
rect 78916 218016 78922 218028
rect 79962 218016 79968 218028
rect 80020 218016 80026 218068
rect 82170 218016 82176 218068
rect 82228 218056 82234 218068
rect 83458 218056 83464 218068
rect 82228 218028 83464 218056
rect 82228 218016 82234 218028
rect 83458 218016 83464 218028
rect 83516 218016 83522 218068
rect 84654 218016 84660 218068
rect 84712 218056 84718 218068
rect 85298 218056 85304 218068
rect 84712 218028 85304 218056
rect 84712 218016 84718 218028
rect 85298 218016 85304 218028
rect 85356 218016 85362 218068
rect 87138 218016 87144 218068
rect 87196 218056 87202 218068
rect 88242 218056 88248 218068
rect 87196 218028 88248 218056
rect 87196 218016 87202 218028
rect 88242 218016 88248 218028
rect 88300 218016 88306 218068
rect 88794 218016 88800 218068
rect 88852 218056 88858 218068
rect 89438 218056 89444 218068
rect 88852 218028 89444 218056
rect 88852 218016 88858 218028
rect 89438 218016 89444 218028
rect 89496 218016 89502 218068
rect 92934 218016 92940 218068
rect 92992 218056 92998 218068
rect 93762 218056 93768 218068
rect 92992 218028 93768 218056
rect 92992 218016 92998 218028
rect 93762 218016 93768 218028
rect 93820 218016 93826 218068
rect 95418 218016 95424 218068
rect 95476 218056 95482 218068
rect 96246 218056 96252 218068
rect 95476 218028 96252 218056
rect 95476 218016 95482 218028
rect 96246 218016 96252 218028
rect 96304 218016 96310 218068
rect 98730 218016 98736 218068
rect 98788 218056 98794 218068
rect 99282 218056 99288 218068
rect 98788 218028 99288 218056
rect 98788 218016 98794 218028
rect 99282 218016 99288 218028
rect 99340 218016 99346 218068
rect 99558 218016 99564 218068
rect 99616 218056 99622 218068
rect 100662 218056 100668 218068
rect 99616 218028 100668 218056
rect 99616 218016 99622 218028
rect 100662 218016 100668 218028
rect 100720 218016 100726 218068
rect 100864 217988 100892 218164
rect 117774 218152 117780 218204
rect 117832 218192 117838 218204
rect 118694 218192 118700 218204
rect 117832 218164 118700 218192
rect 117832 218152 117838 218164
rect 118694 218152 118700 218164
rect 118752 218152 118758 218204
rect 129568 218192 129596 218232
rect 132494 218192 132500 218204
rect 129568 218164 132500 218192
rect 132494 218152 132500 218164
rect 132552 218152 132558 218204
rect 140130 218152 140136 218204
rect 140188 218192 140194 218204
rect 175918 218192 175924 218204
rect 140188 218164 175924 218192
rect 140188 218152 140194 218164
rect 175918 218152 175924 218164
rect 175976 218152 175982 218204
rect 178678 218192 178684 218204
rect 176120 218164 178684 218192
rect 102870 218084 102876 218136
rect 102928 218124 102934 218136
rect 103422 218124 103428 218136
rect 102928 218096 103428 218124
rect 102928 218084 102934 218096
rect 103422 218084 103428 218096
rect 103480 218084 103486 218136
rect 103698 218084 103704 218136
rect 103756 218124 103762 218136
rect 104802 218124 104808 218136
rect 103756 218096 104808 218124
rect 103756 218084 103762 218096
rect 104802 218084 104808 218096
rect 104860 218084 104866 218136
rect 105354 218084 105360 218136
rect 105412 218124 105418 218136
rect 105998 218124 106004 218136
rect 105412 218096 106004 218124
rect 105412 218084 105418 218096
rect 105998 218084 106004 218096
rect 106056 218084 106062 218136
rect 111978 218084 111984 218136
rect 112036 218124 112042 218136
rect 112806 218124 112812 218136
rect 112036 218096 112812 218124
rect 112036 218084 112042 218096
rect 112806 218084 112812 218096
rect 112864 218084 112870 218136
rect 116118 218084 116124 218136
rect 116176 218124 116182 218136
rect 117222 218124 117228 218136
rect 116176 218096 117228 218124
rect 116176 218084 116182 218096
rect 117222 218084 117228 218096
rect 117280 218084 117286 218136
rect 119430 218084 119436 218136
rect 119488 218124 119494 218136
rect 119982 218124 119988 218136
rect 119488 218096 119988 218124
rect 119488 218084 119494 218096
rect 119982 218084 119988 218096
rect 120040 218084 120046 218136
rect 121914 218084 121920 218136
rect 121972 218124 121978 218136
rect 122558 218124 122564 218136
rect 121972 218096 122564 218124
rect 121972 218084 121978 218096
rect 122558 218084 122564 218096
rect 122616 218084 122622 218136
rect 126054 218084 126060 218136
rect 126112 218124 126118 218136
rect 126698 218124 126704 218136
rect 126112 218096 126704 218124
rect 126112 218084 126118 218096
rect 126698 218084 126704 218096
rect 126756 218084 126762 218136
rect 127710 218084 127716 218136
rect 127768 218124 127774 218136
rect 128262 218124 128268 218136
rect 127768 218096 128268 218124
rect 127768 218084 127774 218096
rect 128262 218084 128268 218096
rect 128320 218084 128326 218136
rect 128538 218084 128544 218136
rect 128596 218124 128602 218136
rect 129366 218124 129372 218136
rect 128596 218096 129372 218124
rect 128596 218084 128602 218096
rect 129366 218084 129372 218096
rect 129424 218084 129430 218136
rect 132678 218084 132684 218136
rect 132736 218124 132742 218136
rect 133506 218124 133512 218136
rect 132736 218096 133512 218124
rect 132736 218084 132742 218096
rect 133506 218084 133512 218096
rect 133564 218084 133570 218136
rect 135990 218084 135996 218136
rect 136048 218124 136054 218136
rect 136542 218124 136548 218136
rect 136048 218096 136548 218124
rect 136048 218084 136054 218096
rect 136542 218084 136548 218096
rect 136600 218084 136606 218136
rect 161658 218016 161664 218068
rect 161716 218056 161722 218068
rect 162762 218056 162768 218068
rect 161716 218028 162768 218056
rect 161716 218016 161722 218028
rect 162762 218016 162768 218028
rect 162820 218016 162826 218068
rect 163314 218016 163320 218068
rect 163372 218056 163378 218068
rect 163958 218056 163964 218068
rect 163372 218028 163964 218056
rect 163372 218016 163378 218028
rect 163958 218016 163964 218028
rect 164016 218016 164022 218068
rect 164970 218016 164976 218068
rect 165028 218056 165034 218068
rect 165522 218056 165528 218068
rect 165028 218028 165528 218056
rect 165028 218016 165034 218028
rect 165522 218016 165528 218028
rect 165580 218016 165586 218068
rect 169110 218016 169116 218068
rect 169168 218056 169174 218068
rect 169570 218056 169576 218068
rect 169168 218028 169576 218056
rect 169168 218016 169174 218028
rect 169570 218016 169576 218028
rect 169628 218016 169634 218068
rect 169938 218016 169944 218068
rect 169996 218056 170002 218068
rect 170766 218056 170772 218068
rect 169996 218028 170772 218056
rect 169996 218016 170002 218028
rect 170766 218016 170772 218028
rect 170824 218016 170830 218068
rect 172422 218016 172428 218068
rect 172480 218056 172486 218068
rect 173158 218056 173164 218068
rect 172480 218028 173164 218056
rect 172480 218016 172486 218028
rect 173158 218016 173164 218028
rect 173216 218016 173222 218068
rect 173342 218016 173348 218068
rect 173400 218056 173406 218068
rect 173400 218028 174584 218056
rect 173400 218016 173406 218028
rect 100864 217960 161474 217988
rect 161446 217920 161474 217960
rect 174078 217920 174084 217932
rect 161446 217892 174084 217920
rect 174078 217880 174084 217892
rect 174136 217880 174142 217932
rect 174556 217920 174584 218028
rect 174722 218016 174728 218068
rect 174780 218056 174786 218068
rect 176120 218056 176148 218164
rect 178678 218152 178684 218164
rect 178736 218152 178742 218204
rect 179046 218152 179052 218204
rect 179104 218192 179110 218204
rect 196618 218192 196624 218204
rect 179104 218164 196624 218192
rect 179104 218152 179110 218164
rect 196618 218152 196624 218164
rect 196676 218152 196682 218204
rect 199746 218152 199752 218204
rect 199804 218192 199810 218204
rect 200206 218192 200212 218204
rect 199804 218164 200212 218192
rect 199804 218152 199810 218164
rect 200206 218152 200212 218164
rect 200264 218152 200270 218204
rect 200408 218192 200436 218300
rect 200666 218288 200672 218340
rect 200724 218328 200730 218340
rect 207860 218328 207888 218572
rect 214282 218560 214288 218572
rect 214340 218560 214346 218612
rect 214742 218560 214748 218612
rect 214800 218600 214806 218612
rect 219802 218600 219808 218612
rect 214800 218572 219808 218600
rect 214800 218560 214806 218572
rect 219802 218560 219808 218572
rect 219860 218560 219866 218612
rect 225966 218560 225972 218612
rect 226024 218600 226030 218612
rect 266998 218600 267004 218612
rect 226024 218572 267004 218600
rect 226024 218560 226030 218572
rect 266998 218560 267004 218572
rect 267056 218560 267062 218612
rect 272334 218560 272340 218612
rect 272392 218600 272398 218612
rect 279418 218600 279424 218612
rect 272392 218572 279424 218600
rect 272392 218560 272398 218572
rect 279418 218560 279424 218572
rect 279476 218560 279482 218612
rect 305546 218600 305552 218612
rect 287026 218572 305552 218600
rect 208486 218424 208492 218476
rect 208544 218464 208550 218476
rect 211798 218464 211804 218476
rect 208544 218436 211804 218464
rect 208544 218424 208550 218436
rect 211798 218424 211804 218436
rect 211856 218424 211862 218476
rect 212994 218424 213000 218476
rect 213052 218464 213058 218476
rect 224218 218464 224224 218476
rect 213052 218436 224224 218464
rect 213052 218424 213058 218436
rect 224218 218424 224224 218436
rect 224276 218424 224282 218476
rect 224402 218424 224408 218476
rect 224460 218464 224466 218476
rect 231026 218464 231032 218476
rect 224460 218436 231032 218464
rect 224460 218424 224466 218436
rect 231026 218424 231032 218436
rect 231084 218424 231090 218476
rect 238018 218464 238024 218476
rect 232700 218436 238024 218464
rect 200724 218300 207888 218328
rect 200724 218288 200730 218300
rect 209682 218288 209688 218340
rect 209740 218328 209746 218340
rect 213178 218328 213184 218340
rect 209740 218300 213184 218328
rect 209740 218288 209746 218300
rect 213178 218288 213184 218300
rect 213236 218288 213242 218340
rect 214282 218288 214288 218340
rect 214340 218328 214346 218340
rect 214340 218300 214650 218328
rect 214340 218288 214346 218300
rect 204162 218192 204168 218204
rect 200408 218164 204168 218192
rect 204162 218152 204168 218164
rect 204220 218152 204226 218204
rect 204898 218152 204904 218204
rect 204956 218192 204962 218204
rect 210326 218192 210332 218204
rect 204956 218164 210332 218192
rect 204956 218152 204962 218164
rect 210326 218152 210332 218164
rect 210384 218152 210390 218204
rect 211338 218152 211344 218204
rect 211396 218192 211402 218204
rect 214466 218192 214472 218204
rect 211396 218164 214472 218192
rect 211396 218152 211402 218164
rect 214466 218152 214472 218164
rect 214524 218152 214530 218204
rect 214622 218192 214650 218300
rect 216306 218288 216312 218340
rect 216364 218328 216370 218340
rect 232700 218328 232728 218436
rect 238018 218424 238024 218436
rect 238076 218424 238082 218476
rect 271138 218464 271144 218476
rect 238726 218436 271144 218464
rect 216364 218300 232728 218328
rect 216364 218288 216370 218300
rect 232866 218288 232872 218340
rect 232924 218328 232930 218340
rect 238726 218328 238754 218436
rect 271138 218424 271144 218436
rect 271196 218424 271202 218476
rect 279234 218424 279240 218476
rect 279292 218464 279298 218476
rect 287026 218464 287054 218572
rect 305546 218560 305552 218572
rect 305604 218560 305610 218612
rect 398466 218560 398472 218612
rect 398524 218600 398530 218612
rect 407758 218600 407764 218612
rect 398524 218572 407764 218600
rect 398524 218560 398530 218572
rect 407758 218560 407764 218572
rect 407816 218560 407822 218612
rect 469858 218560 469864 218612
rect 469916 218600 469922 218612
rect 471238 218600 471244 218612
rect 469916 218572 471244 218600
rect 469916 218560 469922 218572
rect 471238 218560 471244 218572
rect 471296 218560 471302 218612
rect 475562 218560 475568 218612
rect 475620 218600 475626 218612
rect 482830 218600 482836 218612
rect 475620 218572 482836 218600
rect 475620 218560 475626 218572
rect 482830 218560 482836 218572
rect 482888 218560 482894 218612
rect 507670 218560 507676 218612
rect 507728 218600 507734 218612
rect 563192 218600 563198 218612
rect 507728 218572 563198 218600
rect 507728 218560 507734 218572
rect 563192 218560 563198 218572
rect 563250 218560 563256 218612
rect 572806 218560 572812 218612
rect 572864 218600 572870 218612
rect 610710 218600 610716 218612
rect 572864 218572 610716 218600
rect 572864 218560 572870 218572
rect 610710 218560 610716 218572
rect 610768 218560 610774 218612
rect 568298 218492 568304 218544
rect 568356 218532 568362 218544
rect 572438 218532 572444 218544
rect 568356 218504 572444 218532
rect 568356 218492 568362 218504
rect 572438 218492 572444 218504
rect 572496 218492 572502 218544
rect 279292 218436 287054 218464
rect 279292 218424 279298 218436
rect 294138 218424 294144 218476
rect 294196 218464 294202 218476
rect 316678 218464 316684 218476
rect 294196 218436 316684 218464
rect 294196 218424 294202 218436
rect 316678 218424 316684 218436
rect 316736 218424 316742 218476
rect 502794 218424 502800 218476
rect 502852 218464 502858 218476
rect 503162 218464 503168 218476
rect 502852 218436 503168 218464
rect 502852 218424 502858 218436
rect 503162 218424 503168 218436
rect 503220 218464 503226 218476
rect 507854 218464 507860 218476
rect 503220 218436 507860 218464
rect 503220 218424 503226 218436
rect 507854 218424 507860 218436
rect 507912 218424 507918 218476
rect 508038 218424 508044 218476
rect 508096 218464 508102 218476
rect 508096 218436 567976 218464
rect 508096 218424 508102 218436
rect 458174 218356 458180 218408
rect 458232 218396 458238 218408
rect 567948 218396 567976 218436
rect 574922 218424 574928 218476
rect 574980 218464 574986 218476
rect 604454 218464 604460 218476
rect 574980 218436 604460 218464
rect 574980 218424 574986 218436
rect 604454 218424 604460 218436
rect 604512 218424 604518 218476
rect 572070 218396 572076 218408
rect 458232 218368 460934 218396
rect 567948 218368 572076 218396
rect 458232 218356 458238 218368
rect 232924 218300 238754 218328
rect 232924 218288 232930 218300
rect 241606 218288 241612 218340
rect 241664 218328 241670 218340
rect 246298 218328 246304 218340
rect 241664 218300 246304 218328
rect 241664 218288 241670 218300
rect 246298 218288 246304 218300
rect 246356 218288 246362 218340
rect 249426 218288 249432 218340
rect 249484 218328 249490 218340
rect 251726 218328 251732 218340
rect 249484 218300 251732 218328
rect 249484 218288 249490 218300
rect 251726 218288 251732 218300
rect 251784 218288 251790 218340
rect 253014 218288 253020 218340
rect 253072 218328 253078 218340
rect 258074 218328 258080 218340
rect 253072 218300 258080 218328
rect 253072 218288 253078 218300
rect 258074 218288 258080 218300
rect 258132 218288 258138 218340
rect 426618 218288 426624 218340
rect 426676 218328 426682 218340
rect 429378 218328 429384 218340
rect 426676 218300 429384 218328
rect 426676 218288 426682 218300
rect 429378 218288 429384 218300
rect 429436 218288 429442 218340
rect 450722 218288 450728 218340
rect 450780 218328 450786 218340
rect 453850 218328 453856 218340
rect 450780 218300 453856 218328
rect 450780 218288 450786 218300
rect 453850 218288 453856 218300
rect 453908 218288 453914 218340
rect 460906 218328 460934 218368
rect 572070 218356 572076 218368
rect 572128 218356 572134 218408
rect 461302 218328 461308 218340
rect 460906 218300 461308 218328
rect 461302 218288 461308 218300
rect 461360 218288 461366 218340
rect 497458 218288 497464 218340
rect 497516 218328 497522 218340
rect 497516 218300 567884 218328
rect 497516 218288 497522 218300
rect 567856 218260 567884 218300
rect 572806 218288 572812 218340
rect 572864 218328 572870 218340
rect 594794 218328 594800 218340
rect 572864 218300 594800 218328
rect 572864 218288 572870 218300
rect 594794 218288 594800 218300
rect 594852 218288 594858 218340
rect 668394 218288 668400 218340
rect 668452 218328 668458 218340
rect 669498 218328 669504 218340
rect 668452 218300 669504 218328
rect 668452 218288 668458 218300
rect 669498 218288 669504 218300
rect 669556 218288 669562 218340
rect 572530 218260 572536 218272
rect 567856 218232 572536 218260
rect 572530 218220 572536 218232
rect 572588 218220 572594 218272
rect 214622 218164 216720 218192
rect 176654 218056 176660 218068
rect 174780 218028 176148 218056
rect 176212 218028 176660 218056
rect 174780 218016 174786 218028
rect 176212 217920 176240 218028
rect 176654 218016 176660 218028
rect 176712 218016 176718 218068
rect 178218 218016 178224 218068
rect 178276 218056 178282 218068
rect 179322 218056 179328 218068
rect 178276 218028 179328 218056
rect 178276 218016 178282 218028
rect 179322 218016 179328 218028
rect 179380 218016 179386 218068
rect 179506 218016 179512 218068
rect 179564 218056 179570 218068
rect 183830 218056 183836 218068
rect 179564 218028 183836 218056
rect 179564 218016 179570 218028
rect 183830 218016 183836 218028
rect 183888 218016 183894 218068
rect 184014 218016 184020 218068
rect 184072 218056 184078 218068
rect 184658 218056 184664 218068
rect 184072 218028 184664 218056
rect 184072 218016 184078 218028
rect 184658 218016 184664 218028
rect 184716 218016 184722 218068
rect 185670 218016 185676 218068
rect 185728 218056 185734 218068
rect 186130 218056 186136 218068
rect 185728 218028 186136 218056
rect 185728 218016 185734 218028
rect 186130 218016 186136 218028
rect 186188 218016 186194 218068
rect 188154 218016 188160 218068
rect 188212 218056 188218 218068
rect 188890 218056 188896 218068
rect 188212 218028 188896 218056
rect 188212 218016 188218 218028
rect 188890 218016 188896 218028
rect 188948 218016 188954 218068
rect 192294 218016 192300 218068
rect 192352 218056 192358 218068
rect 193030 218056 193036 218068
rect 192352 218028 193036 218056
rect 192352 218016 192358 218028
rect 193030 218016 193036 218028
rect 193088 218016 193094 218068
rect 193950 218016 193956 218068
rect 194008 218056 194014 218068
rect 194502 218056 194508 218068
rect 194008 218028 194508 218056
rect 194008 218016 194014 218028
rect 194502 218016 194508 218028
rect 194560 218016 194566 218068
rect 194778 218016 194784 218068
rect 194836 218056 194842 218068
rect 195882 218056 195888 218068
rect 194836 218028 195888 218056
rect 194836 218016 194842 218028
rect 195882 218016 195888 218028
rect 195940 218016 195946 218068
rect 196434 218016 196440 218068
rect 196492 218056 196498 218068
rect 200390 218056 200396 218068
rect 196492 218028 200396 218056
rect 196492 218016 196498 218028
rect 200390 218016 200396 218028
rect 200448 218016 200454 218068
rect 200574 218016 200580 218068
rect 200632 218056 200638 218068
rect 201494 218056 201500 218068
rect 200632 218028 201500 218056
rect 200632 218016 200638 218028
rect 201494 218016 201500 218028
rect 201552 218016 201558 218068
rect 203058 218016 203064 218068
rect 203116 218056 203122 218068
rect 206278 218056 206284 218068
rect 203116 218028 206284 218056
rect 203116 218016 203122 218028
rect 206278 218016 206284 218028
rect 206336 218016 206342 218068
rect 207198 218016 207204 218068
rect 207256 218056 207262 218068
rect 208118 218056 208124 218068
rect 207256 218028 208124 218056
rect 207256 218016 207262 218028
rect 208118 218016 208124 218028
rect 208176 218016 208182 218068
rect 214650 218016 214656 218068
rect 214708 218056 214714 218068
rect 215202 218056 215208 218068
rect 214708 218028 215208 218056
rect 214708 218016 214714 218028
rect 215202 218016 215208 218028
rect 215260 218016 215266 218068
rect 215478 218016 215484 218068
rect 215536 218056 215542 218068
rect 216490 218056 216496 218068
rect 215536 218028 216496 218056
rect 215536 218016 215542 218028
rect 216490 218016 216496 218028
rect 216548 218016 216554 218068
rect 216692 218056 216720 218164
rect 217962 218152 217968 218204
rect 218020 218192 218026 218204
rect 222746 218192 222752 218204
rect 218020 218164 222752 218192
rect 218020 218152 218026 218164
rect 222746 218152 222752 218164
rect 222804 218152 222810 218204
rect 222930 218152 222936 218204
rect 222988 218192 222994 218204
rect 225598 218192 225604 218204
rect 222988 218164 225604 218192
rect 222988 218152 222994 218164
rect 225598 218152 225604 218164
rect 225656 218152 225662 218204
rect 246114 218152 246120 218204
rect 246172 218192 246178 218204
rect 253198 218192 253204 218204
rect 246172 218164 253204 218192
rect 246172 218152 246178 218164
rect 253198 218152 253204 218164
rect 253256 218152 253262 218204
rect 328914 218152 328920 218204
rect 328972 218192 328978 218204
rect 330478 218192 330484 218204
rect 328972 218164 330484 218192
rect 328972 218152 328978 218164
rect 330478 218152 330484 218164
rect 330536 218152 330542 218204
rect 365346 218152 365352 218204
rect 365404 218192 365410 218204
rect 371786 218192 371792 218204
rect 365404 218164 371792 218192
rect 365404 218152 365410 218164
rect 371786 218152 371792 218164
rect 371844 218152 371850 218204
rect 374454 218152 374460 218204
rect 374512 218192 374518 218204
rect 376018 218192 376024 218204
rect 374512 218164 376024 218192
rect 374512 218152 374518 218164
rect 376018 218152 376024 218164
rect 376076 218152 376082 218204
rect 381906 218152 381912 218204
rect 381964 218192 381970 218204
rect 382918 218192 382924 218204
rect 381964 218164 382924 218192
rect 381964 218152 381970 218164
rect 382918 218152 382924 218164
rect 382976 218152 382982 218204
rect 401778 218152 401784 218204
rect 401836 218192 401842 218204
rect 402790 218192 402796 218204
rect 401836 218164 402796 218192
rect 401836 218152 401842 218164
rect 402790 218152 402796 218164
rect 402848 218152 402854 218204
rect 407574 218152 407580 218204
rect 407632 218192 407638 218204
rect 411898 218192 411904 218204
rect 407632 218164 411904 218192
rect 407632 218152 407638 218164
rect 411898 218152 411904 218164
rect 411956 218152 411962 218204
rect 422478 218152 422484 218204
rect 422536 218192 422542 218204
rect 425422 218192 425428 218204
rect 422536 218164 425428 218192
rect 422536 218152 422542 218164
rect 425422 218152 425428 218164
rect 425480 218152 425486 218204
rect 425790 218152 425796 218204
rect 425848 218192 425854 218204
rect 427906 218192 427912 218204
rect 425848 218164 427912 218192
rect 425848 218152 425854 218164
rect 427906 218152 427912 218164
rect 427964 218152 427970 218204
rect 433242 218152 433248 218204
rect 433300 218192 433306 218204
rect 434714 218192 434720 218204
rect 433300 218164 434720 218192
rect 433300 218152 433306 218164
rect 434714 218152 434720 218164
rect 434772 218152 434778 218204
rect 434898 218152 434904 218204
rect 434956 218192 434962 218204
rect 436830 218192 436836 218204
rect 434956 218164 436836 218192
rect 434956 218152 434962 218164
rect 436830 218152 436836 218164
rect 436888 218152 436894 218204
rect 461946 218152 461952 218204
rect 462004 218192 462010 218204
rect 466270 218192 466276 218204
rect 462004 218164 466276 218192
rect 462004 218152 462010 218164
rect 466270 218152 466276 218164
rect 466328 218152 466334 218204
rect 491938 218152 491944 218204
rect 491996 218192 492002 218204
rect 502242 218192 502248 218204
rect 491996 218164 502248 218192
rect 491996 218152 492002 218164
rect 502242 218152 502248 218164
rect 502300 218152 502306 218204
rect 507118 218152 507124 218204
rect 507176 218192 507182 218204
rect 507670 218192 507676 218204
rect 507176 218164 507676 218192
rect 507176 218152 507182 218164
rect 507670 218152 507676 218164
rect 507728 218152 507734 218204
rect 507854 218152 507860 218204
rect 507912 218192 507918 218204
rect 562870 218192 562876 218204
rect 507912 218164 562876 218192
rect 507912 218152 507918 218164
rect 562870 218152 562876 218164
rect 562928 218152 562934 218204
rect 572990 218152 572996 218204
rect 573048 218192 573054 218204
rect 573048 218164 613884 218192
rect 573048 218152 573054 218164
rect 563210 218096 572852 218124
rect 220078 218056 220084 218068
rect 216692 218028 220084 218056
rect 220078 218016 220084 218028
rect 220136 218016 220142 218068
rect 221274 218016 221280 218068
rect 221332 218056 221338 218068
rect 221826 218056 221832 218068
rect 221332 218028 221832 218056
rect 221332 218016 221338 218028
rect 221826 218016 221832 218028
rect 221884 218016 221890 218068
rect 223758 218016 223764 218068
rect 223816 218056 223822 218068
rect 224586 218056 224592 218068
rect 223816 218028 224592 218056
rect 223816 218016 223822 218028
rect 224586 218016 224592 218028
rect 224644 218016 224650 218068
rect 225414 218016 225420 218068
rect 225472 218056 225478 218068
rect 226150 218056 226156 218068
rect 225472 218028 226156 218056
rect 225472 218016 225478 218028
rect 226150 218016 226156 218028
rect 226208 218016 226214 218068
rect 231210 218016 231216 218068
rect 231268 218056 231274 218068
rect 231670 218056 231676 218068
rect 231268 218028 231676 218056
rect 231268 218016 231274 218028
rect 231670 218016 231676 218028
rect 231728 218016 231734 218068
rect 232038 218016 232044 218068
rect 232096 218056 232102 218068
rect 233142 218056 233148 218068
rect 232096 218028 233148 218056
rect 232096 218016 232102 218028
rect 233142 218016 233148 218028
rect 233200 218016 233206 218068
rect 235350 218016 235356 218068
rect 235408 218056 235414 218068
rect 235810 218056 235816 218068
rect 235408 218028 235816 218056
rect 235408 218016 235414 218028
rect 235810 218016 235816 218028
rect 235868 218016 235874 218068
rect 236178 218016 236184 218068
rect 236236 218056 236242 218068
rect 237282 218056 237288 218068
rect 236236 218028 237288 218056
rect 236236 218016 236242 218028
rect 237282 218016 237288 218028
rect 237340 218016 237346 218068
rect 240318 218016 240324 218068
rect 240376 218056 240382 218068
rect 241330 218056 241336 218068
rect 240376 218028 241336 218056
rect 240376 218016 240382 218028
rect 241330 218016 241336 218028
rect 241388 218016 241394 218068
rect 243630 218016 243636 218068
rect 243688 218056 243694 218068
rect 244090 218056 244096 218068
rect 243688 218028 244096 218056
rect 243688 218016 243694 218028
rect 244090 218016 244096 218028
rect 244148 218016 244154 218068
rect 247770 218016 247776 218068
rect 247828 218056 247834 218068
rect 248230 218056 248236 218068
rect 247828 218028 248236 218056
rect 247828 218016 247834 218028
rect 248230 218016 248236 218028
rect 248288 218016 248294 218068
rect 248598 218016 248604 218068
rect 248656 218056 248662 218068
rect 249610 218056 249616 218068
rect 248656 218028 249616 218056
rect 248656 218016 248662 218028
rect 249610 218016 249616 218028
rect 249668 218016 249674 218068
rect 250254 218016 250260 218068
rect 250312 218056 250318 218068
rect 250898 218056 250904 218068
rect 250312 218028 250904 218056
rect 250312 218016 250318 218028
rect 250898 218016 250904 218028
rect 250956 218016 250962 218068
rect 251910 218016 251916 218068
rect 251968 218056 251974 218068
rect 252462 218056 252468 218068
rect 251968 218028 252468 218056
rect 251968 218016 251974 218028
rect 252462 218016 252468 218028
rect 252520 218016 252526 218068
rect 254394 218016 254400 218068
rect 254452 218056 254458 218068
rect 255038 218056 255044 218068
rect 254452 218028 255044 218056
rect 254452 218016 254458 218028
rect 255038 218016 255044 218028
rect 255096 218016 255102 218068
rect 256050 218016 256056 218068
rect 256108 218056 256114 218068
rect 256510 218056 256516 218068
rect 256108 218028 256516 218056
rect 256108 218016 256114 218028
rect 256510 218016 256516 218028
rect 256568 218016 256574 218068
rect 256878 218016 256884 218068
rect 256936 218056 256942 218068
rect 257522 218056 257528 218068
rect 256936 218028 257528 218056
rect 256936 218016 256942 218028
rect 257522 218016 257528 218028
rect 257580 218016 257586 218068
rect 258534 218016 258540 218068
rect 258592 218056 258598 218068
rect 259270 218056 259276 218068
rect 258592 218028 259276 218056
rect 258592 218016 258598 218028
rect 259270 218016 259276 218028
rect 259328 218016 259334 218068
rect 262674 218016 262680 218068
rect 262732 218056 262738 218068
rect 263594 218056 263600 218068
rect 262732 218028 263600 218056
rect 262732 218016 262738 218028
rect 263594 218016 263600 218028
rect 263652 218016 263658 218068
rect 264330 218016 264336 218068
rect 264388 218056 264394 218068
rect 264790 218056 264796 218068
rect 264388 218028 264796 218056
rect 264388 218016 264394 218028
rect 264790 218016 264796 218028
rect 264848 218016 264854 218068
rect 265158 218016 265164 218068
rect 265216 218056 265222 218068
rect 266170 218056 266176 218068
rect 265216 218028 266176 218056
rect 265216 218016 265222 218028
rect 266170 218016 266176 218028
rect 266228 218016 266234 218068
rect 268470 218016 268476 218068
rect 268528 218056 268534 218068
rect 268930 218056 268936 218068
rect 268528 218028 268936 218056
rect 268528 218016 268534 218028
rect 268930 218016 268936 218028
rect 268988 218016 268994 218068
rect 269298 218016 269304 218068
rect 269356 218056 269362 218068
rect 270034 218056 270040 218068
rect 269356 218028 270040 218056
rect 269356 218016 269362 218028
rect 270034 218016 270040 218028
rect 270092 218016 270098 218068
rect 270954 218016 270960 218068
rect 271012 218056 271018 218068
rect 272518 218056 272524 218068
rect 271012 218028 272524 218056
rect 271012 218016 271018 218028
rect 272518 218016 272524 218028
rect 272576 218016 272582 218068
rect 276750 218016 276756 218068
rect 276808 218056 276814 218068
rect 277210 218056 277216 218068
rect 276808 218028 277216 218056
rect 276808 218016 276814 218028
rect 277210 218016 277216 218028
rect 277268 218016 277274 218068
rect 277578 218016 277584 218068
rect 277636 218056 277642 218068
rect 278590 218056 278596 218068
rect 277636 218028 278596 218056
rect 277636 218016 277642 218028
rect 278590 218016 278596 218028
rect 278648 218016 278654 218068
rect 280890 218016 280896 218068
rect 280948 218056 280954 218068
rect 281442 218056 281448 218068
rect 280948 218028 281448 218056
rect 280948 218016 280954 218028
rect 281442 218016 281448 218028
rect 281500 218016 281506 218068
rect 281718 218016 281724 218068
rect 281776 218056 281782 218068
rect 282454 218056 282460 218068
rect 281776 218028 282460 218056
rect 281776 218016 281782 218028
rect 282454 218016 282460 218028
rect 282512 218016 282518 218068
rect 285030 218016 285036 218068
rect 285088 218056 285094 218068
rect 285490 218056 285496 218068
rect 285088 218028 285496 218056
rect 285088 218016 285094 218028
rect 285490 218016 285496 218028
rect 285548 218016 285554 218068
rect 287514 218016 287520 218068
rect 287572 218056 287578 218068
rect 288710 218056 288716 218068
rect 287572 218028 288716 218056
rect 287572 218016 287578 218028
rect 288710 218016 288716 218028
rect 288768 218016 288774 218068
rect 289170 218016 289176 218068
rect 289228 218056 289234 218068
rect 289722 218056 289728 218068
rect 289228 218028 289728 218056
rect 289228 218016 289234 218028
rect 289722 218016 289728 218028
rect 289780 218016 289786 218068
rect 289998 218016 290004 218068
rect 290056 218056 290062 218068
rect 291102 218056 291108 218068
rect 290056 218028 291108 218056
rect 290056 218016 290062 218028
rect 291102 218016 291108 218028
rect 291160 218016 291166 218068
rect 293310 218016 293316 218068
rect 293368 218056 293374 218068
rect 293770 218056 293776 218068
rect 293368 218028 293776 218056
rect 293368 218016 293374 218028
rect 293770 218016 293776 218028
rect 293828 218016 293834 218068
rect 297450 218016 297456 218068
rect 297508 218056 297514 218068
rect 297910 218056 297916 218068
rect 297508 218028 297916 218056
rect 297508 218016 297514 218028
rect 297910 218016 297916 218028
rect 297968 218016 297974 218068
rect 298278 218016 298284 218068
rect 298336 218056 298342 218068
rect 299106 218056 299112 218068
rect 298336 218028 299112 218056
rect 298336 218016 298342 218028
rect 299106 218016 299112 218028
rect 299164 218016 299170 218068
rect 299934 218016 299940 218068
rect 299992 218056 299998 218068
rect 300670 218056 300676 218068
rect 299992 218028 300676 218056
rect 299992 218016 299998 218028
rect 300670 218016 300676 218028
rect 300728 218016 300734 218068
rect 301590 218016 301596 218068
rect 301648 218056 301654 218068
rect 302142 218056 302148 218068
rect 301648 218028 302148 218056
rect 301648 218016 301654 218028
rect 302142 218016 302148 218028
rect 302200 218016 302206 218068
rect 304074 218016 304080 218068
rect 304132 218056 304138 218068
rect 304718 218056 304724 218068
rect 304132 218028 304724 218056
rect 304132 218016 304138 218028
rect 304718 218016 304724 218028
rect 304776 218016 304782 218068
rect 305730 218016 305736 218068
rect 305788 218056 305794 218068
rect 306190 218056 306196 218068
rect 305788 218028 306196 218056
rect 305788 218016 305794 218028
rect 306190 218016 306196 218028
rect 306248 218016 306254 218068
rect 306558 218016 306564 218068
rect 306616 218056 306622 218068
rect 307662 218056 307668 218068
rect 306616 218028 307668 218056
rect 306616 218016 306622 218028
rect 307662 218016 307668 218028
rect 307720 218016 307726 218068
rect 309870 218016 309876 218068
rect 309928 218056 309934 218068
rect 310422 218056 310428 218068
rect 309928 218028 310428 218056
rect 309928 218016 309934 218028
rect 310422 218016 310428 218028
rect 310480 218016 310486 218068
rect 312354 218016 312360 218068
rect 312412 218056 312418 218068
rect 312906 218056 312912 218068
rect 312412 218028 312912 218056
rect 312412 218016 312418 218028
rect 312906 218016 312912 218028
rect 312964 218016 312970 218068
rect 317322 218016 317328 218068
rect 317380 218056 317386 218068
rect 317966 218056 317972 218068
rect 317380 218028 317972 218056
rect 317380 218016 317386 218028
rect 317966 218016 317972 218028
rect 318024 218016 318030 218068
rect 318978 218016 318984 218068
rect 319036 218056 319042 218068
rect 319806 218056 319812 218068
rect 319036 218028 319812 218056
rect 319036 218016 319042 218028
rect 319806 218016 319812 218028
rect 319864 218016 319870 218068
rect 322290 218016 322296 218068
rect 322348 218056 322354 218068
rect 322842 218056 322848 218068
rect 322348 218028 322848 218056
rect 322348 218016 322354 218028
rect 322842 218016 322848 218028
rect 322900 218016 322906 218068
rect 323118 218016 323124 218068
rect 323176 218056 323182 218068
rect 324130 218056 324136 218068
rect 323176 218028 324136 218056
rect 323176 218016 323182 218028
rect 324130 218016 324136 218028
rect 324188 218016 324194 218068
rect 324774 218016 324780 218068
rect 324832 218056 324838 218068
rect 325418 218056 325424 218068
rect 324832 218028 325424 218056
rect 324832 218016 324838 218028
rect 325418 218016 325424 218028
rect 325476 218016 325482 218068
rect 326430 218016 326436 218068
rect 326488 218056 326494 218068
rect 326890 218056 326896 218068
rect 326488 218028 326896 218056
rect 326488 218016 326494 218028
rect 326890 218016 326896 218028
rect 326948 218016 326954 218068
rect 330570 218016 330576 218068
rect 330628 218056 330634 218068
rect 331030 218056 331036 218068
rect 330628 218028 331036 218056
rect 330628 218016 330634 218028
rect 331030 218016 331036 218028
rect 331088 218016 331094 218068
rect 333054 218016 333060 218068
rect 333112 218056 333118 218068
rect 333882 218056 333888 218068
rect 333112 218028 333888 218056
rect 333112 218016 333118 218028
rect 333882 218016 333888 218028
rect 333940 218016 333946 218068
rect 334710 218016 334716 218068
rect 334768 218056 334774 218068
rect 335170 218056 335176 218068
rect 334768 218028 335176 218056
rect 334768 218016 334774 218028
rect 335170 218016 335176 218028
rect 335228 218016 335234 218068
rect 335538 218016 335544 218068
rect 335596 218056 335602 218068
rect 338666 218056 338672 218068
rect 335596 218028 338672 218056
rect 335596 218016 335602 218028
rect 338666 218016 338672 218028
rect 338724 218016 338730 218068
rect 338850 218016 338856 218068
rect 338908 218056 338914 218068
rect 339402 218056 339408 218068
rect 338908 218028 339408 218056
rect 338908 218016 338914 218028
rect 339402 218016 339408 218028
rect 339460 218016 339466 218068
rect 339678 218016 339684 218068
rect 339736 218056 339742 218068
rect 340690 218056 340696 218068
rect 339736 218028 340696 218056
rect 339736 218016 339742 218028
rect 340690 218016 340696 218028
rect 340748 218016 340754 218068
rect 345474 218016 345480 218068
rect 345532 218056 345538 218068
rect 347038 218056 347044 218068
rect 345532 218028 347044 218056
rect 345532 218016 345538 218028
rect 347038 218016 347044 218028
rect 347096 218016 347102 218068
rect 347958 218016 347964 218068
rect 348016 218056 348022 218068
rect 349062 218056 349068 218068
rect 348016 218028 349068 218056
rect 348016 218016 348022 218028
rect 349062 218016 349068 218028
rect 349120 218016 349126 218068
rect 355410 218016 355416 218068
rect 355468 218056 355474 218068
rect 355870 218056 355876 218068
rect 355468 218028 355876 218056
rect 355468 218016 355474 218028
rect 355870 218016 355876 218028
rect 355928 218016 355934 218068
rect 356238 218016 356244 218068
rect 356296 218056 356302 218068
rect 356974 218056 356980 218068
rect 356296 218028 356980 218056
rect 356296 218016 356302 218028
rect 356974 218016 356980 218028
rect 357032 218016 357038 218068
rect 359550 218016 359556 218068
rect 359608 218056 359614 218068
rect 360102 218056 360108 218068
rect 359608 218028 360108 218056
rect 359608 218016 359614 218028
rect 360102 218016 360108 218028
rect 360160 218016 360166 218068
rect 360378 218016 360384 218068
rect 360436 218056 360442 218068
rect 361022 218056 361028 218068
rect 360436 218028 361028 218056
rect 360436 218016 360442 218028
rect 361022 218016 361028 218028
rect 361080 218016 361086 218068
rect 364518 218016 364524 218068
rect 364576 218056 364582 218068
rect 365530 218056 365536 218068
rect 364576 218028 365536 218056
rect 364576 218016 364582 218028
rect 365530 218016 365536 218028
rect 365588 218016 365594 218068
rect 366174 218016 366180 218068
rect 366232 218056 366238 218068
rect 366726 218056 366732 218068
rect 366232 218028 366732 218056
rect 366232 218016 366238 218028
rect 366726 218016 366732 218028
rect 366784 218016 366790 218068
rect 367830 218016 367836 218068
rect 367888 218056 367894 218068
rect 368382 218056 368388 218068
rect 367888 218028 368388 218056
rect 367888 218016 367894 218028
rect 368382 218016 368388 218028
rect 368440 218016 368446 218068
rect 371970 218016 371976 218068
rect 372028 218056 372034 218068
rect 372522 218056 372528 218068
rect 372028 218028 372528 218056
rect 372028 218016 372034 218028
rect 372522 218016 372528 218028
rect 372580 218016 372586 218068
rect 372798 218016 372804 218068
rect 372856 218056 372862 218068
rect 373442 218056 373448 218068
rect 372856 218028 373448 218056
rect 372856 218016 372862 218028
rect 373442 218016 373448 218028
rect 373500 218016 373506 218068
rect 376110 218016 376116 218068
rect 376168 218056 376174 218068
rect 376662 218056 376668 218068
rect 376168 218028 376668 218056
rect 376168 218016 376174 218028
rect 376662 218016 376668 218028
rect 376720 218016 376726 218068
rect 378594 218016 378600 218068
rect 378652 218056 378658 218068
rect 379238 218056 379244 218068
rect 378652 218028 379244 218056
rect 378652 218016 378658 218028
rect 379238 218016 379244 218028
rect 379296 218016 379302 218068
rect 381078 218016 381084 218068
rect 381136 218056 381142 218068
rect 382090 218056 382096 218068
rect 381136 218028 382096 218056
rect 381136 218016 381142 218028
rect 382090 218016 382096 218028
rect 382148 218016 382154 218068
rect 389358 218016 389364 218068
rect 389416 218056 389422 218068
rect 390002 218056 390008 218068
rect 389416 218028 390008 218056
rect 389416 218016 389422 218028
rect 390002 218016 390008 218028
rect 390060 218016 390066 218068
rect 392670 218016 392676 218068
rect 392728 218056 392734 218068
rect 393130 218056 393136 218068
rect 392728 218028 393136 218056
rect 392728 218016 392734 218028
rect 393130 218016 393136 218028
rect 393188 218016 393194 218068
rect 393498 218016 393504 218068
rect 393556 218056 393562 218068
rect 394510 218056 394516 218068
rect 393556 218028 394516 218056
rect 393556 218016 393562 218028
rect 394510 218016 394516 218028
rect 394568 218016 394574 218068
rect 395154 218016 395160 218068
rect 395212 218056 395218 218068
rect 395798 218056 395804 218068
rect 395212 218028 395804 218056
rect 395212 218016 395218 218028
rect 395798 218016 395804 218028
rect 395856 218016 395862 218068
rect 397638 218016 397644 218068
rect 397696 218056 397702 218068
rect 400674 218056 400680 218068
rect 397696 218028 400680 218056
rect 397696 218016 397702 218028
rect 400674 218016 400680 218028
rect 400732 218016 400738 218068
rect 400950 218016 400956 218068
rect 401008 218056 401014 218068
rect 402238 218056 402244 218068
rect 401008 218028 402244 218056
rect 401008 218016 401014 218028
rect 402238 218016 402244 218028
rect 402296 218016 402302 218068
rect 403434 218016 403440 218068
rect 403492 218056 403498 218068
rect 403986 218056 403992 218068
rect 403492 218028 403992 218056
rect 403492 218016 403498 218028
rect 403986 218016 403992 218028
rect 404044 218016 404050 218068
rect 405090 218016 405096 218068
rect 405148 218056 405154 218068
rect 405550 218056 405556 218068
rect 405148 218028 405556 218056
rect 405148 218016 405154 218028
rect 405550 218016 405556 218028
rect 405608 218016 405614 218068
rect 409230 218016 409236 218068
rect 409288 218056 409294 218068
rect 409782 218056 409788 218068
rect 409288 218028 409788 218056
rect 409288 218016 409294 218028
rect 409782 218016 409788 218028
rect 409840 218016 409846 218068
rect 410058 218016 410064 218068
rect 410116 218056 410122 218068
rect 410702 218056 410708 218068
rect 410116 218028 410708 218056
rect 410116 218016 410122 218028
rect 410702 218016 410708 218028
rect 410760 218016 410766 218068
rect 413370 218016 413376 218068
rect 413428 218056 413434 218068
rect 413830 218056 413836 218068
rect 413428 218028 413836 218056
rect 413428 218016 413434 218028
rect 413830 218016 413836 218028
rect 413888 218016 413894 218068
rect 419994 218016 420000 218068
rect 420052 218056 420058 218068
rect 420914 218056 420920 218068
rect 420052 218028 420920 218056
rect 420052 218016 420058 218028
rect 420914 218016 420920 218028
rect 420972 218016 420978 218068
rect 424134 218016 424140 218068
rect 424192 218056 424198 218068
rect 426986 218056 426992 218068
rect 424192 218028 426992 218056
rect 424192 218016 424198 218028
rect 426986 218016 426992 218028
rect 427044 218016 427050 218068
rect 427446 218016 427452 218068
rect 427504 218056 427510 218068
rect 428458 218056 428464 218068
rect 427504 218028 428464 218056
rect 427504 218016 427510 218028
rect 428458 218016 428464 218028
rect 428516 218016 428522 218068
rect 429102 218016 429108 218068
rect 429160 218056 429166 218068
rect 430574 218056 430580 218068
rect 429160 218028 430580 218056
rect 429160 218016 429166 218028
rect 430574 218016 430580 218028
rect 430632 218016 430638 218068
rect 432414 218016 432420 218068
rect 432472 218056 432478 218068
rect 433794 218056 433800 218068
rect 432472 218028 433800 218056
rect 432472 218016 432478 218028
rect 433794 218016 433800 218028
rect 433852 218016 433858 218068
rect 435726 218016 435732 218068
rect 435784 218056 435790 218068
rect 436278 218056 436284 218068
rect 435784 218028 436284 218056
rect 435784 218016 435790 218028
rect 436278 218016 436284 218028
rect 436336 218016 436342 218068
rect 436462 218016 436468 218068
rect 436520 218056 436526 218068
rect 437750 218056 437756 218068
rect 436520 218028 437756 218056
rect 436520 218016 436526 218028
rect 437750 218016 437756 218028
rect 437808 218016 437814 218068
rect 453298 218016 453304 218068
rect 453356 218056 453362 218068
rect 455414 218056 455420 218068
rect 453356 218028 455420 218056
rect 453356 218016 453362 218028
rect 455414 218016 455420 218028
rect 455472 218016 455478 218068
rect 455598 218016 455604 218068
rect 455656 218056 455662 218068
rect 457162 218056 457168 218068
rect 455656 218028 457168 218056
rect 455656 218016 455662 218028
rect 457162 218016 457168 218028
rect 457220 218016 457226 218068
rect 463142 218016 463148 218068
rect 463200 218056 463206 218068
rect 464614 218056 464620 218068
rect 463200 218028 464620 218056
rect 463200 218016 463206 218028
rect 464614 218016 464620 218028
rect 464672 218016 464678 218068
rect 467282 218016 467288 218068
rect 467340 218056 467346 218068
rect 467926 218056 467932 218068
rect 467340 218028 467932 218056
rect 467340 218016 467346 218028
rect 467926 218016 467932 218028
rect 467984 218016 467990 218068
rect 471422 218016 471428 218068
rect 471480 218056 471486 218068
rect 472894 218056 472900 218068
rect 471480 218028 472900 218056
rect 471480 218016 471486 218028
rect 472894 218016 472900 218028
rect 472952 218016 472958 218068
rect 490374 218016 490380 218068
rect 490432 218056 490438 218068
rect 490432 218028 496860 218056
rect 490432 218016 490438 218028
rect 174556 217892 176240 217920
rect 496832 217920 496860 218028
rect 496998 218016 497004 218068
rect 497056 218056 497062 218068
rect 497458 218056 497464 218068
rect 497056 218028 497464 218056
rect 497056 218016 497062 218028
rect 497458 218016 497464 218028
rect 497516 218016 497522 218068
rect 497660 218028 563100 218056
rect 497660 217920 497688 218028
rect 563072 217988 563100 218028
rect 563210 217988 563238 218096
rect 572824 218056 572852 218096
rect 572824 218028 605834 218056
rect 563072 217960 563238 217988
rect 563606 217948 563612 218000
rect 563664 217988 563670 218000
rect 571886 217988 571892 218000
rect 563664 217960 571892 217988
rect 563664 217948 563670 217960
rect 571886 217948 571892 217960
rect 571944 217948 571950 218000
rect 605806 217988 605834 218028
rect 612274 217988 612280 218000
rect 605806 217960 612280 217988
rect 612274 217948 612280 217960
rect 612332 217948 612338 218000
rect 613856 217988 613884 218164
rect 614482 217988 614488 218000
rect 613856 217960 614488 217988
rect 614482 217948 614488 217960
rect 614540 217948 614546 218000
rect 496832 217892 497688 217920
rect 451366 217812 451372 217864
rect 451424 217852 451430 217864
rect 452194 217852 452200 217864
rect 451424 217824 452200 217852
rect 451424 217812 451430 217824
rect 452194 217812 452200 217824
rect 452252 217812 452258 217864
rect 523034 217812 523040 217864
rect 523092 217852 523098 217864
rect 524230 217852 524236 217864
rect 523092 217824 524236 217852
rect 523092 217812 523098 217824
rect 524230 217812 524236 217824
rect 524288 217812 524294 217864
rect 536374 217812 536380 217864
rect 536432 217852 536438 217864
rect 603994 217852 604000 217864
rect 536432 217824 604000 217852
rect 536432 217812 536438 217824
rect 603994 217812 604000 217824
rect 604052 217812 604058 217864
rect 527818 217676 527824 217728
rect 527876 217716 527882 217728
rect 528370 217716 528376 217728
rect 527876 217688 528376 217716
rect 527876 217676 527882 217688
rect 528370 217676 528376 217688
rect 528428 217716 528434 217728
rect 603258 217716 603264 217728
rect 528428 217688 603264 217716
rect 528428 217676 528434 217688
rect 603258 217676 603264 217688
rect 603316 217676 603322 217728
rect 604454 217676 604460 217728
rect 604512 217716 604518 217728
rect 614298 217716 614304 217728
rect 604512 217688 614304 217716
rect 604512 217676 604518 217688
rect 614298 217676 614304 217688
rect 614356 217676 614362 217728
rect 116946 217540 116952 217592
rect 117004 217580 117010 217592
rect 189166 217580 189172 217592
rect 117004 217552 189172 217580
rect 117004 217540 117010 217552
rect 189166 217540 189172 217552
rect 189224 217540 189230 217592
rect 533430 217540 533436 217592
rect 533488 217580 533494 217592
rect 536374 217580 536380 217592
rect 533488 217552 536380 217580
rect 533488 217540 533494 217552
rect 536374 217540 536380 217552
rect 536432 217540 536438 217592
rect 542354 217540 542360 217592
rect 542412 217580 542418 217592
rect 543274 217580 543280 217592
rect 542412 217552 543280 217580
rect 542412 217540 542418 217552
rect 543274 217540 543280 217552
rect 543332 217580 543338 217592
rect 606202 217580 606208 217592
rect 543332 217552 606208 217580
rect 543332 217540 543338 217552
rect 606202 217540 606208 217552
rect 606260 217540 606266 217592
rect 614114 217540 614120 217592
rect 614172 217580 614178 217592
rect 626626 217580 626632 217592
rect 614172 217552 626632 217580
rect 614172 217540 614178 217552
rect 626626 217540 626632 217552
rect 626684 217540 626690 217592
rect 669866 217472 669872 217524
rect 669924 217472 669930 217524
rect 115290 217404 115296 217456
rect 115348 217444 115354 217456
rect 187970 217444 187976 217456
rect 115348 217416 187976 217444
rect 115348 217404 115354 217416
rect 187970 217404 187976 217416
rect 188028 217404 188034 217456
rect 530946 217404 530952 217456
rect 531004 217444 531010 217456
rect 531004 217416 598704 217444
rect 531004 217404 531010 217416
rect 168558 217308 168564 217320
rect 93826 217280 168564 217308
rect 90404 217200 90410 217252
rect 90462 217240 90468 217252
rect 93826 217240 93854 217280
rect 168558 217268 168564 217280
rect 168616 217268 168622 217320
rect 508590 217268 508596 217320
rect 508648 217308 508654 217320
rect 563008 217308 563014 217320
rect 508648 217280 563014 217308
rect 508648 217268 508654 217280
rect 563008 217268 563014 217280
rect 563066 217268 563072 217320
rect 563146 217268 563152 217320
rect 563204 217308 563210 217320
rect 572530 217308 572536 217320
rect 563204 217280 572536 217308
rect 563204 217268 563210 217280
rect 572530 217268 572536 217280
rect 572588 217268 572594 217320
rect 572714 217268 572720 217320
rect 572772 217308 572778 217320
rect 598474 217308 598480 217320
rect 572772 217280 598480 217308
rect 572772 217268 572778 217280
rect 598474 217268 598480 217280
rect 598532 217268 598538 217320
rect 90462 217212 93854 217240
rect 90462 217200 90468 217212
rect 447134 217200 447140 217252
rect 447192 217240 447198 217252
rect 448100 217240 448106 217252
rect 447192 217212 448106 217240
rect 447192 217200 447198 217212
rect 448100 217200 448106 217212
rect 448158 217200 448164 217252
rect 448606 217200 448612 217252
rect 448664 217240 448670 217252
rect 449756 217240 449762 217252
rect 448664 217212 449762 217240
rect 448664 217200 448670 217212
rect 449756 217200 449762 217212
rect 449814 217200 449820 217252
rect 469306 217200 469312 217252
rect 469364 217240 469370 217252
rect 470456 217240 470462 217252
rect 469364 217212 470462 217240
rect 469364 217200 469370 217212
rect 470456 217200 470462 217212
rect 470514 217200 470520 217252
rect 498194 217200 498200 217252
rect 498252 217240 498258 217252
rect 499436 217240 499442 217252
rect 498252 217212 499442 217240
rect 498252 217200 498258 217212
rect 499436 217200 499442 217212
rect 499494 217200 499500 217252
rect 506060 217132 506066 217184
rect 506118 217172 506124 217184
rect 597922 217172 597928 217184
rect 506118 217144 597928 217172
rect 506118 217132 506124 217144
rect 597922 217132 597928 217144
rect 597980 217132 597986 217184
rect 598676 217172 598704 217416
rect 603074 217404 603080 217456
rect 603132 217444 603138 217456
rect 628282 217444 628288 217456
rect 603132 217416 628288 217444
rect 603132 217404 603138 217416
rect 628282 217404 628288 217416
rect 628340 217404 628346 217456
rect 598842 217268 598848 217320
rect 598900 217308 598906 217320
rect 622394 217308 622400 217320
rect 598900 217280 622400 217308
rect 598900 217268 598906 217280
rect 622394 217268 622400 217280
rect 622452 217268 622458 217320
rect 603442 217172 603448 217184
rect 598676 217144 603448 217172
rect 603442 217132 603448 217144
rect 603500 217132 603506 217184
rect 669884 217116 669912 217472
rect 498608 217064 498614 217116
rect 498666 217104 498672 217116
rect 498666 217076 499574 217104
rect 498666 217064 498672 217076
rect 499546 217036 499574 217076
rect 669866 217064 669872 217116
rect 669924 217064 669930 217116
rect 499546 217008 574048 217036
rect 574020 216900 574048 217008
rect 574186 216996 574192 217048
rect 574244 217036 574250 217048
rect 610066 217036 610072 217048
rect 574244 217008 610072 217036
rect 574244 216996 574250 217008
rect 610066 216996 610072 217008
rect 610124 216996 610130 217048
rect 596358 216900 596364 216912
rect 574020 216872 596364 216900
rect 596358 216860 596364 216872
rect 596416 216860 596422 216912
rect 613378 216900 613384 216912
rect 605806 216872 613384 216900
rect 594794 216724 594800 216776
rect 594852 216764 594858 216776
rect 605806 216764 605834 216872
rect 613378 216860 613384 216872
rect 613436 216860 613442 216912
rect 594852 216736 605834 216764
rect 594852 216724 594858 216736
rect 610710 216724 610716 216776
rect 610768 216764 610774 216776
rect 615678 216764 615684 216776
rect 610768 216736 615684 216764
rect 610768 216724 610774 216736
rect 615678 216724 615684 216736
rect 615736 216724 615742 216776
rect 648246 216656 648252 216708
rect 648304 216696 648310 216708
rect 650638 216696 650644 216708
rect 648304 216668 650644 216696
rect 648304 216656 648310 216668
rect 650638 216656 650644 216668
rect 650696 216656 650702 216708
rect 644934 215908 644940 215960
rect 644992 215948 644998 215960
rect 658918 215948 658924 215960
rect 644992 215920 658924 215948
rect 644992 215908 644998 215920
rect 658918 215908 658924 215920
rect 658976 215908 658982 215960
rect 675846 215160 675852 215212
rect 675904 215200 675910 215212
rect 676766 215200 676772 215212
rect 675904 215172 676772 215200
rect 675904 215160 675910 215172
rect 676766 215160 676772 215172
rect 676824 215160 676830 215212
rect 574738 214820 574744 214872
rect 574796 214860 574802 214872
rect 616874 214860 616880 214872
rect 574796 214832 616880 214860
rect 574796 214820 574802 214832
rect 616874 214820 616880 214832
rect 616932 214820 616938 214872
rect 574554 214684 574560 214736
rect 574612 214724 574618 214736
rect 623314 214724 623320 214736
rect 574612 214696 623320 214724
rect 574612 214684 574618 214696
rect 623314 214684 623320 214696
rect 623372 214684 623378 214736
rect 658182 214684 658188 214736
rect 658240 214724 658246 214736
rect 665818 214724 665824 214736
rect 658240 214696 665824 214724
rect 658240 214684 658246 214696
rect 665818 214684 665824 214696
rect 665876 214684 665882 214736
rect 574370 214548 574376 214600
rect 574428 214588 574434 214600
rect 574428 214560 605834 214588
rect 574428 214548 574434 214560
rect 600498 214412 600504 214464
rect 600556 214452 600562 214464
rect 601234 214452 601240 214464
rect 600556 214424 601240 214452
rect 600556 214412 600562 214424
rect 601234 214412 601240 214424
rect 601292 214412 601298 214464
rect 605806 214452 605834 214560
rect 618254 214548 618260 214600
rect 618312 214588 618318 214600
rect 618898 214588 618904 214600
rect 618312 214560 618904 214588
rect 618312 214548 618318 214560
rect 618898 214548 618904 214560
rect 618956 214548 618962 214600
rect 619910 214548 619916 214600
rect 619968 214588 619974 214600
rect 620554 214588 620560 214600
rect 619968 214560 620560 214588
rect 619968 214548 619974 214560
rect 620554 214548 620560 214560
rect 620612 214548 620618 214600
rect 623958 214548 623964 214600
rect 624016 214588 624022 214600
rect 624016 214560 625154 214588
rect 624016 214548 624022 214560
rect 624418 214452 624424 214464
rect 605806 214424 624424 214452
rect 624418 214412 624424 214424
rect 624476 214412 624482 214464
rect 625126 214452 625154 214560
rect 625246 214548 625252 214600
rect 625304 214588 625310 214600
rect 626074 214588 626080 214600
rect 625304 214560 626080 214588
rect 625304 214548 625310 214560
rect 626074 214548 626080 214560
rect 626132 214548 626138 214600
rect 630030 214548 630036 214600
rect 630088 214588 630094 214600
rect 632882 214588 632888 214600
rect 630088 214560 632888 214588
rect 630088 214548 630094 214560
rect 632882 214548 632888 214560
rect 632940 214548 632946 214600
rect 646314 214548 646320 214600
rect 646372 214588 646378 214600
rect 656158 214588 656164 214600
rect 646372 214560 656164 214588
rect 646372 214548 646378 214560
rect 656158 214548 656164 214560
rect 656216 214548 656222 214600
rect 629386 214452 629392 214464
rect 625126 214424 629392 214452
rect 629386 214412 629392 214424
rect 629444 214412 629450 214464
rect 35802 214072 35808 214124
rect 35860 214112 35866 214124
rect 39758 214112 39764 214124
rect 35860 214084 39764 214112
rect 35860 214072 35866 214084
rect 39758 214072 39764 214084
rect 39816 214072 39822 214124
rect 645854 213868 645860 213920
rect 645912 213908 645918 213920
rect 646498 213908 646504 213920
rect 645912 213880 646504 213908
rect 645912 213868 645918 213880
rect 646498 213868 646504 213880
rect 646556 213868 646562 213920
rect 654594 213868 654600 213920
rect 654652 213908 654658 213920
rect 657538 213908 657544 213920
rect 654652 213880 657544 213908
rect 654652 213868 654658 213880
rect 657538 213868 657544 213880
rect 657596 213868 657602 213920
rect 663150 213868 663156 213920
rect 663208 213908 663214 213920
rect 663702 213908 663708 213920
rect 663208 213880 663708 213908
rect 663208 213868 663214 213880
rect 663702 213868 663708 213880
rect 663760 213868 663766 213920
rect 653214 213732 653220 213784
rect 653272 213772 653278 213784
rect 654778 213772 654784 213784
rect 653272 213744 654784 213772
rect 653272 213732 653278 213744
rect 654778 213732 654784 213744
rect 654836 213732 654842 213784
rect 648614 213392 648620 213444
rect 648672 213432 648678 213444
rect 649258 213432 649264 213444
rect 648672 213404 649264 213432
rect 648672 213392 648678 213404
rect 649258 213392 649264 213404
rect 649316 213392 649322 213444
rect 654134 213392 654140 213444
rect 654192 213432 654198 213444
rect 654778 213432 654784 213444
rect 654192 213404 654784 213432
rect 654192 213392 654198 213404
rect 654778 213392 654784 213404
rect 654836 213392 654842 213444
rect 656526 213392 656532 213444
rect 656584 213432 656590 213444
rect 664622 213432 664628 213444
rect 656584 213404 664628 213432
rect 656584 213392 656590 213404
rect 664622 213392 664628 213404
rect 664680 213392 664686 213444
rect 643830 213324 643836 213376
rect 643888 213364 643894 213376
rect 643888 213336 644474 213364
rect 643888 213324 643894 213336
rect 644446 213296 644474 213336
rect 653398 213296 653404 213308
rect 644446 213268 653404 213296
rect 653398 213256 653404 213268
rect 653456 213256 653462 213308
rect 575474 213188 575480 213240
rect 575532 213228 575538 213240
rect 594794 213228 594800 213240
rect 575532 213200 594800 213228
rect 575532 213188 575538 213200
rect 594794 213188 594800 213200
rect 594852 213188 594858 213240
rect 660758 213228 660764 213240
rect 654106 213200 660764 213228
rect 645486 213120 645492 213172
rect 645544 213160 645550 213172
rect 654106 213160 654134 213200
rect 660758 213188 660764 213200
rect 660816 213188 660822 213240
rect 645544 213132 654134 213160
rect 645544 213120 645550 213132
rect 632698 212984 632704 213036
rect 632756 213024 632762 213036
rect 634354 213024 634360 213036
rect 632756 212996 634360 213024
rect 632756 212984 632762 212996
rect 634354 212984 634360 212996
rect 634412 212984 634418 213036
rect 650454 212712 650460 212764
rect 650512 212752 650518 212764
rect 651282 212752 651288 212764
rect 650512 212724 651288 212752
rect 650512 212712 650518 212724
rect 651282 212712 651288 212724
rect 651340 212712 651346 212764
rect 664254 212712 664260 212764
rect 664312 212752 664318 212764
rect 665082 212752 665088 212764
rect 664312 212724 665088 212752
rect 664312 212712 664318 212724
rect 665082 212712 665088 212724
rect 665140 212712 665146 212764
rect 35802 212644 35808 212696
rect 35860 212684 35866 212696
rect 39850 212684 39856 212696
rect 35860 212656 39856 212684
rect 35860 212644 35866 212656
rect 39850 212644 39856 212656
rect 39908 212644 39914 212696
rect 592678 212644 592684 212696
rect 592736 212684 592742 212696
rect 641714 212684 641720 212696
rect 592736 212656 641720 212684
rect 592736 212644 592742 212656
rect 641714 212644 641720 212656
rect 641772 212644 641778 212696
rect 591298 212508 591304 212560
rect 591356 212548 591362 212560
rect 639874 212548 639880 212560
rect 591356 212520 639880 212548
rect 591356 212508 591362 212520
rect 639874 212508 639880 212520
rect 639932 212508 639938 212560
rect 35802 211420 35808 211472
rect 35860 211460 35866 211472
rect 40126 211460 40132 211472
rect 35860 211432 40132 211460
rect 35860 211420 35866 211432
rect 40126 211420 40132 211432
rect 40184 211420 40190 211472
rect 35618 211148 35624 211200
rect 35676 211188 35682 211200
rect 40770 211188 40776 211200
rect 35676 211160 40776 211188
rect 35676 211148 35682 211160
rect 40770 211148 40776 211160
rect 40828 211148 40834 211200
rect 578510 211148 578516 211200
rect 578568 211188 578574 211200
rect 580902 211188 580908 211200
rect 578568 211160 580908 211188
rect 578568 211148 578574 211160
rect 580902 211148 580908 211160
rect 580960 211148 580966 211200
rect 600314 210060 600320 210112
rect 600372 210100 600378 210112
rect 600682 210100 600688 210112
rect 600372 210072 600688 210100
rect 600372 210060 600378 210072
rect 600682 210060 600688 210072
rect 600740 210060 600746 210112
rect 35802 209788 35808 209840
rect 35860 209828 35866 209840
rect 39206 209828 39212 209840
rect 35860 209800 39212 209828
rect 35860 209788 35866 209800
rect 39206 209788 39212 209800
rect 39264 209788 39270 209840
rect 579522 209788 579528 209840
rect 579580 209828 579586 209840
rect 582282 209828 582288 209840
rect 579580 209800 582288 209828
rect 579580 209788 579586 209800
rect 582282 209788 582288 209800
rect 582340 209788 582346 209840
rect 632146 209556 632152 209568
rect 625126 209528 632152 209556
rect 35802 208632 35808 208684
rect 35860 208672 35866 208684
rect 39942 208672 39948 208684
rect 35860 208644 39948 208672
rect 35860 208632 35866 208644
rect 39942 208632 39948 208644
rect 40000 208632 40006 208684
rect 581638 208564 581644 208616
rect 581696 208604 581702 208616
rect 625126 208604 625154 209528
rect 632146 209516 632152 209528
rect 632204 209516 632210 209568
rect 652018 209516 652024 209568
rect 652076 209556 652082 209568
rect 652076 209528 654134 209556
rect 652076 209516 652082 209528
rect 654106 209080 654134 209528
rect 667014 209080 667020 209092
rect 654106 209052 667020 209080
rect 667014 209040 667020 209052
rect 667072 209040 667078 209092
rect 581696 208576 625154 208604
rect 581696 208564 581702 208576
rect 35618 208360 35624 208412
rect 35676 208400 35682 208412
rect 40954 208400 40960 208412
rect 35676 208372 40960 208400
rect 35676 208360 35682 208372
rect 40954 208360 40960 208372
rect 41012 208360 41018 208412
rect 578878 208292 578884 208344
rect 578936 208332 578942 208344
rect 589458 208332 589464 208344
rect 578936 208304 589464 208332
rect 578936 208292 578942 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 35802 207136 35808 207188
rect 35860 207176 35866 207188
rect 40954 207176 40960 207188
rect 35860 207148 40960 207176
rect 35860 207136 35866 207148
rect 40954 207136 40960 207148
rect 41012 207136 41018 207188
rect 580902 206864 580908 206916
rect 580960 206904 580966 206916
rect 589458 206904 589464 206916
rect 580960 206876 589464 206904
rect 580960 206864 580966 206876
rect 589458 206864 589464 206876
rect 589516 206864 589522 206916
rect 35802 205776 35808 205828
rect 35860 205816 35866 205828
rect 41690 205816 41696 205828
rect 35860 205788 41696 205816
rect 35860 205776 35866 205788
rect 41690 205776 41696 205788
rect 41748 205776 41754 205828
rect 579522 205776 579528 205828
rect 579580 205816 579586 205828
rect 580994 205816 581000 205828
rect 579580 205788 581000 205816
rect 579580 205776 579586 205788
rect 580994 205776 581000 205788
rect 581052 205776 581058 205828
rect 42058 205504 42064 205556
rect 42116 205544 42122 205556
rect 43346 205544 43352 205556
rect 42116 205516 43352 205544
rect 42116 205504 42122 205516
rect 43346 205504 43352 205516
rect 43404 205504 43410 205556
rect 582282 205504 582288 205556
rect 582340 205544 582346 205556
rect 589458 205544 589464 205556
rect 582340 205516 589464 205544
rect 582340 205504 582346 205516
rect 589458 205504 589464 205516
rect 589516 205504 589522 205556
rect 35802 204620 35808 204672
rect 35860 204660 35866 204672
rect 35860 204620 35894 204660
rect 35866 204592 35894 204620
rect 35866 204564 41414 204592
rect 41386 204524 41414 204564
rect 41690 204524 41696 204536
rect 41386 204496 41696 204524
rect 41690 204484 41696 204496
rect 41748 204484 41754 204536
rect 35802 204280 35808 204332
rect 35860 204320 35866 204332
rect 39390 204320 39396 204332
rect 35860 204292 39396 204320
rect 35860 204280 35866 204292
rect 39390 204280 39396 204292
rect 39448 204280 39454 204332
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 35802 202852 35808 202904
rect 35860 202892 35866 202904
rect 39298 202892 39304 202904
rect 35860 202864 39304 202892
rect 35860 202852 35866 202864
rect 39298 202852 39304 202864
rect 39356 202852 39362 202904
rect 578326 202852 578332 202904
rect 578384 202892 578390 202904
rect 580258 202892 580264 202904
rect 578384 202864 580264 202892
rect 578384 202852 578390 202864
rect 580258 202852 580264 202864
rect 580316 202852 580322 202904
rect 580994 202784 581000 202836
rect 581052 202824 581058 202836
rect 589458 202824 589464 202836
rect 581052 202796 589464 202824
rect 581052 202784 581058 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 578786 200132 578792 200184
rect 578844 200172 578850 200184
rect 590378 200172 590384 200184
rect 578844 200144 590384 200172
rect 578844 200132 578850 200144
rect 590378 200132 590384 200144
rect 590436 200132 590442 200184
rect 580258 199996 580264 200048
rect 580316 200036 580322 200048
rect 589458 200036 589464 200048
rect 580316 200008 589464 200036
rect 580316 199996 580322 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 579522 198704 579528 198756
rect 579580 198744 579586 198756
rect 589458 198744 589464 198756
rect 579580 198716 589464 198744
rect 579580 198704 579586 198716
rect 589458 198704 589464 198716
rect 589516 198704 589522 198756
rect 42702 197072 42708 197124
rect 42760 197112 42766 197124
rect 43346 197112 43352 197124
rect 42760 197084 43352 197112
rect 42760 197072 42766 197084
rect 43346 197072 43352 197084
rect 43404 197072 43410 197124
rect 578510 195984 578516 196036
rect 578568 196024 578574 196036
rect 589274 196024 589280 196036
rect 578568 195996 589280 196024
rect 578568 195984 578574 195996
rect 589274 195984 589280 195996
rect 589332 195984 589338 196036
rect 579522 194556 579528 194608
rect 579580 194596 579586 194608
rect 589458 194596 589464 194608
rect 579580 194568 589464 194596
rect 579580 194556 579586 194568
rect 589458 194556 589464 194568
rect 589516 194556 589522 194608
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 589458 191876 589464 191888
rect 579580 191848 589464 191876
rect 579580 191836 579586 191848
rect 589458 191836 589464 191848
rect 589516 191836 589522 191888
rect 579522 190476 579528 190528
rect 579580 190516 579586 190528
rect 590562 190516 590568 190528
rect 579580 190488 590568 190516
rect 579580 190476 579586 190488
rect 590562 190476 590568 190488
rect 590620 190476 590626 190528
rect 579522 187688 579528 187740
rect 579580 187728 579586 187740
rect 589458 187728 589464 187740
rect 579580 187700 589464 187728
rect 579580 187688 579586 187700
rect 589458 187688 589464 187700
rect 589516 187688 589522 187740
rect 42426 187280 42432 187332
rect 42484 187320 42490 187332
rect 43070 187320 43076 187332
rect 42484 187292 43076 187320
rect 42484 187280 42490 187292
rect 43070 187280 43076 187292
rect 43128 187280 43134 187332
rect 579522 186260 579528 186312
rect 579580 186300 579586 186312
rect 589642 186300 589648 186312
rect 579580 186272 589648 186300
rect 579580 186260 579586 186272
rect 589642 186260 589648 186272
rect 589700 186260 589706 186312
rect 579522 184832 579528 184884
rect 579580 184872 579586 184884
rect 589458 184872 589464 184884
rect 579580 184844 589464 184872
rect 579580 184832 579586 184844
rect 589458 184832 589464 184844
rect 589516 184832 589522 184884
rect 668946 184832 668952 184884
rect 669004 184872 669010 184884
rect 670694 184872 670700 184884
rect 669004 184844 670700 184872
rect 669004 184832 669010 184844
rect 670694 184832 670700 184844
rect 670752 184832 670758 184884
rect 42426 182112 42432 182164
rect 42484 182152 42490 182164
rect 43254 182152 43260 182164
rect 42484 182124 43260 182152
rect 42484 182112 42490 182124
rect 43254 182112 43260 182124
rect 43312 182112 43318 182164
rect 579522 182112 579528 182164
rect 579580 182152 579586 182164
rect 589458 182152 589464 182164
rect 579580 182124 589464 182152
rect 579580 182112 579586 182124
rect 589458 182112 589464 182124
rect 589516 182112 589522 182164
rect 578786 180752 578792 180804
rect 578844 180792 578850 180804
rect 590562 180792 590568 180804
rect 578844 180764 590568 180792
rect 578844 180752 578850 180764
rect 590562 180752 590568 180764
rect 590620 180752 590626 180804
rect 578786 178032 578792 178084
rect 578844 178072 578850 178084
rect 589458 178072 589464 178084
rect 578844 178044 589464 178072
rect 578844 178032 578850 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 668210 177964 668216 178016
rect 668268 178004 668274 178016
rect 670786 178004 670792 178016
rect 668268 177976 670792 178004
rect 668268 177964 668274 177976
rect 670786 177964 670792 177976
rect 670844 177964 670850 178016
rect 579522 177896 579528 177948
rect 579580 177936 579586 177948
rect 589642 177936 589648 177948
rect 579580 177908 589648 177936
rect 579580 177896 579586 177908
rect 589642 177896 589648 177908
rect 589700 177896 589706 177948
rect 589458 175352 589464 175364
rect 586486 175324 589464 175352
rect 579982 175244 579988 175296
rect 580040 175284 580046 175296
rect 586486 175284 586514 175324
rect 589458 175312 589464 175324
rect 589516 175312 589522 175364
rect 580040 175256 586514 175284
rect 580040 175244 580046 175256
rect 668026 175040 668032 175092
rect 668084 175080 668090 175092
rect 670418 175080 670424 175092
rect 668084 175052 670424 175080
rect 668084 175040 668090 175052
rect 670418 175040 670424 175052
rect 670476 175040 670482 175092
rect 578418 174496 578424 174548
rect 578476 174536 578482 174548
rect 589642 174536 589648 174548
rect 578476 174508 589648 174536
rect 578476 174496 578482 174508
rect 589642 174496 589648 174508
rect 589700 174496 589706 174548
rect 578234 172864 578240 172916
rect 578292 172904 578298 172916
rect 579982 172904 579988 172916
rect 578292 172876 579988 172904
rect 578292 172864 578298 172876
rect 579982 172864 579988 172876
rect 580040 172864 580046 172916
rect 580902 172524 580908 172576
rect 580960 172564 580966 172576
rect 589458 172564 589464 172576
rect 580960 172536 589464 172564
rect 580960 172524 580966 172536
rect 589458 172524 589464 172536
rect 589516 172524 589522 172576
rect 580258 171096 580264 171148
rect 580316 171136 580322 171148
rect 589458 171136 589464 171148
rect 580316 171108 589464 171136
rect 580316 171096 580322 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 578694 169736 578700 169788
rect 578752 169776 578758 169788
rect 580902 169776 580908 169788
rect 578752 169748 580908 169776
rect 578752 169736 578758 169748
rect 580902 169736 580908 169748
rect 580960 169736 580966 169788
rect 667934 169668 667940 169720
rect 667992 169708 667998 169720
rect 669682 169708 669688 169720
rect 667992 169680 669688 169708
rect 667992 169668 667998 169680
rect 669682 169668 669688 169680
rect 669740 169668 669746 169720
rect 582374 168376 582380 168428
rect 582432 168416 582438 168428
rect 589458 168416 589464 168428
rect 582432 168388 589464 168416
rect 582432 168376 582438 168388
rect 589458 168376 589464 168388
rect 589516 168376 589522 168428
rect 578234 167288 578240 167340
rect 578292 167328 578298 167340
rect 580258 167328 580264 167340
rect 578292 167300 580264 167328
rect 578292 167288 578298 167300
rect 580258 167288 580264 167300
rect 580316 167288 580322 167340
rect 579982 167016 579988 167068
rect 580040 167056 580046 167068
rect 589458 167056 589464 167068
rect 580040 167028 589464 167056
rect 580040 167016 580046 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 579522 166268 579528 166320
rect 579580 166308 579586 166320
rect 589642 166308 589648 166320
rect 579580 166280 589648 166308
rect 579580 166268 579586 166280
rect 589642 166268 589648 166280
rect 589700 166268 589706 166320
rect 579338 165180 579344 165232
rect 579396 165220 579402 165232
rect 582374 165220 582380 165232
rect 579396 165192 582380 165220
rect 579396 165180 579402 165192
rect 582374 165180 582380 165192
rect 582432 165180 582438 165232
rect 667934 165044 667940 165096
rect 667992 165084 667998 165096
rect 670050 165084 670056 165096
rect 667992 165056 670056 165084
rect 667992 165044 667998 165056
rect 670050 165044 670056 165056
rect 670108 165044 670114 165096
rect 582466 164228 582472 164280
rect 582524 164268 582530 164280
rect 589458 164268 589464 164280
rect 582524 164240 589464 164268
rect 582524 164228 582530 164240
rect 589458 164228 589464 164240
rect 589516 164228 589522 164280
rect 675846 164160 675852 164212
rect 675904 164200 675910 164212
rect 682378 164200 682384 164212
rect 675904 164172 682384 164200
rect 675904 164160 675910 164172
rect 682378 164160 682384 164172
rect 682436 164160 682442 164212
rect 578234 163616 578240 163668
rect 578292 163656 578298 163668
rect 579982 163656 579988 163668
rect 578292 163628 579988 163656
rect 578292 163616 578298 163628
rect 579982 163616 579988 163628
rect 580040 163616 580046 163668
rect 580902 162868 580908 162920
rect 580960 162908 580966 162920
rect 589458 162908 589464 162920
rect 580960 162880 589464 162908
rect 580960 162868 580966 162880
rect 589458 162868 589464 162880
rect 589516 162868 589522 162920
rect 578418 162664 578424 162716
rect 578476 162704 578482 162716
rect 582466 162704 582472 162716
rect 578476 162676 582472 162704
rect 578476 162664 578482 162676
rect 582466 162664 582472 162676
rect 582524 162664 582530 162716
rect 580534 161440 580540 161492
rect 580592 161480 580598 161492
rect 589458 161480 589464 161492
rect 580592 161452 589464 161480
rect 580592 161440 580598 161452
rect 589458 161440 589464 161452
rect 589516 161440 589522 161492
rect 580718 160080 580724 160132
rect 580776 160120 580782 160132
rect 589458 160120 589464 160132
rect 580776 160092 589464 160120
rect 580776 160080 580782 160092
rect 589458 160080 589464 160092
rect 589516 160080 589522 160132
rect 668210 160012 668216 160064
rect 668268 160052 668274 160064
rect 670786 160052 670792 160064
rect 668268 160024 670792 160052
rect 668268 160012 668274 160024
rect 670786 160012 670792 160024
rect 670844 160012 670850 160064
rect 578878 158720 578884 158772
rect 578936 158760 578942 158772
rect 580902 158760 580908 158772
rect 578936 158732 580908 158760
rect 578936 158720 578942 158732
rect 580902 158720 580908 158732
rect 580960 158720 580966 158772
rect 585778 158720 585784 158772
rect 585836 158760 585842 158772
rect 589458 158760 589464 158772
rect 585836 158732 589464 158760
rect 585836 158720 585842 158732
rect 589458 158720 589464 158732
rect 589516 158720 589522 158772
rect 587158 157360 587164 157412
rect 587216 157400 587222 157412
rect 589274 157400 589280 157412
rect 587216 157372 589280 157400
rect 587216 157360 587222 157372
rect 589274 157360 589280 157372
rect 589332 157360 589338 157412
rect 668210 155524 668216 155576
rect 668268 155564 668274 155576
rect 670786 155564 670792 155576
rect 668268 155536 670792 155564
rect 668268 155524 668274 155536
rect 670786 155524 670792 155536
rect 670844 155524 670850 155576
rect 578326 154640 578332 154692
rect 578384 154680 578390 154692
rect 580534 154680 580540 154692
rect 578384 154652 580540 154680
rect 578384 154640 578390 154652
rect 580534 154640 580540 154652
rect 580592 154640 580598 154692
rect 584398 154572 584404 154624
rect 584456 154612 584462 154624
rect 589458 154612 589464 154624
rect 584456 154584 589464 154612
rect 584456 154572 584462 154584
rect 589458 154572 589464 154584
rect 589516 154572 589522 154624
rect 583018 153212 583024 153264
rect 583076 153252 583082 153264
rect 589458 153252 589464 153264
rect 583076 153224 589464 153252
rect 583076 153212 583082 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 578234 152736 578240 152788
rect 578292 152776 578298 152788
rect 580718 152776 580724 152788
rect 578292 152748 580724 152776
rect 578292 152736 578298 152748
rect 580718 152736 580724 152748
rect 580776 152736 580782 152788
rect 580258 151784 580264 151836
rect 580316 151824 580322 151836
rect 589458 151824 589464 151836
rect 580316 151796 589464 151824
rect 580316 151784 580322 151796
rect 589458 151784 589464 151796
rect 589516 151784 589522 151836
rect 578878 150560 578884 150612
rect 578936 150600 578942 150612
rect 585778 150600 585784 150612
rect 578936 150572 585784 150600
rect 578936 150560 578942 150572
rect 585778 150560 585784 150572
rect 585836 150560 585842 150612
rect 585134 149064 585140 149116
rect 585192 149104 585198 149116
rect 589458 149104 589464 149116
rect 585192 149076 589464 149104
rect 585192 149064 585198 149076
rect 589458 149064 589464 149076
rect 589516 149064 589522 149116
rect 579522 148316 579528 148368
rect 579580 148356 579586 148368
rect 587158 148356 587164 148368
rect 579580 148328 587164 148356
rect 579580 148316 579586 148328
rect 587158 148316 587164 148328
rect 587216 148316 587222 148368
rect 578878 146276 578884 146328
rect 578936 146316 578942 146328
rect 585134 146316 585140 146328
rect 578936 146288 585140 146316
rect 578936 146276 578942 146288
rect 585134 146276 585140 146288
rect 585192 146276 585198 146328
rect 668762 145732 668768 145784
rect 668820 145772 668826 145784
rect 670786 145772 670792 145784
rect 668820 145744 670792 145772
rect 668820 145732 668826 145744
rect 670786 145732 670792 145744
rect 670844 145732 670850 145784
rect 584766 144916 584772 144968
rect 584824 144956 584830 144968
rect 589458 144956 589464 144968
rect 584824 144928 589464 144956
rect 584824 144916 584830 144928
rect 589458 144916 589464 144928
rect 589516 144916 589522 144968
rect 579246 144644 579252 144696
rect 579304 144684 579310 144696
rect 584398 144684 584404 144696
rect 579304 144656 584404 144684
rect 579304 144644 579310 144656
rect 584398 144644 584404 144656
rect 584456 144644 584462 144696
rect 585962 143556 585968 143608
rect 586020 143596 586026 143608
rect 589458 143596 589464 143608
rect 586020 143568 589464 143596
rect 586020 143556 586026 143568
rect 589458 143556 589464 143568
rect 589516 143556 589522 143608
rect 579522 143420 579528 143472
rect 579580 143460 579586 143472
rect 583018 143460 583024 143472
rect 579580 143432 583024 143460
rect 579580 143420 579586 143432
rect 583018 143420 583024 143432
rect 583076 143420 583082 143472
rect 587158 142400 587164 142452
rect 587216 142440 587222 142452
rect 589826 142440 589832 142452
rect 587216 142412 589832 142440
rect 587216 142400 587222 142412
rect 589826 142400 589832 142412
rect 589884 142400 589890 142452
rect 580442 140768 580448 140820
rect 580500 140808 580506 140820
rect 589458 140808 589464 140820
rect 580500 140780 589464 140808
rect 580500 140768 580506 140780
rect 589458 140768 589464 140780
rect 589516 140768 589522 140820
rect 578602 140700 578608 140752
rect 578660 140740 578666 140752
rect 580258 140740 580264 140752
rect 578660 140712 580264 140740
rect 578660 140700 578666 140712
rect 580258 140700 580264 140712
rect 580316 140700 580322 140752
rect 583018 139408 583024 139460
rect 583076 139448 583082 139460
rect 589458 139448 589464 139460
rect 583076 139420 589464 139448
rect 583076 139408 583082 139420
rect 589458 139408 589464 139420
rect 589516 139408 589522 139460
rect 578602 139272 578608 139324
rect 578660 139312 578666 139324
rect 589918 139312 589924 139324
rect 578660 139284 589924 139312
rect 578660 139272 578666 139284
rect 589918 139272 589924 139284
rect 589976 139272 589982 139324
rect 579522 138660 579528 138712
rect 579580 138700 579586 138712
rect 588538 138700 588544 138712
rect 579580 138672 588544 138700
rect 579580 138660 579586 138672
rect 588538 138660 588544 138672
rect 588596 138660 588602 138712
rect 579062 137300 579068 137352
rect 579120 137340 579126 137352
rect 584766 137340 584772 137352
rect 579120 137312 584772 137340
rect 579120 137300 579126 137312
rect 584766 137300 584772 137312
rect 584824 137300 584830 137352
rect 584582 136620 584588 136672
rect 584640 136660 584646 136672
rect 589458 136660 589464 136672
rect 584640 136632 589464 136660
rect 584640 136620 584646 136632
rect 589458 136620 589464 136632
rect 589516 136620 589522 136672
rect 580258 134512 580264 134564
rect 580316 134552 580322 134564
rect 589458 134552 589464 134564
rect 580316 134524 589464 134552
rect 580316 134512 580322 134524
rect 589458 134512 589464 134524
rect 589516 134512 589522 134564
rect 675846 133900 675852 133952
rect 675904 133940 675910 133952
rect 676490 133940 676496 133952
rect 675904 133912 676496 133940
rect 675904 133900 675910 133912
rect 676490 133900 676496 133912
rect 676548 133900 676554 133952
rect 667934 133764 667940 133816
rect 667992 133804 667998 133816
rect 669866 133804 669872 133816
rect 667992 133776 669872 133804
rect 667992 133764 667998 133776
rect 669866 133764 669872 133776
rect 669924 133764 669930 133816
rect 585778 132472 585784 132524
rect 585836 132512 585842 132524
rect 589458 132512 589464 132524
rect 585836 132484 589464 132512
rect 585836 132472 585842 132484
rect 589458 132472 589464 132484
rect 589516 132472 589522 132524
rect 581822 131248 581828 131300
rect 581880 131288 581886 131300
rect 589458 131288 589464 131300
rect 581880 131260 589464 131288
rect 581880 131248 581886 131260
rect 589458 131248 589464 131260
rect 589516 131248 589522 131300
rect 578878 131112 578884 131164
rect 578936 131152 578942 131164
rect 585962 131152 585968 131164
rect 578936 131124 585968 131152
rect 578936 131112 578942 131124
rect 585962 131112 585968 131124
rect 586020 131112 586026 131164
rect 668578 130772 668584 130824
rect 668636 130812 668642 130824
rect 670786 130812 670792 130824
rect 668636 130784 670792 130812
rect 668636 130772 668642 130784
rect 670786 130772 670792 130784
rect 670844 130772 670850 130824
rect 668026 129684 668032 129736
rect 668084 129724 668090 129736
rect 670142 129724 670148 129736
rect 668084 129696 670148 129724
rect 668084 129684 668090 129696
rect 670142 129684 670148 129696
rect 670200 129684 670206 129736
rect 583202 129140 583208 129192
rect 583260 129180 583266 129192
rect 590378 129180 590384 129192
rect 583260 129152 590384 129180
rect 583260 129140 583266 129152
rect 590378 129140 590384 129152
rect 590436 129140 590442 129192
rect 579522 129004 579528 129056
rect 579580 129044 579586 129056
rect 587158 129044 587164 129056
rect 579580 129016 587164 129044
rect 579580 129004 579586 129016
rect 587158 129004 587164 129016
rect 587216 129004 587222 129056
rect 579062 126964 579068 127016
rect 579120 127004 579126 127016
rect 589458 127004 589464 127016
rect 579120 126976 589464 127004
rect 579120 126964 579126 126976
rect 589458 126964 589464 126976
rect 589516 126964 589522 127016
rect 578326 125604 578332 125656
rect 578384 125644 578390 125656
rect 580442 125644 580448 125656
rect 578384 125616 580448 125644
rect 578384 125604 578390 125616
rect 580442 125604 580448 125616
rect 580500 125604 580506 125656
rect 675846 125400 675852 125452
rect 675904 125440 675910 125452
rect 676398 125440 676404 125452
rect 675904 125412 676404 125440
rect 675904 125400 675910 125412
rect 676398 125400 676404 125412
rect 676456 125400 676462 125452
rect 580442 124176 580448 124228
rect 580500 124216 580506 124228
rect 589458 124216 589464 124228
rect 580500 124188 589464 124216
rect 580500 124176 580506 124188
rect 589458 124176 589464 124188
rect 589516 124176 589522 124228
rect 578418 123564 578424 123616
rect 578476 123604 578482 123616
rect 583018 123604 583024 123616
rect 578476 123576 583024 123604
rect 578476 123564 578482 123576
rect 583018 123564 583024 123576
rect 583076 123564 583082 123616
rect 584398 122816 584404 122868
rect 584456 122856 584462 122868
rect 589458 122856 589464 122868
rect 584456 122828 589464 122856
rect 584456 122816 584462 122828
rect 589458 122816 589464 122828
rect 589516 122816 589522 122868
rect 578878 122136 578884 122188
rect 578936 122176 578942 122188
rect 584582 122176 584588 122188
rect 578936 122148 584588 122176
rect 578936 122136 578942 122148
rect 584582 122136 584588 122148
rect 584640 122136 584646 122188
rect 580626 122000 580632 122052
rect 580684 122040 580690 122052
rect 589918 122040 589924 122052
rect 580684 122012 589924 122040
rect 580684 122000 580690 122012
rect 589918 122000 589924 122012
rect 589976 122000 589982 122052
rect 587342 118668 587348 118720
rect 587400 118708 587406 118720
rect 590010 118708 590016 118720
rect 587400 118680 590016 118708
rect 587400 118668 587406 118680
rect 590010 118668 590016 118680
rect 590068 118668 590074 118720
rect 675938 118600 675944 118652
rect 675996 118640 676002 118652
rect 679618 118640 679624 118652
rect 675996 118612 679624 118640
rect 675996 118600 676002 118612
rect 679618 118600 679624 118612
rect 679676 118600 679682 118652
rect 578510 118396 578516 118448
rect 578568 118436 578574 118448
rect 580258 118436 580264 118448
rect 578568 118408 580264 118436
rect 578568 118396 578574 118408
rect 580258 118396 580264 118408
rect 580316 118396 580322 118448
rect 579522 116900 579528 116952
rect 579580 116940 579586 116952
rect 583202 116940 583208 116952
rect 579580 116912 583208 116940
rect 579580 116900 579586 116912
rect 583202 116900 583208 116912
rect 583260 116900 583266 116952
rect 668762 116696 668768 116748
rect 668820 116736 668826 116748
rect 670418 116736 670424 116748
rect 668820 116708 670424 116736
rect 668820 116696 668826 116708
rect 670418 116696 670424 116708
rect 670476 116696 670482 116748
rect 586146 115948 586152 116000
rect 586204 115988 586210 116000
rect 589458 115988 589464 116000
rect 586204 115960 589464 115988
rect 586204 115948 586210 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 583202 115200 583208 115252
rect 583260 115240 583266 115252
rect 589642 115240 589648 115252
rect 583260 115212 589648 115240
rect 583260 115200 583266 115212
rect 589642 115200 589648 115212
rect 589700 115200 589706 115252
rect 579246 114452 579252 114504
rect 579304 114492 579310 114504
rect 581638 114492 581644 114504
rect 579304 114464 581644 114492
rect 579304 114452 579310 114464
rect 581638 114452 581644 114464
rect 581696 114452 581702 114504
rect 583018 113160 583024 113212
rect 583076 113200 583082 113212
rect 589458 113200 589464 113212
rect 583076 113172 589464 113200
rect 583076 113160 583082 113172
rect 589458 113160 589464 113172
rect 589516 113160 589522 113212
rect 579522 112820 579528 112872
rect 579580 112860 579586 112872
rect 585778 112860 585784 112872
rect 579580 112832 585784 112860
rect 579580 112820 579586 112832
rect 585778 112820 585784 112832
rect 585836 112820 585842 112872
rect 585962 112412 585968 112464
rect 586020 112452 586026 112464
rect 590102 112452 590108 112464
rect 586020 112424 590108 112452
rect 586020 112412 586026 112424
rect 590102 112412 590108 112424
rect 590160 112412 590166 112464
rect 581638 110440 581644 110492
rect 581696 110480 581702 110492
rect 589458 110480 589464 110492
rect 581696 110452 589464 110480
rect 581696 110440 581702 110452
rect 589458 110440 589464 110452
rect 589516 110440 589522 110492
rect 579338 110100 579344 110152
rect 579396 110140 579402 110152
rect 581822 110140 581828 110152
rect 579396 110112 581828 110140
rect 579396 110100 579402 110112
rect 581822 110100 581828 110112
rect 581880 110100 581886 110152
rect 584582 109012 584588 109064
rect 584640 109052 584646 109064
rect 589274 109052 589280 109064
rect 584640 109024 589280 109052
rect 584640 109012 584646 109024
rect 589274 109012 589280 109024
rect 589332 109012 589338 109064
rect 667934 108808 667940 108860
rect 667992 108848 667998 108860
rect 669958 108848 669964 108860
rect 667992 108820 669964 108848
rect 667992 108808 667998 108820
rect 669958 108808 669964 108820
rect 670016 108808 670022 108860
rect 578326 108672 578332 108724
rect 578384 108712 578390 108724
rect 580626 108712 580632 108724
rect 578384 108684 580632 108712
rect 578384 108672 578390 108684
rect 580626 108672 580632 108684
rect 580684 108672 580690 108724
rect 589458 107692 589464 107704
rect 579632 107664 589464 107692
rect 578878 107584 578884 107636
rect 578936 107624 578942 107636
rect 579632 107624 579660 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 578936 107596 579660 107624
rect 578936 107584 578942 107596
rect 587158 106292 587164 106344
rect 587216 106332 587222 106344
rect 589826 106332 589832 106344
rect 587216 106304 589832 106332
rect 587216 106292 587222 106304
rect 589826 106292 589832 106304
rect 589884 106292 589890 106344
rect 668394 106156 668400 106208
rect 668452 106196 668458 106208
rect 670786 106196 670792 106208
rect 668452 106168 670792 106196
rect 668452 106156 668458 106168
rect 670786 106156 670792 106168
rect 670844 106156 670850 106208
rect 580258 104864 580264 104916
rect 580316 104904 580322 104916
rect 589458 104904 589464 104916
rect 580316 104876 589464 104904
rect 580316 104864 580322 104876
rect 589458 104864 589464 104876
rect 589516 104864 589522 104916
rect 668762 104660 668768 104712
rect 668820 104700 668826 104712
rect 670786 104700 670792 104712
rect 668820 104672 670792 104700
rect 668820 104660 668826 104672
rect 670786 104660 670792 104672
rect 670844 104660 670850 104712
rect 579522 103436 579528 103488
rect 579580 103476 579586 103488
rect 588538 103476 588544 103488
rect 579580 103448 588544 103476
rect 579580 103436 579586 103448
rect 588538 103436 588544 103448
rect 588596 103436 588602 103488
rect 579522 101804 579528 101856
rect 579580 101844 579586 101856
rect 584398 101844 584404 101856
rect 579580 101816 584404 101844
rect 579580 101804 579586 101816
rect 584398 101804 584404 101816
rect 584456 101804 584462 101856
rect 584398 100104 584404 100156
rect 584456 100144 584462 100156
rect 589458 100144 589464 100156
rect 584456 100116 589464 100144
rect 584456 100104 584462 100116
rect 589458 100104 589464 100116
rect 589516 100104 589522 100156
rect 579062 99356 579068 99408
rect 579120 99396 579126 99408
rect 586146 99396 586152 99408
rect 579120 99368 586152 99396
rect 579120 99356 579126 99368
rect 586146 99356 586152 99368
rect 586204 99356 586210 99408
rect 622302 99288 622308 99340
rect 622360 99328 622366 99340
rect 630766 99328 630772 99340
rect 622360 99300 630772 99328
rect 622360 99288 622366 99300
rect 630766 99288 630772 99300
rect 630824 99288 630830 99340
rect 578602 99220 578608 99272
rect 578660 99260 578666 99272
rect 580442 99260 580448 99272
rect 578660 99232 580448 99260
rect 578660 99220 578666 99232
rect 580442 99220 580448 99232
rect 580500 99220 580506 99272
rect 623682 99152 623688 99204
rect 623740 99192 623746 99204
rect 633434 99192 633440 99204
rect 623740 99164 633440 99192
rect 623740 99152 623746 99164
rect 633434 99152 633440 99164
rect 633492 99152 633498 99204
rect 577498 99084 577504 99136
rect 577556 99124 577562 99136
rect 595254 99124 595260 99136
rect 577556 99096 595260 99124
rect 577556 99084 577562 99096
rect 595254 99084 595260 99096
rect 595312 99084 595318 99136
rect 625062 99016 625068 99068
rect 625120 99056 625126 99068
rect 636286 99056 636292 99068
rect 625120 99028 636292 99056
rect 625120 99016 625126 99028
rect 636286 99016 636292 99028
rect 636344 99016 636350 99068
rect 628282 98880 628288 98932
rect 628340 98920 628346 98932
rect 642174 98920 642180 98932
rect 628340 98892 642180 98920
rect 628340 98880 628346 98892
rect 642174 98880 642180 98892
rect 642232 98880 642238 98932
rect 629018 98744 629024 98796
rect 629076 98784 629082 98796
rect 643646 98784 643652 98796
rect 629076 98756 643652 98784
rect 629076 98744 629082 98756
rect 643646 98744 643652 98756
rect 643704 98744 643710 98796
rect 647142 98744 647148 98796
rect 647200 98784 647206 98796
rect 661954 98784 661960 98796
rect 647200 98756 661960 98784
rect 647200 98744 647206 98756
rect 661954 98744 661960 98756
rect 662012 98744 662018 98796
rect 630490 98608 630496 98660
rect 630548 98648 630554 98660
rect 646590 98648 646596 98660
rect 630548 98620 646596 98648
rect 630548 98608 630554 98620
rect 646590 98608 646596 98620
rect 646648 98608 646654 98660
rect 645302 98240 645308 98252
rect 631980 98212 645308 98240
rect 578326 97928 578332 97980
rect 578384 97968 578390 97980
rect 587342 97968 587348 97980
rect 578384 97940 587348 97968
rect 578384 97928 578390 97940
rect 587342 97928 587348 97940
rect 587400 97928 587406 97980
rect 620186 97928 620192 97980
rect 620244 97968 620250 97980
rect 626258 97968 626264 97980
rect 620244 97940 626264 97968
rect 620244 97928 620250 97940
rect 626258 97928 626264 97940
rect 626316 97928 626322 97980
rect 629754 97928 629760 97980
rect 629812 97968 629818 97980
rect 631980 97968 632008 98212
rect 645302 98200 645308 98212
rect 645360 98200 645366 98252
rect 640702 98036 640708 98048
rect 629812 97940 632008 97968
rect 632072 98008 640708 98036
rect 629812 97928 629818 97940
rect 618714 97792 618720 97844
rect 618772 97832 618778 97844
rect 625798 97832 625804 97844
rect 618772 97804 625804 97832
rect 618772 97792 618778 97804
rect 625798 97792 625804 97804
rect 625856 97792 625862 97844
rect 627546 97792 627552 97844
rect 627604 97832 627610 97844
rect 632072 97832 632100 98008
rect 640702 97996 640708 98008
rect 640760 97996 640766 98048
rect 659930 97928 659936 97980
rect 659988 97968 659994 97980
rect 665542 97968 665548 97980
rect 659988 97940 665548 97968
rect 659988 97928 659994 97940
rect 665542 97928 665548 97940
rect 665600 97928 665606 97980
rect 627604 97804 632100 97832
rect 627604 97792 627610 97804
rect 632698 97792 632704 97844
rect 632756 97832 632762 97844
rect 648246 97832 648252 97844
rect 632756 97804 648252 97832
rect 632756 97792 632762 97804
rect 648246 97792 648252 97804
rect 648304 97792 648310 97844
rect 655422 97792 655428 97844
rect 655480 97832 655486 97844
rect 662506 97832 662512 97844
rect 655480 97804 662512 97832
rect 655480 97792 655486 97804
rect 662506 97792 662512 97804
rect 662564 97792 662570 97844
rect 631962 97656 631968 97708
rect 632020 97696 632026 97708
rect 647510 97696 647516 97708
rect 632020 97668 647516 97696
rect 632020 97656 632026 97668
rect 647510 97656 647516 97668
rect 647568 97656 647574 97708
rect 650362 97656 650368 97708
rect 650420 97696 650426 97708
rect 658274 97696 658280 97708
rect 650420 97668 658280 97696
rect 650420 97656 650426 97668
rect 658274 97656 658280 97668
rect 658332 97656 658338 97708
rect 659838 97696 659844 97708
rect 659028 97668 659844 97696
rect 621658 97520 621664 97572
rect 621716 97560 621722 97572
rect 629294 97560 629300 97572
rect 621716 97532 629300 97560
rect 621716 97520 621722 97532
rect 629294 97520 629300 97532
rect 629352 97520 629358 97572
rect 634170 97520 634176 97572
rect 634228 97560 634234 97572
rect 650546 97560 650552 97572
rect 634228 97532 650552 97560
rect 634228 97520 634234 97532
rect 650546 97520 650552 97532
rect 650604 97520 650610 97572
rect 656618 97520 656624 97572
rect 656676 97560 656682 97572
rect 659028 97560 659056 97668
rect 659838 97656 659844 97668
rect 659896 97656 659902 97708
rect 656676 97532 659056 97560
rect 656676 97520 656682 97532
rect 659194 97520 659200 97572
rect 659252 97560 659258 97572
rect 664162 97560 664168 97572
rect 659252 97532 664168 97560
rect 659252 97520 659258 97532
rect 664162 97520 664168 97532
rect 664220 97520 664226 97572
rect 612642 97384 612648 97436
rect 612700 97424 612706 97436
rect 618898 97424 618904 97436
rect 612700 97396 618904 97424
rect 612700 97384 612706 97396
rect 618898 97384 618904 97396
rect 618956 97384 618962 97436
rect 623130 97384 623136 97436
rect 623188 97424 623194 97436
rect 632054 97424 632060 97436
rect 623188 97396 632060 97424
rect 623188 97384 623194 97396
rect 632054 97384 632060 97396
rect 632112 97384 632118 97436
rect 633250 97384 633256 97436
rect 633308 97424 633314 97436
rect 648614 97424 648620 97436
rect 633308 97396 648620 97424
rect 633308 97384 633314 97396
rect 648614 97384 648620 97396
rect 648672 97384 648678 97436
rect 651834 97384 651840 97436
rect 651892 97424 651898 97436
rect 659562 97424 659568 97436
rect 651892 97396 659568 97424
rect 651892 97384 651898 97396
rect 659562 97384 659568 97396
rect 659620 97384 659626 97436
rect 605466 97248 605472 97300
rect 605524 97288 605530 97300
rect 611906 97288 611912 97300
rect 605524 97260 611912 97288
rect 605524 97248 605530 97260
rect 611906 97248 611912 97260
rect 611964 97248 611970 97300
rect 626810 97248 626816 97300
rect 626868 97288 626874 97300
rect 639230 97288 639236 97300
rect 626868 97260 639236 97288
rect 626868 97248 626874 97260
rect 639230 97248 639236 97260
rect 639288 97248 639294 97300
rect 643002 97248 643008 97300
rect 643060 97288 643066 97300
rect 656618 97288 656624 97300
rect 643060 97260 656624 97288
rect 643060 97248 643066 97260
rect 656618 97248 656624 97260
rect 656676 97248 656682 97300
rect 656802 97248 656808 97300
rect 656860 97288 656866 97300
rect 661402 97288 661408 97300
rect 656860 97260 661408 97288
rect 656860 97248 656866 97260
rect 661402 97248 661408 97260
rect 661460 97248 661466 97300
rect 626074 97112 626080 97164
rect 626132 97152 626138 97164
rect 637758 97152 637764 97164
rect 626132 97124 637764 97152
rect 626132 97112 626138 97124
rect 637758 97112 637764 97124
rect 637816 97112 637822 97164
rect 644290 97112 644296 97164
rect 644348 97152 644354 97164
rect 658826 97152 658832 97164
rect 644348 97124 658832 97152
rect 644348 97112 644354 97124
rect 658826 97112 658832 97124
rect 658884 97112 658890 97164
rect 624602 96976 624608 97028
rect 624660 97016 624666 97028
rect 634998 97016 635004 97028
rect 624660 96988 635004 97016
rect 624660 96976 624666 96988
rect 634998 96976 635004 96988
rect 635056 96976 635062 97028
rect 635550 96976 635556 97028
rect 635608 97016 635614 97028
rect 647694 97016 647700 97028
rect 635608 96988 647700 97016
rect 635608 96976 635614 96988
rect 647694 96976 647700 96988
rect 647752 96976 647758 97028
rect 596174 96908 596180 96960
rect 596232 96948 596238 96960
rect 596726 96948 596732 96960
rect 596232 96920 596732 96948
rect 596232 96908 596238 96920
rect 596726 96908 596732 96920
rect 596784 96908 596790 96960
rect 597646 96908 597652 96960
rect 597704 96948 597710 96960
rect 598198 96948 598204 96960
rect 597704 96920 598204 96948
rect 597704 96908 597710 96920
rect 598198 96908 598204 96920
rect 598256 96908 598262 96960
rect 600314 96908 600320 96960
rect 600372 96948 600378 96960
rect 601142 96948 601148 96960
rect 600372 96920 601148 96948
rect 600372 96908 600378 96920
rect 601142 96908 601148 96920
rect 601200 96908 601206 96960
rect 601694 96908 601700 96960
rect 601752 96948 601758 96960
rect 602614 96948 602620 96960
rect 601752 96920 602620 96948
rect 601752 96908 601758 96920
rect 602614 96908 602620 96920
rect 602672 96908 602678 96960
rect 606202 96908 606208 96960
rect 606260 96948 606266 96960
rect 607122 96948 607128 96960
rect 606260 96920 607128 96948
rect 606260 96908 606266 96920
rect 607122 96908 607128 96920
rect 607180 96908 607186 96960
rect 613562 96908 613568 96960
rect 613620 96948 613626 96960
rect 613930 96948 613936 96960
rect 613620 96920 613936 96948
rect 613620 96908 613626 96920
rect 613930 96908 613936 96920
rect 613988 96908 613994 96960
rect 615770 96908 615776 96960
rect 615828 96948 615834 96960
rect 616782 96948 616788 96960
rect 615828 96920 616788 96948
rect 615828 96908 615834 96920
rect 616782 96908 616788 96920
rect 616840 96908 616846 96960
rect 656710 96908 656716 96960
rect 656768 96948 656774 96960
rect 660114 96948 660120 96960
rect 656768 96920 660120 96948
rect 656768 96908 656774 96920
rect 660114 96908 660120 96920
rect 660172 96908 660178 96960
rect 612090 96840 612096 96892
rect 612148 96880 612154 96892
rect 612642 96880 612648 96892
rect 612148 96852 612648 96880
rect 612148 96840 612154 96852
rect 612642 96840 612648 96852
rect 612700 96840 612706 96892
rect 634722 96840 634728 96892
rect 634780 96880 634786 96892
rect 650362 96880 650368 96892
rect 634780 96852 650368 96880
rect 634780 96840 634786 96852
rect 650362 96840 650368 96852
rect 650420 96840 650426 96892
rect 653950 96840 653956 96892
rect 654008 96880 654014 96892
rect 654594 96880 654600 96892
rect 654008 96852 654600 96880
rect 654008 96840 654014 96852
rect 654594 96840 654600 96852
rect 654652 96840 654658 96892
rect 654778 96840 654784 96892
rect 654836 96880 654842 96892
rect 655422 96880 655428 96892
rect 654836 96852 655428 96880
rect 654836 96840 654842 96852
rect 655422 96840 655428 96852
rect 655480 96840 655486 96892
rect 658090 96772 658096 96824
rect 658148 96812 658154 96824
rect 663058 96812 663064 96824
rect 658148 96784 663064 96812
rect 658148 96772 658154 96784
rect 663058 96772 663064 96784
rect 663116 96772 663122 96824
rect 610618 96704 610624 96756
rect 610676 96744 610682 96756
rect 611262 96744 611268 96756
rect 610676 96716 611268 96744
rect 610676 96704 610682 96716
rect 611262 96704 611268 96716
rect 611320 96704 611326 96756
rect 617242 96704 617248 96756
rect 617300 96744 617306 96756
rect 618070 96744 618076 96756
rect 617300 96716 618076 96744
rect 617300 96704 617306 96716
rect 618070 96704 618076 96716
rect 618128 96704 618134 96756
rect 647878 96744 647884 96756
rect 645596 96716 647884 96744
rect 640518 96568 640524 96620
rect 640576 96608 640582 96620
rect 645596 96608 645624 96716
rect 647878 96704 647884 96716
rect 647936 96704 647942 96756
rect 640576 96580 645624 96608
rect 640576 96568 640582 96580
rect 645762 96568 645768 96620
rect 645820 96608 645826 96620
rect 656342 96608 656348 96620
rect 645820 96580 656348 96608
rect 645820 96568 645826 96580
rect 656342 96568 656348 96580
rect 656400 96568 656406 96620
rect 639046 96432 639052 96484
rect 639104 96472 639110 96484
rect 645118 96472 645124 96484
rect 639104 96444 645124 96472
rect 639104 96432 639110 96444
rect 645118 96432 645124 96444
rect 645176 96432 645182 96484
rect 646406 96432 646412 96484
rect 646464 96472 646470 96484
rect 652018 96472 652024 96484
rect 646464 96444 652024 96472
rect 646464 96432 646470 96444
rect 652018 96432 652024 96444
rect 652076 96432 652082 96484
rect 652570 96432 652576 96484
rect 652628 96472 652634 96484
rect 665358 96472 665364 96484
rect 652628 96444 665364 96472
rect 652628 96432 652634 96444
rect 665358 96432 665364 96444
rect 665416 96432 665422 96484
rect 631226 96296 631232 96348
rect 631284 96336 631290 96348
rect 647142 96336 647148 96348
rect 631284 96308 647148 96336
rect 631284 96296 631290 96308
rect 647142 96296 647148 96308
rect 647200 96296 647206 96348
rect 648890 96296 648896 96348
rect 648948 96336 648954 96348
rect 664346 96336 664352 96348
rect 648948 96308 664352 96336
rect 648948 96296 648954 96308
rect 664346 96296 664352 96308
rect 664404 96296 664410 96348
rect 637574 96160 637580 96212
rect 637632 96200 637638 96212
rect 660666 96200 660672 96212
rect 637632 96172 660672 96200
rect 637632 96160 637638 96172
rect 660666 96160 660672 96172
rect 660724 96160 660730 96212
rect 611078 96024 611084 96076
rect 611136 96064 611142 96076
rect 622302 96064 622308 96076
rect 611136 96036 622308 96064
rect 611136 96024 611142 96036
rect 622302 96024 622308 96036
rect 622360 96024 622366 96076
rect 649902 96024 649908 96076
rect 649960 96064 649966 96076
rect 663794 96064 663800 96076
rect 649960 96036 663800 96064
rect 649960 96024 649966 96036
rect 663794 96024 663800 96036
rect 663852 96024 663858 96076
rect 644934 95956 644940 96008
rect 644992 95996 644998 96008
rect 649534 95996 649540 96008
rect 644992 95968 649540 95996
rect 644992 95956 644998 95968
rect 649534 95956 649540 95968
rect 649592 95956 649598 96008
rect 607674 95888 607680 95940
rect 607732 95928 607738 95940
rect 624970 95928 624976 95940
rect 607732 95900 624976 95928
rect 607732 95888 607738 95900
rect 624970 95888 624976 95900
rect 625028 95888 625034 95940
rect 665174 95928 665180 95940
rect 656866 95900 665180 95928
rect 643462 95820 643468 95872
rect 643520 95860 643526 95872
rect 649258 95860 649264 95872
rect 643520 95832 649264 95860
rect 643520 95820 643526 95832
rect 649258 95820 649264 95832
rect 649316 95820 649322 95872
rect 656866 95860 656894 95900
rect 665174 95888 665180 95900
rect 665232 95888 665238 95940
rect 649460 95832 656894 95860
rect 638586 95684 638592 95736
rect 638644 95724 638650 95736
rect 647326 95724 647332 95736
rect 638644 95696 647332 95724
rect 638644 95684 638650 95696
rect 647326 95684 647332 95696
rect 647384 95684 647390 95736
rect 647878 95684 647884 95736
rect 647936 95724 647942 95736
rect 649460 95724 649488 95832
rect 647936 95696 649488 95724
rect 647936 95684 647942 95696
rect 653306 95616 653312 95668
rect 653364 95656 653370 95668
rect 663978 95656 663984 95668
rect 653364 95628 663984 95656
rect 653364 95616 653370 95628
rect 663978 95616 663984 95628
rect 664036 95616 664042 95668
rect 640058 95548 640064 95600
rect 640116 95588 640122 95600
rect 647878 95588 647884 95600
rect 640116 95560 647884 95588
rect 640116 95548 640122 95560
rect 647878 95548 647884 95560
rect 647936 95548 647942 95600
rect 641530 95412 641536 95464
rect 641588 95412 641594 95464
rect 645118 95412 645124 95464
rect 645176 95452 645182 95464
rect 651834 95452 651840 95464
rect 645176 95424 651840 95452
rect 645176 95412 645182 95424
rect 651834 95412 651840 95424
rect 651892 95412 651898 95464
rect 641548 95316 641576 95412
rect 649902 95316 649908 95328
rect 641548 95288 649908 95316
rect 649902 95276 649908 95288
rect 649960 95276 649966 95328
rect 620922 95140 620928 95192
rect 620980 95180 620986 95192
rect 626442 95180 626448 95192
rect 620980 95152 626448 95180
rect 620980 95140 620986 95152
rect 626442 95140 626448 95152
rect 626500 95140 626506 95192
rect 647694 95072 647700 95124
rect 647752 95112 647758 95124
rect 648798 95112 648804 95124
rect 647752 95084 648804 95112
rect 647752 95072 647758 95084
rect 648798 95072 648804 95084
rect 648856 95072 648862 95124
rect 579522 95004 579528 95056
rect 579580 95044 579586 95056
rect 583202 95044 583208 95056
rect 579580 95016 583208 95044
rect 579580 95004 579586 95016
rect 583202 95004 583208 95016
rect 583260 95004 583266 95056
rect 616506 95004 616512 95056
rect 616564 95044 616570 95056
rect 622946 95044 622952 95056
rect 616564 95016 622952 95044
rect 616564 95004 616570 95016
rect 622946 95004 622952 95016
rect 623004 95004 623010 95056
rect 609146 94460 609152 94512
rect 609204 94500 609210 94512
rect 620278 94500 620284 94512
rect 609204 94472 620284 94500
rect 609204 94460 609210 94472
rect 620278 94460 620284 94472
rect 620336 94460 620342 94512
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626442 93820 626448 93832
rect 619600 93792 626448 93820
rect 619600 93780 619606 93792
rect 626442 93780 626448 93792
rect 626500 93780 626506 93832
rect 651282 93508 651288 93560
rect 651340 93548 651346 93560
rect 655422 93548 655428 93560
rect 651340 93520 655428 93548
rect 651340 93508 651346 93520
rect 655422 93508 655428 93520
rect 655480 93508 655486 93560
rect 578510 93440 578516 93492
rect 578568 93480 578574 93492
rect 585962 93480 585968 93492
rect 578568 93452 585968 93480
rect 578568 93440 578574 93452
rect 585962 93440 585968 93452
rect 586020 93440 586026 93492
rect 611262 93100 611268 93152
rect 611320 93140 611326 93152
rect 619266 93140 619272 93152
rect 611320 93112 619272 93140
rect 611320 93100 611326 93112
rect 619266 93100 619272 93112
rect 619324 93100 619330 93152
rect 649534 92964 649540 93016
rect 649592 93004 649598 93016
rect 656158 93004 656164 93016
rect 649592 92976 656164 93004
rect 649592 92964 649598 92976
rect 656158 92964 656164 92976
rect 656216 92964 656222 93016
rect 606938 92828 606944 92880
rect 606996 92868 607002 92880
rect 610066 92868 610072 92880
rect 606996 92840 610072 92868
rect 606996 92828 607002 92840
rect 610066 92828 610072 92840
rect 610124 92828 610130 92880
rect 648614 92488 648620 92540
rect 648672 92528 648678 92540
rect 649994 92528 650000 92540
rect 648672 92500 650000 92528
rect 648672 92488 648678 92500
rect 649994 92488 650000 92500
rect 650052 92488 650058 92540
rect 617886 92420 617892 92472
rect 617944 92460 617950 92472
rect 626442 92460 626448 92472
rect 617944 92432 626448 92460
rect 617944 92420 617950 92432
rect 626442 92420 626448 92432
rect 626500 92420 626506 92472
rect 647326 92352 647332 92404
rect 647384 92392 647390 92404
rect 654318 92392 654324 92404
rect 647384 92364 654324 92392
rect 647384 92352 647390 92364
rect 654318 92352 654324 92364
rect 654376 92352 654382 92404
rect 579338 91060 579344 91112
rect 579396 91100 579402 91112
rect 584582 91100 584588 91112
rect 579396 91072 584588 91100
rect 579396 91060 579402 91072
rect 584582 91060 584588 91072
rect 584640 91060 584646 91112
rect 618070 90992 618076 91044
rect 618128 91032 618134 91044
rect 626442 91032 626448 91044
rect 618128 91004 626448 91032
rect 618128 90992 618134 91004
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 651834 90652 651840 90704
rect 651892 90692 651898 90704
rect 655422 90692 655428 90704
rect 651892 90664 655428 90692
rect 651892 90652 651898 90664
rect 655422 90652 655428 90664
rect 655480 90652 655486 90704
rect 622946 89632 622952 89684
rect 623004 89672 623010 89684
rect 623004 89644 625154 89672
rect 623004 89632 623010 89644
rect 625126 89604 625154 89644
rect 626442 89604 626448 89616
rect 625126 89576 626448 89604
rect 626442 89564 626448 89576
rect 626500 89564 626506 89616
rect 585134 88952 585140 89004
rect 585192 88992 585198 89004
rect 589918 88992 589924 89004
rect 585192 88964 589924 88992
rect 585192 88952 585198 88964
rect 589918 88952 589924 88964
rect 589976 88952 589982 89004
rect 649718 88748 649724 88800
rect 649776 88788 649782 88800
rect 658550 88788 658556 88800
rect 649776 88760 658556 88788
rect 649776 88748 649782 88760
rect 658550 88748 658556 88760
rect 658608 88748 658614 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 664162 88788 664168 88800
rect 662380 88760 664168 88788
rect 662380 88748 662386 88760
rect 664162 88748 664168 88760
rect 664220 88748 664226 88800
rect 656342 88612 656348 88664
rect 656400 88652 656406 88664
rect 657446 88652 657452 88664
rect 656400 88624 657452 88652
rect 656400 88612 656406 88624
rect 657446 88612 657452 88624
rect 657504 88612 657510 88664
rect 610066 88272 610072 88324
rect 610124 88312 610130 88324
rect 626442 88312 626448 88324
rect 610124 88284 626448 88312
rect 610124 88272 610130 88284
rect 626442 88272 626448 88284
rect 626500 88272 626506 88324
rect 655238 88272 655244 88324
rect 655296 88312 655302 88324
rect 658458 88312 658464 88324
rect 655296 88284 658464 88312
rect 655296 88272 655302 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 622302 88136 622308 88188
rect 622360 88176 622366 88188
rect 626258 88176 626264 88188
rect 622360 88148 626264 88176
rect 622360 88136 622366 88148
rect 626258 88136 626264 88148
rect 626316 88136 626322 88188
rect 579522 88068 579528 88120
rect 579580 88108 579586 88120
rect 585134 88108 585140 88120
rect 579580 88080 585140 88108
rect 579580 88068 579586 88080
rect 585134 88068 585140 88080
rect 585192 88068 585198 88120
rect 648430 86980 648436 87032
rect 648488 87020 648494 87032
rect 662506 87020 662512 87032
rect 648488 86992 662512 87020
rect 648488 86980 648494 86992
rect 662506 86980 662512 86992
rect 662564 86980 662570 87032
rect 656710 86844 656716 86896
rect 656768 86884 656774 86896
rect 659562 86884 659568 86896
rect 656768 86856 659568 86884
rect 656768 86844 656774 86856
rect 659562 86844 659568 86856
rect 659620 86844 659626 86896
rect 656158 86708 656164 86760
rect 656216 86748 656222 86760
rect 660666 86748 660672 86760
rect 656216 86720 660672 86748
rect 656216 86708 656222 86720
rect 660666 86708 660672 86720
rect 660724 86708 660730 86760
rect 649258 86572 649264 86624
rect 649316 86612 649322 86624
rect 661402 86612 661408 86624
rect 649316 86584 661408 86612
rect 649316 86572 649322 86584
rect 661402 86572 661408 86584
rect 661460 86572 661466 86624
rect 652018 86436 652024 86488
rect 652076 86476 652082 86488
rect 657170 86476 657176 86488
rect 652076 86448 657176 86476
rect 652076 86436 652082 86448
rect 657170 86436 657176 86448
rect 657228 86436 657234 86488
rect 619266 86300 619272 86352
rect 619324 86340 619330 86352
rect 626442 86340 626448 86352
rect 619324 86312 626448 86340
rect 619324 86300 619330 86312
rect 626442 86300 626448 86312
rect 626500 86300 626506 86352
rect 647878 86164 647884 86216
rect 647936 86204 647942 86216
rect 660114 86204 660120 86216
rect 647936 86176 660120 86204
rect 647936 86164 647942 86176
rect 660114 86164 660120 86176
rect 660172 86164 660178 86216
rect 609882 85484 609888 85536
rect 609940 85524 609946 85536
rect 626442 85524 626448 85536
rect 609940 85496 626448 85524
rect 609940 85484 609946 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 620278 85348 620284 85400
rect 620336 85388 620342 85400
rect 625246 85388 625252 85400
rect 620336 85360 625252 85388
rect 620336 85348 620342 85360
rect 625246 85348 625252 85360
rect 625304 85348 625310 85400
rect 579154 84124 579160 84176
rect 579212 84164 579218 84176
rect 581638 84164 581644 84176
rect 579212 84136 581644 84164
rect 579212 84124 579218 84136
rect 581638 84124 581644 84136
rect 581696 84124 581702 84176
rect 608502 84124 608508 84176
rect 608560 84164 608566 84176
rect 625798 84164 625804 84176
rect 608560 84136 625804 84164
rect 608560 84124 608566 84136
rect 625798 84124 625804 84136
rect 625856 84124 625862 84176
rect 579062 82356 579068 82408
rect 579120 82396 579126 82408
rect 583018 82396 583024 82408
rect 579120 82368 583024 82396
rect 579120 82356 579126 82368
rect 583018 82356 583024 82368
rect 583076 82356 583082 82408
rect 579522 82084 579528 82136
rect 579580 82124 579586 82136
rect 587158 82124 587164 82136
rect 579580 82096 587164 82124
rect 579580 82084 579586 82096
rect 587158 82084 587164 82096
rect 587216 82084 587222 82136
rect 628742 80928 628748 80980
rect 628800 80968 628806 80980
rect 642450 80968 642456 80980
rect 628800 80940 642456 80968
rect 628800 80928 628806 80940
rect 642450 80928 642456 80940
rect 642508 80928 642514 80980
rect 612642 80792 612648 80844
rect 612700 80832 612706 80844
rect 647418 80832 647424 80844
rect 612700 80804 647424 80832
rect 612700 80792 612706 80804
rect 647418 80792 647424 80804
rect 647476 80792 647482 80844
rect 595438 80656 595444 80708
rect 595496 80696 595502 80708
rect 636746 80696 636752 80708
rect 595496 80668 636752 80696
rect 595496 80656 595502 80668
rect 636746 80656 636752 80668
rect 636804 80656 636810 80708
rect 629202 79976 629208 80028
rect 629260 80016 629266 80028
rect 633434 80016 633440 80028
rect 629260 79988 633440 80016
rect 629260 79976 629266 79988
rect 633434 79976 633440 79988
rect 633492 79976 633498 80028
rect 613746 79432 613752 79484
rect 613804 79472 613810 79484
rect 646038 79472 646044 79484
rect 613804 79444 646044 79472
rect 613804 79432 613810 79444
rect 646038 79432 646044 79444
rect 646096 79432 646102 79484
rect 579062 79296 579068 79348
rect 579120 79336 579126 79348
rect 588722 79336 588728 79348
rect 579120 79308 588728 79336
rect 579120 79296 579126 79308
rect 588722 79296 588728 79308
rect 588780 79296 588786 79348
rect 613930 79296 613936 79348
rect 613988 79336 613994 79348
rect 646498 79336 646504 79348
rect 613988 79308 646504 79336
rect 613988 79296 613994 79308
rect 646498 79296 646504 79308
rect 646556 79296 646562 79348
rect 633434 78072 633440 78124
rect 633492 78112 633498 78124
rect 645302 78112 645308 78124
rect 633492 78084 645308 78112
rect 633492 78072 633498 78084
rect 645302 78072 645308 78084
rect 645360 78072 645366 78124
rect 631042 77936 631048 77988
rect 631100 77976 631106 77988
rect 643094 77976 643100 77988
rect 631100 77948 643100 77976
rect 631100 77936 631106 77948
rect 643094 77936 643100 77948
rect 643152 77936 643158 77988
rect 628466 77732 628472 77784
rect 628524 77772 628530 77784
rect 632790 77772 632796 77784
rect 628524 77744 632796 77772
rect 628524 77732 628530 77744
rect 632790 77732 632796 77744
rect 632848 77732 632854 77784
rect 625798 77256 625804 77308
rect 625856 77296 625862 77308
rect 631042 77296 631048 77308
rect 625856 77268 631048 77296
rect 625856 77256 625862 77268
rect 631042 77256 631048 77268
rect 631100 77256 631106 77308
rect 616782 76644 616788 76696
rect 616840 76684 616846 76696
rect 646682 76684 646688 76696
rect 616840 76656 646688 76684
rect 616840 76644 616846 76656
rect 646682 76644 646688 76656
rect 646740 76644 646746 76696
rect 611998 76508 612004 76560
rect 612056 76548 612062 76560
rect 662414 76548 662420 76560
rect 612056 76520 662420 76548
rect 612056 76508 612062 76520
rect 662414 76508 662420 76520
rect 662472 76508 662478 76560
rect 578234 75828 578240 75880
rect 578292 75868 578298 75880
rect 580258 75868 580264 75880
rect 578292 75840 580264 75868
rect 578292 75828 578298 75840
rect 580258 75828 580264 75840
rect 580316 75828 580322 75880
rect 618898 75420 618904 75472
rect 618956 75460 618962 75472
rect 648614 75460 648620 75472
rect 618956 75432 648620 75460
rect 618956 75420 618962 75432
rect 648614 75420 648620 75432
rect 648672 75420 648678 75472
rect 615402 75284 615408 75336
rect 615460 75324 615466 75336
rect 646866 75324 646872 75336
rect 615460 75296 646872 75324
rect 615460 75284 615466 75296
rect 646866 75284 646872 75296
rect 646924 75284 646930 75336
rect 607122 75148 607128 75200
rect 607180 75188 607186 75200
rect 646222 75188 646228 75200
rect 607180 75160 646228 75188
rect 607180 75148 607186 75160
rect 646222 75148 646228 75160
rect 646280 75148 646286 75200
rect 578878 72428 578884 72480
rect 578936 72468 578942 72480
rect 601878 72468 601884 72480
rect 578936 72440 601884 72468
rect 578936 72428 578942 72440
rect 601878 72428 601884 72440
rect 601936 72428 601942 72480
rect 579062 71340 579068 71392
rect 579120 71380 579126 71392
rect 584398 71380 584404 71392
rect 579120 71352 584404 71380
rect 579120 71340 579126 71352
rect 584398 71340 584404 71352
rect 584456 71340 584462 71392
rect 580258 68280 580264 68332
rect 580316 68320 580322 68332
rect 604454 68320 604460 68332
rect 580316 68292 604460 68320
rect 580316 68280 580322 68292
rect 604454 68280 604460 68292
rect 604512 68280 604518 68332
rect 577498 59984 577504 60036
rect 577556 60024 577562 60036
rect 603074 60024 603080 60036
rect 577556 59996 603080 60024
rect 577556 59984 577562 59996
rect 603074 59984 603080 59996
rect 603132 59984 603138 60036
rect 576118 58624 576124 58676
rect 576176 58664 576182 58676
rect 601694 58664 601700 58676
rect 576176 58636 601700 58664
rect 576176 58624 576182 58636
rect 601694 58624 601700 58636
rect 601752 58624 601758 58676
rect 574922 57196 574928 57248
rect 574980 57236 574986 57248
rect 600314 57236 600320 57248
rect 574980 57208 600320 57236
rect 574980 57196 574986 57208
rect 600314 57196 600320 57208
rect 600372 57196 600378 57248
rect 574554 55972 574560 56024
rect 574612 56012 574618 56024
rect 599118 56012 599124 56024
rect 574612 55984 599124 56012
rect 574612 55972 574618 55984
rect 599118 55972 599124 55984
rect 599176 55972 599182 56024
rect 574738 55836 574744 55888
rect 574796 55876 574802 55888
rect 600498 55876 600504 55888
rect 574796 55848 600504 55876
rect 574796 55836 574802 55848
rect 600498 55836 600504 55848
rect 600556 55836 600562 55888
rect 462976 55576 478874 55604
rect 462976 53644 463004 55576
rect 463298 55236 469214 55264
rect 463298 53644 463326 55236
rect 469186 55060 469214 55236
rect 478846 55196 478874 55576
rect 596450 55196 596456 55208
rect 478846 55168 596456 55196
rect 596450 55156 596456 55168
rect 596508 55156 596514 55208
rect 597830 55060 597836 55072
rect 469186 55032 597836 55060
rect 597830 55020 597836 55032
rect 597888 55020 597894 55072
rect 597646 54924 597652 54936
rect 469186 54896 597652 54924
rect 469186 54720 469214 54896
rect 597646 54884 597652 54896
rect 597704 54884 597710 54936
rect 598934 54788 598940 54800
rect 463528 54692 469214 54720
rect 474016 54760 598940 54788
rect 463528 53644 463556 54692
rect 474016 54584 474044 54760
rect 598934 54748 598940 54760
rect 598992 54748 598998 54800
rect 624418 54652 624424 54664
rect 463712 54556 474044 54584
rect 476500 54624 624424 54652
rect 463712 53644 463740 54556
rect 464448 54420 476252 54448
rect 464448 53644 464476 54420
rect 476224 53644 476252 54420
rect 476500 53768 476528 54624
rect 624418 54612 624424 54624
rect 624476 54612 624482 54664
rect 625798 54516 625804 54528
rect 476408 53740 476528 53768
rect 476592 54488 625804 54516
rect 476408 53644 476436 53740
rect 476592 53644 476620 54488
rect 625798 54476 625804 54488
rect 625856 54476 625862 54528
rect 596174 54380 596180 54392
rect 477052 54352 596180 54380
rect 477052 53644 477080 54352
rect 596174 54340 596180 54352
rect 596232 54340 596238 54392
rect 581638 54244 581644 54256
rect 479628 54216 581644 54244
rect 479628 53972 479656 54216
rect 581638 54204 581644 54216
rect 581696 54204 581702 54256
rect 574738 54108 574744 54120
rect 479260 53944 479656 53972
rect 480226 54080 574744 54108
rect 479260 53768 479288 53944
rect 480226 53768 480254 54080
rect 574738 54068 574744 54080
rect 574796 54068 574802 54120
rect 574554 53972 574560 53984
rect 479076 53740 479288 53768
rect 479444 53740 480254 53768
rect 481606 53944 574560 53972
rect 479076 53644 479104 53740
rect 479444 53644 479472 53740
rect 462958 53592 462964 53644
rect 463016 53592 463022 53644
rect 463234 53592 463240 53644
rect 463292 53604 463326 53644
rect 463292 53592 463298 53604
rect 463510 53592 463516 53644
rect 463568 53592 463574 53644
rect 463694 53592 463700 53644
rect 463752 53592 463758 53644
rect 464430 53592 464436 53644
rect 464488 53592 464494 53644
rect 464706 53592 464712 53644
rect 464764 53632 464770 53644
rect 476022 53632 476028 53644
rect 464764 53604 476028 53632
rect 464764 53592 464770 53604
rect 476022 53592 476028 53604
rect 476080 53592 476086 53644
rect 476206 53592 476212 53644
rect 476264 53592 476270 53644
rect 476390 53592 476396 53644
rect 476448 53592 476454 53644
rect 476574 53592 476580 53644
rect 476632 53592 476638 53644
rect 477034 53592 477040 53644
rect 477092 53592 477098 53644
rect 479058 53592 479064 53644
rect 479116 53592 479122 53644
rect 479426 53592 479432 53644
rect 479484 53592 479490 53644
rect 481606 53632 481634 53944
rect 574554 53932 574560 53944
rect 574612 53932 574618 53984
rect 574922 53836 574928 53848
rect 480226 53604 481634 53632
rect 482986 53808 574928 53836
rect 479610 53524 479616 53576
rect 479668 53564 479674 53576
rect 480226 53564 480254 53604
rect 479668 53536 480254 53564
rect 479668 53524 479674 53536
rect 462222 53456 462228 53508
rect 462280 53496 462286 53508
rect 479426 53496 479432 53508
rect 462280 53468 479432 53496
rect 462280 53456 462286 53468
rect 479426 53456 479432 53468
rect 479484 53456 479490 53508
rect 463142 53320 463148 53372
rect 463200 53360 463206 53372
rect 482986 53360 483014 53808
rect 574922 53796 574928 53808
rect 574980 53796 574986 53848
rect 463200 53332 483014 53360
rect 463200 53320 463206 53332
rect 48958 53184 48964 53236
rect 49016 53224 49022 53236
rect 130378 53224 130384 53236
rect 49016 53196 130384 53224
rect 49016 53184 49022 53196
rect 130378 53184 130384 53196
rect 130436 53184 130442 53236
rect 461302 53184 461308 53236
rect 461360 53224 461366 53236
rect 479610 53224 479616 53236
rect 461360 53196 479616 53224
rect 461360 53184 461366 53196
rect 479610 53184 479616 53196
rect 479668 53184 479674 53236
rect 312354 53116 312360 53168
rect 312412 53156 312418 53168
rect 313734 53156 313740 53168
rect 312412 53128 313740 53156
rect 312412 53116 312418 53128
rect 313734 53116 313740 53128
rect 313792 53116 313798 53168
rect 316310 53116 316316 53168
rect 316368 53156 316374 53168
rect 317690 53156 317696 53168
rect 316368 53128 317696 53156
rect 316368 53116 316374 53128
rect 317690 53116 317696 53128
rect 317748 53116 317754 53168
rect 45462 53048 45468 53100
rect 45520 53088 45526 53100
rect 128998 53088 129004 53100
rect 45520 53060 129004 53088
rect 45520 53048 45526 53060
rect 128998 53048 129004 53060
rect 129056 53048 129062 53100
rect 459462 53048 459468 53100
rect 459520 53088 459526 53100
rect 463694 53088 463700 53100
rect 459520 53060 463700 53088
rect 459520 53048 459526 53060
rect 463694 53048 463700 53060
rect 463752 53048 463758 53100
rect 465442 53048 465448 53100
rect 465500 53088 465506 53100
rect 479058 53088 479064 53100
rect 465500 53060 479064 53088
rect 465500 53048 465506 53060
rect 479058 53048 479064 53060
rect 479116 53048 479122 53100
rect 462958 52912 462964 52964
rect 463016 52952 463022 52964
rect 464522 52952 464528 52964
rect 463016 52924 464528 52952
rect 463016 52912 463022 52924
rect 464522 52912 464528 52924
rect 464580 52912 464586 52964
rect 460060 52776 460066 52828
rect 460118 52816 460124 52828
rect 464706 52816 464712 52828
rect 460118 52788 464712 52816
rect 460118 52776 460124 52788
rect 464706 52776 464712 52788
rect 464764 52776 464770 52828
rect 465580 52776 465586 52828
rect 465638 52816 465644 52828
rect 476390 52816 476396 52828
rect 465638 52788 476396 52816
rect 465638 52776 465644 52788
rect 476390 52776 476396 52788
rect 476448 52776 476454 52828
rect 47578 51960 47584 52012
rect 47636 52000 47642 52012
rect 130562 52000 130568 52012
rect 47636 51972 130568 52000
rect 47636 51960 47642 51972
rect 130562 51960 130568 51972
rect 130620 51960 130626 52012
rect 50338 51824 50344 51876
rect 50396 51864 50402 51876
rect 129182 51864 129188 51876
rect 50396 51836 129188 51864
rect 50396 51824 50402 51836
rect 129182 51824 129188 51836
rect 129240 51824 129246 51876
rect 129550 51824 129556 51876
rect 129608 51864 129614 51876
rect 591298 51864 591304 51876
rect 129608 51836 591304 51864
rect 129608 51824 129614 51836
rect 591298 51824 591304 51836
rect 591356 51824 591362 51876
rect 128814 51688 128820 51740
rect 128872 51728 128878 51740
rect 592678 51728 592684 51740
rect 128872 51700 592684 51728
rect 128872 51688 128878 51700
rect 592678 51688 592684 51700
rect 592736 51688 592742 51740
rect 318334 50464 318340 50516
rect 318392 50504 318398 50516
rect 458174 50504 458180 50516
rect 318392 50476 458180 50504
rect 318392 50464 318398 50476
rect 458174 50464 458180 50476
rect 458232 50464 458238 50516
rect 47762 50328 47768 50380
rect 47820 50368 47826 50380
rect 130838 50368 130844 50380
rect 47820 50340 130844 50368
rect 47820 50328 47826 50340
rect 130838 50328 130844 50340
rect 130896 50328 130902 50380
rect 314010 50328 314016 50380
rect 314068 50368 314074 50380
rect 458358 50368 458364 50380
rect 314068 50340 458364 50368
rect 314068 50328 314074 50340
rect 458358 50328 458364 50340
rect 458416 50328 458422 50380
rect 522942 50328 522948 50380
rect 523000 50368 523006 50380
rect 544010 50368 544016 50380
rect 523000 50340 544016 50368
rect 523000 50328 523006 50340
rect 544010 50328 544016 50340
rect 544068 50328 544074 50380
rect 49142 49104 49148 49156
rect 49200 49144 49206 49156
rect 129366 49144 129372 49156
rect 49200 49116 129372 49144
rect 49200 49104 49206 49116
rect 129366 49104 129372 49116
rect 129424 49104 129430 49156
rect 46198 48968 46204 49020
rect 46256 49008 46262 49020
rect 131022 49008 131028 49020
rect 46256 48980 131028 49008
rect 46256 48968 46262 48980
rect 131022 48968 131028 48980
rect 131080 48968 131086 49020
rect 130562 46044 130568 46096
rect 130620 46084 130626 46096
rect 132862 46084 132868 46096
rect 130620 46056 132868 46084
rect 130620 46044 130626 46056
rect 132862 46044 132868 46056
rect 132920 46044 132926 46096
rect 130378 45908 130384 45960
rect 130436 45948 130442 45960
rect 132586 45948 132592 45960
rect 130436 45920 132592 45948
rect 130436 45908 130442 45920
rect 132586 45908 132592 45920
rect 132644 45908 132650 45960
rect 128998 45364 129004 45416
rect 129056 45404 129062 45416
rect 129056 45376 131390 45404
rect 129056 45364 129062 45376
rect 131362 45090 131390 45376
rect 129550 45024 129556 45076
rect 129608 45064 129614 45076
rect 129608 45036 131068 45064
rect 129608 45024 129614 45036
rect 131040 45020 131068 45036
rect 131040 44992 131330 45020
rect 129366 44888 129372 44940
rect 129424 44928 129430 44940
rect 129424 44900 131620 44928
rect 129424 44888 129430 44900
rect 131684 44824 131790 44852
rect 128814 44752 128820 44804
rect 128872 44792 128878 44804
rect 131684 44792 131712 44824
rect 128872 44764 131712 44792
rect 128872 44752 128878 44764
rect 131776 44740 131974 44768
rect 131574 44644 131580 44696
rect 131632 44684 131638 44696
rect 131776 44684 131804 44740
rect 131632 44656 131804 44684
rect 132144 44656 132172 44670
rect 131632 44644 131638 44656
rect 131868 44628 132172 44656
rect 129182 44548 129188 44600
rect 129240 44588 129246 44600
rect 131868 44588 131896 44628
rect 129240 44560 131896 44588
rect 132236 44560 132402 44588
rect 129240 44548 129246 44560
rect 132236 44520 132264 44560
rect 132144 44492 132264 44520
rect 50522 44276 50528 44328
rect 50580 44316 50586 44328
rect 131574 44316 131580 44328
rect 50580 44288 131580 44316
rect 50580 44276 50586 44288
rect 131574 44276 131580 44288
rect 131632 44276 131638 44328
rect 43438 44140 43444 44192
rect 43496 44180 43502 44192
rect 132144 44180 132172 44492
rect 132604 44396 132632 44502
rect 132586 44344 132592 44396
rect 132644 44344 132650 44396
rect 132862 44364 132868 44416
rect 132920 44364 132926 44416
rect 132770 44252 132776 44304
rect 132828 44292 132834 44304
rect 132828 44264 132986 44292
rect 132828 44252 132834 44264
rect 43496 44152 132172 44180
rect 132466 44152 133170 44180
rect 43496 44140 43502 44152
rect 131022 44004 131028 44056
rect 131080 44044 131086 44056
rect 132466 44044 132494 44152
rect 131080 44016 132494 44044
rect 131080 44004 131086 44016
rect 440234 43800 440240 43852
rect 440292 43840 440298 43852
rect 441062 43840 441068 43852
rect 440292 43812 441068 43840
rect 440292 43800 440298 43812
rect 441062 43800 441068 43812
rect 441120 43800 441126 43852
rect 187326 42780 187332 42832
rect 187384 42820 187390 42832
rect 255866 42820 255872 42832
rect 187384 42792 255872 42820
rect 187384 42780 187390 42792
rect 255866 42780 255872 42792
rect 255924 42780 255930 42832
rect 307294 42712 307300 42764
rect 307352 42752 307358 42764
rect 431218 42752 431224 42764
rect 307352 42724 431224 42752
rect 307352 42712 307358 42724
rect 431218 42712 431224 42724
rect 431276 42712 431282 42764
rect 441062 42712 441068 42764
rect 441120 42752 441126 42764
rect 449158 42752 449164 42764
rect 441120 42724 449164 42752
rect 441120 42712 441126 42724
rect 449158 42712 449164 42724
rect 449216 42712 449222 42764
rect 453574 42712 453580 42764
rect 453632 42752 453638 42764
rect 464154 42752 464160 42764
rect 453632 42724 464160 42752
rect 453632 42712 453638 42724
rect 464154 42712 464160 42724
rect 464212 42712 464218 42764
rect 310422 42576 310428 42628
rect 310480 42616 310486 42628
rect 427078 42616 427084 42628
rect 310480 42588 427084 42616
rect 310480 42576 310486 42588
rect 427078 42576 427084 42588
rect 427136 42576 427142 42628
rect 441246 42576 441252 42628
rect 441304 42616 441310 42628
rect 446398 42616 446404 42628
rect 441304 42588 446404 42616
rect 441304 42576 441310 42588
rect 446398 42576 446404 42588
rect 446456 42576 446462 42628
rect 454494 42440 454500 42492
rect 454552 42480 454558 42492
rect 463050 42480 463056 42492
rect 454552 42452 463056 42480
rect 454552 42440 454558 42452
rect 463050 42440 463056 42452
rect 463108 42440 463114 42492
rect 404446 42304 404452 42356
rect 404504 42344 404510 42356
rect 405182 42344 405188 42356
rect 404504 42316 405188 42344
rect 404504 42304 404510 42316
rect 405182 42304 405188 42316
rect 405240 42304 405246 42356
rect 420730 42304 420736 42356
rect 420788 42344 420794 42356
rect 426894 42344 426900 42356
rect 420788 42316 426900 42344
rect 420788 42304 420794 42316
rect 426894 42304 426900 42316
rect 426952 42304 426958 42356
rect 661402 42129 661408 42181
rect 661460 42129 661466 42181
rect 427078 41964 427084 42016
rect 427136 42004 427142 42016
rect 427136 41976 427814 42004
rect 427136 41964 427142 41976
rect 427786 41868 427814 41976
rect 431218 41964 431224 42016
rect 431276 42004 431282 42016
rect 441062 42004 441068 42016
rect 431276 41976 441068 42004
rect 431276 41964 431282 41976
rect 441062 41964 441068 41976
rect 441120 41964 441126 42016
rect 446398 41964 446404 42016
rect 446456 42004 446462 42016
rect 454494 42004 454500 42016
rect 446456 41976 454500 42004
rect 446456 41964 446462 41976
rect 454494 41964 454500 41976
rect 454552 41964 454558 42016
rect 441246 41868 441252 41880
rect 427786 41840 441252 41868
rect 441246 41828 441252 41840
rect 441304 41828 441310 41880
rect 449158 41828 449164 41880
rect 449216 41868 449222 41880
rect 453574 41868 453580 41880
rect 449216 41840 453580 41868
rect 449216 41828 449222 41840
rect 453574 41828 453580 41840
rect 453632 41828 453638 41880
rect 404446 41420 404452 41472
rect 404504 41460 404510 41472
rect 420730 41460 420736 41472
rect 404504 41432 420736 41460
rect 404504 41420 404510 41432
rect 420730 41420 420736 41432
rect 420788 41420 420794 41472
rect 426894 41420 426900 41472
rect 426952 41460 426958 41472
rect 459186 41460 459192 41472
rect 426952 41432 459192 41460
rect 426952 41420 426958 41432
rect 459186 41420 459192 41432
rect 459244 41420 459250 41472
<< via1 >>
rect 132500 1001920 132552 1001972
rect 133696 1001920 133748 1001972
rect 401692 992196 401744 992248
rect 404360 992196 404412 992248
rect 396080 990836 396132 990888
rect 400220 990836 400272 990888
rect 242256 989068 242308 989120
rect 245660 989068 245712 989120
rect 293960 988184 294012 988236
rect 298100 988184 298152 988236
rect 389180 987504 389232 987556
rect 391940 987504 391992 987556
rect 399760 986348 399812 986400
rect 401692 986348 401744 986400
rect 238668 985940 238720 985992
rect 242256 985940 242308 985992
rect 289728 985396 289780 985448
rect 293960 985396 294012 985448
rect 394424 983492 394476 983544
rect 396080 983492 396132 983544
rect 483020 982472 483072 982524
rect 483848 982472 483900 982524
rect 651380 959080 651432 959132
rect 677416 959080 677468 959132
rect 30104 954932 30156 954984
rect 63408 954932 63460 954984
rect 656164 896996 656216 897048
rect 676036 897064 676088 897116
rect 672724 895772 672776 895824
rect 676036 895772 676088 895824
rect 654784 895636 654836 895688
rect 675852 895636 675904 895688
rect 671896 894412 671948 894464
rect 676036 894412 676088 894464
rect 671068 894276 671120 894328
rect 675852 894276 675904 894328
rect 673276 892984 673328 893036
rect 675852 892984 675904 893036
rect 672264 892848 672316 892900
rect 676036 892848 676088 892900
rect 674840 890332 674892 890384
rect 676036 890332 676088 890384
rect 676220 890128 676272 890180
rect 676864 890128 676916 890180
rect 674380 888904 674432 888956
rect 676036 888904 676088 888956
rect 675024 888700 675076 888752
rect 675852 888700 675904 888752
rect 676220 888700 676272 888752
rect 677048 888700 677100 888752
rect 674656 888496 674708 888548
rect 676036 888496 676088 888548
rect 674196 887272 674248 887324
rect 676036 887272 676088 887324
rect 670884 886864 670936 886916
rect 676036 886864 676088 886916
rect 675576 886592 675628 886644
rect 676404 886592 676456 886644
rect 653404 880472 653456 880524
rect 667296 880472 667348 880524
rect 675392 880336 675444 880388
rect 679624 880404 679676 880456
rect 667296 879588 667348 879640
rect 675576 879588 675628 879640
rect 675760 879316 675812 879368
rect 676864 879316 676916 879368
rect 675944 879180 675996 879232
rect 678244 879180 678296 879232
rect 674012 878976 674064 879028
rect 677048 879044 677100 879096
rect 675760 878364 675812 878416
rect 675484 877208 675536 877260
rect 674840 874896 674892 874948
rect 675392 874896 675444 874948
rect 674012 873672 674064 873724
rect 675392 873672 675444 873724
rect 674196 871972 674248 872024
rect 674656 871972 674708 872024
rect 657544 869388 657596 869440
rect 674656 869388 674708 869440
rect 651472 868844 651524 868896
rect 654784 868844 654836 868896
rect 654140 868028 654192 868080
rect 674840 868028 674892 868080
rect 651472 867892 651524 867944
rect 656164 867892 656216 867944
rect 674656 867892 674708 867944
rect 675208 867892 675260 867944
rect 651472 866600 651524 866652
rect 672724 866600 672776 866652
rect 651380 865172 651432 865224
rect 653404 865172 653456 865224
rect 651472 863812 651524 863864
rect 657544 863812 657596 863864
rect 651472 862452 651524 862504
rect 654140 862452 654192 862504
rect 35808 816960 35860 817012
rect 58624 816960 58676 817012
rect 35808 815736 35860 815788
rect 43444 815736 43496 815788
rect 35624 815600 35676 815652
rect 61384 815600 61436 815652
rect 35440 814852 35492 814904
rect 62764 814852 62816 814904
rect 35624 814376 35676 814428
rect 42892 814376 42944 814428
rect 35808 814240 35860 814292
rect 44732 814240 44784 814292
rect 41328 812812 41380 812864
rect 44180 812812 44232 812864
rect 41328 811724 41380 811776
rect 43076 811724 43128 811776
rect 40960 810704 41012 810756
rect 42616 810704 42668 810756
rect 41328 808596 41380 808648
rect 42248 808596 42300 808648
rect 41328 807440 41380 807492
rect 43260 807440 43312 807492
rect 41144 807304 41196 807356
rect 44364 807304 44416 807356
rect 41328 806080 41380 806132
rect 50344 806080 50396 806132
rect 41144 805944 41196 805996
rect 64144 805944 64196 805996
rect 34520 802408 34572 802460
rect 42156 802408 42208 802460
rect 37924 801728 37976 801780
rect 41972 801728 42024 801780
rect 36544 801252 36596 801304
rect 42616 801252 42668 801304
rect 41972 801116 42024 801168
rect 42708 801116 42760 801168
rect 31024 801048 31076 801100
rect 42800 800980 42852 801032
rect 43628 799076 43680 799128
rect 53104 799076 53156 799128
rect 43812 797648 43864 797700
rect 62948 797648 63000 797700
rect 42248 795608 42300 795660
rect 43812 795608 43864 795660
rect 44364 794860 44416 794912
rect 42340 794316 42392 794368
rect 653404 790780 653456 790832
rect 675392 790780 675444 790832
rect 53104 790712 53156 790764
rect 62212 790712 62264 790764
rect 42156 790100 42208 790152
rect 42708 790100 42760 790152
rect 61384 788604 61436 788656
rect 62948 788604 63000 788656
rect 42616 787992 42668 788044
rect 43076 787992 43128 788044
rect 42708 786632 42760 786684
rect 62120 786632 62172 786684
rect 58624 786496 58676 786548
rect 62120 786496 62172 786548
rect 670608 784252 670660 784304
rect 675116 784252 675168 784304
rect 669228 784116 669280 784168
rect 675392 784116 675444 784168
rect 673920 782620 673972 782672
rect 675116 782620 675168 782672
rect 669044 782484 669096 782536
rect 675300 782484 675352 782536
rect 655520 781056 655572 781108
rect 675208 781056 675260 781108
rect 655060 778336 655112 778388
rect 674932 778336 674984 778388
rect 651472 777588 651524 777640
rect 660304 777588 660356 777640
rect 670424 776976 670476 777028
rect 675300 776976 675352 777028
rect 672724 775616 672776 775668
rect 674932 775616 674984 775668
rect 651472 775548 651524 775600
rect 669964 775548 670016 775600
rect 651380 775276 651432 775328
rect 653404 775276 653456 775328
rect 35808 774188 35860 774240
rect 41696 774188 41748 774240
rect 42064 774188 42116 774240
rect 58624 774188 58676 774240
rect 651472 774120 651524 774172
rect 655520 774120 655572 774172
rect 651472 773780 651524 773832
rect 655060 773780 655112 773832
rect 671436 773372 671488 773424
rect 675300 773372 675352 773424
rect 35808 773304 35860 773356
rect 40316 773304 40368 773356
rect 35808 773100 35860 773152
rect 39580 773100 39632 773152
rect 35624 772964 35676 773016
rect 41696 772964 41748 773016
rect 42064 772964 42116 773016
rect 44548 772964 44600 773016
rect 35440 772828 35492 772880
rect 41696 772828 41748 772880
rect 42064 772828 42116 772880
rect 61384 772828 61436 772880
rect 35624 771808 35676 771860
rect 40776 771808 40828 771860
rect 35808 771536 35860 771588
rect 41696 771604 41748 771656
rect 42064 771604 42116 771656
rect 44732 771604 44784 771656
rect 35440 771400 35492 771452
rect 41696 771400 41748 771452
rect 42064 771400 42116 771452
rect 44364 771400 44416 771452
rect 35808 770448 35860 770500
rect 40500 770448 40552 770500
rect 35440 770176 35492 770228
rect 39948 770244 40000 770296
rect 35624 770040 35676 770092
rect 41696 770040 41748 770092
rect 42064 770040 42116 770092
rect 44180 770040 44232 770092
rect 652024 768884 652076 768936
rect 656164 768884 656216 768936
rect 35624 768816 35676 768868
rect 41696 768816 41748 768868
rect 35808 768680 35860 768732
rect 40040 768680 40092 768732
rect 35808 767592 35860 767644
rect 36544 767592 36596 767644
rect 35808 765892 35860 765944
rect 39764 765892 39816 765944
rect 40040 765280 40092 765332
rect 41696 765280 41748 765332
rect 42064 765144 42116 765196
rect 42524 765144 42576 765196
rect 35808 764804 35860 764856
rect 39212 764804 39264 764856
rect 35808 764532 35860 764584
rect 39764 764532 39816 764584
rect 35624 763444 35676 763496
rect 41696 763444 41748 763496
rect 35808 763172 35860 763224
rect 41696 763104 41748 763156
rect 57244 763172 57296 763224
rect 42616 763036 42668 763088
rect 42064 761880 42116 761932
rect 48964 761880 49016 761932
rect 35808 761812 35860 761864
rect 41696 761812 41748 761864
rect 35164 759772 35216 759824
rect 41696 759772 41748 759824
rect 32404 759636 32456 759688
rect 41604 759636 41656 759688
rect 33784 758276 33836 758328
rect 39304 758276 39356 758328
rect 42432 758072 42484 758124
rect 42800 758072 42852 758124
rect 42064 757936 42116 757988
rect 42432 757936 42484 757988
rect 45100 755488 45152 755540
rect 62764 755488 62816 755540
rect 42892 754876 42944 754928
rect 44732 754876 44784 754928
rect 42248 754264 42300 754316
rect 45100 754264 45152 754316
rect 44180 753516 44232 753568
rect 42248 753380 42300 753432
rect 42340 749980 42392 750032
rect 42340 749300 42392 749352
rect 61384 747124 61436 747176
rect 63040 747124 63092 747176
rect 653404 746580 653456 746632
rect 675392 746580 675444 746632
rect 45100 746512 45152 746564
rect 62120 746512 62172 746564
rect 42156 745424 42208 745476
rect 42708 745424 42760 745476
rect 42800 744064 42852 744116
rect 62120 743860 62172 743912
rect 671712 743860 671764 743912
rect 675116 743860 675168 743912
rect 46204 743724 46256 743776
rect 62120 743724 62172 743776
rect 58624 742364 58676 742416
rect 62120 742364 62172 742416
rect 671804 742160 671856 742212
rect 675484 742160 675536 742212
rect 674840 739780 674892 739832
rect 675392 739780 675444 739832
rect 672448 739100 672500 739152
rect 675300 739100 675352 739152
rect 673460 738624 673512 738676
rect 675392 738624 675444 738676
rect 669596 738284 669648 738336
rect 675300 737944 675352 737996
rect 657544 735564 657596 735616
rect 675208 735700 675260 735752
rect 654784 734136 654836 734188
rect 675300 734136 675352 734188
rect 675300 733660 675352 733712
rect 651472 733388 651524 733440
rect 668584 733388 668636 733440
rect 675300 733320 675352 733372
rect 651472 731416 651524 731468
rect 658924 731416 658976 731468
rect 651380 731076 651432 731128
rect 653404 731076 653456 731128
rect 652668 730668 652720 730720
rect 661684 730668 661736 730720
rect 673828 730464 673880 730516
rect 674656 730464 674708 730516
rect 675300 730464 675352 730516
rect 43628 730328 43680 730380
rect 58624 730328 58676 730380
rect 651472 729988 651524 730040
rect 657544 729988 657596 730040
rect 675024 729852 675076 729904
rect 42432 729308 42484 729360
rect 62764 729308 62816 729360
rect 41328 728764 41380 728816
rect 41696 728764 41748 728816
rect 42064 728764 42116 728816
rect 44364 728764 44416 728816
rect 41328 728628 41380 728680
rect 41696 728628 41748 728680
rect 42064 728628 42116 728680
rect 44548 728628 44600 728680
rect 651472 728492 651524 728544
rect 654784 728492 654836 728544
rect 673092 728288 673144 728340
rect 670884 728084 670936 728136
rect 40684 727404 40736 727456
rect 41696 727404 41748 727456
rect 42064 727404 42116 727456
rect 43444 727404 43496 727456
rect 40868 727268 40920 727320
rect 41696 727268 41748 727320
rect 42064 727268 42116 727320
rect 43444 727268 43496 727320
rect 674748 727200 674800 727252
rect 681004 727200 681056 727252
rect 674472 726656 674524 726708
rect 684132 726656 684184 726708
rect 674288 726452 674340 726504
rect 683488 726384 683540 726436
rect 41144 726044 41196 726096
rect 41604 726044 41656 726096
rect 40960 725908 41012 725960
rect 41420 725908 41472 725960
rect 673828 724344 673880 724396
rect 673368 724208 673420 724260
rect 675300 721692 675352 721744
rect 675300 721216 675352 721268
rect 675300 720808 675352 720860
rect 675300 720468 675352 720520
rect 42800 718972 42852 719024
rect 61384 718972 61436 719024
rect 32404 716864 32456 716916
rect 40224 716864 40276 716916
rect 674288 716456 674340 716508
rect 676036 716456 676088 716508
rect 656164 716252 656216 716304
rect 674012 716252 674064 716304
rect 669964 715708 670016 715760
rect 674012 715708 674064 715760
rect 35164 715640 35216 715692
rect 41512 715640 41564 715692
rect 31668 715504 31720 715556
rect 40592 715504 40644 715556
rect 671068 715436 671120 715488
rect 674012 715436 674064 715488
rect 674288 715436 674340 715488
rect 675852 715436 675904 715488
rect 674288 715300 674340 715352
rect 676036 715300 676088 715352
rect 42064 715028 42116 715080
rect 42432 715028 42484 715080
rect 660304 714824 660356 714876
rect 674012 714892 674064 714944
rect 39304 714756 39356 714808
rect 41696 714756 41748 714808
rect 671896 714484 671948 714536
rect 674012 714484 674064 714536
rect 671068 713192 671120 713244
rect 674012 713192 674064 713244
rect 672264 712852 672316 712904
rect 674012 712852 674064 712904
rect 671896 712376 671948 712428
rect 674012 712376 674064 712428
rect 43812 712240 43864 712292
rect 51724 712240 51776 712292
rect 42340 711084 42392 711136
rect 43812 711084 43864 711136
rect 43812 710948 43864 711000
rect 44732 710948 44784 711000
rect 42340 710404 42392 710456
rect 42800 710404 42852 710456
rect 671436 709996 671488 710048
rect 674012 709996 674064 710048
rect 674288 709452 674340 709504
rect 676036 709452 676088 709504
rect 669044 709316 669096 709368
rect 674012 709316 674064 709368
rect 670608 709180 670660 709232
rect 674012 709180 674064 709232
rect 674656 707548 674708 707600
rect 676036 707548 676088 707600
rect 670424 705916 670476 705968
rect 674012 705916 674064 705968
rect 674288 705780 674340 705832
rect 676036 705780 676088 705832
rect 674472 705304 674524 705356
rect 683120 705304 683172 705356
rect 669228 705168 669280 705220
rect 674012 705168 674064 705220
rect 51724 705100 51776 705152
rect 62120 705100 62172 705152
rect 674288 704012 674340 704064
rect 676036 704012 676088 704064
rect 667848 703808 667900 703860
rect 674012 703808 674064 703860
rect 44732 703740 44784 703792
rect 62120 703740 62172 703792
rect 654784 701156 654836 701208
rect 674012 701156 674064 701208
rect 674288 701088 674340 701140
rect 675392 701088 675444 701140
rect 42800 701020 42852 701072
rect 62212 701020 62264 701072
rect 666468 701020 666520 701072
rect 674012 701020 674064 701072
rect 46204 700272 46256 700324
rect 62120 700272 62172 700324
rect 58624 699524 58676 699576
rect 62304 699524 62356 699576
rect 666284 696940 666336 696992
rect 674012 696940 674064 696992
rect 674288 696940 674340 696992
rect 675116 696940 675168 696992
rect 674288 693132 674340 693184
rect 675116 693132 675168 693184
rect 668952 693064 669004 693116
rect 674012 693064 674064 693116
rect 674288 692996 674340 693048
rect 675392 692996 675444 693048
rect 656440 690072 656492 690124
rect 674012 690072 674064 690124
rect 674472 690004 674524 690056
rect 675116 690004 675168 690056
rect 674748 688984 674800 689036
rect 675208 688984 675260 689036
rect 652760 688780 652812 688832
rect 674012 688780 674064 688832
rect 651472 688644 651524 688696
rect 657544 688644 657596 688696
rect 35808 687488 35860 687540
rect 41696 687488 41748 687540
rect 35440 687216 35492 687268
rect 651472 687216 651524 687268
rect 669964 687216 670016 687268
rect 41696 687148 41748 687200
rect 651472 687012 651524 687064
rect 654784 687012 654836 687064
rect 42064 686468 42116 686520
rect 63408 686468 63460 686520
rect 651656 686468 651708 686520
rect 667204 686468 667256 686520
rect 35624 686400 35676 686452
rect 41696 686400 41748 686452
rect 35808 686264 35860 686316
rect 41696 686264 41748 686316
rect 42064 686264 42116 686316
rect 43812 686264 43864 686316
rect 42064 686060 42116 686112
rect 44548 686060 44600 686112
rect 35808 685992 35860 686044
rect 41696 685992 41748 686044
rect 670884 685924 670936 685976
rect 673000 685924 673052 685976
rect 35440 685856 35492 685908
rect 41696 685856 41748 685908
rect 42064 685856 42116 685908
rect 44272 685856 44324 685908
rect 651472 685516 651524 685568
rect 656440 685516 656492 685568
rect 35808 684972 35860 685024
rect 42064 684904 42116 684956
rect 45100 684904 45152 684956
rect 41328 684768 41380 684820
rect 35624 684632 35676 684684
rect 41512 684632 41564 684684
rect 35808 684496 35860 684548
rect 41696 684496 41748 684548
rect 35808 683408 35860 683460
rect 41696 683408 41748 683460
rect 35624 683272 35676 683324
rect 41512 683272 41564 683324
rect 35440 683136 35492 683188
rect 41696 683136 41748 683188
rect 42064 683136 42116 683188
rect 44364 683136 44416 683188
rect 674840 682524 674892 682576
rect 683212 682524 683264 682576
rect 674840 682388 674892 682440
rect 683488 682388 683540 682440
rect 35624 681844 35676 681896
rect 41604 681844 41656 681896
rect 35808 681708 35860 681760
rect 41420 681708 41472 681760
rect 42064 681708 42116 681760
rect 42616 681708 42668 681760
rect 35808 680620 35860 680672
rect 41696 680620 41748 680672
rect 35808 679396 35860 679448
rect 41696 679396 41748 679448
rect 35624 679124 35676 679176
rect 41696 679192 41748 679244
rect 42064 679192 42116 679244
rect 44180 679192 44232 679244
rect 35440 678988 35492 679040
rect 41696 678988 41748 679040
rect 42064 678988 42116 679040
rect 44640 678988 44692 679040
rect 40776 677696 40828 677748
rect 41604 677696 41656 677748
rect 42800 676200 42852 676252
rect 55864 676200 55916 676252
rect 33048 674092 33100 674144
rect 41512 674092 41564 674144
rect 35164 672868 35216 672920
rect 39580 672868 39632 672920
rect 31024 672732 31076 672784
rect 41696 672596 41748 672648
rect 42064 672528 42116 672580
rect 42800 672528 42852 672580
rect 42616 672392 42668 672444
rect 42800 672188 42852 672240
rect 673736 671304 673788 671356
rect 668584 671100 668636 671152
rect 673736 671100 673788 671152
rect 661684 670692 661736 670744
rect 674840 669808 674892 669860
rect 676496 669808 676548 669860
rect 658924 669468 658976 669520
rect 673736 669468 673788 669520
rect 45836 669400 45888 669452
rect 53104 669332 53156 669384
rect 670240 669332 670292 669384
rect 673368 669332 673420 669384
rect 673736 668652 673788 668704
rect 671068 668516 671120 668568
rect 673736 668516 673788 668568
rect 671436 668176 671488 668228
rect 45652 667904 45704 667956
rect 58624 667904 58676 667956
rect 671068 667904 671120 667956
rect 673736 667904 673788 667956
rect 673736 667292 673788 667344
rect 671620 667156 671672 667208
rect 673736 667156 673788 667208
rect 42248 666884 42300 666936
rect 44180 666884 44232 666936
rect 671896 666884 671948 666936
rect 44640 666544 44692 666596
rect 671896 666544 671948 666596
rect 673736 666544 673788 666596
rect 42340 665660 42392 665712
rect 669596 665252 669648 665304
rect 673736 665252 673788 665304
rect 672448 665116 672500 665168
rect 673368 665116 673420 665168
rect 671712 664368 671764 664420
rect 673736 664368 673788 664420
rect 669412 663892 669464 663944
rect 673736 663892 673788 663944
rect 674840 663756 674892 663808
rect 676036 663756 676088 663808
rect 672080 663416 672132 663468
rect 673368 663416 673420 663468
rect 42248 663008 42300 663060
rect 43996 663008 44048 663060
rect 42432 662872 42484 662924
rect 45560 662872 45612 662924
rect 671252 661580 671304 661632
rect 673736 661580 673788 661632
rect 668216 661104 668268 661156
rect 673736 661104 673788 661156
rect 53104 660900 53156 660952
rect 62120 660900 62172 660952
rect 668768 660084 668820 660136
rect 673736 660084 673788 660136
rect 674840 659812 674892 659864
rect 683120 659812 683172 659864
rect 58624 659540 58676 659592
rect 62120 659540 62172 659592
rect 45376 658928 45428 658980
rect 62304 658928 62356 658980
rect 42524 657500 42576 657552
rect 62120 657500 62172 657552
rect 46204 656820 46256 656872
rect 62120 656820 62172 656872
rect 653404 655528 653456 655580
rect 673736 655528 673788 655580
rect 655520 645872 655572 645924
rect 673736 645872 673788 645924
rect 35808 644444 35860 644496
rect 39764 644444 39816 644496
rect 35808 643492 35860 643544
rect 40224 643492 40276 643544
rect 35532 643220 35584 643272
rect 41696 643288 41748 643340
rect 42064 643288 42116 643340
rect 43812 643288 43864 643340
rect 35348 643084 35400 643136
rect 41696 643084 41748 643136
rect 42064 643084 42116 643136
rect 58624 643084 58676 643136
rect 655336 643084 655388 643136
rect 673736 643084 673788 643136
rect 38568 642472 38620 642524
rect 41696 642472 41748 642524
rect 42064 642336 42116 642388
rect 62948 642336 63000 642388
rect 651472 642336 651524 642388
rect 660304 642336 660356 642388
rect 35808 642132 35860 642184
rect 39580 642132 39632 642184
rect 35808 641860 35860 641912
rect 40776 641996 40828 642048
rect 35624 641724 35676 641776
rect 41696 641724 41748 641776
rect 42064 641724 42116 641776
rect 45284 641724 45336 641776
rect 35808 640772 35860 640824
rect 39304 640704 39356 640756
rect 35808 640432 35860 640484
rect 40408 640500 40460 640552
rect 674840 640364 674892 640416
rect 35624 640296 35676 640348
rect 40868 640296 40920 640348
rect 651472 640296 651524 640348
rect 668584 640296 668636 640348
rect 675300 640228 675352 640280
rect 651380 640092 651432 640144
rect 653404 640092 653456 640144
rect 35808 639208 35860 639260
rect 41696 639208 41748 639260
rect 35532 638936 35584 638988
rect 39304 638936 39356 638988
rect 651656 638868 651708 638920
rect 655336 638868 655388 638920
rect 651472 638732 651524 638784
rect 655520 638732 655572 638784
rect 34428 638188 34480 638240
rect 41696 638188 41748 638240
rect 35808 637848 35860 637900
rect 36544 637848 36596 637900
rect 674472 636964 674524 637016
rect 683212 636964 683264 637016
rect 35624 636896 35676 636948
rect 40592 636896 40644 636948
rect 674288 636828 674340 636880
rect 683396 636828 683448 636880
rect 35808 636692 35860 636744
rect 40132 636624 40184 636676
rect 35808 636352 35860 636404
rect 40776 636420 40828 636472
rect 35532 636216 35584 636268
rect 40592 636216 40644 636268
rect 671988 636148 672040 636200
rect 672172 636148 672224 636200
rect 651840 635468 651892 635520
rect 661684 635468 661736 635520
rect 674932 635468 674984 635520
rect 675668 635468 675720 635520
rect 35808 634788 35860 634840
rect 39948 634788 40000 634840
rect 35808 633836 35860 633888
rect 40500 633700 40552 633752
rect 35808 633428 35860 633480
rect 41512 633428 41564 633480
rect 42156 633428 42208 633480
rect 63408 633428 63460 633480
rect 671528 632952 671580 633004
rect 671344 632884 671396 632936
rect 671344 632748 671396 632800
rect 671528 632612 671580 632664
rect 36544 630572 36596 630624
rect 41604 630504 41656 630556
rect 671896 630028 671948 630080
rect 672080 629348 672132 629400
rect 35164 628532 35216 628584
rect 39672 628532 39724 628584
rect 667204 626084 667256 626136
rect 672816 626084 672868 626136
rect 44180 625812 44232 625864
rect 63132 625812 63184 625864
rect 669964 625540 670016 625592
rect 672172 625540 672224 625592
rect 42340 625132 42392 625184
rect 44364 625132 44416 625184
rect 657544 625132 657596 625184
rect 672816 625132 672868 625184
rect 670240 624996 670292 625048
rect 672816 624996 672868 625048
rect 670424 624656 670476 624708
rect 672816 624656 672868 624708
rect 671436 624316 671488 624368
rect 672816 624316 672868 624368
rect 670240 623840 670292 623892
rect 672816 623840 672868 623892
rect 44088 623772 44140 623824
rect 671068 623500 671120 623552
rect 672816 623500 672868 623552
rect 42340 623364 42392 623416
rect 669412 623024 669464 623076
rect 672816 623024 672868 623076
rect 674656 623024 674708 623076
rect 683396 623024 683448 623076
rect 42432 621460 42484 621512
rect 42616 621188 42668 621240
rect 666468 621052 666520 621104
rect 672816 621052 672868 621104
rect 674288 620984 674340 621036
rect 676220 620984 676272 621036
rect 668952 620236 669004 620288
rect 672816 620236 672868 620288
rect 670884 619964 670936 620016
rect 672816 619964 672868 620016
rect 666284 619692 666336 619744
rect 672816 619692 672868 619744
rect 674380 619692 674432 619744
rect 676036 619692 676088 619744
rect 42248 619624 42300 619676
rect 42892 619624 42944 619676
rect 42708 618876 42760 618928
rect 43904 618876 43956 618928
rect 674288 618468 674340 618520
rect 676220 618468 676272 618520
rect 674288 617992 674340 618044
rect 676496 617992 676548 618044
rect 674288 617856 674340 617908
rect 676220 617856 676272 617908
rect 670608 617448 670660 617500
rect 674012 617448 674064 617500
rect 674288 617448 674340 617500
rect 676220 617448 676272 617500
rect 42156 617108 42208 617160
rect 42708 617108 42760 617160
rect 668400 616836 668452 616888
rect 674012 616836 674064 616888
rect 44180 616768 44232 616820
rect 62120 616768 62172 616820
rect 669780 615612 669832 615664
rect 674012 615612 674064 615664
rect 674288 615476 674340 615528
rect 683120 615476 683172 615528
rect 674288 614592 674340 614644
rect 676220 614592 676272 614644
rect 42800 614116 42852 614168
rect 62120 614116 62172 614168
rect 670608 614116 670660 614168
rect 674012 614116 674064 614168
rect 58624 613980 58676 614032
rect 62120 613980 62172 614032
rect 46204 613368 46256 613420
rect 62120 613368 62172 613420
rect 43076 612824 43128 612876
rect 43904 612688 43956 612740
rect 43260 612620 43312 612672
rect 42248 612348 42300 612400
rect 53104 612552 53156 612604
rect 44916 611940 44968 611992
rect 46204 611668 46256 611720
rect 44088 611532 44140 611584
rect 653404 611328 653456 611380
rect 674012 611328 674064 611380
rect 674288 611328 674340 611380
rect 675392 611328 675444 611380
rect 50160 611260 50212 611312
rect 44318 611124 44370 611176
rect 44732 610716 44784 610768
rect 50160 610104 50212 610156
rect 58624 610104 58676 610156
rect 64328 609968 64380 610020
rect 669044 608608 669096 608660
rect 674012 608608 674064 608660
rect 674288 608608 674340 608660
rect 675116 608608 675168 608660
rect 673552 607248 673604 607300
rect 673552 607044 673604 607096
rect 673276 603508 673328 603560
rect 674012 603508 674064 603560
rect 674288 603236 674340 603288
rect 675116 603236 675168 603288
rect 657544 600312 657596 600364
rect 674012 600312 674064 600364
rect 654784 598952 654836 599004
rect 674012 599360 674064 599412
rect 674564 598952 674616 599004
rect 675300 598952 675352 599004
rect 674472 598340 674524 598392
rect 675300 598340 675352 598392
rect 651472 597524 651524 597576
rect 669964 597524 670016 597576
rect 43076 597388 43128 597440
rect 43076 596980 43128 597032
rect 651472 596164 651524 596216
rect 667204 596164 667256 596216
rect 40132 595756 40184 595808
rect 41696 595756 41748 595808
rect 651656 595484 651708 595536
rect 653404 595484 653456 595536
rect 41328 594804 41380 594856
rect 41696 594804 41748 594856
rect 651472 594804 651524 594856
rect 658924 594804 658976 594856
rect 39948 594668 40000 594720
rect 41696 594668 41748 594720
rect 651472 594668 651524 594720
rect 657544 594668 657596 594720
rect 651472 593240 651524 593292
rect 654784 593240 654836 593292
rect 674748 592560 674800 592612
rect 683396 592628 683448 592680
rect 39304 591404 39356 591456
rect 41420 591404 41472 591456
rect 35808 590928 35860 590980
rect 40776 590928 40828 590980
rect 35624 590656 35676 590708
rect 41696 590724 41748 590776
rect 42064 590656 42116 590708
rect 43260 590656 43312 590708
rect 674840 590588 674892 590640
rect 682384 590588 682436 590640
rect 675300 590384 675352 590436
rect 675116 590180 675168 590232
rect 674472 588548 674524 588600
rect 684040 588548 684092 588600
rect 33048 587120 33100 587172
rect 41512 587120 41564 587172
rect 37924 585828 37976 585880
rect 41696 585828 41748 585880
rect 42064 585828 42116 585880
rect 42616 585828 42668 585880
rect 31024 585692 31076 585744
rect 41696 585692 41748 585744
rect 42064 585624 42116 585676
rect 42708 585624 42760 585676
rect 672264 584400 672316 584452
rect 672632 584400 672684 584452
rect 42432 582428 42484 582480
rect 42248 582088 42300 582140
rect 661684 581000 661736 581052
rect 673644 581000 673696 581052
rect 42432 580592 42484 580644
rect 43260 580592 43312 580644
rect 668584 580252 668636 580304
rect 673644 580252 673696 580304
rect 42248 580048 42300 580100
rect 42248 579912 42300 579964
rect 670424 579844 670476 579896
rect 673644 579844 673696 579896
rect 660304 579640 660356 579692
rect 673092 579640 673144 579692
rect 670792 579368 670844 579420
rect 673644 579368 673696 579420
rect 670240 579028 670292 579080
rect 673644 579028 673696 579080
rect 671160 578552 671212 578604
rect 673644 578552 673696 578604
rect 669412 578144 669464 578196
rect 673644 578144 673696 578196
rect 670240 577736 670292 577788
rect 673644 577736 673696 577788
rect 671436 577396 671488 577448
rect 673644 577396 673696 577448
rect 669412 576920 669464 576972
rect 673644 576920 673696 576972
rect 45100 575424 45152 575476
rect 62120 575424 62172 575476
rect 671620 574540 671672 574592
rect 673644 574540 673696 574592
rect 671988 574132 672040 574184
rect 673644 574132 673696 574184
rect 51724 573996 51776 574048
rect 62120 573996 62172 574048
rect 672264 573996 672316 574048
rect 673092 573996 673144 574048
rect 42248 573452 42300 573504
rect 42708 573452 42760 573504
rect 669596 572228 669648 572280
rect 673644 572228 673696 572280
rect 674472 571548 674524 571600
rect 676220 571548 676272 571600
rect 671804 571412 671856 571464
rect 673644 571412 673696 571464
rect 42064 570936 42116 570988
rect 42616 570936 42668 570988
rect 674840 570460 674892 570512
rect 675484 570460 675536 570512
rect 683120 570460 683172 570512
rect 671344 570392 671396 570444
rect 671988 570120 672040 570172
rect 673644 570120 673696 570172
rect 673644 569916 673696 569968
rect 669780 568556 669832 568608
rect 673644 568556 673696 568608
rect 653404 565836 653456 565888
rect 673644 565836 673696 565888
rect 665088 564544 665140 564596
rect 673644 564544 673696 564596
rect 661040 554752 661092 554804
rect 673644 554752 673696 554804
rect 655152 553392 655204 553444
rect 673644 553392 673696 553444
rect 651472 552644 651524 552696
rect 665824 552644 665876 552696
rect 675208 552576 675260 552628
rect 675208 552304 675260 552356
rect 674656 550604 674708 550656
rect 674840 550604 674892 550656
rect 40960 550468 41012 550520
rect 41696 550468 41748 550520
rect 675208 550468 675260 550520
rect 651656 550332 651708 550384
rect 653404 550332 653456 550384
rect 651472 549856 651524 549908
rect 664444 549856 664496 549908
rect 675300 549788 675352 549840
rect 651472 549176 651524 549228
rect 661040 549176 661092 549228
rect 651472 548836 651524 548888
rect 655152 548836 655204 548888
rect 41328 547952 41380 548004
rect 41696 547884 41748 547936
rect 42064 547884 42116 547936
rect 43260 547884 43312 547936
rect 29644 547136 29696 547188
rect 41696 547136 41748 547188
rect 675576 547136 675628 547188
rect 683212 547136 683264 547188
rect 674840 545980 674892 546032
rect 682384 545844 682436 545896
rect 667204 535916 667256 535968
rect 672632 535916 672684 535968
rect 669964 535644 670016 535696
rect 672632 535644 672684 535696
rect 670792 534828 670844 534880
rect 672632 534828 672684 534880
rect 671160 534556 671212 534608
rect 672632 534556 672684 534608
rect 658924 534216 658976 534268
rect 672632 534216 672684 534268
rect 674288 534080 674340 534132
rect 676036 534080 676088 534132
rect 670240 533332 670292 533384
rect 672448 533332 672500 533384
rect 674288 533332 674340 533384
rect 683580 533332 683632 533384
rect 42432 532720 42484 532772
rect 43076 532720 43128 532772
rect 669412 532516 669464 532568
rect 672448 532516 672500 532568
rect 673828 532176 673880 532228
rect 675484 531972 675536 532024
rect 676220 531972 676272 532024
rect 673828 531768 673880 531820
rect 51724 531224 51776 531276
rect 62120 531224 62172 531276
rect 45284 531088 45336 531140
rect 62120 531088 62172 531140
rect 673276 530884 673328 530936
rect 674012 530884 674064 530936
rect 674288 530816 674340 530868
rect 676036 530816 676088 530868
rect 667388 529932 667440 529984
rect 674012 529932 674064 529984
rect 674288 529932 674340 529984
rect 676036 529932 676088 529984
rect 42156 529456 42208 529508
rect 42616 529456 42668 529508
rect 670976 529252 671028 529304
rect 674012 529252 674064 529304
rect 674288 529184 674340 529236
rect 676036 529184 676088 529236
rect 674288 528980 674340 529032
rect 676220 528980 676272 529032
rect 45284 528572 45336 528624
rect 62120 528572 62172 528624
rect 668860 528572 668912 528624
rect 674012 528572 674064 528624
rect 54484 527076 54536 527128
rect 62120 527076 62172 527128
rect 42064 527008 42116 527060
rect 42616 527008 42668 527060
rect 674656 526736 674708 526788
rect 676036 526736 676088 526788
rect 674288 526328 674340 526380
rect 676036 526328 676088 526380
rect 667572 524424 667624 524476
rect 674012 524424 674064 524476
rect 674288 524424 674340 524476
rect 683120 524424 683172 524476
rect 663800 521568 663852 521620
rect 667572 521568 667624 521620
rect 675484 520208 675536 520260
rect 678980 520208 679032 520260
rect 675668 518780 675720 518832
rect 677876 518780 677928 518832
rect 656348 514020 656400 514072
rect 663800 514020 663852 514072
rect 653404 510620 653456 510672
rect 656348 510620 656400 510672
rect 675116 503616 675168 503668
rect 679624 503616 679676 503668
rect 675300 503480 675352 503532
rect 681004 503480 681056 503532
rect 674840 500896 674892 500948
rect 681188 500896 681240 500948
rect 652024 500216 652076 500268
rect 669964 500216 670016 500268
rect 650644 494708 650696 494760
rect 653404 494708 653456 494760
rect 674288 491988 674340 492040
rect 674656 491988 674708 492040
rect 669964 491852 670016 491904
rect 674012 491852 674064 491904
rect 674288 491784 674340 491836
rect 675852 491784 675904 491836
rect 674288 491648 674340 491700
rect 676036 491648 676088 491700
rect 665824 491444 665876 491496
rect 674012 491444 674064 491496
rect 664444 491308 664496 491360
rect 673828 491308 673880 491360
rect 670792 490900 670844 490952
rect 674012 490900 674064 490952
rect 672448 490424 672500 490476
rect 674012 490424 674064 490476
rect 672632 490084 672684 490136
rect 674012 490084 674064 490136
rect 672632 489608 672684 489660
rect 674012 489608 674064 489660
rect 671620 489268 671672 489320
rect 674012 489268 674064 489320
rect 671160 488452 671212 488504
rect 674012 488452 674064 488504
rect 674288 486140 674340 486192
rect 676036 486140 676088 486192
rect 672264 486004 672316 486056
rect 673828 486004 673880 486056
rect 665088 485800 665140 485852
rect 674012 485800 674064 485852
rect 674288 485120 674340 485172
rect 676036 485120 676088 485172
rect 667020 484372 667072 484424
rect 674012 484372 674064 484424
rect 674472 483964 674524 484016
rect 676036 483964 676088 484016
rect 671804 483148 671856 483200
rect 674012 483148 674064 483200
rect 676220 482944 676272 482996
rect 677416 482944 677468 482996
rect 669964 480700 670016 480752
rect 670424 480700 670476 480752
rect 674012 480700 674064 480752
rect 674288 480360 674340 480412
rect 683120 480360 683172 480412
rect 676036 476076 676088 476128
rect 680360 476076 680412 476128
rect 657544 467100 657596 467152
rect 669964 467100 670016 467152
rect 653404 460164 653456 460216
rect 657544 460164 657596 460216
rect 667848 456560 667900 456612
rect 669228 455948 669280 456000
rect 673368 455812 673420 455864
rect 668216 455608 668268 455660
rect 673276 455336 673328 455388
rect 673388 455200 673440 455252
rect 673506 455200 673558 455252
rect 674288 454860 674340 454912
rect 675852 454860 675904 454912
rect 672080 454792 672132 454844
rect 673046 454588 673098 454640
rect 674288 454588 674340 454640
rect 675484 454588 675536 454640
rect 672816 454452 672868 454504
rect 672954 454316 673006 454368
rect 674288 454316 674340 454368
rect 675668 454316 675720 454368
rect 672264 453908 672316 453960
rect 674288 453908 674340 453960
rect 676036 453908 676088 453960
rect 44824 451392 44876 451444
rect 47768 451392 47820 451444
rect 35808 429156 35860 429208
rect 41328 429156 41380 429208
rect 35808 427932 35860 427984
rect 41604 427932 41656 427984
rect 41144 424328 41196 424380
rect 41696 424328 41748 424380
rect 33048 417392 33100 417444
rect 41696 417392 41748 417444
rect 42064 417256 42116 417308
rect 42524 417256 42576 417308
rect 34520 416032 34572 416084
rect 41604 416032 41656 416084
rect 42248 409776 42300 409828
rect 42708 409776 42760 409828
rect 42248 407668 42300 407720
rect 42616 407668 42668 407720
rect 51080 404268 51132 404320
rect 62120 404268 62172 404320
rect 674564 403248 674616 403300
rect 676220 403248 676272 403300
rect 51448 402908 51500 402960
rect 62120 402908 62172 402960
rect 51080 400188 51132 400240
rect 62120 400188 62172 400240
rect 44824 400052 44876 400104
rect 62120 400052 62172 400104
rect 674932 398828 674984 398880
rect 676036 398828 676088 398880
rect 54484 398760 54536 398812
rect 62120 398760 62172 398812
rect 675024 395700 675076 395752
rect 676220 395700 676272 395752
rect 674380 395496 674432 395548
rect 676220 395496 676272 395548
rect 674472 394272 674524 394324
rect 676220 394272 676272 394324
rect 41328 386384 41380 386436
rect 41604 386384 41656 386436
rect 679624 386724 679676 386776
rect 674840 386112 674892 386164
rect 675300 386112 675352 386164
rect 675484 385976 675536 386028
rect 41328 382508 41380 382560
rect 41604 382508 41656 382560
rect 35808 379516 35860 379568
rect 40408 379516 40460 379568
rect 674472 378088 674524 378140
rect 675116 378088 675168 378140
rect 35808 376728 35860 376780
rect 41696 376728 41748 376780
rect 674380 375300 674432 375352
rect 675116 375300 675168 375352
rect 651472 373940 651524 373992
rect 663064 373940 663116 373992
rect 33968 373260 34020 373312
rect 41696 373260 41748 373312
rect 39304 371628 39356 371680
rect 41696 371628 41748 371680
rect 42064 371560 42116 371612
rect 42524 371560 42576 371612
rect 651472 370948 651524 371000
rect 654784 370948 654836 371000
rect 42248 365304 42300 365356
rect 43076 365304 43128 365356
rect 662420 364352 662472 364404
rect 666468 364352 666520 364404
rect 42248 362856 42300 362908
rect 42248 362584 42300 362636
rect 44732 361496 44784 361548
rect 62120 361496 62172 361548
rect 657544 360204 657596 360256
rect 662420 360204 662472 360256
rect 51080 360136 51132 360188
rect 62120 360136 62172 360188
rect 42156 359932 42208 359984
rect 42892 359932 42944 359984
rect 54484 356668 54536 356720
rect 62120 356668 62172 356720
rect 44640 354968 44692 355020
rect 44640 354832 44692 354884
rect 44640 354492 44692 354544
rect 44732 354356 44784 354408
rect 45652 353812 45704 353864
rect 45836 353676 45888 353728
rect 45652 353404 45704 353456
rect 46020 353200 46072 353252
rect 652024 348372 652076 348424
rect 657544 348372 657596 348424
rect 35808 343748 35860 343800
rect 40224 343748 40276 343800
rect 35532 343612 35584 343664
rect 40040 343612 40092 343664
rect 35808 341300 35860 341352
rect 39856 341300 39908 341352
rect 35808 341164 35860 341216
rect 40224 341164 40276 341216
rect 35532 341028 35584 341080
rect 40040 341028 40092 341080
rect 35808 339600 35860 339652
rect 37924 339600 37976 339652
rect 35532 339464 35584 339516
rect 38936 339464 38988 339516
rect 35808 335316 35860 335368
rect 40224 335316 40276 335368
rect 35808 334092 35860 334144
rect 39764 334092 39816 334144
rect 674472 331032 674524 331084
rect 675116 331032 675168 331084
rect 651472 328244 651524 328296
rect 654784 328244 654836 328296
rect 651748 325592 651800 325644
rect 653588 325592 653640 325644
rect 650828 322940 650880 322992
rect 653404 322940 653456 322992
rect 42248 320220 42300 320272
rect 42616 319948 42668 320000
rect 53840 317364 53892 317416
rect 62120 317364 62172 317416
rect 53840 314712 53892 314764
rect 62120 314712 62172 314764
rect 674380 311992 674432 312044
rect 675484 311992 675536 312044
rect 676220 306348 676272 306400
rect 676864 306348 676916 306400
rect 50528 305600 50580 305652
rect 58808 305600 58860 305652
rect 675852 304852 675904 304904
rect 676404 304852 676456 304904
rect 651380 303356 651432 303408
rect 653404 303356 653456 303408
rect 651472 300772 651524 300824
rect 658924 300772 658976 300824
rect 41144 299072 41196 299124
rect 41696 299072 41748 299124
rect 651472 298120 651524 298172
rect 660580 298120 660632 298172
rect 675852 298052 675904 298104
rect 678244 298052 678296 298104
rect 651656 296760 651708 296812
rect 658924 296692 658976 296744
rect 675484 296352 675536 296404
rect 675300 296148 675352 296200
rect 675300 295400 675352 295452
rect 675484 295196 675536 295248
rect 41328 294584 41380 294636
rect 41696 294584 41748 294636
rect 42064 294448 42116 294500
rect 42524 294448 42576 294500
rect 57428 294040 57480 294092
rect 62120 294040 62172 294092
rect 651472 293972 651524 294024
rect 664444 293972 664496 294024
rect 47584 293904 47636 293956
rect 50528 293904 50580 293956
rect 40592 292544 40644 292596
rect 41604 292544 41656 292596
rect 56048 292544 56100 292596
rect 62764 292544 62816 292596
rect 651472 292544 651524 292596
rect 660304 292544 660356 292596
rect 54484 292408 54536 292460
rect 62120 292408 62172 292460
rect 35808 291320 35860 291372
rect 41604 291320 41656 291372
rect 51724 291116 51776 291168
rect 62120 291116 62172 291168
rect 649264 290776 649316 290828
rect 651748 290776 651800 290828
rect 651472 289824 651524 289876
rect 663064 289824 663116 289876
rect 51724 288464 51776 288516
rect 62120 288464 62172 288516
rect 651472 288396 651524 288448
rect 672172 288396 672224 288448
rect 33048 287648 33100 287700
rect 41512 287648 41564 287700
rect 651472 287036 651524 287088
rect 667756 287036 667808 287088
rect 674380 286628 674432 286680
rect 675300 286628 675352 286680
rect 35164 286288 35216 286340
rect 41696 286288 41748 286340
rect 42248 286288 42300 286340
rect 42616 286288 42668 286340
rect 46388 285676 46440 285728
rect 62120 285676 62172 285728
rect 651472 285676 651524 285728
rect 667572 285676 667624 285728
rect 47768 284928 47820 284980
rect 60004 284928 60056 284980
rect 45560 284316 45612 284368
rect 62948 284316 63000 284368
rect 651472 284316 651524 284368
rect 672356 284316 672408 284368
rect 651472 282888 651524 282940
rect 667204 282888 667256 282940
rect 54484 280372 54536 280424
rect 62120 280372 62172 280424
rect 53288 280168 53340 280220
rect 62304 280168 62356 280220
rect 651472 280168 651524 280220
rect 667388 280168 667440 280220
rect 62580 278672 62632 278724
rect 671344 278672 671396 278724
rect 63316 278536 63368 278588
rect 671712 278468 671764 278520
rect 58808 278400 58860 278452
rect 650828 278400 650880 278452
rect 50528 278264 50580 278316
rect 69204 278264 69256 278316
rect 60004 278128 60056 278180
rect 649264 278264 649316 278316
rect 69204 277992 69256 278044
rect 650644 278128 650696 278180
rect 45468 277380 45520 277432
rect 637856 277380 637908 277432
rect 42248 277312 42300 277364
rect 43352 277312 43404 277364
rect 487988 277176 488040 277228
rect 565820 277176 565872 277228
rect 497924 277040 497976 277092
rect 579988 277040 580040 277092
rect 511632 276904 511684 276956
rect 600136 276904 600188 276956
rect 42248 276768 42300 276820
rect 42616 276768 42668 276820
rect 514484 276768 514536 276820
rect 603632 276768 603684 276820
rect 518348 276632 518400 276684
rect 609612 276632 609664 276684
rect 479984 276496 480036 276548
rect 555240 276496 555292 276548
rect 482836 276360 482888 276412
rect 557540 276360 557592 276412
rect 477040 276224 477092 276276
rect 550456 276224 550508 276276
rect 471612 276088 471664 276140
rect 543372 276088 543424 276140
rect 107200 275952 107252 276004
rect 163504 275952 163556 276004
rect 167552 275952 167604 276004
rect 178684 275952 178736 276004
rect 185216 275952 185268 276004
rect 221280 275952 221332 276004
rect 232504 275952 232556 276004
rect 240048 275952 240100 276004
rect 410800 275952 410852 276004
rect 455880 275952 455932 276004
rect 456064 275952 456116 276004
rect 509056 275952 509108 276004
rect 513196 275952 513248 276004
rect 601332 275952 601384 276004
rect 139124 275816 139176 275868
rect 174268 275816 174320 275868
rect 178132 275816 178184 275868
rect 216680 275816 216732 275868
rect 224224 275816 224276 275868
rect 232688 275816 232740 275868
rect 236092 275816 236144 275868
rect 250444 275816 250496 275868
rect 284576 275816 284628 275868
rect 290096 275816 290148 275868
rect 430212 275816 430264 275868
rect 484308 275816 484360 275868
rect 490564 275816 490616 275868
rect 505560 275816 505612 275868
rect 522764 275816 522816 275868
rect 615500 275816 615552 275868
rect 260932 275748 260984 275800
rect 266360 275748 266412 275800
rect 93032 275680 93084 275732
rect 152832 275680 152884 275732
rect 160468 275680 160520 275732
rect 199568 275680 199620 275732
rect 217140 275680 217192 275732
rect 224224 275680 224276 275732
rect 229008 275680 229060 275732
rect 243728 275680 243780 275732
rect 250260 275680 250312 275732
rect 259368 275680 259420 275732
rect 286876 275680 286928 275732
rect 291844 275680 291896 275732
rect 445024 275680 445076 275732
rect 498476 275680 498528 275732
rect 498844 275680 498896 275732
rect 512644 275680 512696 275732
rect 528192 275680 528244 275732
rect 622584 275680 622636 275732
rect 76472 275544 76524 275596
rect 86224 275544 86276 275596
rect 90732 275544 90784 275596
rect 154764 275544 154816 275596
rect 171048 275544 171100 275596
rect 211436 275544 211488 275596
rect 218336 275544 218388 275596
rect 233884 275544 233936 275596
rect 239588 275544 239640 275596
rect 255964 275544 256016 275596
rect 257344 275544 257396 275596
rect 262312 275544 262364 275596
rect 266820 275544 266872 275596
rect 276480 275544 276532 275596
rect 363880 275544 363932 275596
rect 388536 275544 388588 275596
rect 416412 275544 416464 275596
rect 462964 275544 463016 275596
rect 463148 275544 463200 275596
rect 516232 275544 516284 275596
rect 516784 275544 516836 275596
rect 526812 275544 526864 275596
rect 532332 275544 532384 275596
rect 629668 275544 629720 275596
rect 277492 275476 277544 275528
rect 285128 275476 285180 275528
rect 100116 275408 100168 275460
rect 71780 275272 71832 275324
rect 141056 275272 141108 275324
rect 156880 275408 156932 275460
rect 159456 275272 159508 275324
rect 163964 275408 164016 275460
rect 206376 275408 206428 275460
rect 221924 275408 221976 275460
rect 243544 275408 243596 275460
rect 256148 275408 256200 275460
rect 270132 275408 270184 275460
rect 358636 275408 358688 275460
rect 381452 275408 381504 275460
rect 386052 275408 386104 275460
rect 420460 275408 420512 275460
rect 435640 275408 435692 275460
rect 481732 275408 481784 275460
rect 483664 275408 483716 275460
rect 530400 275408 530452 275460
rect 537668 275408 537720 275460
rect 636752 275408 636804 275460
rect 297548 275340 297600 275392
rect 299572 275340 299624 275392
rect 299940 275340 299992 275392
rect 301136 275340 301188 275392
rect 201040 275272 201092 275324
rect 214840 275272 214892 275324
rect 239404 275272 239456 275324
rect 243176 275272 243228 275324
rect 256700 275272 256752 275324
rect 263232 275272 263284 275324
rect 273260 275272 273312 275324
rect 276296 275272 276348 275324
rect 283104 275272 283156 275324
rect 285680 275272 285732 275324
rect 291292 275272 291344 275324
rect 291660 275272 291712 275324
rect 295340 275272 295392 275324
rect 326436 275272 326488 275324
rect 335360 275272 335412 275324
rect 371056 275272 371108 275324
rect 399208 275272 399260 275324
rect 418804 275272 418856 275324
rect 466552 275272 466604 275324
rect 467564 275272 467616 275324
rect 537484 275272 537536 275324
rect 542268 275272 542320 275324
rect 643836 275272 643888 275324
rect 298744 275204 298796 275256
rect 300032 275204 300084 275256
rect 96620 275136 96672 275188
rect 149612 275136 149664 275188
rect 153384 275136 153436 275188
rect 169024 275136 169076 275188
rect 190000 275136 190052 275188
rect 222936 275136 222988 275188
rect 292856 275136 292908 275188
rect 295800 275136 295852 275188
rect 427084 275136 427136 275188
rect 477224 275136 477276 275188
rect 481732 275136 481784 275188
rect 491392 275136 491444 275188
rect 507492 275136 507544 275188
rect 594248 275136 594300 275188
rect 269212 275068 269264 275120
rect 274640 275068 274692 275120
rect 136824 275000 136876 275052
rect 137652 275000 137704 275052
rect 146208 275000 146260 275052
rect 185308 275000 185360 275052
rect 288072 275000 288124 275052
rect 292856 275000 292908 275052
rect 420552 275000 420604 275052
rect 470140 275000 470192 275052
rect 503444 275000 503496 275052
rect 587072 275000 587124 275052
rect 81256 274932 81308 274984
rect 293960 274932 294012 274984
rect 296812 274932 296864 274984
rect 145288 274864 145340 274916
rect 149796 274864 149848 274916
rect 189080 274864 189132 274916
rect 289268 274864 289320 274916
rect 292672 274864 292724 274916
rect 473084 274864 473136 274916
rect 544568 274864 544620 274916
rect 295156 274796 295208 274848
rect 297456 274796 297508 274848
rect 128544 274728 128596 274780
rect 168288 274728 168340 274780
rect 207756 274728 207808 274780
rect 210700 274728 210752 274780
rect 476764 274728 476816 274780
rect 523316 274728 523368 274780
rect 523684 274728 523736 274780
rect 533896 274728 533948 274780
rect 534724 274728 534776 274780
rect 540980 274728 541032 274780
rect 74172 274660 74224 274712
rect 76840 274660 76892 274712
rect 85948 274660 86000 274712
rect 90364 274660 90416 274712
rect 103704 274660 103756 274712
rect 104808 274660 104860 274712
rect 110788 274660 110840 274712
rect 111708 274660 111760 274712
rect 253848 274660 253900 274712
rect 256884 274660 256936 274712
rect 275100 274660 275152 274712
rect 278044 274660 278096 274712
rect 283380 274660 283432 274712
rect 289176 274660 289228 274712
rect 290464 274660 290516 274712
rect 294144 274660 294196 274712
rect 296352 274660 296404 274712
rect 298376 274660 298428 274712
rect 303436 274660 303488 274712
rect 303988 274660 304040 274712
rect 321192 274660 321244 274712
rect 328276 274660 328328 274712
rect 114376 274592 114428 274644
rect 171600 274592 171652 274644
rect 179328 274592 179380 274644
rect 214564 274592 214616 274644
rect 409788 274592 409840 274644
rect 453580 274592 453632 274644
rect 457444 274592 457496 274644
rect 480720 274592 480772 274644
rect 486792 274592 486844 274644
rect 563428 274592 563480 274644
rect 101312 274456 101364 274508
rect 160928 274456 160980 274508
rect 168748 274456 168800 274508
rect 208400 274456 208452 274508
rect 381544 274456 381596 274508
rect 392124 274456 392176 274508
rect 413836 274456 413888 274508
rect 460664 274456 460716 274508
rect 463240 274456 463292 274508
rect 483664 274456 483716 274508
rect 488356 274456 488408 274508
rect 567016 274456 567068 274508
rect 95424 274320 95476 274372
rect 157616 274320 157668 274372
rect 159272 274320 159324 274372
rect 202328 274320 202380 274372
rect 223120 274320 223172 274372
rect 247224 274320 247276 274372
rect 369124 274320 369176 274372
rect 387340 274320 387392 274372
rect 419080 274320 419132 274372
rect 467748 274320 467800 274372
rect 506204 274320 506256 274372
rect 591856 274320 591908 274372
rect 331956 274252 332008 274304
rect 337752 274252 337804 274304
rect 67088 274184 67140 274236
rect 130384 274184 130436 274236
rect 130844 274184 130896 274236
rect 182456 274184 182508 274236
rect 192392 274184 192444 274236
rect 224960 274184 225012 274236
rect 240048 274184 240100 274236
rect 253940 274184 253992 274236
rect 359464 274184 359516 274236
rect 380256 274184 380308 274236
rect 388996 274184 389048 274236
rect 425152 274184 425204 274236
rect 425704 274184 425756 274236
rect 474832 274184 474884 274236
rect 511816 274184 511868 274236
rect 598940 274184 598992 274236
rect 77668 274048 77720 274100
rect 144920 274048 144972 274100
rect 154488 274048 154540 274100
rect 198096 274048 198148 274100
rect 210056 274048 210108 274100
rect 237840 274048 237892 274100
rect 249064 274048 249116 274100
rect 265256 274048 265308 274100
rect 266360 274048 266412 274100
rect 273536 274048 273588 274100
rect 278596 274048 278648 274100
rect 285864 274048 285916 274100
rect 337752 274048 337804 274100
rect 351920 274048 351972 274100
rect 353944 274048 353996 274100
rect 369584 274048 369636 274100
rect 373264 274048 373316 274100
rect 400312 274048 400364 274100
rect 401508 274048 401560 274100
rect 442908 274048 442960 274100
rect 451188 274048 451240 274100
rect 513840 274048 513892 274100
rect 536748 274048 536800 274100
rect 634360 274048 634412 274100
rect 69388 273912 69440 273964
rect 139400 273912 139452 273964
rect 148600 273912 148652 273964
rect 194784 273912 194836 273964
rect 208860 273912 208912 273964
rect 237472 273912 237524 273964
rect 238484 273912 238536 273964
rect 88340 273776 88392 273828
rect 119344 273776 119396 273828
rect 120264 273776 120316 273828
rect 175280 273776 175332 273828
rect 193496 273776 193548 273828
rect 226432 273776 226484 273828
rect 271512 273912 271564 273964
rect 280344 273912 280396 273964
rect 322756 273912 322808 273964
rect 330576 273912 330628 273964
rect 335268 273912 335320 273964
rect 348332 273912 348384 273964
rect 350356 273912 350408 273964
rect 368480 273912 368532 273964
rect 377680 273912 377732 273964
rect 408592 273912 408644 273964
rect 422116 273912 422168 273964
rect 472440 273912 472492 273964
rect 474648 273912 474700 273964
rect 545764 273912 545816 273964
rect 545948 273912 546000 273964
rect 639144 273912 639196 273964
rect 258080 273776 258132 273828
rect 397000 273776 397052 273828
rect 435824 273776 435876 273828
rect 438124 273776 438176 273828
rect 473636 273776 473688 273828
rect 481364 273776 481416 273828
rect 556344 273776 556396 273828
rect 556804 273776 556856 273828
rect 590660 273776 590712 273828
rect 119068 273640 119120 273692
rect 173256 273640 173308 273692
rect 447784 273640 447836 273692
rect 481916 273640 481968 273692
rect 484216 273640 484268 273692
rect 559932 273640 559984 273692
rect 132040 273504 132092 273556
rect 153844 273504 153896 273556
rect 259368 273504 259420 273556
rect 266360 273504 266412 273556
rect 440884 273504 440936 273556
rect 471244 273504 471296 273556
rect 478696 273504 478748 273556
rect 552848 273504 552900 273556
rect 145288 273368 145340 273420
rect 147864 273368 147916 273420
rect 476028 273368 476080 273420
rect 549260 273368 549312 273420
rect 549904 273368 549956 273420
rect 583576 273368 583628 273420
rect 460020 273300 460072 273352
rect 461400 273300 461452 273352
rect 327724 273232 327776 273284
rect 329472 273232 329524 273284
rect 42432 273164 42484 273216
rect 42984 273164 43036 273216
rect 108396 273164 108448 273216
rect 165896 273164 165948 273216
rect 186412 273164 186464 273216
rect 218704 273164 218756 273216
rect 362776 273164 362828 273216
rect 385868 273164 385920 273216
rect 400036 273164 400088 273216
rect 439320 273164 439372 273216
rect 444012 273164 444064 273216
rect 503168 273164 503220 273216
rect 504180 273164 504232 273216
rect 511448 273164 511500 273216
rect 515404 273164 515456 273216
rect 519728 273164 519780 273216
rect 521476 273164 521528 273216
rect 614304 273164 614356 273216
rect 102508 273028 102560 273080
rect 162860 273028 162912 273080
rect 172244 273028 172296 273080
rect 209780 273028 209832 273080
rect 219532 273028 219584 273080
rect 244556 273028 244608 273080
rect 280988 273028 281040 273080
rect 286324 273028 286376 273080
rect 361212 273028 361264 273080
rect 384948 273028 385000 273080
rect 385684 273028 385736 273080
rect 395620 273028 395672 273080
rect 404176 273028 404228 273080
rect 446496 273028 446548 273080
rect 446864 273028 446916 273080
rect 507952 273028 508004 273080
rect 94228 272892 94280 272944
rect 155960 272892 156012 272944
rect 166356 272892 166408 272944
rect 207296 272892 207348 272944
rect 211252 272892 211304 272944
rect 220084 272892 220136 272944
rect 220728 272892 220780 272944
rect 245752 272892 245804 272944
rect 247868 272892 247920 272944
rect 264244 272892 264296 272944
rect 333796 272892 333848 272944
rect 345940 272892 345992 272944
rect 348424 272892 348476 272944
rect 362500 272892 362552 272944
rect 365444 272892 365496 272944
rect 390928 272892 390980 272944
rect 405556 272892 405608 272944
rect 448796 272892 448848 272944
rect 455328 272892 455380 272944
rect 457260 272892 457312 272944
rect 457996 272892 458048 272944
rect 465908 272892 465960 272944
rect 466092 272892 466144 272944
rect 518532 273028 518584 273080
rect 518716 273028 518768 273080
rect 569408 273028 569460 273080
rect 82452 272756 82504 272808
rect 148416 272756 148468 272808
rect 155684 272756 155736 272808
rect 200120 272756 200172 272808
rect 205364 272756 205416 272808
rect 234804 272756 234856 272808
rect 245384 272756 245436 272808
rect 72976 272620 73028 272672
rect 142160 272620 142212 272672
rect 142712 272620 142764 272672
rect 145564 272620 145616 272672
rect 147404 272620 147456 272672
rect 193220 272620 193272 272672
rect 197084 272620 197136 272672
rect 229100 272620 229152 272672
rect 233700 272620 233752 272672
rect 254400 272620 254452 272672
rect 262312 272756 262364 272808
rect 270960 272756 271012 272808
rect 273904 272756 273956 272808
rect 282920 272756 282972 272808
rect 325332 272756 325384 272808
rect 332968 272756 333020 272808
rect 344652 272756 344704 272808
rect 361396 272756 361448 272808
rect 362224 272756 362276 272808
rect 370320 272756 370372 272808
rect 370504 272756 370556 272808
rect 396816 272756 396868 272808
rect 406844 272756 406896 272808
rect 449992 272756 450044 272808
rect 452292 272756 452344 272808
rect 515036 272892 515088 272944
rect 532516 272892 532568 272944
rect 513748 272756 513800 272808
rect 525616 272756 525668 272808
rect 529848 272756 529900 272808
rect 532884 272756 532936 272808
rect 533712 272756 533764 272808
rect 538680 272756 538732 272808
rect 539048 272892 539100 272944
rect 624976 272892 625028 272944
rect 628472 272756 628524 272808
rect 262680 272620 262732 272672
rect 264428 272620 264480 272672
rect 276020 272620 276072 272672
rect 324044 272620 324096 272672
rect 331772 272620 331824 272672
rect 332324 272620 332376 272672
rect 343640 272620 343692 272672
rect 346216 272620 346268 272672
rect 363696 272620 363748 272672
rect 376116 272620 376168 272672
rect 406292 272620 406344 272672
rect 412272 272620 412324 272672
rect 457076 272620 457128 272672
rect 457260 272620 457312 272672
rect 460020 272620 460072 272672
rect 460204 272620 460256 272672
rect 319076 272552 319128 272604
rect 319628 272552 319680 272604
rect 65892 272484 65944 272536
rect 136824 272484 136876 272536
rect 137928 272484 137980 272536
rect 116676 272348 116728 272400
rect 172520 272348 172572 272400
rect 181720 272484 181772 272536
rect 186964 272484 187016 272536
rect 195888 272484 195940 272536
rect 227904 272484 227956 272536
rect 228088 272484 228140 272536
rect 249064 272484 249116 272536
rect 254952 272484 255004 272536
rect 269304 272484 269356 272536
rect 270316 272484 270368 272536
rect 280528 272484 280580 272536
rect 329748 272484 329800 272536
rect 338856 272484 338908 272536
rect 339224 272484 339276 272536
rect 354220 272484 354272 272536
rect 354496 272484 354548 272536
rect 375564 272484 375616 272536
rect 379428 272484 379480 272536
rect 410984 272484 411036 272536
rect 416596 272484 416648 272536
rect 460848 272484 460900 272536
rect 461400 272484 461452 272536
rect 465540 272484 465592 272536
rect 465908 272620 465960 272672
rect 522120 272620 522172 272672
rect 526812 272620 526864 272672
rect 621388 272620 621440 272672
rect 470554 272484 470606 272536
rect 470692 272484 470744 272536
rect 532700 272484 532752 272536
rect 532884 272484 532936 272536
rect 538496 272484 538548 272536
rect 538680 272484 538732 272536
rect 632060 272892 632112 272944
rect 318708 272416 318760 272468
rect 324688 272416 324740 272468
rect 187700 272348 187752 272400
rect 194968 272348 195020 272400
rect 227168 272348 227220 272400
rect 395988 272348 396040 272400
rect 434628 272348 434680 272400
rect 449716 272348 449768 272400
rect 504180 272348 504232 272400
rect 504364 272348 504416 272400
rect 513748 272348 513800 272400
rect 517428 272348 517480 272400
rect 600780 272348 600832 272400
rect 600964 272348 601016 272400
rect 635556 272756 635608 272808
rect 634084 272620 634136 272672
rect 640340 272620 640392 272672
rect 127348 272212 127400 272264
rect 179880 272212 179932 272264
rect 189080 272212 189132 272264
rect 196440 272212 196492 272264
rect 391848 272212 391900 272264
rect 428740 272212 428792 272264
rect 450544 272212 450596 272264
rect 510252 272212 510304 272264
rect 510436 272212 510488 272264
rect 518716 272212 518768 272264
rect 520096 272212 520148 272264
rect 610716 272212 610768 272264
rect 145104 272076 145156 272128
rect 192392 272076 192444 272128
rect 384948 272076 385000 272128
rect 418068 272076 418120 272128
rect 428464 272076 428516 272128
rect 470554 272076 470606 272128
rect 470784 272076 470836 272128
rect 124956 271940 125008 271992
rect 151084 271940 151136 271992
rect 431684 271940 431736 271992
rect 106004 271804 106056 271856
rect 164976 271804 165028 271856
rect 174268 271804 174320 271856
rect 189172 271804 189224 271856
rect 202972 271804 203024 271856
rect 233240 271804 233292 271856
rect 274640 271804 274692 271856
rect 279240 271804 279292 271856
rect 355324 271804 355376 271856
rect 356612 271804 356664 271856
rect 375288 271804 375340 271856
rect 403900 271804 403952 271856
rect 433156 271804 433208 271856
rect 480168 271804 480220 271856
rect 480536 271940 480588 271992
rect 485044 271940 485096 271992
rect 485412 272076 485464 272128
rect 547512 272076 547564 272128
rect 547696 272076 547748 272128
rect 504364 271940 504416 271992
rect 504548 271940 504600 271992
rect 562324 271940 562376 271992
rect 600780 272076 600832 272128
rect 607220 272076 607272 272128
rect 600964 271940 601016 271992
rect 484676 271804 484728 271856
rect 494704 271804 494756 271856
rect 501420 271804 501472 271856
rect 504364 271804 504416 271856
rect 578516 271804 578568 271856
rect 578884 271804 578936 271856
rect 604828 271804 604880 271856
rect 97816 271668 97868 271720
rect 158812 271668 158864 271720
rect 169852 271668 169904 271720
rect 209964 271668 210016 271720
rect 225420 271668 225472 271720
rect 228364 271668 228416 271720
rect 351184 271668 351236 271720
rect 366088 271668 366140 271720
rect 382004 271668 382056 271720
rect 414572 271668 414624 271720
rect 87144 271532 87196 271584
rect 152004 271532 152056 271584
rect 165160 271532 165212 271584
rect 205640 271532 205692 271584
rect 215944 271532 215996 271584
rect 242072 271532 242124 271584
rect 337936 271532 337988 271584
rect 350724 271532 350776 271584
rect 360844 271532 360896 271584
rect 377864 271532 377916 271584
rect 387708 271532 387760 271584
rect 421656 271668 421708 271720
rect 430396 271668 430448 271720
rect 483204 271668 483256 271720
rect 499304 271668 499356 271720
rect 582380 271668 582432 271720
rect 583024 271668 583076 271720
rect 611912 271668 611964 271720
rect 420184 271532 420236 271584
rect 431132 271532 431184 271584
rect 437204 271532 437256 271584
rect 493692 271532 493744 271584
rect 75368 271396 75420 271448
rect 142712 271396 142764 271448
rect 162676 271396 162728 271448
rect 204720 271396 204772 271448
rect 213644 271396 213696 271448
rect 240416 271396 240468 271448
rect 240784 271396 240836 271448
rect 259644 271396 259696 271448
rect 259828 271396 259880 271448
rect 272616 271396 272668 271448
rect 325516 271396 325568 271448
rect 334164 271396 334216 271448
rect 347688 271396 347740 271448
rect 364892 271396 364944 271448
rect 366364 271396 366416 271448
rect 383844 271396 383896 271448
rect 384764 271396 384816 271448
rect 419264 271396 419316 271448
rect 76840 271260 76892 271312
rect 143540 271260 143592 271312
rect 152188 271260 152240 271312
rect 197360 271260 197412 271312
rect 198280 271260 198332 271312
rect 229560 271260 229612 271312
rect 235264 271260 235316 271312
rect 255320 271260 255372 271312
rect 256700 271260 256752 271312
rect 261024 271260 261076 271312
rect 262036 271260 262088 271312
rect 274640 271260 274692 271312
rect 329564 271260 329616 271312
rect 340052 271260 340104 271312
rect 340604 271260 340656 271312
rect 355140 271260 355192 271312
rect 357164 271260 357216 271312
rect 379060 271260 379112 271312
rect 390284 271260 390336 271312
rect 426348 271396 426400 271448
rect 439964 271396 440016 271448
rect 497280 271532 497332 271584
rect 501972 271532 502024 271584
rect 585968 271532 586020 271584
rect 612004 271532 612056 271584
rect 618996 271532 619048 271584
rect 496544 271396 496596 271448
rect 504364 271396 504416 271448
rect 505008 271396 505060 271448
rect 589464 271396 589516 271448
rect 589924 271396 589976 271448
rect 633256 271396 633308 271448
rect 68192 271124 68244 271176
rect 138480 271124 138532 271176
rect 141516 271124 141568 271176
rect 189816 271124 189868 271176
rect 191196 271124 191248 271176
rect 225144 271124 225196 271176
rect 230204 271124 230256 271176
rect 252008 271124 252060 271176
rect 268016 271124 268068 271176
rect 278780 271124 278832 271176
rect 279792 271124 279844 271176
rect 287060 271124 287112 271176
rect 331128 271124 331180 271176
rect 342444 271124 342496 271176
rect 343548 271124 343600 271176
rect 360200 271124 360252 271176
rect 364156 271124 364208 271176
rect 389732 271124 389784 271176
rect 394332 271124 394384 271176
rect 432236 271260 432288 271312
rect 442908 271260 442960 271312
rect 500868 271260 500920 271312
rect 507676 271260 507728 271312
rect 593052 271260 593104 271312
rect 598204 271260 598256 271312
rect 645032 271260 645084 271312
rect 113456 270988 113508 271040
rect 169944 270988 169996 271040
rect 187424 270988 187476 271040
rect 215944 270988 215996 271040
rect 251456 270988 251508 271040
rect 266912 270988 266964 271040
rect 417424 270988 417476 271040
rect 437940 271124 437992 271176
rect 441344 271124 441396 271176
rect 445024 271124 445076 271176
rect 445668 271124 445720 271176
rect 503996 271124 504048 271176
rect 524052 271124 524104 271176
rect 617340 271124 617392 271176
rect 617524 271124 617576 271176
rect 626080 271124 626132 271176
rect 427452 270988 427504 271040
rect 479156 270988 479208 271040
rect 485044 270988 485096 271040
rect 494704 270988 494756 271040
rect 495072 270988 495124 271040
rect 575296 270988 575348 271040
rect 123760 270852 123812 270904
rect 177488 270852 177540 270904
rect 407764 270852 407816 270904
rect 440516 270852 440568 270904
rect 449164 270852 449216 270904
rect 490196 270852 490248 270904
rect 492588 270852 492640 270904
rect 571708 270852 571760 270904
rect 134432 270716 134484 270768
rect 185124 270716 185176 270768
rect 321376 270716 321428 270768
rect 327080 270716 327132 270768
rect 414664 270716 414716 270768
rect 450820 270716 450872 270768
rect 480260 270716 480312 270768
rect 486608 270716 486660 270768
rect 486976 270716 487028 270768
rect 564624 270716 564676 270768
rect 567844 270716 567896 270768
rect 597744 270716 597796 270768
rect 121460 270580 121512 270632
rect 168104 270580 168156 270632
rect 403624 270580 403676 270632
rect 433432 270580 433484 270632
rect 453304 270580 453356 270632
rect 487804 270580 487856 270632
rect 489644 270580 489696 270632
rect 568212 270580 568264 270632
rect 84108 270444 84160 270496
rect 137468 270444 137520 270496
rect 137652 270444 137704 270496
rect 186136 270444 186188 270496
rect 201040 270444 201092 270496
rect 201868 270444 201920 270496
rect 206836 270444 206888 270496
rect 235816 270444 235868 270496
rect 278044 270444 278096 270496
rect 283840 270444 283892 270496
rect 400864 270444 400916 270496
rect 441620 270444 441672 270496
rect 456432 270444 456484 270496
rect 520280 270444 520332 270496
rect 523132 270444 523184 270496
rect 532792 270444 532844 270496
rect 619640 270444 619692 270496
rect 78864 270308 78916 270360
rect 132500 270308 132552 270360
rect 133788 270308 133840 270360
rect 183652 270308 183704 270360
rect 185308 270308 185360 270360
rect 194416 270308 194468 270360
rect 199936 270308 199988 270360
rect 230848 270308 230900 270360
rect 232688 270308 232740 270360
rect 248236 270308 248288 270360
rect 283104 270308 283156 270360
rect 284668 270308 284720 270360
rect 355048 270308 355100 270360
rect 376760 270308 376812 270360
rect 380532 270308 380584 270360
rect 404360 270308 404412 270360
rect 415032 270308 415084 270360
rect 461216 270308 461268 270360
rect 461400 270308 461452 270360
rect 111984 270172 112036 270224
rect 168748 270172 168800 270224
rect 184848 270172 184900 270224
rect 219348 270172 219400 270224
rect 244372 270172 244424 270224
rect 262312 270172 262364 270224
rect 334348 270172 334400 270224
rect 346400 270172 346452 270224
rect 372252 270172 372304 270224
rect 397460 270172 397512 270224
rect 409604 270172 409656 270224
rect 454040 270172 454092 270224
rect 458824 270172 458876 270224
rect 524420 270172 524472 270224
rect 525616 270308 525668 270360
rect 533528 270308 533580 270360
rect 626540 270308 626592 270360
rect 527180 270172 527232 270224
rect 528376 270172 528428 270224
rect 533252 270172 533304 270224
rect 533528 270172 533580 270224
rect 623964 270172 624016 270224
rect 89628 270036 89680 270088
rect 153016 270036 153068 270088
rect 176568 270036 176620 270088
rect 211160 270036 211212 270088
rect 212448 270036 212500 270088
rect 239956 270036 240008 270088
rect 241888 270036 241940 270088
rect 260656 270036 260708 270088
rect 266176 270036 266228 270088
rect 277216 270036 277268 270088
rect 345296 270036 345348 270088
rect 358820 270036 358872 270088
rect 366640 270036 366692 270088
rect 393320 270036 393372 270088
rect 394700 270036 394752 270088
rect 408776 270036 408828 270088
rect 412456 270036 412508 270088
rect 458180 270036 458232 270088
rect 463516 270036 463568 270088
rect 530768 270036 530820 270088
rect 530952 270036 531004 270088
rect 532976 270036 533028 270088
rect 85488 269900 85540 269952
rect 149428 269900 149480 269952
rect 152832 269900 152884 269952
rect 157156 269900 157208 269952
rect 173808 269900 173860 269952
rect 212632 269900 212684 269952
rect 226616 269900 226668 269952
rect 249892 269900 249944 269952
rect 256884 269900 256936 269952
rect 268936 269900 268988 269952
rect 330208 269900 330260 269952
rect 340880 269900 340932 269952
rect 341800 269900 341852 269952
rect 357440 269900 357492 269952
rect 359188 269900 359240 269952
rect 382280 269900 382332 269952
rect 383016 269900 383068 269952
rect 411260 269900 411312 269952
rect 419632 269900 419684 269952
rect 468024 269900 468076 269952
rect 468484 269900 468536 269952
rect 538312 270036 538364 270088
rect 533988 269900 534040 269952
rect 630680 270036 630732 270088
rect 539048 269900 539100 269952
rect 541532 269900 541584 269952
rect 70584 269764 70636 269816
rect 79324 269764 79376 269816
rect 80060 269764 80112 269816
rect 146392 269764 146444 269816
rect 158628 269764 158680 269816
rect 201040 269764 201092 269816
rect 201684 269764 201736 269816
rect 232504 269764 232556 269816
rect 237288 269764 237340 269816
rect 257344 269764 257396 269816
rect 258540 269764 258592 269816
rect 272248 269764 272300 269816
rect 273076 269764 273128 269816
rect 282184 269764 282236 269816
rect 326896 269764 326948 269816
rect 335544 269764 335596 269816
rect 336004 269764 336056 269816
rect 349160 269764 349212 269816
rect 351736 269764 351788 269816
rect 371240 269764 371292 269816
rect 376576 269764 376628 269816
rect 407120 269764 407172 269816
rect 417148 269764 417200 269816
rect 465080 269764 465132 269816
rect 466000 269764 466052 269816
rect 532240 269764 532292 269816
rect 122748 269628 122800 269680
rect 176200 269628 176252 269680
rect 183468 269628 183520 269680
rect 205456 269628 205508 269680
rect 392032 269628 392084 269680
rect 401692 269628 401744 269680
rect 404360 269628 404412 269680
rect 423680 269628 423732 269680
rect 423956 269628 424008 269680
rect 451372 269628 451424 269680
rect 453580 269628 453632 269680
rect 509240 269628 509292 269680
rect 538864 269764 538916 269816
rect 540520 269764 540572 269816
rect 640524 269900 640576 269952
rect 542452 269764 542504 269816
rect 637672 269764 637724 269816
rect 129648 269492 129700 269544
rect 181168 269492 181220 269544
rect 204168 269492 204220 269544
rect 223488 269492 223540 269544
rect 398748 269492 398800 269544
rect 412640 269492 412692 269544
rect 424600 269492 424652 269544
rect 475016 269492 475068 269544
rect 495256 269492 495308 269544
rect 532792 269628 532844 269680
rect 616420 269628 616472 269680
rect 509884 269492 509936 269544
rect 596180 269492 596232 269544
rect 126888 269356 126940 269408
rect 178316 269356 178368 269408
rect 408316 269356 408368 269408
rect 426532 269356 426584 269408
rect 441620 269356 441672 269408
rect 458456 269356 458508 269408
rect 470968 269356 471020 269408
rect 538680 269356 538732 269408
rect 538864 269356 538916 269408
rect 575480 269356 575532 269408
rect 143908 269220 143960 269272
rect 191104 269220 191156 269272
rect 282736 269220 282788 269272
rect 288808 269220 288860 269272
rect 401692 269220 401744 269272
rect 416780 269220 416832 269272
rect 474280 269220 474332 269272
rect 546500 269220 546552 269272
rect 319444 269084 319496 269136
rect 325700 269084 325752 269136
rect 118608 269016 118660 269068
rect 174544 269016 174596 269068
rect 175096 269016 175148 269068
rect 177672 269016 177724 269068
rect 273260 269016 273312 269068
rect 275560 269016 275612 269068
rect 436560 269016 436612 269068
rect 491668 269016 491720 269068
rect 495808 269016 495860 269068
rect 576860 269016 576912 269068
rect 115848 268880 115900 268932
rect 171232 268880 171284 268932
rect 382372 268880 382424 268932
rect 415400 268880 415452 268932
rect 433708 268880 433760 268932
rect 488540 268880 488592 268932
rect 498292 268880 498344 268932
rect 581000 268880 581052 268932
rect 110328 268744 110380 268796
rect 167920 268744 167972 268796
rect 168288 268744 168340 268796
rect 181996 268744 182048 268796
rect 188896 268744 188948 268796
rect 190460 268744 190512 268796
rect 200580 268744 200632 268796
rect 231308 268744 231360 268796
rect 387340 268744 387392 268796
rect 422300 268744 422352 268796
rect 438676 268744 438728 268796
rect 495440 268744 495492 268796
rect 500776 268744 500828 268796
rect 583760 268744 583812 268796
rect 104992 268608 105044 268660
rect 163780 268608 163832 268660
rect 176936 268608 176988 268660
rect 215116 268608 215168 268660
rect 224224 268608 224276 268660
rect 243268 268608 243320 268660
rect 352564 268608 352616 268660
rect 372620 268608 372672 268660
rect 393688 268608 393740 268660
rect 429200 268608 429252 268660
rect 441160 268608 441212 268660
rect 499580 268608 499632 268660
rect 503260 268608 503312 268660
rect 587900 268608 587952 268660
rect 99288 268472 99340 268524
rect 160468 268472 160520 268524
rect 180708 268472 180760 268524
rect 217600 268472 217652 268524
rect 231676 268472 231728 268524
rect 253204 268472 253256 268524
rect 338488 268472 338540 268524
rect 352104 268472 352156 268524
rect 367468 268472 367520 268524
rect 393504 268472 393556 268524
rect 397276 268472 397328 268524
rect 436100 268472 436152 268524
rect 446128 268472 446180 268524
rect 506480 268472 506532 268524
rect 508228 268472 508280 268524
rect 594800 268472 594852 268524
rect 92388 268336 92440 268388
rect 155500 268336 155552 268388
rect 161572 268336 161624 268388
rect 203524 268336 203576 268388
rect 210700 268336 210752 268388
rect 236644 268336 236696 268388
rect 252652 268336 252704 268388
rect 268108 268336 268160 268388
rect 348792 268336 348844 268388
rect 367100 268336 367152 268388
rect 372436 268336 372488 268388
rect 400496 268336 400548 268388
rect 402244 268336 402296 268388
rect 443092 268336 443144 268388
rect 461860 268336 461912 268388
rect 528560 268336 528612 268388
rect 541348 268336 541400 268388
rect 641720 268336 641772 268388
rect 135628 268200 135680 268252
rect 140688 268200 140740 268252
rect 140872 268200 140924 268252
rect 188620 268200 188672 268252
rect 416228 268200 416280 268252
rect 447140 268200 447192 268252
rect 493324 268200 493376 268252
rect 574100 268200 574152 268252
rect 151728 268064 151780 268116
rect 196072 268064 196124 268116
rect 422300 268064 422352 268116
rect 444380 268064 444432 268116
rect 448428 268064 448480 268116
rect 494060 268064 494112 268116
rect 527180 268064 527232 268116
rect 607404 268064 607456 268116
rect 490840 267928 490892 267980
rect 569960 267928 570012 267980
rect 276480 267724 276532 267776
rect 278044 267724 278096 267776
rect 119344 267656 119396 267708
rect 153476 267656 153528 267708
rect 111708 267520 111760 267572
rect 169576 267656 169628 267708
rect 178684 267656 178736 267708
rect 209320 267656 209372 267708
rect 390652 267656 390704 267708
rect 408316 267656 408368 267708
rect 422944 267656 422996 267708
rect 438124 267656 438176 267708
rect 445300 267656 445352 267708
rect 490564 267656 490616 267708
rect 509884 267656 509936 267708
rect 567844 267656 567896 267708
rect 169024 267520 169076 267572
rect 199384 267520 199436 267572
rect 215944 267520 215996 267572
rect 222568 267520 222620 267572
rect 362500 267520 362552 267572
rect 369124 267520 369176 267572
rect 380716 267520 380768 267572
rect 398748 267520 398800 267572
rect 404728 267520 404780 267572
rect 416228 267520 416280 267572
rect 421288 267520 421340 267572
rect 440884 267520 440936 267572
rect 450268 267520 450320 267572
rect 498844 267520 498896 267572
rect 514852 267520 514904 267572
rect 578884 267520 578936 267572
rect 86224 267384 86276 267436
rect 144736 267384 144788 267436
rect 145564 267384 145616 267436
rect 191932 267384 191984 267436
rect 199568 267384 199620 267436
rect 204352 267384 204404 267436
rect 205456 267384 205508 267436
rect 218428 267384 218480 267436
rect 233884 267384 233936 267436
rect 104808 267248 104860 267300
rect 164608 267248 164660 267300
rect 186964 267248 187016 267300
rect 219256 267248 219308 267300
rect 223488 267248 223540 267300
rect 234160 267248 234212 267300
rect 243728 267384 243780 267436
rect 251548 267384 251600 267436
rect 315304 267384 315356 267436
rect 319076 267384 319128 267436
rect 340972 267384 341024 267436
rect 355324 267384 355376 267436
rect 365812 267384 365864 267436
rect 381544 267384 381596 267436
rect 383200 267384 383252 267436
rect 401692 267384 401744 267436
rect 403072 267384 403124 267436
rect 422300 267384 422352 267436
rect 428740 267384 428792 267436
rect 447784 267384 447836 267436
rect 460480 267384 460532 267436
rect 516784 267384 516836 267436
rect 519820 267384 519872 267436
rect 583024 267384 583076 267436
rect 244096 267248 244148 267300
rect 321928 267248 321980 267300
rect 327724 267248 327776 267300
rect 350908 267248 350960 267300
rect 362224 267248 362276 267300
rect 90364 267112 90416 267164
rect 151360 267112 151412 267164
rect 159456 267112 159508 267164
rect 162124 267112 162176 267164
rect 168104 267112 168156 267164
rect 177028 267112 177080 267164
rect 177672 267112 177724 267164
rect 214288 267112 214340 267164
rect 220084 267112 220136 267164
rect 239128 267112 239180 267164
rect 246948 267112 247000 267164
rect 263968 267112 264020 267164
rect 314476 267112 314528 267164
rect 319260 267112 319312 267164
rect 360016 267112 360068 267164
rect 366364 267112 366416 267164
rect 79324 266976 79376 267028
rect 140228 266976 140280 267028
rect 140688 266976 140740 267028
rect 186964 266976 187016 267028
rect 190460 266976 190512 267028
rect 224224 266976 224276 267028
rect 228364 266976 228416 267028
rect 248788 266976 248840 267028
rect 255964 266976 256016 267028
rect 259000 266976 259052 267028
rect 286324 266976 286376 267028
rect 287980 266976 288032 267028
rect 313648 266976 313700 267028
rect 317420 266976 317472 267028
rect 353392 266976 353444 267028
rect 374460 267248 374512 267300
rect 378784 267248 378836 267300
rect 385684 267248 385736 267300
rect 398104 267248 398156 267300
rect 417424 267248 417476 267300
rect 432880 267248 432932 267300
rect 453304 267248 453356 267300
rect 373632 267112 373684 267164
rect 392032 267112 392084 267164
rect 399760 267112 399812 267164
rect 407764 267112 407816 267164
rect 413008 267112 413060 267164
rect 441620 267112 441672 267164
rect 447140 267112 447192 267164
rect 448428 267112 448480 267164
rect 452752 267112 452804 267164
rect 462964 267248 463016 267300
rect 465172 267248 465224 267300
rect 523684 267248 523736 267300
rect 524788 267248 524840 267300
rect 612004 267248 612056 267300
rect 455144 267112 455196 267164
rect 515404 267112 515456 267164
rect 517244 267112 517296 267164
rect 527180 267112 527232 267164
rect 529664 267112 529716 267164
rect 617524 267112 617576 267164
rect 393136 266976 393188 267028
rect 420184 266976 420236 267028
rect 132500 266840 132552 266892
rect 147220 266840 147272 266892
rect 153844 266840 153896 266892
rect 184480 266840 184532 266892
rect 218704 266840 218756 266892
rect 220912 266840 220964 266892
rect 312820 266840 312872 266892
rect 316040 266840 316092 266892
rect 332692 266840 332744 266892
rect 343824 266840 343876 266892
rect 374920 266840 374972 266892
rect 380532 266840 380584 266892
rect 388168 266840 388220 266892
rect 317788 266772 317840 266824
rect 322940 266772 322992 266824
rect 137468 266704 137520 266756
rect 150532 266704 150584 266756
rect 151084 266704 151136 266756
rect 179512 266704 179564 266756
rect 368296 266704 368348 266756
rect 378784 266704 378836 266756
rect 308680 266636 308732 266688
rect 310612 266636 310664 266688
rect 316960 266636 317012 266688
rect 321560 266636 321612 266688
rect 347504 266636 347556 266688
rect 351184 266636 351236 266688
rect 130384 266568 130436 266620
rect 138112 266568 138164 266620
rect 149612 266568 149664 266620
rect 159640 266568 159692 266620
rect 378232 266568 378284 266620
rect 394700 266704 394752 266756
rect 427912 266840 427964 266892
rect 457444 266976 457496 267028
rect 470140 266976 470192 267028
rect 534724 266976 534776 267028
rect 535552 266976 535604 267028
rect 536748 266976 536800 267028
rect 539692 266976 539744 267028
rect 634084 266976 634136 267028
rect 442724 266840 442776 266892
rect 485044 266840 485096 266892
rect 499948 266840 500000 266892
rect 507860 266840 507912 266892
rect 534724 266840 534776 266892
rect 589924 266840 589976 266892
rect 404360 266704 404412 266756
rect 408040 266704 408092 266756
rect 423956 266704 424008 266756
rect 434536 266704 434588 266756
rect 449164 266704 449216 266756
rect 457720 266704 457772 266756
rect 476764 266704 476816 266756
rect 485044 266704 485096 266756
rect 394792 266568 394844 266620
rect 403624 266568 403676 266620
rect 407212 266568 407264 266620
rect 414664 266568 414716 266620
rect 437848 266568 437900 266620
rect 447140 266568 447192 266620
rect 490012 266704 490064 266756
rect 509700 266704 509752 266756
rect 510712 266704 510764 266756
rect 511816 266704 511868 266756
rect 512368 266704 512420 266756
rect 513196 266704 513248 266756
rect 516508 266704 516560 266756
rect 517428 266704 517480 266756
rect 518992 266704 519044 266756
rect 520096 266704 520148 266756
rect 527272 266704 527324 266756
rect 528192 266704 528244 266756
rect 528928 266704 528980 266756
rect 529848 266704 529900 266756
rect 531412 266704 531464 266756
rect 532608 266704 532660 266756
rect 533068 266704 533120 266756
rect 533988 266704 534040 266756
rect 543004 266704 543056 266756
rect 598204 266704 598256 266756
rect 501604 266568 501656 266620
rect 504824 266568 504876 266620
rect 556804 266568 556856 266620
rect 250444 266500 250496 266552
rect 256516 266500 256568 266552
rect 310336 266500 310388 266552
rect 311900 266500 311952 266552
rect 312360 266500 312412 266552
rect 314660 266500 314712 266552
rect 316132 266500 316184 266552
rect 320180 266500 320232 266552
rect 327724 266500 327776 266552
rect 331956 266500 332008 266552
rect 345112 266500 345164 266552
rect 348424 266500 348476 266552
rect 350080 266500 350132 266552
rect 353944 266500 353996 266552
rect 355876 266500 355928 266552
rect 360844 266500 360896 266552
rect 369952 266500 370004 266552
rect 372252 266500 372304 266552
rect 423772 266500 423824 266552
rect 425704 266500 425756 266552
rect 426256 266500 426308 266552
rect 428464 266500 428516 266552
rect 447784 266500 447836 266552
rect 456064 266500 456116 266552
rect 491668 266432 491720 266484
rect 492588 266432 492640 266484
rect 494152 266432 494204 266484
rect 495072 266432 495124 266484
rect 502432 266432 502484 266484
rect 503444 266432 503496 266484
rect 504088 266432 504140 266484
rect 505008 266432 505060 266484
rect 506572 266432 506624 266484
rect 507676 266432 507728 266484
rect 507860 266432 507912 266484
rect 549904 266432 549956 266484
rect 163504 266364 163556 266416
rect 167092 266364 167144 266416
rect 211160 266364 211212 266416
rect 213460 266364 213512 266416
rect 214564 266364 214616 266416
rect 215944 266364 215996 266416
rect 239404 266364 239456 266416
rect 241612 266364 241664 266416
rect 243544 266364 243596 266416
rect 246580 266364 246632 266416
rect 249064 266364 249116 266416
rect 250720 266364 250772 266416
rect 300952 266364 301004 266416
rect 302056 266364 302108 266416
rect 303712 266364 303764 266416
rect 304540 266364 304592 266416
rect 307852 266364 307904 266416
rect 309140 266364 309192 266416
rect 309508 266364 309560 266416
rect 310796 266364 310848 266416
rect 311164 266364 311216 266416
rect 313280 266364 313332 266416
rect 320272 266364 320324 266416
rect 321376 266364 321428 266416
rect 324412 266364 324464 266416
rect 325332 266364 325384 266416
rect 328552 266364 328604 266416
rect 329748 266364 329800 266416
rect 336832 266364 336884 266416
rect 337936 266364 337988 266416
rect 342628 266364 342680 266416
rect 345296 266364 345348 266416
rect 346768 266364 346820 266416
rect 347688 266364 347740 266416
rect 349252 266364 349304 266416
rect 350356 266364 350408 266416
rect 357532 266364 357584 266416
rect 359464 266364 359516 266416
rect 361672 266364 361724 266416
rect 362776 266364 362828 266416
rect 369124 266364 369176 266416
rect 370504 266364 370556 266416
rect 371608 266364 371660 266416
rect 373264 266364 373316 266416
rect 374092 266364 374144 266416
rect 375288 266364 375340 266416
rect 379888 266364 379940 266416
rect 383016 266364 383068 266416
rect 384028 266364 384080 266416
rect 384948 266364 385000 266416
rect 386512 266364 386564 266416
rect 387708 266364 387760 266416
rect 392308 266364 392360 266416
rect 393688 266364 393740 266416
rect 398932 266364 398984 266416
rect 400036 266364 400088 266416
rect 408868 266364 408920 266416
rect 409788 266364 409840 266416
rect 411352 266364 411404 266416
rect 412272 266364 412324 266416
rect 415492 266364 415544 266416
rect 416412 266364 416464 266416
rect 417976 266364 418028 266416
rect 418804 266364 418856 266416
rect 425428 266364 425480 266416
rect 427084 266364 427136 266416
rect 429568 266364 429620 266416
rect 430396 266364 430448 266416
rect 432052 266364 432104 266416
rect 433156 266364 433208 266416
rect 440332 266364 440384 266416
rect 441344 266364 441396 266416
rect 441988 266364 442040 266416
rect 442908 266364 442960 266416
rect 444472 266364 444524 266416
rect 445668 266364 445720 266416
rect 448612 266364 448664 266416
rect 450544 266364 450596 266416
rect 454408 266364 454460 266416
rect 455328 266364 455380 266416
rect 456892 266364 456944 266416
rect 457996 266364 458048 266416
rect 459376 266364 459428 266416
rect 460204 266364 460256 266416
rect 473452 266364 473504 266416
rect 474648 266364 474700 266416
rect 475108 266364 475160 266416
rect 479524 266364 479576 266416
rect 481732 266364 481784 266416
rect 482836 266364 482888 266416
rect 483388 266364 483440 266416
rect 484216 266364 484268 266416
rect 485872 266364 485924 266416
rect 486792 266364 486844 266416
rect 487160 266296 487212 266348
rect 557724 266296 557776 266348
rect 484216 266160 484268 266212
rect 560300 266160 560352 266212
rect 482560 266024 482612 266076
rect 487160 266024 487212 266076
rect 492496 266024 492548 266076
rect 572720 266024 572772 266076
rect 513196 265888 513248 265940
rect 601700 265888 601752 265940
rect 515680 265752 515732 265804
rect 605840 265752 605892 265804
rect 209780 265616 209832 265668
rect 210700 265616 210752 265668
rect 224960 265616 225012 265668
rect 225604 265616 225656 265668
rect 280344 265616 280396 265668
rect 280988 265616 281040 265668
rect 292672 265616 292724 265668
rect 293500 265616 293552 265668
rect 520648 265616 520700 265668
rect 612740 265616 612792 265668
rect 479248 265480 479300 265532
rect 553400 265480 553452 265532
rect 477592 265344 477644 265396
rect 550640 265344 550692 265396
rect 469312 265208 469364 265260
rect 539968 265208 540020 265260
rect 466828 265072 466880 265124
rect 535736 265072 535788 265124
rect 58624 264460 58676 264512
rect 669136 264460 669188 264512
rect 53104 264324 53156 264376
rect 668216 264324 668268 264376
rect 46204 264188 46256 264240
rect 668952 264188 669004 264240
rect 570604 261468 570656 261520
rect 645860 261468 645912 261520
rect 554412 260856 554464 260908
rect 568580 260856 568632 260908
rect 554320 259428 554372 259480
rect 563704 259428 563756 259480
rect 675852 259428 675904 259480
rect 676404 259428 676456 259480
rect 35808 256776 35860 256828
rect 39580 256776 39632 256828
rect 553952 256708 554004 256760
rect 560944 256708 560996 256760
rect 554504 255552 554556 255604
rect 558184 255552 558236 255604
rect 35808 255416 35860 255468
rect 40500 255416 40552 255468
rect 35624 255280 35676 255332
rect 41696 255280 41748 255332
rect 42064 255280 42116 255332
rect 42800 255280 42852 255332
rect 35808 254328 35860 254380
rect 40684 254328 40736 254380
rect 35808 254056 35860 254108
rect 41512 254056 41564 254108
rect 35624 253920 35676 253972
rect 39948 253920 40000 253972
rect 675852 253104 675904 253156
rect 679624 253104 679676 253156
rect 35808 252696 35860 252748
rect 41328 252696 41380 252748
rect 35624 252560 35676 252612
rect 41696 252560 41748 252612
rect 42064 252560 42116 252612
rect 42708 252560 42760 252612
rect 554412 252560 554464 252612
rect 562324 252560 562376 252612
rect 35808 251200 35860 251252
rect 37924 251200 37976 251252
rect 554136 251200 554188 251252
rect 556804 251200 556856 251252
rect 35808 249908 35860 249960
rect 40316 249908 40368 249960
rect 675392 249568 675444 249620
rect 675392 248480 675444 248532
rect 559564 246304 559616 246356
rect 647240 246304 647292 246356
rect 553860 245624 553912 245676
rect 596824 245624 596876 245676
rect 553492 244264 553544 244316
rect 555424 244264 555476 244316
rect 674656 243652 674708 243704
rect 675208 243652 675260 243704
rect 674840 243176 674892 243228
rect 675208 242904 675260 242956
rect 37924 242836 37976 242888
rect 41696 242836 41748 242888
rect 576124 242156 576176 242208
rect 648620 242156 648672 242208
rect 553676 241476 553728 241528
rect 629944 241476 629996 241528
rect 554504 240116 554556 240168
rect 577504 240116 577556 240168
rect 554320 238688 554372 238740
rect 576124 238688 576176 238740
rect 672172 237056 672224 237108
rect 553768 236784 553820 236836
rect 559564 236784 559616 236836
rect 671160 236580 671212 236632
rect 672954 236648 673006 236700
rect 671988 236444 672040 236496
rect 673184 236240 673236 236292
rect 670976 235900 671028 235952
rect 672908 235900 672960 235952
rect 673000 235696 673052 235748
rect 673184 235492 673236 235544
rect 671988 235288 672040 235340
rect 673874 235084 673926 235136
rect 669688 234812 669740 234864
rect 554412 234540 554464 234592
rect 570604 234540 570656 234592
rect 672172 234472 672224 234524
rect 673552 234472 673604 234524
rect 671344 234336 671396 234388
rect 670332 234132 670384 234184
rect 652208 233860 652260 233912
rect 675484 233860 675536 233912
rect 675852 233860 675904 233912
rect 678244 233860 678296 233912
rect 673000 233384 673052 233436
rect 42340 233248 42392 233300
rect 42708 233248 42760 233300
rect 670884 233180 670936 233232
rect 670056 232840 670108 232892
rect 671988 232840 672040 232892
rect 663064 232636 663116 232688
rect 675484 232636 675536 232688
rect 675852 232636 675904 232688
rect 683120 232636 683172 232688
rect 660304 232500 660356 232552
rect 675484 232500 675536 232552
rect 675852 232500 675904 232552
rect 683304 232500 683356 232552
rect 155132 231752 155184 231804
rect 156972 231752 157024 231804
rect 134892 231616 134944 231668
rect 142068 231616 142120 231668
rect 155500 231616 155552 231668
rect 162676 231616 162728 231668
rect 92388 231480 92440 231532
rect 170772 231480 170824 231532
rect 662512 231480 662564 231532
rect 668584 231480 668636 231532
rect 128268 231344 128320 231396
rect 195888 231344 195940 231396
rect 64328 231208 64380 231260
rect 668032 231208 668084 231260
rect 57244 231072 57296 231124
rect 674840 231276 674892 231328
rect 665088 230936 665140 230988
rect 672172 230936 672224 230988
rect 94504 230868 94556 230920
rect 171416 230868 171468 230920
rect 668584 230800 668636 230852
rect 104808 230732 104860 230784
rect 179144 230732 179196 230784
rect 118608 230596 118660 230648
rect 188160 230596 188212 230648
rect 665272 230596 665324 230648
rect 439320 230528 439372 230580
rect 142160 230460 142212 230512
rect 201040 230460 201092 230512
rect 42340 230392 42392 230444
rect 43076 230392 43128 230444
rect 126888 230392 126940 230444
rect 141976 230392 142028 230444
rect 213092 230392 213144 230444
rect 261576 230392 261628 230444
rect 311992 230392 312044 230444
rect 313096 230392 313148 230444
rect 374644 230392 374696 230444
rect 376208 230392 376260 230444
rect 440700 230392 440752 230444
rect 441896 230392 441948 230444
rect 443460 230392 443512 230444
rect 444472 230392 444524 230444
rect 447600 230392 447652 230444
rect 451556 230392 451608 230444
rect 453304 230392 453356 230444
rect 476120 230392 476172 230444
rect 478604 230392 478656 230444
rect 387432 230324 387484 230376
rect 388444 230324 388496 230376
rect 398104 230324 398156 230376
rect 399392 230324 399444 230376
rect 438676 230324 438728 230376
rect 439320 230324 439372 230376
rect 455420 230324 455472 230376
rect 457168 230324 457220 230376
rect 470876 230324 470928 230376
rect 471888 230324 471940 230376
rect 493416 230324 493468 230376
rect 496360 230324 496412 230376
rect 497280 230324 497332 230376
rect 498108 230324 498160 230376
rect 510804 230324 510856 230376
rect 511908 230324 511960 230376
rect 521108 230324 521160 230376
rect 526444 230324 526496 230376
rect 530124 230324 530176 230376
rect 531136 230324 531188 230376
rect 133788 230256 133840 230308
rect 202328 230256 202380 230308
rect 206284 230256 206336 230308
rect 256424 230256 256476 230308
rect 256608 230256 256660 230308
rect 297640 230256 297692 230308
rect 297824 230256 297876 230308
rect 323400 230256 323452 230308
rect 443828 230188 443880 230240
rect 444656 230188 444708 230240
rect 452844 230188 452896 230240
rect 454316 230188 454368 230240
rect 468300 230188 468352 230240
rect 469128 230188 469180 230240
rect 487620 230188 487672 230240
rect 488448 230188 488500 230240
rect 95240 230120 95292 230172
rect 86224 229984 86276 230036
rect 157156 229984 157208 230036
rect 157432 230120 157484 230172
rect 161112 230120 161164 230172
rect 161296 230120 161348 230172
rect 166264 230120 166316 230172
rect 176476 230120 176528 230172
rect 235816 230120 235868 230172
rect 240324 230120 240376 230172
rect 282184 230120 282236 230172
rect 282644 230120 282696 230172
rect 307944 230120 307996 230172
rect 308128 230120 308180 230172
rect 334992 230120 335044 230172
rect 335176 230120 335228 230172
rect 350448 230120 350500 230172
rect 454132 230052 454184 230104
rect 455328 230052 455380 230104
rect 157800 229984 157852 230036
rect 157984 229984 158036 230036
rect 163688 229984 163740 230036
rect 170956 229984 171008 230036
rect 230664 229984 230716 230036
rect 130384 229848 130436 229900
rect 68284 229712 68336 229764
rect 142160 229712 142212 229764
rect 142620 229848 142672 229900
rect 195060 229848 195112 229900
rect 195428 229848 195480 229900
rect 145012 229712 145064 229764
rect 146944 229712 146996 229764
rect 82084 229576 82136 229628
rect 147772 229576 147824 229628
rect 148140 229712 148192 229764
rect 155960 229712 156012 229764
rect 156328 229712 156380 229764
rect 157294 229712 157346 229764
rect 157432 229712 157484 229764
rect 162584 229712 162636 229764
rect 164056 229712 164108 229764
rect 225512 229712 225564 229764
rect 230480 229848 230532 229900
rect 277032 229984 277084 230036
rect 277216 229984 277268 230036
rect 302792 229984 302844 230036
rect 303252 229984 303304 230036
rect 329840 229984 329892 230036
rect 330944 229984 330996 230036
rect 355600 229984 355652 230036
rect 476672 229984 476724 230036
rect 481640 229984 481692 230036
rect 484400 229984 484452 230036
rect 495164 230188 495216 230240
rect 511448 230188 511500 230240
rect 517520 230188 517572 230240
rect 530768 230188 530820 230240
rect 539600 230392 539652 230444
rect 674676 230392 674728 230444
rect 533528 230256 533580 230308
rect 538312 230256 538364 230308
rect 673092 230188 673144 230240
rect 532700 230120 532752 230172
rect 547144 230120 547196 230172
rect 491484 230052 491536 230104
rect 492496 230052 492548 230104
rect 560944 230052 560996 230104
rect 568120 230052 568172 230104
rect 517244 229984 517296 230036
rect 524604 229984 524656 230036
rect 528836 229984 528888 230036
rect 533528 229984 533580 230036
rect 534632 229984 534684 230036
rect 549260 229984 549312 230036
rect 673276 229984 673328 230036
rect 453488 229916 453540 229968
rect 455788 229916 455840 229968
rect 233700 229848 233752 229900
rect 271880 229848 271932 229900
rect 275652 229848 275704 229900
rect 311992 229848 312044 229900
rect 312636 229848 312688 229900
rect 340144 229848 340196 229900
rect 345664 229848 345716 229900
rect 360752 229848 360804 229900
rect 361212 229848 361264 229900
rect 378784 229848 378836 229900
rect 410892 229848 410944 229900
rect 417424 229848 417476 229900
rect 449624 229848 449676 229900
rect 450544 229848 450596 229900
rect 457352 229848 457404 229900
rect 464068 229848 464120 229900
rect 469588 229848 469640 229900
rect 476764 229848 476816 229900
rect 481824 229848 481876 229900
rect 493692 229848 493744 229900
rect 495992 229848 496044 229900
rect 506388 229848 506440 229900
rect 507584 229848 507636 229900
rect 516784 229848 516836 229900
rect 519176 229848 519228 229900
rect 528560 229848 528612 229900
rect 536564 229848 536616 229900
rect 559564 229848 559616 229900
rect 433524 229780 433576 229832
rect 434168 229780 434220 229832
rect 673874 229780 673926 229832
rect 246120 229712 246172 229764
rect 246488 229712 246540 229764
rect 287336 229712 287388 229764
rect 287704 229712 287756 229764
rect 318248 229712 318300 229764
rect 153384 229576 153436 229628
rect 153844 229576 153896 229628
rect 158536 229576 158588 229628
rect 158720 229576 158772 229628
rect 161756 229576 161808 229628
rect 161940 229576 161992 229628
rect 220360 229576 220412 229628
rect 102140 229440 102192 229492
rect 145656 229440 145708 229492
rect 145840 229440 145892 229492
rect 210056 229440 210108 229492
rect 220268 229440 220320 229492
rect 251272 229576 251324 229628
rect 251732 229576 251784 229628
rect 292488 229576 292540 229628
rect 318064 229576 318116 229628
rect 345296 229712 345348 229764
rect 351736 229712 351788 229764
rect 371056 229712 371108 229764
rect 377680 229712 377732 229764
rect 389088 229712 389140 229764
rect 399852 229712 399904 229764
rect 409696 229712 409748 229764
rect 467012 229712 467064 229764
rect 474004 229712 474056 229764
rect 479248 229712 479300 229764
rect 489920 229712 489972 229764
rect 492128 229712 492180 229764
rect 507124 229712 507176 229764
rect 523040 229712 523092 229764
rect 534724 229712 534776 229764
rect 538496 229712 538548 229764
rect 566832 229712 566884 229764
rect 662328 229712 662380 229764
rect 672172 229712 672224 229764
rect 509516 229644 509568 229696
rect 515496 229644 515548 229696
rect 388628 229576 388680 229628
rect 398748 229576 398800 229628
rect 463792 229576 463844 229628
rect 465724 229576 465776 229628
rect 526904 229576 526956 229628
rect 536104 229576 536156 229628
rect 660948 229576 661000 229628
rect 662512 229576 662564 229628
rect 672908 229576 672960 229628
rect 448980 229508 449032 229560
rect 451372 229508 451424 229560
rect 225604 229440 225656 229492
rect 233700 229440 233752 229492
rect 465448 229440 465500 229492
rect 467472 229440 467524 229492
rect 446404 229372 446456 229424
rect 448980 229372 449032 229424
rect 450912 229372 450964 229424
rect 452660 229372 452712 229424
rect 673460 229372 673512 229424
rect 110144 229304 110196 229356
rect 144644 229304 144696 229356
rect 144828 229304 144880 229356
rect 151452 229304 151504 229356
rect 151636 229304 151688 229356
rect 123484 229168 123536 229220
rect 146944 229168 146996 229220
rect 148324 229168 148376 229220
rect 154028 229168 154080 229220
rect 154396 229304 154448 229356
rect 157156 229304 157208 229356
rect 157340 229304 157392 229356
rect 215208 229304 215260 229356
rect 413836 229304 413888 229356
rect 420000 229304 420052 229356
rect 472164 229304 472216 229356
rect 472992 229304 473044 229356
rect 450268 229236 450320 229288
rect 451740 229236 451792 229288
rect 495348 229236 495400 229288
rect 500224 229236 500276 229288
rect 505652 229236 505704 229288
rect 510620 229236 510672 229288
rect 513380 229236 513432 229288
rect 519084 229236 519136 229288
rect 156328 229168 156380 229220
rect 162584 229168 162636 229220
rect 180432 229168 180484 229220
rect 183376 229168 183428 229220
rect 240968 229168 241020 229220
rect 423496 229100 423548 229152
rect 427728 229100 427780 229152
rect 441252 229100 441304 229152
rect 442080 229100 442132 229152
rect 503720 229100 503772 229152
rect 509884 229100 509936 229152
rect 515312 229100 515364 229152
rect 520924 229100 520976 229152
rect 524972 229100 525024 229152
rect 529940 229100 529992 229152
rect 673874 229100 673926 229152
rect 100668 229032 100720 229084
rect 167368 229032 167420 229084
rect 167552 229032 167604 229084
rect 169484 229032 169536 229084
rect 106188 228896 106240 228948
rect 179788 229032 179840 229084
rect 180064 229032 180116 229084
rect 185584 229032 185636 229084
rect 189724 229032 189776 229084
rect 93768 228760 93820 228812
rect 166356 228760 166408 228812
rect 184940 228896 184992 228948
rect 185400 228896 185452 228948
rect 190092 228896 190144 228948
rect 192484 229032 192536 229084
rect 200396 229032 200448 229084
rect 201408 229032 201460 229084
rect 252560 229032 252612 229084
rect 255228 229032 255280 229084
rect 295708 229032 295760 229084
rect 305552 229032 305604 229084
rect 315672 229032 315724 229084
rect 326896 229032 326948 229084
rect 351092 229032 351144 229084
rect 195244 228896 195296 228948
rect 195612 228896 195664 228948
rect 246764 228896 246816 228948
rect 248236 228896 248288 228948
rect 291844 228896 291896 228948
rect 302148 228896 302200 228948
rect 331220 228896 331272 228948
rect 506388 228896 506440 228948
rect 512736 228896 512788 228948
rect 526444 228896 526496 228948
rect 544016 228896 544068 228948
rect 67548 228624 67600 228676
rect 146024 228624 146076 228676
rect 173164 228760 173216 228812
rect 231308 228760 231360 228812
rect 238576 228760 238628 228812
rect 282828 228760 282880 228812
rect 291844 228760 291896 228812
rect 300216 228760 300268 228812
rect 300676 228760 300728 228812
rect 330484 228760 330536 228812
rect 376024 228760 376076 228812
rect 387800 228760 387852 228812
rect 478880 228760 478932 228812
rect 490380 228760 490432 228812
rect 499856 228760 499908 228812
rect 518164 228760 518216 228812
rect 518532 228760 518584 228812
rect 541624 228760 541676 228812
rect 61384 228488 61436 228540
rect 57244 228352 57296 228404
rect 136824 228352 136876 228404
rect 137376 228488 137428 228540
rect 166954 228624 167006 228676
rect 181444 228624 181496 228676
rect 181628 228624 181680 228676
rect 185400 228624 185452 228676
rect 185584 228624 185636 228676
rect 226156 228624 226208 228676
rect 226340 228624 226392 228676
rect 272524 228624 272576 228676
rect 296628 228624 296680 228676
rect 329196 228624 329248 228676
rect 336464 228624 336516 228676
rect 358820 228624 358872 228676
rect 359924 228624 359976 228676
rect 376852 228624 376904 228676
rect 485688 228624 485740 228676
rect 498292 228624 498344 228676
rect 498568 228624 498620 228676
rect 515772 228624 515824 228676
rect 517888 228624 517940 228676
rect 539416 228624 539468 228676
rect 539600 228624 539652 228676
rect 557172 228624 557224 228676
rect 147128 228488 147180 228540
rect 200120 228488 200172 228540
rect 200304 228488 200356 228540
rect 221004 228488 221056 228540
rect 112996 228216 113048 228268
rect 137192 228216 137244 228268
rect 139308 228352 139360 228404
rect 143080 228216 143132 228268
rect 143448 228216 143500 228268
rect 145840 228216 145892 228268
rect 146024 228216 146076 228268
rect 148876 228216 148928 228268
rect 153108 228352 153160 228404
rect 215852 228352 215904 228404
rect 216496 228352 216548 228404
rect 264796 228488 264848 228540
rect 272524 228488 272576 228540
rect 309876 228488 309928 228540
rect 313924 228488 313976 228540
rect 320824 228488 320876 228540
rect 325424 228488 325476 228540
rect 349160 228488 349212 228540
rect 350448 228488 350500 228540
rect 369124 228488 369176 228540
rect 371056 228488 371108 228540
rect 385224 228488 385276 228540
rect 386052 228488 386104 228540
rect 397460 228488 397512 228540
rect 224776 228352 224828 228404
rect 273812 228352 273864 228404
rect 285496 228352 285548 228404
rect 318892 228352 318944 228404
rect 330484 228352 330536 228404
rect 354956 228352 355008 228404
rect 355324 228352 355376 228404
rect 372988 228352 373040 228404
rect 373448 228352 373500 228404
rect 387156 228352 387208 228404
rect 390008 228352 390060 228404
rect 400036 228352 400088 228404
rect 205548 228216 205600 228268
rect 205732 228216 205784 228268
rect 257068 228216 257120 228268
rect 257620 228216 257672 228268
rect 296352 228216 296404 228268
rect 407764 228488 407816 228540
rect 409788 228488 409840 228540
rect 415492 228488 415544 228540
rect 485044 228488 485096 228540
rect 498660 228488 498712 228540
rect 502432 228488 502484 228540
rect 521108 228488 521160 228540
rect 527548 228488 527600 228540
rect 553308 228488 553360 228540
rect 556804 228488 556856 228540
rect 570604 228488 570656 228540
rect 402796 228352 402848 228404
rect 411628 228352 411680 228404
rect 474464 228352 474516 228404
rect 484492 228352 484544 228404
rect 490196 228352 490248 228404
rect 505192 228352 505244 228404
rect 512092 228352 512144 228404
rect 533528 228352 533580 228404
rect 537208 228352 537260 228404
rect 565636 228352 565688 228404
rect 672494 228352 672546 228404
rect 673092 228352 673144 228404
rect 539416 228216 539468 228268
rect 540796 228216 540848 228268
rect 119988 228080 120040 228132
rect 181260 228080 181312 228132
rect 181444 228080 181496 228132
rect 126704 227944 126756 227996
rect 195244 228080 195296 228132
rect 239036 228080 239088 228132
rect 246304 228080 246356 228132
rect 253848 228080 253900 228132
rect 268936 228080 268988 228132
rect 306012 228080 306064 228132
rect 400128 228080 400180 228132
rect 415032 228012 415084 228064
rect 421932 228012 421984 228064
rect 88248 227808 88300 227860
rect 95240 227808 95292 227860
rect 133512 227808 133564 227860
rect 136640 227808 136692 227860
rect 136824 227808 136876 227860
rect 141148 227808 141200 227860
rect 141516 227808 141568 227860
rect 192484 227808 192536 227860
rect 200304 227944 200356 227996
rect 210424 227944 210476 227996
rect 238392 227944 238444 227996
rect 416688 227876 416740 227928
rect 420644 227876 420696 227928
rect 447048 227876 447100 227928
rect 450544 227876 450596 227928
rect 195060 227808 195112 227860
rect 200120 227808 200172 227860
rect 210240 227808 210292 227860
rect 409052 227740 409104 227792
rect 410340 227740 410392 227792
rect 411904 227740 411956 227792
rect 413560 227740 413612 227792
rect 420644 227740 420696 227792
rect 423864 227740 423916 227792
rect 471520 227740 471572 227792
rect 479524 227740 479576 227792
rect 75184 227672 75236 227724
rect 146300 227672 146352 227724
rect 150072 227672 150124 227724
rect 213368 227672 213420 227724
rect 213828 227672 213880 227724
rect 262864 227672 262916 227724
rect 263508 227672 263560 227724
rect 277216 227672 277268 227724
rect 64788 227536 64840 227588
rect 110144 227536 110196 227588
rect 110328 227536 110380 227588
rect 182364 227536 182416 227588
rect 185400 227536 185452 227588
rect 192668 227536 192720 227588
rect 200028 227536 200080 227588
rect 205640 227536 205692 227588
rect 214564 227536 214616 227588
rect 214748 227536 214800 227588
rect 262220 227536 262272 227588
rect 277216 227536 277268 227588
rect 311808 227672 311860 227724
rect 465908 227604 465960 227656
rect 469864 227604 469916 227656
rect 282184 227536 282236 227588
rect 308588 227536 308640 227588
rect 524604 227536 524656 227588
rect 539968 227536 540020 227588
rect 60648 227400 60700 227452
rect 102140 227400 102192 227452
rect 103428 227400 103480 227452
rect 177212 227400 177264 227452
rect 181260 227400 181312 227452
rect 96528 227264 96580 227316
rect 169392 227264 169444 227316
rect 169576 227264 169628 227316
rect 172060 227264 172112 227316
rect 185584 227264 185636 227316
rect 186136 227400 186188 227452
rect 204812 227400 204864 227452
rect 251916 227400 251968 227452
rect 259276 227400 259328 227452
rect 298284 227400 298336 227452
rect 304908 227400 304960 227452
rect 333704 227400 333756 227452
rect 333888 227400 333940 227452
rect 356244 227400 356296 227452
rect 357072 227400 357124 227452
rect 374276 227400 374328 227452
rect 514024 227400 514076 227452
rect 535736 227400 535788 227452
rect 538312 227400 538364 227452
rect 556068 227400 556120 227452
rect 219164 227264 219216 227316
rect 220084 227264 220136 227316
rect 241612 227264 241664 227316
rect 257804 227264 257856 227316
rect 299572 227264 299624 227316
rect 310428 227264 310480 227316
rect 338212 227264 338264 227316
rect 340696 227264 340748 227316
rect 361396 227264 361448 227316
rect 89628 227128 89680 227180
rect 157294 227128 157346 227180
rect 157432 227128 157484 227180
rect 171508 227128 171560 227180
rect 56508 226992 56560 227044
rect 142436 226992 142488 227044
rect 143264 226992 143316 227044
rect 208124 226992 208176 227044
rect 214564 226992 214616 227044
rect 220084 226992 220136 227044
rect 220452 226992 220504 227044
rect 222936 226992 222988 227044
rect 235816 227128 235868 227180
rect 280252 227128 280304 227180
rect 306196 227128 306248 227180
rect 336924 227128 336976 227180
rect 338672 227128 338724 227180
rect 360108 227128 360160 227180
rect 362776 227128 362828 227180
rect 379428 227128 379480 227180
rect 382096 227128 382148 227180
rect 392952 227128 393004 227180
rect 393136 227128 393188 227180
rect 402612 227264 402664 227316
rect 494704 227264 494756 227316
rect 402244 227128 402296 227180
rect 408408 227128 408460 227180
rect 478604 227128 478656 227180
rect 486792 227128 486844 227180
rect 489552 227128 489604 227180
rect 504180 227128 504232 227180
rect 228732 226992 228784 227044
rect 228916 226992 228968 227044
rect 271236 226992 271288 227044
rect 271788 226992 271840 227044
rect 282184 226992 282236 227044
rect 122748 226856 122800 226908
rect 185400 226856 185452 226908
rect 185584 226856 185636 226908
rect 218428 226856 218480 226908
rect 219348 226856 219400 226908
rect 267372 226856 267424 226908
rect 281356 226856 281408 226908
rect 317604 226992 317656 227044
rect 322848 226992 322900 227044
rect 349804 226992 349856 227044
rect 355876 226992 355928 227044
rect 375564 226992 375616 227044
rect 376668 226992 376720 227044
rect 389732 226992 389784 227044
rect 391848 226992 391900 227044
rect 403532 226992 403584 227044
rect 412548 226992 412600 227044
rect 419356 226992 419408 227044
rect 486976 226992 487028 227044
rect 500960 226992 501012 227044
rect 293776 226856 293828 226908
rect 324964 226856 325016 226908
rect 510620 227264 510672 227316
rect 524420 227264 524472 227316
rect 526260 227264 526312 227316
rect 551560 227264 551612 227316
rect 506204 227128 506256 227180
rect 525984 227128 526036 227180
rect 533344 227128 533396 227180
rect 560944 227128 560996 227180
rect 669228 227128 669280 227180
rect 669872 227128 669924 227180
rect 505008 226992 505060 227044
rect 523040 226992 523092 227044
rect 523684 226992 523736 227044
rect 548340 226992 548392 227044
rect 555424 226992 555476 227044
rect 633716 226992 633768 227044
rect 510988 226856 511040 226908
rect 117228 226720 117280 226772
rect 187516 226720 187568 226772
rect 190000 226720 190052 226772
rect 233884 226720 233936 226772
rect 249616 226720 249668 226772
rect 290556 226720 290608 226772
rect 668400 226720 668452 226772
rect 672540 226992 672592 227044
rect 243452 226652 243504 226704
rect 248696 226652 248748 226704
rect 129556 226584 129608 226636
rect 197360 226584 197412 226636
rect 203524 226584 203576 226636
rect 136548 226448 136600 226500
rect 141792 226448 141844 226500
rect 142252 226448 142304 226500
rect 202972 226448 203024 226500
rect 212172 226448 212224 226500
rect 214748 226448 214800 226500
rect 219164 226584 219216 226636
rect 223580 226584 223632 226636
rect 231032 226584 231084 226636
rect 243268 226584 243320 226636
rect 264152 226584 264204 226636
rect 269304 226584 269356 226636
rect 669872 226584 669924 226636
rect 670516 226584 670568 226636
rect 673276 226516 673328 226568
rect 220452 226448 220504 226500
rect 221832 226448 221884 226500
rect 228916 226448 228968 226500
rect 351092 226448 351144 226500
rect 353024 226448 353076 226500
rect 403992 226448 404044 226500
rect 412272 226448 412324 226500
rect 474740 226448 474792 226500
rect 482744 226448 482796 226500
rect 141976 226380 142028 226432
rect 142114 226380 142166 226432
rect 271144 226380 271196 226432
rect 279608 226380 279660 226432
rect 672724 226380 672776 226432
rect 350264 226312 350316 226364
rect 351736 226312 351788 226364
rect 388536 226312 388588 226364
rect 391664 226312 391716 226364
rect 407764 226312 407816 226364
rect 408684 226312 408736 226364
rect 481640 226312 481692 226364
rect 487804 226312 487856 226364
rect 663432 226312 663484 226364
rect 665272 226312 665324 226364
rect 58992 226244 59044 226296
rect 130384 226244 130436 226296
rect 135076 226244 135128 226296
rect 204260 226244 204312 226296
rect 208124 226244 208176 226296
rect 257436 226244 257488 226296
rect 267004 226244 267056 226296
rect 274456 226244 274508 226296
rect 286324 226244 286376 226296
rect 289912 226244 289964 226296
rect 291016 226244 291068 226296
rect 322112 226244 322164 226296
rect 458640 226244 458692 226296
rect 462964 226244 463016 226296
rect 127440 226108 127492 226160
rect 142114 226108 142166 226160
rect 142252 226108 142304 226160
rect 209412 226108 209464 226160
rect 209688 226108 209740 226160
rect 259644 226108 259696 226160
rect 261852 226108 261904 226160
rect 300860 226108 300912 226160
rect 309048 226108 309100 226160
rect 336280 226108 336332 226160
rect 528560 226108 528612 226160
rect 542636 226108 542688 226160
rect 672604 226108 672656 226160
rect 66168 225972 66220 226024
rect 142620 225972 142672 226024
rect 142804 225972 142856 226024
rect 147588 225972 147640 226024
rect 147772 225972 147824 226024
rect 83464 225836 83516 225888
rect 155500 225836 155552 225888
rect 157340 225972 157392 226024
rect 217140 225972 217192 226024
rect 222016 225972 222068 226024
rect 269948 225972 270000 226024
rect 278412 225972 278464 226024
rect 313280 225972 313332 226024
rect 329748 225972 329800 226024
rect 353668 225972 353720 226024
rect 354588 225972 354640 226024
rect 372344 225972 372396 226024
rect 498108 225972 498160 226024
rect 514300 225972 514352 226024
rect 516600 225972 516652 226024
rect 538680 225972 538732 226024
rect 672494 225904 672546 225956
rect 198004 225836 198056 225888
rect 249340 225836 249392 225888
rect 252468 225836 252520 225888
rect 293132 225836 293184 225888
rect 296444 225836 296496 225888
rect 327540 225836 327592 225888
rect 332232 225836 332284 225888
rect 357532 225836 357584 225888
rect 373816 225836 373868 225888
rect 377680 225836 377732 225888
rect 377864 225836 377916 225888
rect 390376 225836 390428 225888
rect 394332 225836 394384 225888
rect 403256 225836 403308 225888
rect 483756 225836 483808 225888
rect 497280 225836 497332 225888
rect 501144 225836 501196 225888
rect 519268 225836 519320 225888
rect 521752 225836 521804 225888
rect 545764 225836 545816 225888
rect 558184 225836 558236 225888
rect 572260 225836 572312 225888
rect 672172 225836 672224 225888
rect 76564 225700 76616 225752
rect 184020 225700 184072 225752
rect 184204 225700 184256 225752
rect 212632 225700 212684 225752
rect 237288 225700 237340 225752
rect 240324 225700 240376 225752
rect 255044 225700 255096 225752
rect 296996 225700 297048 225752
rect 315672 225700 315724 225752
rect 344652 225700 344704 225752
rect 352932 225700 352984 225752
rect 371608 225700 371660 225752
rect 371792 225700 371844 225752
rect 382740 225700 382792 225752
rect 382924 225700 382976 225752
rect 396172 225700 396224 225752
rect 488908 225700 488960 225752
rect 503628 225700 503680 225752
rect 508872 225700 508924 225752
rect 529204 225700 529256 225752
rect 535920 225700 535972 225752
rect 563980 225700 564032 225752
rect 156604 225632 156656 225684
rect 72424 225564 72476 225616
rect 142114 225564 142166 225616
rect 142252 225564 142304 225616
rect 147680 225564 147732 225616
rect 157340 225564 157392 225616
rect 214380 225564 214432 225616
rect 215208 225564 215260 225616
rect 266084 225564 266136 225616
rect 270040 225564 270092 225616
rect 282644 225564 282696 225616
rect 284116 225564 284168 225616
rect 320180 225564 320232 225616
rect 321376 225564 321428 225616
rect 346584 225564 346636 225616
rect 347044 225564 347096 225616
rect 367836 225564 367888 225616
rect 372528 225564 372580 225616
rect 387432 225564 387484 225616
rect 390192 225564 390244 225616
rect 401968 225564 402020 225616
rect 410984 225564 411036 225616
rect 416136 225564 416188 225616
rect 467656 225564 467708 225616
rect 476580 225564 476632 225616
rect 477316 225564 477368 225616
rect 488816 225564 488868 225616
rect 494060 225564 494112 225616
rect 509700 225564 509752 225616
rect 510160 225564 510212 225616
rect 530952 225564 531004 225616
rect 531412 225564 531464 225616
rect 558276 225564 558328 225616
rect 672264 225496 672316 225548
rect 110144 225428 110196 225480
rect 127440 225428 127492 225480
rect 122564 225156 122616 225208
rect 193588 225428 193640 225480
rect 193772 225428 193824 225480
rect 244188 225428 244240 225480
rect 463148 225360 463200 225412
rect 467288 225360 467340 225412
rect 672156 225360 672208 225412
rect 125232 225020 125284 225072
rect 196164 225292 196216 225344
rect 196624 225292 196676 225344
rect 236460 225292 236512 225344
rect 241152 225292 241204 225344
rect 286692 225292 286744 225344
rect 129372 225156 129424 225208
rect 199108 225156 199160 225208
rect 242716 225156 242768 225208
rect 285036 225156 285088 225208
rect 132408 225020 132460 225072
rect 201684 225020 201736 225072
rect 202236 225020 202288 225072
rect 254492 225020 254544 225072
rect 297272 224952 297324 225004
rect 305368 224952 305420 225004
rect 327724 224952 327776 225004
rect 332048 224952 332100 225004
rect 369124 224952 369176 225004
rect 373632 224952 373684 225004
rect 404176 224952 404228 225004
rect 410616 224952 410668 225004
rect 416504 224952 416556 225004
rect 422208 224952 422260 225004
rect 493692 224952 493744 225004
rect 494704 224952 494756 225004
rect 495164 224952 495216 225004
rect 567016 225088 567068 225140
rect 571432 225088 571484 225140
rect 563704 224952 563756 225004
rect 672034 225224 672086 225276
rect 666468 225156 666520 225208
rect 96068 224884 96120 224936
rect 172980 224884 173032 224936
rect 174912 224884 174964 224936
rect 185584 224884 185636 224936
rect 185768 224884 185820 224936
rect 195244 224884 195296 224936
rect 195612 224884 195664 224936
rect 242900 224884 242952 224936
rect 266176 224884 266228 224936
rect 630864 224952 630916 225004
rect 568948 224884 569000 224936
rect 303436 224816 303488 224868
rect 549260 224816 549312 224868
rect 554780 224816 554832 224868
rect 610992 224816 611044 224868
rect 614948 224816 615000 224868
rect 102048 224748 102100 224800
rect 178500 224748 178552 224800
rect 178684 224748 178736 224800
rect 204536 224748 204588 224800
rect 204720 224748 204772 224800
rect 79968 224612 80020 224664
rect 160468 224612 160520 224664
rect 162768 224612 162820 224664
rect 224040 224612 224092 224664
rect 224592 224748 224644 224800
rect 237748 224612 237800 224664
rect 245292 224748 245344 224800
rect 287980 224748 288032 224800
rect 311532 224748 311584 224800
rect 338856 224748 338908 224800
rect 462504 224748 462556 224800
rect 469312 224748 469364 224800
rect 506940 224748 506992 224800
rect 526720 224748 526772 224800
rect 529940 224748 529992 224800
rect 549076 224748 549128 224800
rect 554964 224748 555016 224800
rect 555792 224748 555844 224800
rect 555976 224748 556028 224800
rect 562140 224748 562192 224800
rect 562324 224748 562376 224800
rect 567016 224748 567068 224800
rect 567844 224748 567896 224800
rect 610808 224748 610860 224800
rect 670516 224748 670568 224800
rect 270592 224612 270644 224664
rect 274272 224612 274324 224664
rect 312452 224612 312504 224664
rect 319996 224612 320048 224664
rect 345940 224612 345992 224664
rect 346216 224612 346268 224664
rect 366548 224612 366600 224664
rect 505192 224612 505244 224664
rect 610440 224612 610492 224664
rect 610624 224612 610676 224664
rect 616052 224612 616104 224664
rect 668584 224612 668636 224664
rect 85488 224476 85540 224528
rect 165620 224476 165672 224528
rect 179328 224476 179380 224528
rect 185400 224476 185452 224528
rect 185584 224476 185636 224528
rect 235172 224476 235224 224528
rect 251088 224476 251140 224528
rect 294420 224476 294472 224528
rect 299296 224476 299348 224528
rect 331772 224476 331824 224528
rect 335176 224476 335228 224528
rect 356888 224476 356940 224528
rect 366732 224476 366784 224528
rect 381636 224476 381688 224528
rect 456064 224476 456116 224528
rect 459744 224476 459796 224528
rect 491300 224476 491352 224528
rect 506020 224476 506072 224528
rect 515956 224476 516008 224528
rect 538312 224476 538364 224528
rect 538864 224476 538916 224528
rect 73712 224340 73764 224392
rect 155316 224340 155368 224392
rect 157248 224340 157300 224392
rect 161940 224340 161992 224392
rect 165528 224340 165580 224392
rect 227444 224340 227496 224392
rect 228732 224340 228784 224392
rect 274916 224340 274968 224392
rect 275100 224340 275152 224392
rect 311164 224340 311216 224392
rect 319812 224340 319864 224392
rect 347228 224340 347280 224392
rect 361212 224340 361264 224392
rect 377496 224340 377548 224392
rect 387708 224340 387760 224392
rect 397828 224340 397880 224392
rect 480536 224340 480588 224392
rect 492772 224340 492824 224392
rect 499212 224340 499264 224392
rect 516784 224340 516836 224392
rect 525616 224340 525668 224392
rect 550824 224340 550876 224392
rect 552848 224476 552900 224528
rect 625436 224476 625488 224528
rect 68928 224204 68980 224256
rect 96252 224204 96304 224256
rect 89444 224068 89496 224120
rect 167828 224204 167880 224256
rect 168288 224204 168340 224256
rect 230020 224204 230072 224256
rect 231676 224204 231728 224256
rect 278964 224204 279016 224256
rect 290832 224204 290884 224256
rect 323676 224204 323728 224256
rect 323952 224204 324004 224256
rect 334992 224204 335044 224256
rect 339408 224204 339460 224256
rect 362316 224204 362368 224256
rect 363604 224204 363656 224256
rect 368480 224204 368532 224256
rect 379244 224204 379296 224256
rect 393596 224204 393648 224256
rect 394516 224204 394568 224256
rect 404544 224204 404596 224256
rect 405556 224204 405608 224256
rect 414204 224204 414256 224256
rect 470232 224204 470284 224256
rect 480444 224204 480496 224256
rect 486608 224204 486660 224256
rect 500408 224204 500460 224256
rect 504364 224204 504416 224256
rect 523500 224204 523552 224256
rect 524420 224204 524472 224256
rect 525064 224204 525116 224256
rect 538864 224204 538916 224256
rect 539324 224204 539376 224256
rect 555976 224204 556028 224256
rect 556344 224340 556396 224392
rect 625252 224340 625304 224392
rect 671596 224340 671648 224392
rect 671482 224272 671534 224324
rect 619640 224204 619692 224256
rect 96252 223932 96304 223984
rect 137974 224068 138026 224120
rect 138112 224068 138164 224120
rect 194600 224068 194652 224120
rect 195244 224068 195296 224120
rect 204720 224068 204772 224120
rect 204904 224068 204956 224120
rect 250628 224068 250680 224120
rect 286692 224068 286744 224120
rect 319536 224068 319588 224120
rect 358084 224068 358136 224120
rect 363236 224068 363288 224120
rect 509700 224068 509752 224120
rect 510160 224068 510212 224120
rect 610624 224068 610676 224120
rect 377404 224000 377456 224052
rect 385868 224000 385920 224052
rect 610808 224000 610860 224052
rect 623780 224000 623832 224052
rect 106004 223932 106056 223984
rect 181076 223932 181128 223984
rect 201224 223932 201276 223984
rect 255780 223932 255832 223984
rect 279424 223932 279476 223984
rect 284760 223932 284812 223984
rect 519084 223932 519136 223984
rect 108672 223796 108724 223848
rect 183836 223796 183888 223848
rect 112812 223660 112864 223712
rect 185952 223796 186004 223848
rect 186964 223796 187016 223848
rect 217784 223796 217836 223848
rect 233148 223796 233200 223848
rect 277676 223796 277728 223848
rect 535276 223932 535328 223984
rect 539324 223932 539376 223984
rect 539968 223864 540020 223916
rect 622676 223864 622728 223916
rect 535092 223728 535144 223780
rect 621572 223728 621624 223780
rect 184848 223660 184900 223712
rect 195612 223660 195664 223712
rect 195888 223660 195940 223712
rect 204904 223660 204956 223712
rect 238024 223660 238076 223712
rect 266728 223660 266780 223712
rect 460572 223660 460624 223712
rect 463148 223660 463200 223712
rect 520464 223592 520516 223644
rect 543832 223592 543884 223644
rect 544016 223592 544068 223644
rect 544936 223592 544988 223644
rect 567844 223592 567896 223644
rect 81348 223524 81400 223576
rect 159824 223524 159876 223576
rect 162124 223524 162176 223576
rect 186596 223524 186648 223576
rect 187332 223524 187384 223576
rect 242256 223524 242308 223576
rect 250904 223524 250956 223576
rect 291200 223524 291252 223576
rect 297916 223524 297968 223576
rect 303252 223524 303304 223576
rect 307668 223524 307720 223576
rect 335636 223524 335688 223576
rect 406752 223524 406804 223576
rect 414848 223524 414900 223576
rect 454868 223524 454920 223576
rect 460480 223524 460532 223576
rect 473452 223524 473504 223576
rect 475568 223524 475620 223576
rect 75828 223388 75880 223440
rect 154672 223388 154724 223440
rect 159364 223388 159416 223440
rect 175924 223388 175976 223440
rect 184664 223388 184716 223440
rect 239680 223388 239732 223440
rect 244096 223388 244148 223440
rect 286048 223388 286100 223440
rect 312912 223388 312964 223440
rect 342076 223456 342128 223508
rect 566832 223456 566884 223508
rect 628748 223592 628800 223644
rect 342812 223388 342864 223440
rect 347872 223388 347924 223440
rect 493048 223388 493100 223440
rect 508596 223388 508648 223440
rect 517520 223388 517572 223440
rect 531504 223388 531556 223440
rect 534724 223388 534776 223440
rect 547420 223388 547472 223440
rect 336004 223320 336056 223372
rect 342260 223320 342312 223372
rect 69572 223252 69624 223304
rect 66904 223116 66956 223168
rect 142528 223116 142580 223168
rect 143816 223252 143868 223304
rect 152096 223252 152148 223304
rect 156420 223252 156472 223304
rect 162400 223252 162452 223304
rect 171784 223252 171836 223304
rect 199752 223252 199804 223304
rect 204720 223252 204772 223304
rect 51908 222980 51960 223032
rect 63132 222980 63184 223032
rect 71412 222980 71464 223032
rect 139860 222980 139912 223032
rect 143632 223116 143684 223168
rect 146576 223116 146628 223168
rect 146760 223116 146812 223168
rect 173348 223116 173400 223168
rect 173532 223116 173584 223168
rect 185768 223116 185820 223168
rect 194508 223116 194560 223168
rect 204904 223116 204956 223168
rect 211436 223252 211488 223304
rect 214380 223252 214432 223304
rect 211620 223116 211672 223168
rect 149520 222980 149572 223032
rect 62764 222844 62816 222896
rect 144000 222844 144052 222896
rect 145104 222844 145156 222896
rect 166264 222980 166316 223032
rect 166448 222980 166500 223032
rect 219532 223252 219584 223304
rect 246856 223252 246908 223304
rect 288624 223252 288676 223304
rect 289728 223252 289780 223304
rect 297732 223252 297784 223304
rect 299112 223252 299164 223304
rect 328552 223252 328604 223304
rect 347228 223252 347280 223304
rect 357900 223252 357952 223304
rect 483112 223252 483164 223304
rect 496084 223252 496136 223304
rect 514668 223252 514720 223304
rect 536656 223252 536708 223304
rect 564624 223252 564676 223304
rect 154212 222844 154264 222896
rect 211436 222844 211488 222896
rect 211804 222844 211856 222896
rect 228088 223116 228140 223168
rect 241336 223116 241388 223168
rect 283472 223116 283524 223168
rect 288256 223116 288308 223168
rect 321100 223116 321152 223168
rect 344652 223116 344704 223168
rect 364616 223116 364668 223168
rect 365536 223116 365588 223168
rect 379612 223116 379664 223168
rect 380072 223116 380124 223168
rect 386512 223116 386564 223168
rect 488632 223116 488684 223168
rect 503168 223116 503220 223168
rect 503352 223116 503404 223168
rect 521752 223116 521804 223168
rect 532056 223116 532108 223168
rect 559012 223116 559064 223168
rect 561680 223116 561732 223168
rect 562416 223116 562468 223168
rect 564808 223116 564860 223168
rect 214840 222980 214892 223032
rect 216220 222980 216272 223032
rect 230204 222980 230256 223032
rect 275468 222980 275520 223032
rect 278596 222980 278648 223032
rect 315028 222980 315080 223032
rect 316684 222980 316736 223032
rect 327264 222980 327316 223032
rect 328092 222980 328144 223032
rect 351460 222980 351512 223032
rect 353944 222980 353996 223032
rect 365904 222980 365956 223032
rect 366916 222980 366968 223032
rect 383936 222980 383988 223032
rect 384304 222980 384356 223032
rect 393964 222980 394016 223032
rect 482744 222980 482796 223032
rect 593972 222980 594024 223032
rect 620652 223116 620704 223168
rect 669228 224000 669280 224052
rect 670516 224000 670568 224052
rect 669228 223728 669280 223780
rect 670056 223728 670108 223780
rect 669872 223592 669924 223644
rect 669688 223524 669740 223576
rect 669596 223388 669648 223440
rect 669872 223116 669924 223168
rect 620284 222980 620336 223032
rect 625620 222980 625672 223032
rect 669688 223048 669740 223100
rect 669872 222912 669924 222964
rect 215944 222844 215996 222896
rect 233332 222844 233384 222896
rect 234528 222844 234580 222896
rect 281540 222844 281592 222896
rect 282460 222844 282512 222896
rect 316316 222844 316368 222896
rect 324136 222844 324188 222896
rect 348516 222844 348568 222896
rect 349068 222844 349120 222896
rect 367192 222844 367244 222896
rect 368388 222844 368440 222896
rect 382372 222844 382424 222896
rect 383476 222844 383528 222896
rect 394884 222844 394936 222896
rect 395804 222844 395856 222896
rect 406476 222844 406528 222896
rect 420828 222844 420880 222896
rect 425152 222844 425204 222896
rect 459928 222844 459980 222896
rect 467104 222844 467156 222896
rect 467472 222844 467524 222896
rect 473728 222844 473780 222896
rect 479892 222844 479944 222896
rect 491944 222844 491996 222896
rect 500776 222844 500828 222896
rect 517520 222844 517572 222896
rect 519820 222844 519872 222896
rect 542360 222844 542412 222896
rect 554044 222844 554096 222896
rect 632704 222844 632756 222896
rect 651288 222844 651340 222896
rect 666468 222844 666520 222896
rect 670056 222844 670108 222896
rect 78588 222708 78640 222760
rect 155132 222708 155184 222760
rect 155684 222708 155736 222760
rect 87972 222572 88024 222624
rect 164976 222572 165028 222624
rect 166264 222708 166316 222760
rect 173532 222708 173584 222760
rect 166448 222572 166500 222624
rect 166632 222572 166684 222624
rect 173900 222572 173952 222624
rect 175556 222572 175608 222624
rect 175924 222572 175976 222624
rect 181812 222572 181864 222624
rect 185768 222708 185820 222760
rect 204720 222708 204772 222760
rect 204904 222708 204956 222760
rect 247408 222708 247460 222760
rect 264796 222708 264848 222760
rect 304356 222708 304408 222760
rect 508228 222708 508280 222760
rect 527824 222708 527876 222760
rect 552480 222708 552532 222760
rect 555700 222708 555752 222760
rect 558184 222708 558236 222760
rect 620284 222708 620336 222760
rect 620468 222708 620520 222760
rect 627092 222708 627144 222760
rect 304724 222640 304776 222692
rect 308128 222640 308180 222692
rect 670516 223116 670568 223168
rect 670516 222640 670568 222692
rect 192024 222572 192076 222624
rect 197176 222572 197228 222624
rect 249984 222572 250036 222624
rect 529848 222572 529900 222624
rect 619916 222572 619968 222624
rect 426440 222504 426492 222556
rect 426992 222504 427044 222556
rect 85304 222436 85356 222488
rect 156420 222436 156472 222488
rect 156604 222436 156656 222488
rect 99288 222300 99340 222352
rect 118424 222164 118476 222216
rect 156604 222164 156656 222216
rect 173348 222300 173400 222352
rect 175740 222300 175792 222352
rect 176108 222436 176160 222488
rect 207480 222436 207532 222488
rect 207664 222436 207716 222488
rect 258356 222436 258408 222488
rect 489920 222436 489972 222488
rect 491116 222436 491168 222488
rect 173900 222164 173952 222216
rect 188896 222300 188948 222352
rect 245108 222300 245160 222352
rect 287888 222300 287940 222352
rect 295064 222300 295116 222352
rect 484492 222300 484544 222352
rect 504364 222436 504416 222488
rect 523684 222436 523736 222488
rect 529480 222436 529532 222488
rect 552480 222436 552532 222488
rect 552664 222436 552716 222488
rect 564624 222436 564676 222488
rect 564808 222436 564860 222488
rect 627920 222436 627972 222488
rect 191012 222164 191064 222216
rect 629852 222300 629904 222352
rect 504364 222164 504416 222216
rect 523684 222164 523736 222216
rect 552664 222164 552716 222216
rect 552848 222164 552900 222216
rect 558184 222164 558236 222216
rect 558552 222164 558604 222216
rect 559932 222164 559984 222216
rect 620468 222164 620520 222216
rect 620652 222164 620704 222216
rect 631508 222164 631560 222216
rect 160836 222096 160888 222148
rect 166080 222096 166132 222148
rect 97908 221960 97960 222012
rect 172704 222096 172756 222148
rect 174360 222096 174412 222148
rect 167460 221960 167512 222012
rect 175924 221960 175976 222012
rect 181444 222096 181496 222148
rect 182640 222096 182692 222148
rect 191472 222096 191524 222148
rect 247592 222096 247644 222148
rect 258080 222096 258132 222148
rect 263692 222096 263744 222148
rect 270224 222096 270276 222148
rect 306564 222096 306616 222148
rect 310704 222096 310756 222148
rect 312636 222096 312688 222148
rect 331404 222096 331456 222148
rect 353760 222096 353812 222148
rect 452476 222096 452528 222148
rect 455604 222096 455656 222148
rect 462136 222096 462188 222148
rect 468760 222096 468812 222148
rect 471888 222096 471940 222148
rect 477868 222096 477920 222148
rect 495164 222028 495216 222080
rect 497740 222028 497792 222080
rect 515496 222028 515548 222080
rect 529848 222028 529900 222080
rect 533988 222028 534040 222080
rect 536104 222028 536156 222080
rect 539600 222028 539652 222080
rect 539784 222028 539836 222080
rect 232136 221960 232188 222012
rect 233700 221960 233752 222012
rect 277952 221960 278004 222012
rect 280068 221960 280120 222012
rect 313740 221960 313792 222012
rect 318248 221960 318300 222012
rect 343824 221960 343876 222012
rect 367652 221960 367704 222012
rect 380256 221960 380308 222012
rect 424968 221892 425020 221944
rect 429200 221892 429252 221944
rect 559380 221892 559432 221944
rect 559564 221892 559616 221944
rect 564808 221892 564860 221944
rect 104532 221824 104584 221876
rect 173348 221824 173400 221876
rect 173532 221824 173584 221876
rect 181444 221824 181496 221876
rect 181628 221824 181680 221876
rect 240140 221824 240192 221876
rect 263324 221824 263376 221876
rect 301136 221824 301188 221876
rect 301964 221824 302016 221876
rect 310888 221824 310940 221876
rect 313188 221824 313240 221876
rect 340420 221824 340472 221876
rect 351276 221824 351328 221876
rect 369308 221824 369360 221876
rect 509884 221824 509936 221876
rect 522580 221824 522632 221876
rect 596640 221960 596692 222012
rect 605012 221960 605064 222012
rect 600780 221824 600832 221876
rect 600964 221824 601016 221876
rect 606668 221824 606720 221876
rect 80520 221688 80572 221740
rect 86224 221688 86276 221740
rect 94688 221688 94740 221740
rect 161434 221688 161486 221740
rect 161572 221688 161624 221740
rect 167184 221688 167236 221740
rect 167644 221688 167696 221740
rect 169760 221688 169812 221740
rect 171600 221688 171652 221740
rect 232320 221688 232372 221740
rect 239312 221688 239364 221740
rect 283656 221688 283708 221740
rect 303252 221688 303304 221740
rect 332784 221688 332836 221740
rect 357164 221688 357216 221740
rect 374644 221688 374696 221740
rect 391020 221688 391072 221740
rect 400312 221688 400364 221740
rect 475936 221688 475988 221740
rect 486148 221688 486200 221740
rect 496268 221688 496320 221740
rect 513564 221688 513616 221740
rect 524236 221688 524288 221740
rect 539324 221756 539376 221808
rect 539600 221756 539652 221808
rect 547834 221756 547886 221808
rect 547972 221756 548024 221808
rect 549076 221756 549128 221808
rect 549260 221756 549312 221808
rect 552112 221756 552164 221808
rect 552848 221756 552900 221808
rect 553308 221756 553360 221808
rect 608600 221688 608652 221740
rect 59360 221552 59412 221604
rect 141332 221552 141384 221604
rect 141516 221552 141568 221604
rect 147404 221552 147456 221604
rect 147588 221552 147640 221604
rect 205916 221552 205968 221604
rect 208400 221552 208452 221604
rect 260840 221552 260892 221604
rect 261024 221552 261076 221604
rect 301780 221552 301832 221604
rect 308864 221552 308916 221604
rect 339684 221552 339736 221604
rect 341340 221552 341392 221604
rect 361764 221552 361816 221604
rect 369492 221552 369544 221604
rect 384120 221552 384172 221604
rect 384488 221552 384540 221604
rect 395160 221552 395212 221604
rect 400680 221552 400732 221604
rect 405832 221552 405884 221604
rect 480812 221552 480864 221604
rect 492956 221552 493008 221604
rect 497464 221552 497516 221604
rect 515128 221552 515180 221604
rect 522856 221552 522908 221604
rect 546592 221620 546644 221672
rect 547144 221620 547196 221672
rect 553952 221620 554004 221672
rect 539324 221484 539376 221536
rect 547834 221484 547886 221536
rect 547972 221484 548024 221536
rect 552296 221484 552348 221536
rect 596640 221552 596692 221604
rect 596824 221552 596876 221604
rect 633440 221552 633492 221604
rect 73896 221416 73948 221468
rect 82084 221416 82136 221468
rect 86316 221416 86368 221468
rect 91284 221280 91336 221332
rect 118148 221280 118200 221332
rect 127440 221280 127492 221332
rect 161434 221280 161486 221332
rect 161756 221416 161808 221468
rect 164332 221280 164384 221332
rect 173532 221280 173584 221332
rect 175924 221416 175976 221468
rect 226524 221416 226576 221468
rect 227904 221416 227956 221468
rect 276112 221416 276164 221468
rect 292488 221416 292540 221468
rect 326252 221416 326304 221468
rect 342168 221416 342220 221468
rect 364800 221416 364852 221468
rect 375288 221416 375340 221468
rect 390744 221416 390796 221468
rect 396816 221416 396868 221468
rect 407304 221416 407356 221468
rect 408408 221416 408460 221468
rect 416872 221416 416924 221468
rect 468944 221416 468996 221468
rect 476212 221416 476264 221468
rect 483756 221416 483808 221468
rect 538496 221416 538548 221468
rect 538680 221348 538732 221400
rect 553124 221348 553176 221400
rect 600964 221416 601016 221468
rect 193404 221280 193456 221332
rect 204168 221280 204220 221332
rect 252744 221280 252796 221332
rect 266820 221280 266872 221332
rect 303804 221280 303856 221332
rect 600872 221280 600924 221332
rect 604644 221280 604696 221332
rect 521108 221212 521160 221264
rect 600504 221212 600556 221264
rect 111156 221008 111208 221060
rect 118148 221008 118200 221060
rect 124404 221008 124456 221060
rect 127256 221008 127308 221060
rect 127440 221008 127492 221060
rect 166080 221144 166132 221196
rect 221280 221144 221332 221196
rect 222752 221144 222804 221196
rect 268292 221144 268344 221196
rect 523500 221076 523552 221128
rect 601792 221076 601844 221128
rect 127900 221008 127952 221060
rect 83004 220872 83056 220924
rect 147634 221008 147686 221060
rect 206468 221008 206520 221060
rect 219808 221008 219860 221060
rect 263048 221008 263100 221060
rect 525984 220940 526036 220992
rect 602252 220940 602304 220992
rect 161434 220872 161486 220924
rect 161572 220872 161624 220924
rect 222292 220872 222344 220924
rect 282644 220872 282696 220924
rect 287704 220872 287756 220924
rect 456708 220872 456760 220924
rect 147220 220804 147272 220856
rect 253848 220804 253900 220856
rect 258632 220804 258684 220856
rect 418344 220804 418396 220856
rect 424048 220804 424100 220856
rect 462136 220804 462188 220856
rect 466092 220804 466144 220856
rect 471428 220804 471480 220856
rect 517520 220804 517572 220856
rect 518532 220804 518584 220856
rect 600320 220804 600372 220856
rect 114284 220736 114336 220788
rect 146760 220736 146812 220788
rect 101220 220600 101272 220652
rect 147036 220600 147088 220652
rect 180754 220736 180806 220788
rect 181076 220736 181128 220788
rect 190368 220736 190420 220788
rect 190552 220736 190604 220788
rect 236644 220736 236696 220788
rect 242624 220736 242676 220788
rect 246488 220736 246540 220788
rect 260196 220736 260248 220788
rect 298560 220736 298612 220788
rect 321560 220736 321612 220788
rect 324504 220736 324556 220788
rect 385224 220736 385276 220788
rect 388720 220736 388772 220788
rect 414204 220736 414256 220788
rect 418160 220736 418212 220788
rect 455328 220736 455380 220788
rect 458824 220736 458876 220788
rect 474004 220736 474056 220788
rect 475384 220736 475436 220788
rect 476764 220736 476816 220788
rect 478696 220736 478748 220788
rect 511816 220736 511868 220788
rect 465724 220668 465776 220720
rect 469588 220668 469640 220720
rect 69756 220464 69808 220516
rect 136916 220464 136968 220516
rect 137100 220464 137152 220516
rect 147680 220600 147732 220652
rect 175280 220600 175332 220652
rect 177396 220600 177448 220652
rect 180754 220600 180806 220652
rect 180892 220600 180944 220652
rect 224224 220600 224276 220652
rect 253572 220600 253624 220652
rect 293316 220600 293368 220652
rect 302424 220600 302476 220652
rect 334072 220600 334124 220652
rect 357900 220600 357952 220652
rect 374460 220600 374512 220652
rect 500224 220600 500276 220652
rect 511816 220600 511868 220652
rect 147588 220464 147640 220516
rect 150716 220464 150768 220516
rect 150900 220464 150952 220516
rect 73068 220328 73120 220380
rect 147220 220328 147272 220380
rect 147404 220328 147456 220380
rect 151544 220328 151596 220380
rect 151912 220464 151964 220516
rect 211252 220464 211304 220516
rect 214104 220464 214156 220516
rect 214288 220464 214340 220516
rect 218704 220464 218756 220516
rect 220452 220464 220504 220516
rect 267924 220464 267976 220516
rect 273444 220464 273496 220516
rect 309232 220464 309284 220516
rect 338028 220464 338080 220516
rect 359004 220464 359056 220516
rect 432236 220464 432288 220516
rect 434812 220464 434864 220516
rect 469128 220464 469180 220516
rect 474556 220464 474608 220516
rect 488448 220464 488500 220516
rect 501880 220464 501932 220516
rect 545764 220668 545816 220720
rect 547972 220668 548024 220720
rect 558736 220668 558788 220720
rect 562968 220668 563020 220720
rect 563152 220668 563204 220720
rect 566464 220668 566516 220720
rect 566832 220668 566884 220720
rect 567292 220668 567344 220720
rect 520924 220600 520976 220652
rect 537484 220600 537536 220652
rect 550824 220600 550876 220652
rect 558552 220600 558604 220652
rect 568580 220600 568632 220652
rect 569776 220600 569828 220652
rect 569960 220600 570012 220652
rect 572444 220600 572496 220652
rect 572628 220600 572680 220652
rect 610532 220600 610584 220652
rect 531688 220464 531740 220516
rect 548340 220464 548392 220516
rect 598572 220464 598624 220516
rect 600964 220464 601016 220516
rect 611452 220464 611504 220516
rect 213644 220328 213696 220380
rect 79692 220192 79744 220244
rect 151728 220192 151780 220244
rect 151912 220192 151964 220244
rect 154028 220192 154080 220244
rect 154396 220192 154448 220244
rect 158904 220192 158956 220244
rect 164240 220192 164292 220244
rect 223764 220192 223816 220244
rect 224408 220328 224460 220380
rect 265164 220328 265216 220380
rect 267648 220328 267700 220380
rect 306932 220328 306984 220380
rect 314844 220328 314896 220380
rect 341064 220328 341116 220380
rect 342996 220328 343048 220380
rect 363420 220328 363472 220380
rect 472992 220328 473044 220380
rect 481180 220328 481232 220380
rect 496452 220328 496504 220380
rect 509332 220328 509384 220380
rect 516968 220328 517020 220380
rect 527548 220328 527600 220380
rect 531136 220328 531188 220380
rect 556528 220328 556580 220380
rect 234160 220192 234212 220244
rect 237012 220192 237064 220244
rect 280436 220192 280488 220244
rect 283380 220192 283432 220244
rect 316316 220192 316368 220244
rect 316500 220192 316552 220244
rect 342628 220192 342680 220244
rect 348792 220192 348844 220244
rect 369952 220192 370004 220244
rect 370504 220192 370556 220244
rect 381084 220192 381136 220244
rect 388720 220192 388772 220244
rect 400956 220192 401008 220244
rect 459468 220192 459520 220244
rect 465448 220192 465500 220244
rect 473176 220192 473228 220244
rect 482008 220192 482060 220244
rect 482928 220192 482980 220244
rect 495256 220192 495308 220244
rect 501328 220192 501380 220244
rect 520188 220192 520240 220244
rect 528376 220192 528428 220244
rect 554044 220192 554096 220244
rect 555700 220192 555752 220244
rect 558000 220192 558052 220244
rect 76380 220056 76432 220108
rect 156144 220056 156196 220108
rect 157524 220056 157576 220108
rect 214288 220056 214340 220108
rect 107844 219920 107896 219972
rect 114284 219920 114336 219972
rect 114468 219920 114520 219972
rect 121092 219784 121144 219836
rect 127624 219920 127676 219972
rect 180754 219920 180806 219972
rect 180892 219920 180944 219972
rect 213644 219920 213696 219972
rect 137100 219784 137152 219836
rect 127624 219648 127676 219700
rect 131028 219648 131080 219700
rect 197636 219784 197688 219836
rect 197820 219784 197872 219836
rect 244280 220056 244332 220108
rect 244464 220056 244516 220108
rect 288532 220056 288584 220108
rect 288716 220056 288768 220108
rect 322388 220056 322440 220108
rect 325608 220056 325660 220108
rect 352104 220056 352156 220108
rect 358820 220056 358872 220108
rect 378324 220056 378376 220108
rect 379428 220056 379480 220108
rect 392124 220056 392176 220108
rect 395988 220056 396040 220108
rect 404820 220056 404872 220108
rect 421656 220056 421708 220108
rect 426716 220056 426768 220108
rect 478328 220056 478380 220108
rect 489460 220056 489512 220108
rect 492496 220056 492548 220108
rect 506848 220056 506900 220108
rect 513104 220056 513156 220108
rect 534172 220056 534224 220108
rect 538128 220056 538180 220108
rect 563198 220328 563250 220380
rect 563336 220328 563388 220380
rect 609428 220328 609480 220380
rect 558368 220192 558420 220244
rect 562876 220192 562928 220244
rect 563060 220192 563112 220244
rect 608876 220192 608928 220244
rect 648620 220192 648672 220244
rect 652760 220192 652812 220244
rect 572674 220056 572726 220108
rect 558368 219988 558420 220040
rect 572536 219988 572588 220040
rect 214748 219920 214800 219972
rect 254768 219920 254820 219972
rect 294972 219920 295024 219972
rect 325884 219920 325936 219972
rect 598572 220056 598624 220108
rect 607312 220056 607364 220108
rect 676220 220056 676272 220108
rect 677324 220056 677376 220108
rect 600964 219920 601016 219972
rect 503628 219852 503680 219904
rect 589280 219852 589332 219904
rect 589464 219852 589516 219904
rect 596732 219852 596784 219904
rect 136916 219512 136968 219564
rect 137652 219512 137704 219564
rect 142712 219512 142764 219564
rect 143080 219648 143132 219700
rect 203156 219648 203208 219700
rect 144092 219512 144144 219564
rect 144276 219512 144328 219564
rect 208584 219648 208636 219700
rect 210516 219648 210568 219700
rect 259920 219784 259972 219836
rect 540796 219716 540848 219768
rect 606024 219716 606076 219768
rect 217140 219648 217192 219700
rect 224408 219648 224460 219700
rect 227076 219648 227128 219700
rect 272708 219648 272760 219700
rect 464988 219580 465040 219632
rect 472072 219580 472124 219632
rect 527548 219580 527600 219632
rect 558368 219580 558420 219632
rect 558552 219580 558604 219632
rect 600872 219580 600924 219632
rect 203892 219512 203944 219564
rect 214748 219512 214800 219564
rect 224224 219512 224276 219564
rect 229284 219512 229336 219564
rect 332692 219512 332744 219564
rect 337200 219512 337252 219564
rect 109500 219376 109552 219428
rect 110420 219376 110472 219428
rect 113640 219376 113692 219428
rect 156512 219376 156564 219428
rect 165804 219376 165856 219428
rect 70584 219240 70636 219292
rect 117780 219240 117832 219292
rect 131856 219240 131908 219292
rect 132408 219240 132460 219292
rect 132592 219240 132644 219292
rect 136180 219240 136232 219292
rect 136364 219240 136416 219292
rect 170956 219240 171008 219292
rect 175740 219376 175792 219428
rect 181444 219376 181496 219428
rect 183836 219376 183888 219428
rect 190000 219376 190052 219428
rect 192300 219376 192352 219428
rect 224408 219376 224460 219428
rect 229560 219376 229612 219428
rect 230480 219376 230532 219428
rect 237840 219376 237892 219428
rect 239312 219376 239364 219428
rect 239496 219376 239548 219428
rect 405924 219444 405976 219496
rect 412732 219444 412784 219496
rect 241796 219376 241848 219428
rect 241980 219376 242032 219428
rect 242900 219376 242952 219428
rect 244924 219376 244976 219428
rect 272340 219376 272392 219428
rect 272708 219376 272760 219428
rect 180064 219240 180116 219292
rect 180248 219240 180300 219292
rect 215944 219240 215996 219292
rect 219624 219240 219676 219292
rect 264152 219240 264204 219292
rect 285864 219376 285916 219428
rect 301964 219240 302016 219292
rect 308220 219376 308272 219428
rect 309140 219376 309192 219428
rect 333704 219376 333756 219428
rect 347228 219376 347280 219428
rect 349620 219376 349672 219428
rect 350540 219376 350592 219428
rect 352104 219376 352156 219428
rect 355324 219376 355376 219428
rect 362040 219376 362092 219428
rect 367652 219376 367704 219428
rect 380256 219376 380308 219428
rect 384212 219376 384264 219428
rect 399300 219376 399352 219428
rect 400220 219376 400272 219428
rect 415860 219376 415912 219428
rect 416780 219376 416832 219428
rect 417516 219376 417568 219428
rect 421012 219444 421064 219496
rect 432052 219512 432104 219564
rect 501144 219512 501196 219564
rect 428280 219376 428332 219428
rect 589096 219444 589148 219496
rect 620100 219580 620152 219632
rect 438216 219376 438268 219428
rect 438860 219376 438912 219428
rect 439872 219376 439924 219428
rect 440332 219376 440384 219428
rect 572674 219308 572726 219360
rect 601240 219444 601292 219496
rect 607496 219444 607548 219496
rect 313924 219240 313976 219292
rect 320640 219240 320692 219292
rect 342812 219240 342864 219292
rect 419172 219240 419224 219292
rect 422668 219240 422720 219292
rect 548156 219240 548208 219292
rect 563060 219240 563112 219292
rect 563244 219240 563296 219292
rect 574376 219172 574428 219224
rect 589280 219172 589332 219224
rect 597560 219172 597612 219224
rect 64604 219104 64656 219156
rect 66904 219104 66956 219156
rect 93584 219104 93636 219156
rect 94412 219104 94464 219156
rect 117964 219104 118016 219156
rect 154672 219104 154724 219156
rect 62304 218968 62356 219020
rect 72424 218968 72476 219020
rect 83832 218968 83884 219020
rect 157984 219104 158036 219156
rect 166632 219104 166684 219156
rect 208492 219104 208544 219156
rect 208860 219104 208912 219156
rect 209688 219104 209740 219156
rect 218796 219104 218848 219156
rect 219348 219104 219400 219156
rect 224224 219104 224276 219156
rect 253020 219104 253072 219156
rect 265992 219104 266044 219156
rect 156512 218968 156564 219020
rect 162124 218968 162176 219020
rect 162492 218968 162544 219020
rect 175740 218968 175792 219020
rect 176660 218968 176712 219020
rect 180248 218968 180300 219020
rect 182364 218968 182416 219020
rect 189724 218968 189776 219020
rect 190644 218968 190696 219020
rect 197820 218968 197872 219020
rect 200212 218968 200264 219020
rect 241612 218968 241664 219020
rect 241796 218968 241848 219020
rect 244924 218968 244976 219020
rect 252744 218968 252796 219020
rect 287888 218968 287940 219020
rect 295800 219104 295852 219156
rect 296720 219104 296772 219156
rect 314016 219104 314068 219156
rect 336004 219104 336056 219156
rect 343824 219104 343876 219156
rect 353944 219104 353996 219156
rect 542636 219104 542688 219156
rect 297272 218968 297324 219020
rect 307392 218968 307444 219020
rect 332692 218968 332744 219020
rect 337200 218968 337252 219020
rect 345664 218968 345716 219020
rect 347228 218968 347280 219020
rect 363604 218968 363656 219020
rect 368664 218968 368716 219020
rect 377404 218968 377456 219020
rect 63132 218832 63184 218884
rect 75184 218832 75236 218884
rect 77208 218832 77260 218884
rect 150440 218832 150492 218884
rect 152372 218832 152424 218884
rect 153844 218832 153896 218884
rect 154672 218832 154724 218884
rect 159364 218832 159416 218884
rect 159824 218832 159876 218884
rect 203524 218832 203576 218884
rect 206468 218832 206520 218884
rect 253848 218832 253900 218884
rect 259092 218832 259144 218884
rect 59820 218696 59872 218748
rect 140044 218696 140096 218748
rect 140964 218696 141016 218748
rect 142068 218696 142120 218748
rect 142620 218696 142672 218748
rect 143264 218696 143316 218748
rect 146760 218696 146812 218748
rect 184204 218696 184256 218748
rect 186504 218696 186556 218748
rect 192300 218696 192352 218748
rect 192852 218696 192904 218748
rect 243452 218696 243504 218748
rect 253204 218696 253256 218748
rect 286324 218696 286376 218748
rect 291660 218832 291712 218884
rect 291844 218696 291896 218748
rect 300492 218832 300544 218884
rect 327724 218832 327776 218884
rect 340512 218832 340564 218884
rect 358084 218832 358136 218884
rect 363696 218832 363748 218884
rect 370504 218832 370556 218884
rect 376944 218832 376996 218884
rect 382740 218832 382792 218884
rect 383476 218832 383528 218884
rect 386880 218968 386932 219020
rect 398104 218968 398156 219020
rect 547420 218968 547472 219020
rect 562876 219104 562928 219156
rect 563520 219104 563572 219156
rect 572076 219104 572128 219156
rect 388536 218832 388588 218884
rect 402612 218832 402664 218884
rect 409052 218832 409104 218884
rect 411720 218832 411772 218884
rect 412548 218832 412600 218884
rect 512736 218832 512788 218884
rect 321560 218696 321612 218748
rect 327264 218696 327316 218748
rect 351092 218696 351144 218748
rect 353760 218696 353812 218748
rect 369124 218696 369176 218748
rect 370320 218696 370372 218748
rect 380072 218696 380124 218748
rect 383568 218696 383620 218748
rect 396264 218696 396316 218748
rect 412548 218696 412600 218748
rect 417148 218696 417200 218748
rect 429936 218696 429988 218748
rect 432696 218696 432748 218748
rect 482744 218696 482796 218748
rect 485320 218696 485372 218748
rect 500408 218696 500460 218748
rect 508044 218696 508096 218748
rect 517704 218696 517756 218748
rect 518164 218696 518216 218748
rect 520004 218696 520056 218748
rect 548156 218832 548208 218884
rect 557356 218968 557408 219020
rect 614120 218968 614172 219020
rect 562692 218832 562744 218884
rect 563612 218832 563664 218884
rect 572076 218832 572128 218884
rect 574744 218832 574796 218884
rect 603080 218832 603132 218884
rect 537484 218696 537536 218748
rect 563336 218696 563388 218748
rect 564164 218696 564216 218748
rect 598848 218696 598900 218748
rect 100392 218560 100444 218612
rect 146576 218560 146628 218612
rect 148416 218560 148468 218612
rect 148876 218560 148928 218612
rect 149244 218560 149296 218612
rect 150072 218560 150124 218612
rect 150440 218560 150492 218612
rect 152372 218560 152424 218612
rect 152556 218560 152608 218612
rect 153108 218560 153160 218612
rect 153384 218560 153436 218612
rect 154488 218560 154540 218612
rect 155040 218560 155092 218612
rect 155684 218560 155736 218612
rect 156696 218560 156748 218612
rect 157248 218560 157300 218612
rect 159180 218560 159232 218612
rect 160008 218560 160060 218612
rect 160192 218560 160244 218612
rect 186964 218560 187016 218612
rect 188712 218560 188764 218612
rect 193588 218560 193640 218612
rect 195612 218560 195664 218612
rect 198004 218560 198056 218612
rect 198924 218560 198976 218612
rect 200028 218560 200080 218612
rect 204720 218560 204772 218612
rect 207664 218560 207716 218612
rect 107016 218424 107068 218476
rect 117964 218424 118016 218476
rect 120264 218424 120316 218476
rect 166264 218424 166316 218476
rect 170956 218424 171008 218476
rect 176292 218424 176344 218476
rect 179880 218424 179932 218476
rect 204904 218424 204956 218476
rect 117780 218288 117832 218340
rect 123484 218288 123536 218340
rect 130200 218288 130252 218340
rect 136364 218288 136416 218340
rect 136824 218288 136876 218340
rect 174728 218288 174780 218340
rect 175740 218288 175792 218340
rect 179512 218288 179564 218340
rect 180708 218288 180760 218340
rect 185952 218288 186004 218340
rect 189816 218288 189868 218340
rect 195244 218288 195296 218340
rect 198096 218288 198148 218340
rect 123668 218220 123720 218272
rect 55680 218152 55732 218204
rect 56508 218152 56560 218204
rect 57428 218152 57480 218204
rect 61384 218152 61436 218204
rect 66444 218152 66496 218204
rect 67548 218152 67600 218204
rect 68100 218152 68152 218204
rect 69572 218152 69624 218204
rect 75552 218152 75604 218204
rect 76564 218152 76616 218204
rect 97080 218152 97132 218204
rect 56508 218016 56560 218068
rect 57244 218016 57296 218068
rect 58164 218016 58216 218068
rect 59360 218016 59412 218068
rect 61476 218016 61528 218068
rect 62764 218016 62816 218068
rect 63960 218016 64012 218068
rect 64788 218016 64840 218068
rect 65616 218016 65668 218068
rect 66168 218016 66220 218068
rect 67272 218016 67324 218068
rect 68284 218016 68336 218068
rect 72240 218016 72292 218068
rect 73712 218016 73764 218068
rect 74724 218016 74776 218068
rect 75828 218016 75880 218068
rect 78036 218016 78088 218068
rect 78588 218016 78640 218068
rect 78864 218016 78916 218068
rect 79968 218016 80020 218068
rect 82176 218016 82228 218068
rect 83464 218016 83516 218068
rect 84660 218016 84712 218068
rect 85304 218016 85356 218068
rect 87144 218016 87196 218068
rect 88248 218016 88300 218068
rect 88800 218016 88852 218068
rect 89444 218016 89496 218068
rect 92940 218016 92992 218068
rect 93768 218016 93820 218068
rect 95424 218016 95476 218068
rect 96252 218016 96304 218068
rect 98736 218016 98788 218068
rect 99288 218016 99340 218068
rect 99564 218016 99616 218068
rect 100668 218016 100720 218068
rect 117780 218152 117832 218204
rect 118700 218152 118752 218204
rect 132500 218152 132552 218204
rect 140136 218152 140188 218204
rect 175924 218152 175976 218204
rect 102876 218084 102928 218136
rect 103428 218084 103480 218136
rect 103704 218084 103756 218136
rect 104808 218084 104860 218136
rect 105360 218084 105412 218136
rect 106004 218084 106056 218136
rect 111984 218084 112036 218136
rect 112812 218084 112864 218136
rect 116124 218084 116176 218136
rect 117228 218084 117280 218136
rect 119436 218084 119488 218136
rect 119988 218084 120040 218136
rect 121920 218084 121972 218136
rect 122564 218084 122616 218136
rect 126060 218084 126112 218136
rect 126704 218084 126756 218136
rect 127716 218084 127768 218136
rect 128268 218084 128320 218136
rect 128544 218084 128596 218136
rect 129372 218084 129424 218136
rect 132684 218084 132736 218136
rect 133512 218084 133564 218136
rect 135996 218084 136048 218136
rect 136548 218084 136600 218136
rect 161664 218016 161716 218068
rect 162768 218016 162820 218068
rect 163320 218016 163372 218068
rect 163964 218016 164016 218068
rect 164976 218016 165028 218068
rect 165528 218016 165580 218068
rect 169116 218016 169168 218068
rect 169576 218016 169628 218068
rect 169944 218016 169996 218068
rect 170772 218016 170824 218068
rect 172428 218016 172480 218068
rect 173164 218016 173216 218068
rect 173348 218016 173400 218068
rect 174084 217880 174136 217932
rect 174728 218016 174780 218068
rect 178684 218152 178736 218204
rect 179052 218152 179104 218204
rect 196624 218152 196676 218204
rect 199752 218152 199804 218204
rect 200212 218152 200264 218204
rect 200672 218288 200724 218340
rect 214288 218560 214340 218612
rect 214748 218560 214800 218612
rect 219808 218560 219860 218612
rect 225972 218560 226024 218612
rect 267004 218560 267056 218612
rect 272340 218560 272392 218612
rect 279424 218560 279476 218612
rect 208492 218424 208544 218476
rect 211804 218424 211856 218476
rect 213000 218424 213052 218476
rect 224224 218424 224276 218476
rect 224408 218424 224460 218476
rect 231032 218424 231084 218476
rect 209688 218288 209740 218340
rect 213184 218288 213236 218340
rect 214288 218288 214340 218340
rect 204168 218152 204220 218204
rect 204904 218152 204956 218204
rect 210332 218152 210384 218204
rect 211344 218152 211396 218204
rect 214472 218152 214524 218204
rect 216312 218288 216364 218340
rect 238024 218424 238076 218476
rect 232872 218288 232924 218340
rect 271144 218424 271196 218476
rect 279240 218424 279292 218476
rect 305552 218560 305604 218612
rect 398472 218560 398524 218612
rect 407764 218560 407816 218612
rect 469864 218560 469916 218612
rect 471244 218560 471296 218612
rect 475568 218560 475620 218612
rect 482836 218560 482888 218612
rect 507676 218560 507728 218612
rect 563198 218560 563250 218612
rect 572812 218560 572864 218612
rect 610716 218560 610768 218612
rect 568304 218492 568356 218544
rect 572444 218492 572496 218544
rect 294144 218424 294196 218476
rect 316684 218424 316736 218476
rect 502800 218424 502852 218476
rect 503168 218424 503220 218476
rect 507860 218424 507912 218476
rect 508044 218424 508096 218476
rect 458180 218356 458232 218408
rect 574928 218424 574980 218476
rect 604460 218424 604512 218476
rect 241612 218288 241664 218340
rect 246304 218288 246356 218340
rect 249432 218288 249484 218340
rect 251732 218288 251784 218340
rect 253020 218288 253072 218340
rect 258080 218288 258132 218340
rect 426624 218288 426676 218340
rect 429384 218288 429436 218340
rect 450728 218288 450780 218340
rect 453856 218288 453908 218340
rect 572076 218356 572128 218408
rect 461308 218288 461360 218340
rect 497464 218288 497516 218340
rect 572812 218288 572864 218340
rect 594800 218288 594852 218340
rect 668400 218288 668452 218340
rect 669504 218288 669556 218340
rect 572536 218220 572588 218272
rect 176660 218016 176712 218068
rect 178224 218016 178276 218068
rect 179328 218016 179380 218068
rect 179512 218016 179564 218068
rect 183836 218016 183888 218068
rect 184020 218016 184072 218068
rect 184664 218016 184716 218068
rect 185676 218016 185728 218068
rect 186136 218016 186188 218068
rect 188160 218016 188212 218068
rect 188896 218016 188948 218068
rect 192300 218016 192352 218068
rect 193036 218016 193088 218068
rect 193956 218016 194008 218068
rect 194508 218016 194560 218068
rect 194784 218016 194836 218068
rect 195888 218016 195940 218068
rect 196440 218016 196492 218068
rect 200396 218016 200448 218068
rect 200580 218016 200632 218068
rect 201500 218016 201552 218068
rect 203064 218016 203116 218068
rect 206284 218016 206336 218068
rect 207204 218016 207256 218068
rect 208124 218016 208176 218068
rect 214656 218016 214708 218068
rect 215208 218016 215260 218068
rect 215484 218016 215536 218068
rect 216496 218016 216548 218068
rect 217968 218152 218020 218204
rect 222752 218152 222804 218204
rect 222936 218152 222988 218204
rect 225604 218152 225656 218204
rect 246120 218152 246172 218204
rect 253204 218152 253256 218204
rect 328920 218152 328972 218204
rect 330484 218152 330536 218204
rect 365352 218152 365404 218204
rect 371792 218152 371844 218204
rect 374460 218152 374512 218204
rect 376024 218152 376076 218204
rect 381912 218152 381964 218204
rect 382924 218152 382976 218204
rect 401784 218152 401836 218204
rect 402796 218152 402848 218204
rect 407580 218152 407632 218204
rect 411904 218152 411956 218204
rect 422484 218152 422536 218204
rect 425428 218152 425480 218204
rect 425796 218152 425848 218204
rect 427912 218152 427964 218204
rect 433248 218152 433300 218204
rect 434720 218152 434772 218204
rect 434904 218152 434956 218204
rect 436836 218152 436888 218204
rect 461952 218152 462004 218204
rect 466276 218152 466328 218204
rect 491944 218152 491996 218204
rect 502248 218152 502300 218204
rect 507124 218152 507176 218204
rect 507676 218152 507728 218204
rect 507860 218152 507912 218204
rect 562876 218152 562928 218204
rect 572996 218152 573048 218204
rect 220084 218016 220136 218068
rect 221280 218016 221332 218068
rect 221832 218016 221884 218068
rect 223764 218016 223816 218068
rect 224592 218016 224644 218068
rect 225420 218016 225472 218068
rect 226156 218016 226208 218068
rect 231216 218016 231268 218068
rect 231676 218016 231728 218068
rect 232044 218016 232096 218068
rect 233148 218016 233200 218068
rect 235356 218016 235408 218068
rect 235816 218016 235868 218068
rect 236184 218016 236236 218068
rect 237288 218016 237340 218068
rect 240324 218016 240376 218068
rect 241336 218016 241388 218068
rect 243636 218016 243688 218068
rect 244096 218016 244148 218068
rect 247776 218016 247828 218068
rect 248236 218016 248288 218068
rect 248604 218016 248656 218068
rect 249616 218016 249668 218068
rect 250260 218016 250312 218068
rect 250904 218016 250956 218068
rect 251916 218016 251968 218068
rect 252468 218016 252520 218068
rect 254400 218016 254452 218068
rect 255044 218016 255096 218068
rect 256056 218016 256108 218068
rect 256516 218016 256568 218068
rect 256884 218016 256936 218068
rect 257528 218016 257580 218068
rect 258540 218016 258592 218068
rect 259276 218016 259328 218068
rect 262680 218016 262732 218068
rect 263600 218016 263652 218068
rect 264336 218016 264388 218068
rect 264796 218016 264848 218068
rect 265164 218016 265216 218068
rect 266176 218016 266228 218068
rect 268476 218016 268528 218068
rect 268936 218016 268988 218068
rect 269304 218016 269356 218068
rect 270040 218016 270092 218068
rect 270960 218016 271012 218068
rect 272524 218016 272576 218068
rect 276756 218016 276808 218068
rect 277216 218016 277268 218068
rect 277584 218016 277636 218068
rect 278596 218016 278648 218068
rect 280896 218016 280948 218068
rect 281448 218016 281500 218068
rect 281724 218016 281776 218068
rect 282460 218016 282512 218068
rect 285036 218016 285088 218068
rect 285496 218016 285548 218068
rect 287520 218016 287572 218068
rect 288716 218016 288768 218068
rect 289176 218016 289228 218068
rect 289728 218016 289780 218068
rect 290004 218016 290056 218068
rect 291108 218016 291160 218068
rect 293316 218016 293368 218068
rect 293776 218016 293828 218068
rect 297456 218016 297508 218068
rect 297916 218016 297968 218068
rect 298284 218016 298336 218068
rect 299112 218016 299164 218068
rect 299940 218016 299992 218068
rect 300676 218016 300728 218068
rect 301596 218016 301648 218068
rect 302148 218016 302200 218068
rect 304080 218016 304132 218068
rect 304724 218016 304776 218068
rect 305736 218016 305788 218068
rect 306196 218016 306248 218068
rect 306564 218016 306616 218068
rect 307668 218016 307720 218068
rect 309876 218016 309928 218068
rect 310428 218016 310480 218068
rect 312360 218016 312412 218068
rect 312912 218016 312964 218068
rect 317328 218016 317380 218068
rect 317972 218016 318024 218068
rect 318984 218016 319036 218068
rect 319812 218016 319864 218068
rect 322296 218016 322348 218068
rect 322848 218016 322900 218068
rect 323124 218016 323176 218068
rect 324136 218016 324188 218068
rect 324780 218016 324832 218068
rect 325424 218016 325476 218068
rect 326436 218016 326488 218068
rect 326896 218016 326948 218068
rect 330576 218016 330628 218068
rect 331036 218016 331088 218068
rect 333060 218016 333112 218068
rect 333888 218016 333940 218068
rect 334716 218016 334768 218068
rect 335176 218016 335228 218068
rect 335544 218016 335596 218068
rect 338672 218016 338724 218068
rect 338856 218016 338908 218068
rect 339408 218016 339460 218068
rect 339684 218016 339736 218068
rect 340696 218016 340748 218068
rect 345480 218016 345532 218068
rect 347044 218016 347096 218068
rect 347964 218016 348016 218068
rect 349068 218016 349120 218068
rect 355416 218016 355468 218068
rect 355876 218016 355928 218068
rect 356244 218016 356296 218068
rect 356980 218016 357032 218068
rect 359556 218016 359608 218068
rect 360108 218016 360160 218068
rect 360384 218016 360436 218068
rect 361028 218016 361080 218068
rect 364524 218016 364576 218068
rect 365536 218016 365588 218068
rect 366180 218016 366232 218068
rect 366732 218016 366784 218068
rect 367836 218016 367888 218068
rect 368388 218016 368440 218068
rect 371976 218016 372028 218068
rect 372528 218016 372580 218068
rect 372804 218016 372856 218068
rect 373448 218016 373500 218068
rect 376116 218016 376168 218068
rect 376668 218016 376720 218068
rect 378600 218016 378652 218068
rect 379244 218016 379296 218068
rect 381084 218016 381136 218068
rect 382096 218016 382148 218068
rect 389364 218016 389416 218068
rect 390008 218016 390060 218068
rect 392676 218016 392728 218068
rect 393136 218016 393188 218068
rect 393504 218016 393556 218068
rect 394516 218016 394568 218068
rect 395160 218016 395212 218068
rect 395804 218016 395856 218068
rect 397644 218016 397696 218068
rect 400680 218016 400732 218068
rect 400956 218016 401008 218068
rect 402244 218016 402296 218068
rect 403440 218016 403492 218068
rect 403992 218016 404044 218068
rect 405096 218016 405148 218068
rect 405556 218016 405608 218068
rect 409236 218016 409288 218068
rect 409788 218016 409840 218068
rect 410064 218016 410116 218068
rect 410708 218016 410760 218068
rect 413376 218016 413428 218068
rect 413836 218016 413888 218068
rect 420000 218016 420052 218068
rect 420920 218016 420972 218068
rect 424140 218016 424192 218068
rect 426992 218016 427044 218068
rect 427452 218016 427504 218068
rect 428464 218016 428516 218068
rect 429108 218016 429160 218068
rect 430580 218016 430632 218068
rect 432420 218016 432472 218068
rect 433800 218016 433852 218068
rect 435732 218016 435784 218068
rect 436284 218016 436336 218068
rect 436468 218016 436520 218068
rect 437756 218016 437808 218068
rect 453304 218016 453356 218068
rect 455420 218016 455472 218068
rect 455604 218016 455656 218068
rect 457168 218016 457220 218068
rect 463148 218016 463200 218068
rect 464620 218016 464672 218068
rect 467288 218016 467340 218068
rect 467932 218016 467984 218068
rect 471428 218016 471480 218068
rect 472900 218016 472952 218068
rect 490380 218016 490432 218068
rect 497004 218016 497056 218068
rect 497464 218016 497516 218068
rect 563612 217948 563664 218000
rect 571892 217948 571944 218000
rect 612280 217948 612332 218000
rect 614488 217948 614540 218000
rect 451372 217812 451424 217864
rect 452200 217812 452252 217864
rect 523040 217812 523092 217864
rect 524236 217812 524288 217864
rect 536380 217812 536432 217864
rect 604000 217812 604052 217864
rect 527824 217676 527876 217728
rect 528376 217676 528428 217728
rect 603264 217676 603316 217728
rect 604460 217676 604512 217728
rect 614304 217676 614356 217728
rect 116952 217540 117004 217592
rect 189172 217540 189224 217592
rect 533436 217540 533488 217592
rect 536380 217540 536432 217592
rect 542360 217540 542412 217592
rect 543280 217540 543332 217592
rect 606208 217540 606260 217592
rect 614120 217540 614172 217592
rect 626632 217540 626684 217592
rect 669872 217472 669924 217524
rect 115296 217404 115348 217456
rect 187976 217404 188028 217456
rect 530952 217404 531004 217456
rect 90410 217200 90462 217252
rect 168564 217268 168616 217320
rect 508596 217268 508648 217320
rect 563014 217268 563066 217320
rect 563152 217268 563204 217320
rect 572536 217268 572588 217320
rect 572720 217268 572772 217320
rect 598480 217268 598532 217320
rect 447140 217200 447192 217252
rect 448106 217200 448158 217252
rect 448612 217200 448664 217252
rect 449762 217200 449814 217252
rect 469312 217200 469364 217252
rect 470462 217200 470514 217252
rect 498200 217200 498252 217252
rect 499442 217200 499494 217252
rect 506066 217132 506118 217184
rect 597928 217132 597980 217184
rect 603080 217404 603132 217456
rect 628288 217404 628340 217456
rect 598848 217268 598900 217320
rect 622400 217268 622452 217320
rect 603448 217132 603500 217184
rect 498614 217064 498666 217116
rect 669872 217064 669924 217116
rect 574192 216996 574244 217048
rect 610072 216996 610124 217048
rect 596364 216860 596416 216912
rect 594800 216724 594852 216776
rect 613384 216860 613436 216912
rect 610716 216724 610768 216776
rect 615684 216724 615736 216776
rect 648252 216656 648304 216708
rect 650644 216656 650696 216708
rect 644940 215908 644992 215960
rect 658924 215908 658976 215960
rect 675852 215160 675904 215212
rect 676772 215160 676824 215212
rect 574744 214820 574796 214872
rect 616880 214820 616932 214872
rect 574560 214684 574612 214736
rect 623320 214684 623372 214736
rect 658188 214684 658240 214736
rect 665824 214684 665876 214736
rect 574376 214548 574428 214600
rect 600504 214412 600556 214464
rect 601240 214412 601292 214464
rect 618260 214548 618312 214600
rect 618904 214548 618956 214600
rect 619916 214548 619968 214600
rect 620560 214548 620612 214600
rect 623964 214548 624016 214600
rect 624424 214412 624476 214464
rect 625252 214548 625304 214600
rect 626080 214548 626132 214600
rect 630036 214548 630088 214600
rect 632888 214548 632940 214600
rect 646320 214548 646372 214600
rect 656164 214548 656216 214600
rect 629392 214412 629444 214464
rect 35808 214072 35860 214124
rect 39764 214072 39816 214124
rect 645860 213868 645912 213920
rect 646504 213868 646556 213920
rect 654600 213868 654652 213920
rect 657544 213868 657596 213920
rect 663156 213868 663208 213920
rect 663708 213868 663760 213920
rect 653220 213732 653272 213784
rect 654784 213732 654836 213784
rect 648620 213392 648672 213444
rect 649264 213392 649316 213444
rect 654140 213392 654192 213444
rect 654784 213392 654836 213444
rect 656532 213392 656584 213444
rect 664628 213392 664680 213444
rect 643836 213324 643888 213376
rect 653404 213256 653456 213308
rect 575480 213188 575532 213240
rect 594800 213188 594852 213240
rect 645492 213120 645544 213172
rect 660764 213188 660816 213240
rect 632704 212984 632756 213036
rect 634360 212984 634412 213036
rect 650460 212712 650512 212764
rect 651288 212712 651340 212764
rect 664260 212712 664312 212764
rect 665088 212712 665140 212764
rect 35808 212644 35860 212696
rect 39856 212644 39908 212696
rect 592684 212644 592736 212696
rect 641720 212644 641772 212696
rect 591304 212508 591356 212560
rect 639880 212508 639932 212560
rect 35808 211420 35860 211472
rect 40132 211420 40184 211472
rect 35624 211148 35676 211200
rect 40776 211148 40828 211200
rect 578516 211148 578568 211200
rect 580908 211148 580960 211200
rect 600320 210060 600372 210112
rect 600688 210060 600740 210112
rect 35808 209788 35860 209840
rect 39212 209788 39264 209840
rect 579528 209788 579580 209840
rect 582288 209788 582340 209840
rect 35808 208632 35860 208684
rect 39948 208632 40000 208684
rect 581644 208564 581696 208616
rect 632152 209516 632204 209568
rect 652024 209516 652076 209568
rect 667020 209040 667072 209092
rect 35624 208360 35676 208412
rect 40960 208360 41012 208412
rect 578884 208292 578936 208344
rect 589464 208292 589516 208344
rect 35808 207136 35860 207188
rect 40960 207136 41012 207188
rect 580908 206864 580960 206916
rect 589464 206864 589516 206916
rect 35808 205776 35860 205828
rect 41696 205776 41748 205828
rect 579528 205776 579580 205828
rect 581000 205776 581052 205828
rect 42064 205504 42116 205556
rect 43352 205504 43404 205556
rect 582288 205504 582340 205556
rect 589464 205504 589516 205556
rect 35808 204620 35860 204672
rect 41696 204484 41748 204536
rect 35808 204280 35860 204332
rect 39396 204280 39448 204332
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 35808 202852 35860 202904
rect 39304 202852 39356 202904
rect 578332 202852 578384 202904
rect 580264 202852 580316 202904
rect 581000 202784 581052 202836
rect 589464 202784 589516 202836
rect 578792 200132 578844 200184
rect 590384 200132 590436 200184
rect 580264 199996 580316 200048
rect 589464 199996 589516 200048
rect 579528 198704 579580 198756
rect 589464 198704 589516 198756
rect 42708 197072 42760 197124
rect 43352 197072 43404 197124
rect 578516 195984 578568 196036
rect 589280 195984 589332 196036
rect 579528 194556 579580 194608
rect 589464 194556 589516 194608
rect 579528 191836 579580 191888
rect 589464 191836 589516 191888
rect 579528 190476 579580 190528
rect 590568 190476 590620 190528
rect 579528 187688 579580 187740
rect 589464 187688 589516 187740
rect 42432 187280 42484 187332
rect 43076 187280 43128 187332
rect 579528 186260 579580 186312
rect 589648 186260 589700 186312
rect 579528 184832 579580 184884
rect 589464 184832 589516 184884
rect 668952 184832 669004 184884
rect 670700 184832 670752 184884
rect 42432 182112 42484 182164
rect 43260 182112 43312 182164
rect 579528 182112 579580 182164
rect 589464 182112 589516 182164
rect 578792 180752 578844 180804
rect 590568 180752 590620 180804
rect 578792 178032 578844 178084
rect 589464 178032 589516 178084
rect 668216 177964 668268 178016
rect 670792 177964 670844 178016
rect 579528 177896 579580 177948
rect 589648 177896 589700 177948
rect 579988 175244 580040 175296
rect 589464 175312 589516 175364
rect 668032 175040 668084 175092
rect 670424 175040 670476 175092
rect 578424 174496 578476 174548
rect 589648 174496 589700 174548
rect 578240 172864 578292 172916
rect 579988 172864 580040 172916
rect 580908 172524 580960 172576
rect 589464 172524 589516 172576
rect 580264 171096 580316 171148
rect 589464 171096 589516 171148
rect 578700 169736 578752 169788
rect 580908 169736 580960 169788
rect 667940 169668 667992 169720
rect 669688 169668 669740 169720
rect 582380 168376 582432 168428
rect 589464 168376 589516 168428
rect 578240 167288 578292 167340
rect 580264 167288 580316 167340
rect 579988 167016 580040 167068
rect 589464 167016 589516 167068
rect 579528 166268 579580 166320
rect 589648 166268 589700 166320
rect 579344 165180 579396 165232
rect 582380 165180 582432 165232
rect 667940 165044 667992 165096
rect 670056 165044 670108 165096
rect 582472 164228 582524 164280
rect 589464 164228 589516 164280
rect 675852 164160 675904 164212
rect 682384 164160 682436 164212
rect 578240 163616 578292 163668
rect 579988 163616 580040 163668
rect 580908 162868 580960 162920
rect 589464 162868 589516 162920
rect 578424 162664 578476 162716
rect 582472 162664 582524 162716
rect 580540 161440 580592 161492
rect 589464 161440 589516 161492
rect 580724 160080 580776 160132
rect 589464 160080 589516 160132
rect 668216 160012 668268 160064
rect 670792 160012 670844 160064
rect 578884 158720 578936 158772
rect 580908 158720 580960 158772
rect 585784 158720 585836 158772
rect 589464 158720 589516 158772
rect 587164 157360 587216 157412
rect 589280 157360 589332 157412
rect 668216 155524 668268 155576
rect 670792 155524 670844 155576
rect 578332 154640 578384 154692
rect 580540 154640 580592 154692
rect 584404 154572 584456 154624
rect 589464 154572 589516 154624
rect 583024 153212 583076 153264
rect 589464 153212 589516 153264
rect 578240 152736 578292 152788
rect 580724 152736 580776 152788
rect 580264 151784 580316 151836
rect 589464 151784 589516 151836
rect 578884 150560 578936 150612
rect 585784 150560 585836 150612
rect 585140 149064 585192 149116
rect 589464 149064 589516 149116
rect 579528 148316 579580 148368
rect 587164 148316 587216 148368
rect 578884 146276 578936 146328
rect 585140 146276 585192 146328
rect 668768 145732 668820 145784
rect 670792 145732 670844 145784
rect 584772 144916 584824 144968
rect 589464 144916 589516 144968
rect 579252 144644 579304 144696
rect 584404 144644 584456 144696
rect 585968 143556 586020 143608
rect 589464 143556 589516 143608
rect 579528 143420 579580 143472
rect 583024 143420 583076 143472
rect 587164 142400 587216 142452
rect 589832 142400 589884 142452
rect 580448 140768 580500 140820
rect 589464 140768 589516 140820
rect 578608 140700 578660 140752
rect 580264 140700 580316 140752
rect 583024 139408 583076 139460
rect 589464 139408 589516 139460
rect 578608 139272 578660 139324
rect 589924 139272 589976 139324
rect 579528 138660 579580 138712
rect 588544 138660 588596 138712
rect 579068 137300 579120 137352
rect 584772 137300 584824 137352
rect 584588 136620 584640 136672
rect 589464 136620 589516 136672
rect 580264 134512 580316 134564
rect 589464 134512 589516 134564
rect 675852 133900 675904 133952
rect 676496 133900 676548 133952
rect 667940 133764 667992 133816
rect 669872 133764 669924 133816
rect 585784 132472 585836 132524
rect 589464 132472 589516 132524
rect 581828 131248 581880 131300
rect 589464 131248 589516 131300
rect 578884 131112 578936 131164
rect 585968 131112 586020 131164
rect 668584 130772 668636 130824
rect 670792 130772 670844 130824
rect 668032 129684 668084 129736
rect 670148 129684 670200 129736
rect 583208 129140 583260 129192
rect 590384 129140 590436 129192
rect 579528 129004 579580 129056
rect 587164 129004 587216 129056
rect 579068 126964 579120 127016
rect 589464 126964 589516 127016
rect 578332 125604 578384 125656
rect 580448 125604 580500 125656
rect 675852 125400 675904 125452
rect 676404 125400 676456 125452
rect 580448 124176 580500 124228
rect 589464 124176 589516 124228
rect 578424 123564 578476 123616
rect 583024 123564 583076 123616
rect 584404 122816 584456 122868
rect 589464 122816 589516 122868
rect 578884 122136 578936 122188
rect 584588 122136 584640 122188
rect 580632 122000 580684 122052
rect 589924 122000 589976 122052
rect 587348 118668 587400 118720
rect 590016 118668 590068 118720
rect 675944 118600 675996 118652
rect 679624 118600 679676 118652
rect 578516 118396 578568 118448
rect 580264 118396 580316 118448
rect 579528 116900 579580 116952
rect 583208 116900 583260 116952
rect 668768 116696 668820 116748
rect 670424 116696 670476 116748
rect 586152 115948 586204 116000
rect 589464 115948 589516 116000
rect 583208 115200 583260 115252
rect 589648 115200 589700 115252
rect 579252 114452 579304 114504
rect 581644 114452 581696 114504
rect 583024 113160 583076 113212
rect 589464 113160 589516 113212
rect 579528 112820 579580 112872
rect 585784 112820 585836 112872
rect 585968 112412 586020 112464
rect 590108 112412 590160 112464
rect 581644 110440 581696 110492
rect 589464 110440 589516 110492
rect 579344 110100 579396 110152
rect 581828 110100 581880 110152
rect 584588 109012 584640 109064
rect 589280 109012 589332 109064
rect 667940 108808 667992 108860
rect 669964 108808 670016 108860
rect 578332 108672 578384 108724
rect 580632 108672 580684 108724
rect 578884 107584 578936 107636
rect 589464 107652 589516 107704
rect 587164 106292 587216 106344
rect 589832 106292 589884 106344
rect 668400 106156 668452 106208
rect 670792 106156 670844 106208
rect 580264 104864 580316 104916
rect 589464 104864 589516 104916
rect 668768 104660 668820 104712
rect 670792 104660 670844 104712
rect 579528 103436 579580 103488
rect 588544 103436 588596 103488
rect 579528 101804 579580 101856
rect 584404 101804 584456 101856
rect 584404 100104 584456 100156
rect 589464 100104 589516 100156
rect 579068 99356 579120 99408
rect 586152 99356 586204 99408
rect 622308 99288 622360 99340
rect 630772 99288 630824 99340
rect 578608 99220 578660 99272
rect 580448 99220 580500 99272
rect 623688 99152 623740 99204
rect 633440 99152 633492 99204
rect 577504 99084 577556 99136
rect 595260 99084 595312 99136
rect 625068 99016 625120 99068
rect 636292 99016 636344 99068
rect 628288 98880 628340 98932
rect 642180 98880 642232 98932
rect 629024 98744 629076 98796
rect 643652 98744 643704 98796
rect 647148 98744 647200 98796
rect 661960 98744 662012 98796
rect 630496 98608 630548 98660
rect 646596 98608 646648 98660
rect 578332 97928 578384 97980
rect 587348 97928 587400 97980
rect 620192 97928 620244 97980
rect 626264 97928 626316 97980
rect 629760 97928 629812 97980
rect 645308 98200 645360 98252
rect 618720 97792 618772 97844
rect 625804 97792 625856 97844
rect 627552 97792 627604 97844
rect 640708 97996 640760 98048
rect 659936 97928 659988 97980
rect 665548 97928 665600 97980
rect 632704 97792 632756 97844
rect 648252 97792 648304 97844
rect 655428 97792 655480 97844
rect 662512 97792 662564 97844
rect 631968 97656 632020 97708
rect 647516 97656 647568 97708
rect 650368 97656 650420 97708
rect 658280 97656 658332 97708
rect 621664 97520 621716 97572
rect 629300 97520 629352 97572
rect 634176 97520 634228 97572
rect 650552 97520 650604 97572
rect 656624 97520 656676 97572
rect 659844 97656 659896 97708
rect 659200 97520 659252 97572
rect 664168 97520 664220 97572
rect 612648 97384 612700 97436
rect 618904 97384 618956 97436
rect 623136 97384 623188 97436
rect 632060 97384 632112 97436
rect 633256 97384 633308 97436
rect 648620 97384 648672 97436
rect 651840 97384 651892 97436
rect 659568 97384 659620 97436
rect 605472 97248 605524 97300
rect 611912 97248 611964 97300
rect 626816 97248 626868 97300
rect 639236 97248 639288 97300
rect 643008 97248 643060 97300
rect 656624 97248 656676 97300
rect 656808 97248 656860 97300
rect 661408 97248 661460 97300
rect 626080 97112 626132 97164
rect 637764 97112 637816 97164
rect 644296 97112 644348 97164
rect 658832 97112 658884 97164
rect 624608 96976 624660 97028
rect 635004 96976 635056 97028
rect 635556 96976 635608 97028
rect 647700 96976 647752 97028
rect 596180 96908 596232 96960
rect 596732 96908 596784 96960
rect 597652 96908 597704 96960
rect 598204 96908 598256 96960
rect 600320 96908 600372 96960
rect 601148 96908 601200 96960
rect 601700 96908 601752 96960
rect 602620 96908 602672 96960
rect 606208 96908 606260 96960
rect 607128 96908 607180 96960
rect 613568 96908 613620 96960
rect 613936 96908 613988 96960
rect 615776 96908 615828 96960
rect 616788 96908 616840 96960
rect 656716 96908 656768 96960
rect 660120 96908 660172 96960
rect 612096 96840 612148 96892
rect 612648 96840 612700 96892
rect 634728 96840 634780 96892
rect 650368 96840 650420 96892
rect 653956 96840 654008 96892
rect 654600 96840 654652 96892
rect 654784 96840 654836 96892
rect 655428 96840 655480 96892
rect 658096 96772 658148 96824
rect 663064 96772 663116 96824
rect 610624 96704 610676 96756
rect 611268 96704 611320 96756
rect 617248 96704 617300 96756
rect 618076 96704 618128 96756
rect 640524 96568 640576 96620
rect 647884 96704 647936 96756
rect 645768 96568 645820 96620
rect 656348 96568 656400 96620
rect 639052 96432 639104 96484
rect 645124 96432 645176 96484
rect 646412 96432 646464 96484
rect 652024 96432 652076 96484
rect 652576 96432 652628 96484
rect 665364 96432 665416 96484
rect 631232 96296 631284 96348
rect 647148 96296 647200 96348
rect 648896 96296 648948 96348
rect 664352 96296 664404 96348
rect 637580 96160 637632 96212
rect 660672 96160 660724 96212
rect 611084 96024 611136 96076
rect 622308 96024 622360 96076
rect 649908 96024 649960 96076
rect 663800 96024 663852 96076
rect 644940 95956 644992 96008
rect 649540 95956 649592 96008
rect 607680 95888 607732 95940
rect 624976 95888 625028 95940
rect 643468 95820 643520 95872
rect 649264 95820 649316 95872
rect 665180 95888 665232 95940
rect 638592 95684 638644 95736
rect 647332 95684 647384 95736
rect 647884 95684 647936 95736
rect 653312 95616 653364 95668
rect 663984 95616 664036 95668
rect 640064 95548 640116 95600
rect 647884 95548 647936 95600
rect 641536 95412 641588 95464
rect 645124 95412 645176 95464
rect 651840 95412 651892 95464
rect 649908 95276 649960 95328
rect 620928 95140 620980 95192
rect 626448 95140 626500 95192
rect 647700 95072 647752 95124
rect 648804 95072 648856 95124
rect 579528 95004 579580 95056
rect 583208 95004 583260 95056
rect 616512 95004 616564 95056
rect 622952 95004 623004 95056
rect 609152 94460 609204 94512
rect 620284 94460 620336 94512
rect 619548 93780 619600 93832
rect 626448 93780 626500 93832
rect 651288 93508 651340 93560
rect 655428 93508 655480 93560
rect 578516 93440 578568 93492
rect 585968 93440 586020 93492
rect 611268 93100 611320 93152
rect 619272 93100 619324 93152
rect 649540 92964 649592 93016
rect 656164 92964 656216 93016
rect 606944 92828 606996 92880
rect 610072 92828 610124 92880
rect 648620 92488 648672 92540
rect 650000 92488 650052 92540
rect 617892 92420 617944 92472
rect 626448 92420 626500 92472
rect 647332 92352 647384 92404
rect 654324 92352 654376 92404
rect 579344 91060 579396 91112
rect 584588 91060 584640 91112
rect 618076 90992 618128 91044
rect 626448 90992 626500 91044
rect 651840 90652 651892 90704
rect 655428 90652 655480 90704
rect 622952 89632 623004 89684
rect 626448 89564 626500 89616
rect 585140 88952 585192 89004
rect 589924 88952 589976 89004
rect 649724 88748 649776 88800
rect 658556 88748 658608 88800
rect 662328 88748 662380 88800
rect 664168 88748 664220 88800
rect 656348 88612 656400 88664
rect 657452 88612 657504 88664
rect 610072 88272 610124 88324
rect 626448 88272 626500 88324
rect 655244 88272 655296 88324
rect 658464 88272 658516 88324
rect 622308 88136 622360 88188
rect 626264 88136 626316 88188
rect 579528 88068 579580 88120
rect 585140 88068 585192 88120
rect 648436 86980 648488 87032
rect 662512 86980 662564 87032
rect 656716 86844 656768 86896
rect 659568 86844 659620 86896
rect 656164 86708 656216 86760
rect 660672 86708 660724 86760
rect 649264 86572 649316 86624
rect 661408 86572 661460 86624
rect 652024 86436 652076 86488
rect 657176 86436 657228 86488
rect 619272 86300 619324 86352
rect 626448 86300 626500 86352
rect 647884 86164 647936 86216
rect 660120 86164 660172 86216
rect 609888 85484 609940 85536
rect 626448 85484 626500 85536
rect 620284 85348 620336 85400
rect 625252 85348 625304 85400
rect 579160 84124 579212 84176
rect 581644 84124 581696 84176
rect 608508 84124 608560 84176
rect 625804 84124 625856 84176
rect 579068 82356 579120 82408
rect 583024 82356 583076 82408
rect 579528 82084 579580 82136
rect 587164 82084 587216 82136
rect 628748 80928 628800 80980
rect 642456 80928 642508 80980
rect 612648 80792 612700 80844
rect 647424 80792 647476 80844
rect 595444 80656 595496 80708
rect 636752 80656 636804 80708
rect 629208 79976 629260 80028
rect 633440 79976 633492 80028
rect 613752 79432 613804 79484
rect 646044 79432 646096 79484
rect 579068 79296 579120 79348
rect 588728 79296 588780 79348
rect 613936 79296 613988 79348
rect 646504 79296 646556 79348
rect 633440 78072 633492 78124
rect 645308 78072 645360 78124
rect 631048 77936 631100 77988
rect 643100 77936 643152 77988
rect 628472 77732 628524 77784
rect 632796 77732 632848 77784
rect 625804 77256 625856 77308
rect 631048 77256 631100 77308
rect 616788 76644 616840 76696
rect 646688 76644 646740 76696
rect 612004 76508 612056 76560
rect 662420 76508 662472 76560
rect 578240 75828 578292 75880
rect 580264 75828 580316 75880
rect 618904 75420 618956 75472
rect 648620 75420 648672 75472
rect 615408 75284 615460 75336
rect 646872 75284 646924 75336
rect 607128 75148 607180 75200
rect 646228 75148 646280 75200
rect 578884 72428 578936 72480
rect 601884 72428 601936 72480
rect 579068 71340 579120 71392
rect 584404 71340 584456 71392
rect 580264 68280 580316 68332
rect 604460 68280 604512 68332
rect 577504 59984 577556 60036
rect 603080 59984 603132 60036
rect 576124 58624 576176 58676
rect 601700 58624 601752 58676
rect 574928 57196 574980 57248
rect 600320 57196 600372 57248
rect 574560 55972 574612 56024
rect 599124 55972 599176 56024
rect 574744 55836 574796 55888
rect 600504 55836 600556 55888
rect 596456 55156 596508 55208
rect 597836 55020 597888 55072
rect 597652 54884 597704 54936
rect 598940 54748 598992 54800
rect 624424 54612 624476 54664
rect 625804 54476 625856 54528
rect 596180 54340 596232 54392
rect 581644 54204 581696 54256
rect 574744 54068 574796 54120
rect 462964 53592 463016 53644
rect 463240 53592 463292 53644
rect 463516 53592 463568 53644
rect 463700 53592 463752 53644
rect 464436 53592 464488 53644
rect 464712 53592 464764 53644
rect 476028 53592 476080 53644
rect 476212 53592 476264 53644
rect 476396 53592 476448 53644
rect 476580 53592 476632 53644
rect 477040 53592 477092 53644
rect 479064 53592 479116 53644
rect 479432 53592 479484 53644
rect 574560 53932 574612 53984
rect 479616 53524 479668 53576
rect 462228 53456 462280 53508
rect 479432 53456 479484 53508
rect 463148 53320 463200 53372
rect 574928 53796 574980 53848
rect 48964 53184 49016 53236
rect 130384 53184 130436 53236
rect 461308 53184 461360 53236
rect 479616 53184 479668 53236
rect 312360 53116 312412 53168
rect 313740 53116 313792 53168
rect 316316 53116 316368 53168
rect 317696 53116 317748 53168
rect 45468 53048 45520 53100
rect 129004 53048 129056 53100
rect 459468 53048 459520 53100
rect 463700 53048 463752 53100
rect 465448 53048 465500 53100
rect 479064 53048 479116 53100
rect 462964 52912 463016 52964
rect 464528 52912 464580 52964
rect 460066 52776 460118 52828
rect 464712 52776 464764 52828
rect 465586 52776 465638 52828
rect 476396 52776 476448 52828
rect 47584 51960 47636 52012
rect 130568 51960 130620 52012
rect 50344 51824 50396 51876
rect 129188 51824 129240 51876
rect 129556 51824 129608 51876
rect 591304 51824 591356 51876
rect 128820 51688 128872 51740
rect 592684 51688 592736 51740
rect 318340 50464 318392 50516
rect 458180 50464 458232 50516
rect 47768 50328 47820 50380
rect 130844 50328 130896 50380
rect 314016 50328 314068 50380
rect 458364 50328 458416 50380
rect 522948 50328 523000 50380
rect 544016 50328 544068 50380
rect 49148 49104 49200 49156
rect 129372 49104 129424 49156
rect 46204 48968 46256 49020
rect 131028 48968 131080 49020
rect 130568 46044 130620 46096
rect 132868 46044 132920 46096
rect 130384 45908 130436 45960
rect 132592 45908 132644 45960
rect 129004 45364 129056 45416
rect 129556 45024 129608 45076
rect 129372 44888 129424 44940
rect 128820 44752 128872 44804
rect 131580 44644 131632 44696
rect 129188 44548 129240 44600
rect 50528 44276 50580 44328
rect 131580 44276 131632 44328
rect 43444 44140 43496 44192
rect 132592 44344 132644 44396
rect 132868 44364 132920 44416
rect 132776 44252 132828 44304
rect 131028 44004 131080 44056
rect 440240 43800 440292 43852
rect 441068 43800 441120 43852
rect 187332 42780 187384 42832
rect 255872 42780 255924 42832
rect 307300 42712 307352 42764
rect 431224 42712 431276 42764
rect 441068 42712 441120 42764
rect 449164 42712 449216 42764
rect 453580 42712 453632 42764
rect 464160 42712 464212 42764
rect 310428 42576 310480 42628
rect 427084 42576 427136 42628
rect 441252 42576 441304 42628
rect 446404 42576 446456 42628
rect 454500 42440 454552 42492
rect 463056 42440 463108 42492
rect 404452 42304 404504 42356
rect 405188 42304 405240 42356
rect 420736 42304 420788 42356
rect 426900 42304 426952 42356
rect 661408 42129 661460 42181
rect 427084 41964 427136 42016
rect 431224 41964 431276 42016
rect 441068 41964 441120 42016
rect 446404 41964 446456 42016
rect 454500 41964 454552 42016
rect 441252 41828 441304 41880
rect 449164 41828 449216 41880
rect 453580 41828 453632 41880
rect 404452 41420 404504 41472
rect 420736 41420 420788 41472
rect 426900 41420 426952 41472
rect 459192 41420 459244 41472
<< metal2 >>
rect 185030 1002144 185086 1002153
rect 185030 1002079 185086 1002088
rect 82174 1002008 82230 1002017
rect 81452 1001966 82174 1001994
rect 81452 997098 81480 1001966
rect 133694 1002008 133750 1002017
rect 82174 1001943 82230 1001952
rect 132500 1001972 132552 1001978
rect 133694 1001943 133696 1001952
rect 132500 1001914 132552 1001920
rect 133748 1001943 133750 1001952
rect 133696 1001914 133748 1001920
rect 81360 997070 81480 997098
rect 81360 983521 81388 997070
rect 81346 983512 81402 983521
rect 81346 983447 81402 983456
rect 132512 982569 132540 1001914
rect 185044 992234 185072 1002079
rect 483018 1002008 483074 1002017
rect 483018 1001943 483074 1001952
rect 534998 1002008 535054 1002017
rect 636198 1002008 636254 1002017
rect 535054 1001966 535500 1001994
rect 534998 1001943 535054 1001952
rect 232976 997393 233004 997628
rect 245226 997614 245700 997642
rect 232962 997384 233018 997393
rect 232962 997319 233018 997328
rect 240138 997248 240194 997257
rect 240138 997183 240194 997192
rect 184952 992206 185072 992234
rect 184952 983521 184980 992206
rect 235906 990992 235962 991001
rect 235906 990927 235962 990936
rect 235920 983793 235948 990927
rect 238668 985992 238720 985998
rect 238668 985934 238720 985940
rect 238680 984065 238708 985934
rect 238666 984056 238722 984065
rect 238666 983991 238722 984000
rect 240152 983793 240180 997183
rect 245672 989126 245700 997614
rect 285416 997393 285444 997628
rect 297850 997614 298140 997642
rect 285402 997384 285458 997393
rect 285402 997319 285458 997328
rect 292578 997384 292634 997393
rect 292578 997319 292634 997328
rect 242256 989120 242308 989126
rect 242256 989062 242308 989068
rect 245660 989120 245712 989126
rect 245660 989062 245712 989068
rect 242268 985998 242296 989062
rect 286966 988000 287022 988009
rect 286966 987935 287022 987944
rect 242256 985992 242308 985998
rect 242256 985934 242308 985940
rect 286980 983793 287008 987935
rect 289728 985448 289780 985454
rect 289728 985390 289780 985396
rect 235906 983784 235962 983793
rect 235906 983719 235962 983728
rect 240138 983784 240194 983793
rect 240138 983719 240194 983728
rect 286966 983784 287022 983793
rect 286966 983719 287022 983728
rect 184938 983512 184994 983521
rect 184938 983447 184994 983456
rect 132498 982560 132554 982569
rect 132498 982495 132554 982504
rect 289740 980937 289768 985390
rect 292592 983793 292620 997319
rect 298112 988242 298140 997614
rect 387536 997393 387564 997628
rect 399602 997614 400260 997642
rect 387522 997384 387578 997393
rect 387522 997319 387578 997328
rect 389178 990992 389234 991001
rect 389178 990927 389234 990936
rect 293960 988236 294012 988242
rect 293960 988178 294012 988184
rect 298100 988236 298152 988242
rect 298100 988178 298152 988184
rect 293972 985454 294000 988178
rect 389192 987562 389220 990927
rect 400232 990894 400260 997614
rect 404358 997384 404414 997393
rect 404358 997319 404414 997328
rect 404372 992254 404400 997319
rect 401692 992248 401744 992254
rect 401692 992190 401744 992196
rect 404360 992248 404412 992254
rect 404360 992190 404412 992196
rect 396080 990888 396132 990894
rect 396080 990830 396132 990836
rect 400220 990888 400272 990894
rect 400220 990830 400272 990836
rect 389180 987556 389232 987562
rect 389180 987498 389232 987504
rect 391940 987556 391992 987562
rect 391940 987498 391992 987504
rect 293960 985448 294012 985454
rect 293960 985390 294012 985396
rect 292578 983784 292634 983793
rect 292578 983719 292634 983728
rect 391952 983521 391980 987498
rect 396092 983550 396120 990830
rect 401704 986406 401732 992190
rect 399760 986400 399812 986406
rect 399760 986342 399812 986348
rect 401692 986400 401744 986406
rect 401692 986342 401744 986348
rect 394424 983544 394476 983550
rect 391938 983512 391994 983521
rect 391938 983447 391994 983456
rect 394422 983512 394424 983521
rect 396080 983544 396132 983550
rect 394476 983512 394478 983521
rect 399772 983521 399800 986342
rect 396080 983486 396132 983492
rect 399758 983512 399814 983521
rect 394422 983447 394478 983456
rect 399758 983447 399814 983456
rect 483032 982530 483060 1001943
rect 535472 983793 535500 1001966
rect 636198 1001943 636254 1001952
rect 636212 983793 636240 1001943
rect 535458 983784 535514 983793
rect 535458 983719 535514 983728
rect 636198 983784 636254 983793
rect 636198 983719 636254 983728
rect 483846 982560 483902 982569
rect 483020 982524 483072 982530
rect 483846 982495 483848 982504
rect 483020 982466 483072 982472
rect 483900 982495 483902 982504
rect 483848 982466 483900 982472
rect 289726 980928 289782 980937
rect 289726 980863 289782 980872
rect 30102 960256 30158 960265
rect 30102 960191 30158 960200
rect 30116 954990 30144 960191
rect 651378 959168 651434 959177
rect 651378 959103 651380 959112
rect 651432 959103 651434 959112
rect 677414 959168 677470 959177
rect 677414 959103 677416 959112
rect 651380 959074 651432 959080
rect 677468 959103 677470 959112
rect 677416 959074 677468 959080
rect 63406 959032 63462 959041
rect 63406 958967 63462 958976
rect 63420 954990 63448 958967
rect 30104 954984 30156 954990
rect 30104 954926 30156 954932
rect 63408 954984 63460 954990
rect 63408 954926 63460 954932
rect 703694 897668 703722 897804
rect 704154 897668 704182 897804
rect 704614 897668 704642 897804
rect 705074 897668 705102 897804
rect 705534 897668 705562 897804
rect 705994 897668 706022 897804
rect 706454 897668 706482 897804
rect 706914 897668 706942 897804
rect 707374 897668 707402 897804
rect 707834 897668 707862 897804
rect 708294 897668 708322 897804
rect 708754 897668 708782 897804
rect 709214 897668 709242 897804
rect 676034 897152 676090 897161
rect 676034 897087 676036 897096
rect 676088 897087 676090 897096
rect 676036 897058 676088 897064
rect 656164 897048 656216 897054
rect 656164 896990 656216 896996
rect 654784 895688 654836 895694
rect 654784 895630 654836 895636
rect 653404 880524 653456 880530
rect 653404 880466 653456 880472
rect 651472 868896 651524 868902
rect 651472 868838 651524 868844
rect 651484 868601 651512 868838
rect 651470 868592 651526 868601
rect 651470 868527 651526 868536
rect 651472 867944 651524 867950
rect 651472 867886 651524 867892
rect 651484 867513 651512 867886
rect 651470 867504 651526 867513
rect 651470 867439 651526 867448
rect 651472 866652 651524 866658
rect 651472 866594 651524 866600
rect 651484 866289 651512 866594
rect 651470 866280 651526 866289
rect 651470 866215 651526 866224
rect 653416 865230 653444 880466
rect 654796 868902 654824 895630
rect 654784 868896 654836 868902
rect 654784 868838 654836 868844
rect 654140 868080 654192 868086
rect 654140 868022 654192 868028
rect 651380 865224 651432 865230
rect 651378 865192 651380 865201
rect 653404 865224 653456 865230
rect 651432 865192 651434 865201
rect 653404 865166 653456 865172
rect 651378 865127 651434 865136
rect 651472 863864 651524 863870
rect 651470 863832 651472 863841
rect 651524 863832 651526 863841
rect 651470 863767 651526 863776
rect 654152 862510 654180 868022
rect 656176 867950 656204 896990
rect 675850 896744 675906 896753
rect 675850 896679 675906 896688
rect 672724 895824 672776 895830
rect 672724 895766 672776 895772
rect 671896 894464 671948 894470
rect 671896 894406 671948 894412
rect 671068 894328 671120 894334
rect 671068 894270 671120 894276
rect 670884 886916 670936 886922
rect 670884 886858 670936 886864
rect 667296 880524 667348 880530
rect 667296 880466 667348 880472
rect 667308 879646 667336 880466
rect 667296 879640 667348 879646
rect 667296 879582 667348 879588
rect 657544 869440 657596 869446
rect 657544 869382 657596 869388
rect 656164 867944 656216 867950
rect 656164 867886 656216 867892
rect 657556 863870 657584 869382
rect 657544 863864 657596 863870
rect 657544 863806 657596 863812
rect 651472 862504 651524 862510
rect 651472 862446 651524 862452
rect 654140 862504 654192 862510
rect 654140 862446 654192 862452
rect 651484 862345 651512 862446
rect 651470 862336 651526 862345
rect 651470 862271 651526 862280
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35806 818000 35862 818009
rect 35806 817935 35862 817944
rect 35438 817320 35494 817329
rect 35438 817255 35494 817264
rect 35452 814910 35480 817255
rect 35820 817018 35848 817935
rect 35808 817012 35860 817018
rect 35808 816954 35860 816960
rect 58624 817012 58676 817018
rect 58624 816954 58676 816960
rect 35622 816912 35678 816921
rect 35622 816847 35678 816856
rect 35636 815658 35664 816847
rect 35806 816096 35862 816105
rect 35806 816031 35862 816040
rect 35820 815794 35848 816031
rect 35808 815788 35860 815794
rect 35808 815730 35860 815736
rect 43444 815788 43496 815794
rect 43444 815730 43496 815736
rect 35624 815652 35676 815658
rect 35624 815594 35676 815600
rect 35622 815280 35678 815289
rect 35622 815215 35678 815224
rect 35440 814904 35492 814910
rect 35440 814846 35492 814852
rect 35636 814434 35664 815215
rect 35806 814464 35862 814473
rect 35624 814428 35676 814434
rect 35806 814399 35862 814408
rect 42892 814428 42944 814434
rect 35624 814370 35676 814376
rect 35820 814298 35848 814399
rect 42892 814370 42944 814376
rect 35808 814292 35860 814298
rect 35808 814234 35860 814240
rect 41326 813648 41382 813657
rect 41326 813583 41382 813592
rect 41340 812870 41368 813583
rect 41328 812864 41380 812870
rect 40958 812832 41014 812841
rect 41328 812806 41380 812812
rect 40958 812767 41014 812776
rect 37922 811608 37978 811617
rect 37922 811543 37978 811552
rect 34518 811200 34574 811209
rect 34518 811135 34574 811144
rect 32586 810792 32642 810801
rect 32586 810727 32642 810736
rect 31022 809976 31078 809985
rect 31022 809911 31078 809920
rect 31036 801106 31064 809911
rect 32600 802505 32628 810727
rect 32586 802496 32642 802505
rect 34532 802466 34560 811135
rect 36542 809568 36598 809577
rect 36542 809503 36598 809512
rect 32586 802431 32642 802440
rect 34520 802460 34572 802466
rect 34520 802402 34572 802408
rect 36556 801310 36584 809503
rect 37936 801786 37964 811543
rect 40972 810762 41000 812767
rect 41326 812424 41382 812433
rect 41326 812359 41382 812368
rect 41142 812016 41198 812025
rect 41142 811951 41198 811960
rect 40960 810756 41012 810762
rect 40960 810698 41012 810704
rect 41156 809962 41184 811951
rect 41340 811782 41368 812359
rect 41328 811776 41380 811782
rect 41328 811718 41380 811724
rect 42616 810756 42668 810762
rect 42616 810698 42668 810704
rect 41970 810384 42026 810393
rect 41970 810319 42026 810328
rect 41786 809976 41842 809985
rect 41156 809934 41786 809962
rect 41786 809911 41842 809920
rect 41326 809160 41382 809169
rect 41326 809095 41382 809104
rect 41340 808654 41368 809095
rect 41786 808752 41842 808761
rect 41786 808687 41842 808696
rect 41328 808648 41380 808654
rect 41328 808590 41380 808596
rect 41142 808344 41198 808353
rect 41142 808279 41198 808288
rect 41156 807362 41184 808279
rect 41326 807528 41382 807537
rect 41326 807463 41328 807472
rect 41380 807463 41382 807472
rect 41328 807434 41380 807440
rect 41144 807356 41196 807362
rect 41144 807298 41196 807304
rect 41142 806712 41198 806721
rect 41142 806647 41198 806656
rect 41156 806002 41184 806647
rect 41326 806304 41382 806313
rect 41326 806239 41382 806248
rect 41340 806138 41368 806239
rect 41328 806132 41380 806138
rect 41328 806074 41380 806080
rect 41144 805996 41196 806002
rect 41144 805938 41196 805944
rect 41800 805225 41828 808687
rect 41984 805633 42012 810319
rect 42628 808694 42656 810698
rect 42444 808666 42656 808694
rect 42904 808694 42932 814370
rect 43076 811776 43128 811782
rect 43076 811718 43128 811724
rect 42904 808666 43024 808694
rect 42248 808648 42300 808654
rect 42300 808596 42380 808602
rect 42248 808590 42380 808596
rect 42260 808574 42380 808590
rect 41970 805624 42026 805633
rect 41970 805559 42026 805568
rect 41786 805216 41842 805225
rect 41786 805151 41842 805160
rect 42156 802460 42208 802466
rect 42156 802402 42208 802408
rect 42168 802346 42196 802402
rect 42168 802318 42288 802346
rect 37924 801780 37976 801786
rect 37924 801722 37976 801728
rect 41972 801780 42024 801786
rect 41972 801722 42024 801728
rect 36544 801304 36596 801310
rect 36544 801246 36596 801252
rect 41984 801174 42012 801722
rect 41972 801168 42024 801174
rect 41972 801110 42024 801116
rect 31024 801100 31076 801106
rect 31024 801042 31076 801048
rect 42260 799459 42288 802318
rect 42182 799431 42288 799459
rect 42154 798144 42210 798153
rect 42352 798130 42380 808574
rect 42210 798102 42380 798130
rect 42154 798079 42210 798088
rect 42444 797994 42472 808666
rect 42616 801304 42668 801310
rect 42352 797966 42472 797994
rect 42536 801252 42616 801258
rect 42536 801246 42668 801252
rect 42536 801230 42656 801246
rect 42352 797858 42380 797966
rect 42260 797830 42380 797858
rect 42260 797619 42288 797830
rect 42536 797722 42564 801230
rect 42708 801168 42760 801174
rect 42182 797591 42288 797619
rect 42352 797694 42564 797722
rect 42628 801116 42708 801122
rect 42628 801110 42760 801116
rect 42628 801094 42748 801110
rect 42062 797328 42118 797337
rect 42062 797263 42118 797272
rect 42076 796960 42104 797263
rect 42352 795779 42380 797694
rect 42182 795751 42380 795779
rect 42248 795660 42300 795666
rect 42248 795602 42300 795608
rect 42260 795138 42288 795602
rect 42182 795110 42288 795138
rect 41786 794880 41842 794889
rect 41786 794815 41842 794824
rect 41800 794580 41828 794815
rect 42154 794472 42210 794481
rect 42154 794407 42210 794416
rect 42168 793900 42196 794407
rect 42340 794368 42392 794374
rect 42340 794310 42392 794316
rect 42352 793778 42380 794310
rect 42168 793750 42380 793778
rect 42168 793288 42196 793750
rect 42628 792962 42656 801094
rect 42800 801032 42852 801038
rect 42720 800980 42800 800986
rect 42720 800974 42852 800980
rect 42720 800958 42840 800974
rect 42720 795682 42748 800958
rect 42720 795654 42932 795682
rect 42904 795138 42932 795654
rect 42260 792934 42656 792962
rect 42720 795110 42932 795138
rect 42260 792758 42288 792934
rect 42182 792730 42288 792758
rect 42430 792024 42486 792033
rect 42430 791959 42486 791968
rect 41786 790664 41842 790673
rect 41786 790599 41842 790608
rect 41800 790228 41828 790599
rect 42156 790152 42208 790158
rect 42156 790094 42208 790100
rect 42168 789616 42196 790094
rect 42444 789374 42472 791959
rect 42720 790158 42748 795110
rect 42996 794894 43024 808666
rect 42904 794866 43024 794894
rect 42708 790152 42760 790158
rect 42708 790094 42760 790100
rect 42260 789346 42472 789374
rect 41786 789304 41842 789313
rect 41786 789239 41842 789248
rect 41800 788936 41828 789239
rect 42260 788406 42288 789346
rect 42182 788378 42288 788406
rect 42430 788352 42486 788361
rect 42430 788287 42486 788296
rect 42444 788202 42472 788287
rect 42168 788174 42472 788202
rect 42168 787930 42196 788174
rect 42430 788080 42486 788089
rect 42430 788015 42486 788024
rect 42616 788044 42668 788050
rect 42168 787902 42288 787930
rect 42260 786978 42288 787902
rect 42168 786950 42288 786978
rect 42168 786556 42196 786950
rect 42444 785958 42472 788015
rect 42616 787986 42668 787992
rect 42628 786842 42656 787986
rect 42168 785890 42196 785944
rect 42260 785930 42472 785958
rect 42536 786814 42656 786842
rect 42260 785890 42288 785930
rect 42168 785862 42288 785890
rect 42536 785278 42564 786814
rect 42708 786684 42760 786690
rect 42708 786626 42760 786632
rect 42182 785250 42564 785278
rect 42720 784802 42748 786626
rect 42536 784774 42748 784802
rect 42536 784734 42564 784774
rect 42182 784706 42564 784734
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 774752 35862 774761
rect 35806 774687 35862 774696
rect 35820 774246 35848 774687
rect 35808 774240 35860 774246
rect 35808 774182 35860 774188
rect 41696 774240 41748 774246
rect 42064 774240 42116 774246
rect 41748 774188 42064 774194
rect 41696 774182 42116 774188
rect 41708 774166 42104 774182
rect 35438 773936 35494 773945
rect 35438 773871 35494 773880
rect 35452 772886 35480 773871
rect 35806 773528 35862 773537
rect 35806 773463 35862 773472
rect 39578 773528 39634 773537
rect 39578 773463 39634 773472
rect 35820 773362 35848 773463
rect 35808 773356 35860 773362
rect 35808 773298 35860 773304
rect 39592 773158 39620 773463
rect 40316 773356 40368 773362
rect 40316 773298 40368 773304
rect 35808 773152 35860 773158
rect 35806 773120 35808 773129
rect 39580 773152 39632 773158
rect 35860 773120 35862 773129
rect 40328 773129 40356 773298
rect 39580 773094 39632 773100
rect 40314 773120 40370 773129
rect 35806 773055 35862 773064
rect 40314 773055 40370 773064
rect 35624 773016 35676 773022
rect 35624 772958 35676 772964
rect 41696 773016 41748 773022
rect 42064 773016 42116 773022
rect 41748 772964 42064 772970
rect 41696 772958 42116 772964
rect 35440 772880 35492 772886
rect 35440 772822 35492 772828
rect 35636 772721 35664 772958
rect 41708 772942 42104 772958
rect 41696 772880 41748 772886
rect 42064 772880 42116 772886
rect 41748 772828 42064 772834
rect 41696 772822 42116 772828
rect 41708 772806 42104 772822
rect 35622 772712 35678 772721
rect 35622 772647 35678 772656
rect 42904 772313 42932 794866
rect 43088 788050 43116 811718
rect 43260 807492 43312 807498
rect 43260 807434 43312 807440
rect 43076 788044 43128 788050
rect 43076 787986 43128 787992
rect 35622 772304 35678 772313
rect 35622 772239 35678 772248
rect 40774 772304 40830 772313
rect 40774 772239 40830 772248
rect 42890 772304 42946 772313
rect 42890 772239 42946 772248
rect 35438 771896 35494 771905
rect 35636 771866 35664 772239
rect 35806 771896 35862 771905
rect 35438 771831 35494 771840
rect 35624 771860 35676 771866
rect 35452 771458 35480 771831
rect 40788 771866 40816 772239
rect 35806 771831 35862 771840
rect 40776 771860 40828 771866
rect 35624 771802 35676 771808
rect 35820 771594 35848 771831
rect 40776 771802 40828 771808
rect 41696 771656 41748 771662
rect 42064 771656 42116 771662
rect 41748 771604 42064 771610
rect 41696 771598 42116 771604
rect 35808 771588 35860 771594
rect 41708 771582 42104 771598
rect 35808 771530 35860 771536
rect 41708 771458 42104 771474
rect 35440 771452 35492 771458
rect 35440 771394 35492 771400
rect 41696 771452 42116 771458
rect 41748 771446 42064 771452
rect 41696 771394 41748 771400
rect 42064 771394 42116 771400
rect 35438 771080 35494 771089
rect 35438 771015 35494 771024
rect 35452 770234 35480 771015
rect 35622 770672 35678 770681
rect 35622 770607 35678 770616
rect 35440 770228 35492 770234
rect 35440 770170 35492 770176
rect 35636 770098 35664 770607
rect 35808 770500 35860 770506
rect 35808 770442 35860 770448
rect 40500 770500 40552 770506
rect 40500 770442 40552 770448
rect 35820 770273 35848 770442
rect 39948 770296 40000 770302
rect 35806 770264 35862 770273
rect 40512 770273 40540 770442
rect 39948 770238 40000 770244
rect 40498 770264 40554 770273
rect 35806 770199 35862 770208
rect 35624 770092 35676 770098
rect 35624 770034 35676 770040
rect 39960 769457 39988 770238
rect 40498 770199 40554 770208
rect 43074 770264 43130 770273
rect 43074 770199 43130 770208
rect 41708 770098 42104 770114
rect 41696 770092 42116 770098
rect 41748 770086 42064 770092
rect 41696 770034 41748 770040
rect 42064 770034 42116 770040
rect 35622 769448 35678 769457
rect 35622 769383 35678 769392
rect 39946 769448 40002 769457
rect 39946 769383 40002 769392
rect 35636 768874 35664 769383
rect 35806 769040 35862 769049
rect 35806 768975 35862 768984
rect 35624 768868 35676 768874
rect 35624 768810 35676 768816
rect 35820 768738 35848 768975
rect 41696 768868 41748 768874
rect 41696 768810 41748 768816
rect 35808 768732 35860 768738
rect 35808 768674 35860 768680
rect 40040 768732 40092 768738
rect 40040 768674 40092 768680
rect 35162 768224 35218 768233
rect 35162 768159 35218 768168
rect 32402 767816 32458 767825
rect 32402 767751 32458 767760
rect 32416 759694 32444 767751
rect 33782 767000 33838 767009
rect 33782 766935 33838 766944
rect 32404 759688 32456 759694
rect 32404 759630 32456 759636
rect 33796 758334 33824 766935
rect 35176 759830 35204 768159
rect 35808 767644 35860 767650
rect 35808 767586 35860 767592
rect 36544 767644 36596 767650
rect 36544 767586 36596 767592
rect 35820 767417 35848 767586
rect 35806 767408 35862 767417
rect 35806 767343 35862 767352
rect 35806 766184 35862 766193
rect 35806 766119 35862 766128
rect 35820 765950 35848 766119
rect 35808 765944 35860 765950
rect 35808 765886 35860 765892
rect 35806 765776 35862 765785
rect 35806 765711 35862 765720
rect 35820 764862 35848 765711
rect 35808 764856 35860 764862
rect 35808 764798 35860 764804
rect 35808 764584 35860 764590
rect 35806 764552 35808 764561
rect 35860 764552 35862 764561
rect 35806 764487 35862 764496
rect 35622 764144 35678 764153
rect 35622 764079 35678 764088
rect 35636 763502 35664 764079
rect 35806 763736 35862 763745
rect 35806 763671 35862 763680
rect 35624 763496 35676 763502
rect 35624 763438 35676 763444
rect 35820 763230 35848 763671
rect 35808 763224 35860 763230
rect 35808 763166 35860 763172
rect 35806 762920 35862 762929
rect 35806 762855 35862 762864
rect 35820 761870 35848 762855
rect 35808 761864 35860 761870
rect 35808 761806 35860 761812
rect 35164 759824 35216 759830
rect 35164 759766 35216 759772
rect 33784 758328 33836 758334
rect 33784 758270 33836 758276
rect 36556 757761 36584 767586
rect 39764 765944 39816 765950
rect 39764 765886 39816 765892
rect 39776 765785 39804 765886
rect 39762 765776 39818 765785
rect 39762 765711 39818 765720
rect 40052 765338 40080 768674
rect 41708 765914 41736 768810
rect 41708 765886 42288 765914
rect 40040 765332 40092 765338
rect 40040 765274 40092 765280
rect 41696 765332 41748 765338
rect 41696 765274 41748 765280
rect 41708 765218 41736 765274
rect 41708 765202 42104 765218
rect 41708 765196 42116 765202
rect 41708 765190 42064 765196
rect 42064 765138 42116 765144
rect 39212 764856 39264 764862
rect 39212 764798 39264 764804
rect 39224 764153 39252 764798
rect 39764 764584 39816 764590
rect 39762 764552 39764 764561
rect 39816 764552 39818 764561
rect 39762 764487 39818 764496
rect 39210 764144 39266 764153
rect 39210 764079 39266 764088
rect 41696 763496 41748 763502
rect 41696 763438 41748 763444
rect 41708 763337 41736 763438
rect 41694 763328 41750 763337
rect 41694 763263 41750 763272
rect 41696 763156 41748 763162
rect 41696 763098 41748 763104
rect 41708 762929 41736 763098
rect 41694 762920 41750 762929
rect 41694 762855 41750 762864
rect 42064 761932 42116 761938
rect 42064 761874 42116 761880
rect 41696 761864 41748 761870
rect 42076 761818 42104 761874
rect 41748 761812 42104 761818
rect 41696 761806 42104 761812
rect 41708 761790 42104 761806
rect 41696 759824 41748 759830
rect 41748 759772 42104 759778
rect 41696 759766 42104 759772
rect 41708 759750 42104 759766
rect 41604 759688 41656 759694
rect 41656 759636 41828 759642
rect 41604 759630 41828 759636
rect 41616 759614 41828 759630
rect 39304 758328 39356 758334
rect 39302 758296 39304 758305
rect 39356 758296 39358 758305
rect 39302 758231 39358 758240
rect 36542 757752 36598 757761
rect 36542 757687 36598 757696
rect 41800 757081 41828 759614
rect 42076 757994 42104 759750
rect 42064 757988 42116 757994
rect 42064 757930 42116 757936
rect 41786 757072 41842 757081
rect 41786 757007 41842 757016
rect 41878 756664 41934 756673
rect 41878 756599 41934 756608
rect 41892 756226 41920 756599
rect 42260 754406 42288 765886
rect 42524 765196 42576 765202
rect 42524 765138 42576 765144
rect 42536 763154 42564 765138
rect 42444 763126 42564 763154
rect 43088 763154 43116 770199
rect 43088 763126 43208 763154
rect 42444 758130 42472 763126
rect 42616 763088 42668 763094
rect 42616 763030 42668 763036
rect 42628 762929 42656 763030
rect 42614 762920 42670 762929
rect 42614 762855 42670 762864
rect 42798 758296 42854 758305
rect 42628 758254 42798 758282
rect 42432 758124 42484 758130
rect 42432 758066 42484 758072
rect 42432 757988 42484 757994
rect 42432 757930 42484 757936
rect 42444 757874 42472 757930
rect 42444 757846 42564 757874
rect 42182 754378 42288 754406
rect 42248 754316 42300 754322
rect 42248 754258 42300 754264
rect 42260 754066 42288 754258
rect 42076 754038 42288 754066
rect 42076 753780 42104 754038
rect 42338 753944 42394 753953
rect 42338 753879 42394 753888
rect 42352 753494 42380 753879
rect 42352 753466 42472 753494
rect 42248 753432 42300 753438
rect 42248 753374 42300 753380
rect 42062 752992 42118 753001
rect 42062 752927 42118 752936
rect 42076 752556 42104 752927
rect 42168 751777 42196 751944
rect 42260 751890 42288 753374
rect 42260 751862 42380 751890
rect 42154 751768 42210 751777
rect 42154 751703 42210 751712
rect 42352 751383 42380 751862
rect 42182 751355 42380 751383
rect 42062 750952 42118 750961
rect 42062 750887 42118 750896
rect 42076 750720 42104 750887
rect 41786 750544 41842 750553
rect 41786 750479 41842 750488
rect 41800 750108 41828 750479
rect 42444 750122 42472 753466
rect 42352 750094 42472 750122
rect 42352 750038 42380 750094
rect 42340 750032 42392 750038
rect 42340 749974 42392 749980
rect 42536 749714 42564 757846
rect 42352 749686 42564 749714
rect 42352 749543 42380 749686
rect 42182 749515 42380 749543
rect 42340 749352 42392 749358
rect 42340 749294 42392 749300
rect 42352 747402 42380 749294
rect 42168 747374 42380 747402
rect 42168 747048 42196 747374
rect 41786 746736 41842 746745
rect 41786 746671 41842 746680
rect 41800 746401 41828 746671
rect 42628 746594 42656 758254
rect 42798 758231 42854 758240
rect 42800 758124 42852 758130
rect 42800 758066 42852 758072
rect 42812 755426 42840 758066
rect 42352 746566 42656 746594
rect 42720 755398 42840 755426
rect 42352 745906 42380 746566
rect 42168 745878 42380 745906
rect 42168 745756 42196 745878
rect 42338 745648 42394 745657
rect 42338 745583 42394 745592
rect 42156 745476 42208 745482
rect 42156 745418 42208 745424
rect 42168 745212 42196 745418
rect 42352 743390 42380 745583
rect 42720 745482 42748 755398
rect 42892 754928 42944 754934
rect 42892 754870 42944 754876
rect 42904 753001 42932 754870
rect 42890 752992 42946 753001
rect 42890 752927 42946 752936
rect 43180 746594 43208 763126
rect 42904 746566 43208 746594
rect 42904 745906 42932 746566
rect 42904 745878 43024 745906
rect 42708 745476 42760 745482
rect 42708 745418 42760 745424
rect 42614 745104 42670 745113
rect 42614 745039 42670 745048
rect 42182 743362 42380 743390
rect 41878 743064 41934 743073
rect 41878 742999 41934 743008
rect 41892 742696 41920 742999
rect 42628 742098 42656 745039
rect 42800 744116 42852 744122
rect 42800 744058 42852 744064
rect 42812 744002 42840 744058
rect 42182 742070 42656 742098
rect 42720 743974 42840 744002
rect 42720 741690 42748 743974
rect 42536 741662 42748 741690
rect 42536 741554 42564 741662
rect 42182 741526 42564 741554
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 42430 730552 42486 730561
rect 42430 730487 42486 730496
rect 42444 729366 42472 730487
rect 42432 729360 42484 729366
rect 41326 729328 41382 729337
rect 42432 729302 42484 729308
rect 41326 729263 41382 729272
rect 41340 728822 41368 729263
rect 41328 728816 41380 728822
rect 41328 728758 41380 728764
rect 41696 728816 41748 728822
rect 42064 728816 42116 728822
rect 41748 728776 42064 728804
rect 41696 728758 41748 728764
rect 42064 728758 42116 728764
rect 40682 728682 40738 728691
rect 40682 728617 40738 728626
rect 41326 728682 41382 728691
rect 41326 728617 41382 728626
rect 41696 728680 41748 728686
rect 42064 728680 42116 728686
rect 41748 728640 42064 728668
rect 41696 728622 41748 728628
rect 42064 728622 42116 728628
rect 40696 727462 40724 728617
rect 40866 728104 40922 728113
rect 40866 728039 40922 728048
rect 40684 727456 40736 727462
rect 40684 727398 40736 727404
rect 40880 727326 40908 728039
rect 42996 727705 43024 745878
rect 42982 727696 43038 727705
rect 42982 727631 43038 727640
rect 41696 727456 41748 727462
rect 42064 727456 42116 727462
rect 41748 727416 42064 727444
rect 41696 727398 41748 727404
rect 42064 727398 42116 727404
rect 40868 727320 40920 727326
rect 40868 727262 40920 727268
rect 41696 727320 41748 727326
rect 42064 727320 42116 727326
rect 41748 727268 42064 727274
rect 41696 727262 42116 727268
rect 42982 727288 43038 727297
rect 41708 727246 42104 727262
rect 42982 727223 43038 727232
rect 41142 726880 41198 726889
rect 41142 726815 41198 726824
rect 40958 726472 41014 726481
rect 40958 726407 41014 726416
rect 40972 725966 41000 726407
rect 41156 726102 41184 726815
rect 41144 726096 41196 726102
rect 41144 726038 41196 726044
rect 41604 726096 41656 726102
rect 41604 726038 41656 726044
rect 40960 725960 41012 725966
rect 40960 725902 41012 725908
rect 41420 725960 41472 725966
rect 41420 725902 41472 725908
rect 40958 725656 41014 725665
rect 40958 725591 41014 725600
rect 32402 725248 32458 725257
rect 32402 725183 32458 725192
rect 31666 724024 31722 724033
rect 31666 723959 31722 723968
rect 31680 715562 31708 723959
rect 32416 716922 32444 725183
rect 35162 724840 35218 724849
rect 35162 724775 35218 724784
rect 32404 716916 32456 716922
rect 32404 716858 32456 716864
rect 35176 715698 35204 724775
rect 37278 724432 37334 724441
rect 37278 724367 37334 724376
rect 37292 716961 37320 724367
rect 39302 723208 39358 723217
rect 39302 723143 39358 723152
rect 37278 716952 37334 716961
rect 37278 716887 37334 716896
rect 35164 715692 35216 715698
rect 35164 715634 35216 715640
rect 31668 715556 31720 715562
rect 31668 715498 31720 715504
rect 39316 714814 39344 723143
rect 40972 719001 41000 725591
rect 41432 725506 41460 725902
rect 41616 725642 41644 726038
rect 41786 725656 41842 725665
rect 41616 725614 41786 725642
rect 41786 725591 41842 725600
rect 41432 725478 41644 725506
rect 41616 719273 41644 725478
rect 41786 722392 41842 722401
rect 41786 722327 41842 722336
rect 41602 719264 41658 719273
rect 41602 719199 41658 719208
rect 40958 718992 41014 719001
rect 40958 718927 41014 718936
rect 41800 718593 41828 722327
rect 42798 720352 42854 720361
rect 42798 720287 42854 720296
rect 42246 719264 42302 719273
rect 42246 719199 42302 719208
rect 42062 718992 42118 719001
rect 42062 718927 42118 718936
rect 41786 718584 41842 718593
rect 41786 718519 41842 718528
rect 40224 716916 40276 716922
rect 40224 716858 40276 716864
rect 40236 715873 40264 716858
rect 40222 715864 40278 715873
rect 40222 715799 40278 715808
rect 41512 715692 41564 715698
rect 41512 715634 41564 715640
rect 40592 715556 40644 715562
rect 40592 715498 40644 715504
rect 40604 715329 40632 715498
rect 40590 715320 40646 715329
rect 40590 715255 40646 715264
rect 39304 714808 39356 714814
rect 39304 714750 39356 714756
rect 41524 714218 41552 715634
rect 42076 715086 42104 718927
rect 42064 715080 42116 715086
rect 42064 715022 42116 715028
rect 42260 714854 42288 719199
rect 42812 719030 42840 720287
rect 42800 719024 42852 719030
rect 42800 718966 42852 718972
rect 42706 715864 42762 715873
rect 42706 715799 42762 715808
rect 42430 715320 42486 715329
rect 42486 715278 42656 715306
rect 42430 715255 42486 715264
rect 42432 715080 42484 715086
rect 42484 715028 42564 715034
rect 42432 715022 42564 715028
rect 42444 715006 42564 715022
rect 42260 714826 42472 714854
rect 41696 714808 41748 714814
rect 41696 714750 41748 714756
rect 41708 714513 41736 714750
rect 41694 714504 41750 714513
rect 41694 714439 41750 714448
rect 41524 714190 42288 714218
rect 42260 713062 42288 714190
rect 42182 713034 42288 713062
rect 42444 711226 42472 714826
rect 42182 711198 42472 711226
rect 42340 711136 42392 711142
rect 42340 711078 42392 711084
rect 42352 710575 42380 711078
rect 42182 710547 42380 710575
rect 42340 710456 42392 710462
rect 42340 710398 42392 710404
rect 42062 709880 42118 709889
rect 42062 709815 42118 709824
rect 42076 709376 42104 709815
rect 42076 708529 42104 708696
rect 41878 708520 41934 708529
rect 41878 708455 41934 708464
rect 42062 708520 42118 708529
rect 42062 708455 42118 708464
rect 41892 708152 41920 708455
rect 42154 707704 42210 707713
rect 42154 707639 42210 707648
rect 42168 707540 42196 707639
rect 41786 707432 41842 707441
rect 41786 707367 41842 707376
rect 41800 706860 41828 707367
rect 42352 706330 42380 710398
rect 42182 706302 42380 706330
rect 42246 706208 42302 706217
rect 42246 706143 42302 706152
rect 42260 704290 42288 706143
rect 42536 705194 42564 715006
rect 42628 710002 42656 715278
rect 42720 714854 42748 715799
rect 42720 714826 42840 714854
rect 42812 710462 42840 714826
rect 42800 710456 42852 710462
rect 42800 710398 42852 710404
rect 42628 709974 42748 710002
rect 42536 705166 42656 705194
rect 42076 704262 42288 704290
rect 42076 703868 42104 704262
rect 42062 703488 42118 703497
rect 42062 703423 42118 703432
rect 42076 703188 42104 703423
rect 42628 703202 42656 705166
rect 42260 703174 42656 703202
rect 42062 703080 42118 703089
rect 42062 703015 42118 703024
rect 42076 702576 42104 703015
rect 42260 702386 42288 703174
rect 42720 703089 42748 709974
rect 42706 703080 42762 703089
rect 42706 703015 42762 703024
rect 42614 702808 42670 702817
rect 42614 702743 42670 702752
rect 42076 702358 42288 702386
rect 42076 702032 42104 702358
rect 42628 702250 42656 702743
rect 42260 702222 42656 702250
rect 42260 700179 42288 702222
rect 42614 702128 42670 702137
rect 42614 702063 42670 702072
rect 42430 701856 42486 701865
rect 42430 701791 42486 701800
rect 42182 700151 42288 700179
rect 42444 699530 42472 701791
rect 42182 699502 42472 699530
rect 42628 698918 42656 702063
rect 42800 701072 42852 701078
rect 42168 698850 42196 698904
rect 42260 698890 42656 698918
rect 42720 701020 42800 701026
rect 42720 701014 42852 701020
rect 42720 700998 42840 701014
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 42720 698339 42748 700998
rect 42182 698311 42748 698339
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 35438 688392 35494 688401
rect 35438 688327 35494 688336
rect 35452 687274 35480 688327
rect 35806 687712 35862 687721
rect 35806 687647 35862 687656
rect 35820 687546 35848 687647
rect 41694 687576 41750 687585
rect 35808 687540 35860 687546
rect 41694 687511 41696 687520
rect 35808 687482 35860 687488
rect 41748 687511 41750 687520
rect 41696 687482 41748 687488
rect 35622 687304 35678 687313
rect 35440 687268 35492 687274
rect 35622 687239 35678 687248
rect 35440 687210 35492 687216
rect 35438 686896 35494 686905
rect 35438 686831 35494 686840
rect 35452 685914 35480 686831
rect 35636 686458 35664 687239
rect 41696 687200 41748 687206
rect 41694 687168 41696 687177
rect 41748 687168 41750 687177
rect 41694 687103 41750 687112
rect 42064 686520 42116 686526
rect 35806 686488 35862 686497
rect 35624 686452 35676 686458
rect 41708 686468 42064 686474
rect 41708 686462 42116 686468
rect 41708 686458 42104 686462
rect 35806 686423 35862 686432
rect 41696 686452 42104 686458
rect 35624 686394 35676 686400
rect 35820 686322 35848 686423
rect 41748 686446 42104 686452
rect 41696 686394 41748 686400
rect 41708 686322 42104 686338
rect 35808 686316 35860 686322
rect 35808 686258 35860 686264
rect 41696 686316 42116 686322
rect 41748 686310 42064 686316
rect 41696 686258 41748 686264
rect 42064 686258 42116 686264
rect 42064 686112 42116 686118
rect 35806 686080 35862 686089
rect 41708 686060 42064 686066
rect 41708 686054 42116 686060
rect 41708 686050 42104 686054
rect 35806 686015 35808 686024
rect 35860 686015 35862 686024
rect 41696 686044 42104 686050
rect 35808 685986 35860 685992
rect 41748 686038 42104 686044
rect 41696 685986 41748 685992
rect 41708 685914 42104 685930
rect 35440 685908 35492 685914
rect 35440 685850 35492 685856
rect 41696 685908 42116 685914
rect 41748 685902 42064 685908
rect 41696 685850 41748 685856
rect 42064 685850 42116 685856
rect 35806 685672 35862 685681
rect 35806 685607 35862 685616
rect 35622 685264 35678 685273
rect 35622 685199 35678 685208
rect 35636 684690 35664 685199
rect 35820 685030 35848 685607
rect 41694 685128 41750 685137
rect 41524 685086 41694 685114
rect 35808 685024 35860 685030
rect 35808 684966 35860 684972
rect 35806 684856 35862 684865
rect 35806 684791 35862 684800
rect 41328 684820 41380 684826
rect 35624 684684 35676 684690
rect 35624 684626 35676 684632
rect 35820 684554 35848 684791
rect 41328 684762 41380 684768
rect 35808 684548 35860 684554
rect 35808 684490 35860 684496
rect 35622 684448 35678 684457
rect 35622 684383 35678 684392
rect 35438 684040 35494 684049
rect 35438 683975 35494 683984
rect 35452 683194 35480 683975
rect 35636 683330 35664 684383
rect 41340 684298 41368 684762
rect 41524 684690 41552 685086
rect 41694 685063 41750 685072
rect 42064 684956 42116 684962
rect 42064 684898 42116 684904
rect 42076 684842 42104 684898
rect 41708 684814 42104 684842
rect 41512 684684 41564 684690
rect 41512 684626 41564 684632
rect 41708 684554 41736 684814
rect 41696 684548 41748 684554
rect 41696 684490 41748 684496
rect 41694 684312 41750 684321
rect 41340 684270 41694 684298
rect 41694 684247 41750 684256
rect 42996 683913 43024 727223
rect 41694 683904 41750 683913
rect 41524 683862 41694 683890
rect 35808 683460 35860 683466
rect 35808 683402 35860 683408
rect 35624 683324 35676 683330
rect 35624 683266 35676 683272
rect 35820 683233 35848 683402
rect 41524 683330 41552 683862
rect 41694 683839 41750 683848
rect 42982 683904 43038 683913
rect 42982 683839 43038 683848
rect 41696 683460 41748 683466
rect 41696 683402 41748 683408
rect 41708 683346 41736 683402
rect 41512 683324 41564 683330
rect 41708 683318 42288 683346
rect 41512 683266 41564 683272
rect 35806 683224 35862 683233
rect 35440 683188 35492 683194
rect 41708 683194 42104 683210
rect 35806 683159 35862 683168
rect 41696 683188 42116 683194
rect 35440 683130 35492 683136
rect 41748 683182 42064 683188
rect 41696 683130 41748 683136
rect 42064 683130 42116 683136
rect 35622 682816 35678 682825
rect 35622 682751 35678 682760
rect 35162 682000 35218 682009
rect 35162 681935 35218 681944
rect 33046 681592 33102 681601
rect 33046 681527 33102 681536
rect 31022 680776 31078 680785
rect 31022 680711 31078 680720
rect 31036 672790 31064 680711
rect 33060 674150 33088 681527
rect 33782 681184 33838 681193
rect 33782 681119 33838 681128
rect 33048 674144 33100 674150
rect 33048 674086 33100 674092
rect 31024 672784 31076 672790
rect 33796 672761 33824 681119
rect 35176 672926 35204 681935
rect 35636 681902 35664 682751
rect 35806 682408 35862 682417
rect 35806 682343 35862 682352
rect 35624 681896 35676 681902
rect 35624 681838 35676 681844
rect 35820 681766 35848 682343
rect 41604 681896 41656 681902
rect 41604 681838 41656 681844
rect 35808 681760 35860 681766
rect 35808 681702 35860 681708
rect 41420 681760 41472 681766
rect 41420 681702 41472 681708
rect 41616 681714 41644 681838
rect 42064 681760 42116 681766
rect 41786 681728 41842 681737
rect 41432 681578 41460 681702
rect 41616 681686 41786 681714
rect 42064 681702 42116 681708
rect 41786 681663 41842 681672
rect 42076 681578 42104 681702
rect 41432 681550 42104 681578
rect 35808 680672 35860 680678
rect 41696 680672 41748 680678
rect 35808 680614 35860 680620
rect 41694 680640 41696 680649
rect 41748 680640 41750 680649
rect 35820 680377 35848 680614
rect 41694 680575 41750 680584
rect 35806 680368 35862 680377
rect 35806 680303 35862 680312
rect 35622 679960 35678 679969
rect 35622 679895 35678 679904
rect 35438 679552 35494 679561
rect 35438 679487 35494 679496
rect 35452 679046 35480 679487
rect 35636 679182 35664 679895
rect 35808 679448 35860 679454
rect 41696 679448 41748 679454
rect 35808 679390 35860 679396
rect 41694 679416 41696 679425
rect 41748 679416 41750 679425
rect 35624 679176 35676 679182
rect 35820 679153 35848 679390
rect 41694 679351 41750 679360
rect 41708 679250 42104 679266
rect 41696 679244 42116 679250
rect 41748 679238 42064 679244
rect 41696 679186 41748 679192
rect 42064 679186 42116 679192
rect 35624 679118 35676 679124
rect 35806 679144 35862 679153
rect 35806 679079 35862 679088
rect 35440 679040 35492 679046
rect 35440 678982 35492 678988
rect 41696 679040 41748 679046
rect 42064 679040 42116 679046
rect 41748 678988 42064 678994
rect 41696 678982 42116 678988
rect 41708 678966 42104 678982
rect 42260 678974 42288 683318
rect 42616 681760 42668 681766
rect 42616 681702 42668 681708
rect 42260 678946 42472 678974
rect 41786 678328 41842 678337
rect 41616 678286 41786 678314
rect 40774 677750 40830 677759
rect 41616 677754 41644 678286
rect 41786 678263 41842 678272
rect 40774 677685 40830 677694
rect 41604 677748 41656 677754
rect 41604 677690 41656 677696
rect 41512 674144 41564 674150
rect 41512 674086 41564 674092
rect 35164 672920 35216 672926
rect 35164 672862 35216 672868
rect 39580 672920 39632 672926
rect 39580 672862 39632 672868
rect 31024 672726 31076 672732
rect 33782 672752 33838 672761
rect 33782 672687 33838 672696
rect 39592 670993 39620 672862
rect 41524 672738 41552 674086
rect 42444 673169 42472 678946
rect 42430 673160 42486 673169
rect 42430 673095 42486 673104
rect 41524 672710 42288 672738
rect 41696 672648 41748 672654
rect 41748 672596 42104 672602
rect 41696 672590 42104 672596
rect 41708 672586 42104 672590
rect 41708 672580 42116 672586
rect 41708 672574 42064 672580
rect 42064 672522 42116 672528
rect 39578 670984 39634 670993
rect 39578 670919 39634 670928
rect 42168 669746 42196 669868
rect 42260 669746 42288 672710
rect 42628 672450 42656 681702
rect 42982 677920 43038 677929
rect 42982 677855 43038 677864
rect 42798 677104 42854 677113
rect 42798 677039 42854 677048
rect 42812 676258 42840 677039
rect 42800 676252 42852 676258
rect 42800 676194 42852 676200
rect 42800 672580 42852 672586
rect 42800 672522 42852 672528
rect 42616 672444 42668 672450
rect 42616 672386 42668 672392
rect 42812 672330 42840 672522
rect 42168 669718 42288 669746
rect 42628 672302 42840 672330
rect 41970 668536 42026 668545
rect 41970 668471 42026 668480
rect 41984 668032 42012 668471
rect 42154 667720 42210 667729
rect 42154 667655 42210 667664
rect 42168 667352 42196 667655
rect 42338 667448 42394 667457
rect 42394 667406 42564 667434
rect 42338 667383 42394 667392
rect 42062 667040 42118 667049
rect 42118 666998 42472 667026
rect 42062 666975 42118 666984
rect 42248 666936 42300 666942
rect 42248 666878 42300 666884
rect 42260 666179 42288 666878
rect 42444 666179 42472 666998
rect 42182 666151 42288 666179
rect 42352 666151 42472 666179
rect 42352 665938 42380 666151
rect 42168 665910 42380 665938
rect 42168 665516 42196 665910
rect 42340 665712 42392 665718
rect 42340 665654 42392 665660
rect 41786 665272 41842 665281
rect 41786 665207 41842 665216
rect 41800 664972 41828 665207
rect 42352 664339 42380 665654
rect 42182 664311 42380 664339
rect 41786 664184 41842 664193
rect 41786 664119 41842 664128
rect 41800 663680 41828 664119
rect 42536 663150 42564 667406
rect 42182 663122 42564 663150
rect 42248 663060 42300 663066
rect 42248 663002 42300 663008
rect 42260 660770 42288 663002
rect 42432 662924 42484 662930
rect 42432 662866 42484 662872
rect 42168 660742 42288 660770
rect 42168 660620 42196 660742
rect 42444 660022 42472 662866
rect 42182 659994 42472 660022
rect 42628 659654 42656 672302
rect 42800 672240 42852 672246
rect 42536 659626 42656 659654
rect 42720 672188 42800 672194
rect 42720 672182 42852 672188
rect 42720 672166 42840 672182
rect 42536 659371 42564 659626
rect 42182 659343 42564 659371
rect 42168 658838 42380 658866
rect 42168 658784 42196 658838
rect 42352 658798 42380 658838
rect 42720 658798 42748 672166
rect 42352 658770 42748 658798
rect 42522 658608 42578 658617
rect 42352 658566 42522 658594
rect 41800 658430 42288 658458
rect 41800 658345 41828 658430
rect 41786 658336 41842 658345
rect 41786 658271 41842 658280
rect 41786 657248 41842 657257
rect 41786 657183 41842 657192
rect 41800 656948 41828 657183
rect 42260 656350 42288 658430
rect 42182 656322 42288 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42352 655670 42380 658566
rect 42522 658543 42578 658552
rect 42524 657552 42576 657558
rect 42524 657494 42576 657500
rect 42260 655642 42380 655670
rect 42536 655126 42564 657494
rect 42182 655098 42564 655126
rect 42996 649994 43024 677855
rect 42996 649966 43116 649994
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 35820 644502 35848 644671
rect 35808 644496 35860 644502
rect 35808 644438 35860 644444
rect 39764 644496 39816 644502
rect 39764 644438 39816 644444
rect 38566 644328 38622 644337
rect 38566 644263 38622 644272
rect 39578 644328 39634 644337
rect 39578 644263 39634 644272
rect 35346 643920 35402 643929
rect 35346 643855 35402 643864
rect 35360 643142 35388 643855
rect 35808 643544 35860 643550
rect 35530 643512 35586 643521
rect 35530 643447 35586 643456
rect 35806 643512 35808 643521
rect 35860 643512 35862 643521
rect 35806 643447 35862 643456
rect 35544 643278 35572 643447
rect 35532 643272 35584 643278
rect 35532 643214 35584 643220
rect 35348 643136 35400 643142
rect 35348 643078 35400 643084
rect 35806 642696 35862 642705
rect 35806 642631 35862 642640
rect 35622 642288 35678 642297
rect 35622 642223 35678 642232
rect 35636 641782 35664 642223
rect 35820 642190 35848 642631
rect 38580 642530 38608 644263
rect 38568 642524 38620 642530
rect 38568 642466 38620 642472
rect 39592 642190 39620 644263
rect 39776 643929 39804 644438
rect 39762 643920 39818 643929
rect 39762 643855 39818 643864
rect 40224 643544 40276 643550
rect 40224 643486 40276 643492
rect 35808 642184 35860 642190
rect 35808 642126 35860 642132
rect 39580 642184 39632 642190
rect 39580 642126 39632 642132
rect 35808 641912 35860 641918
rect 35806 641880 35808 641889
rect 35860 641880 35862 641889
rect 35806 641815 35862 641824
rect 35624 641776 35676 641782
rect 35624 641718 35676 641724
rect 35622 641472 35678 641481
rect 35622 641407 35678 641416
rect 35636 640354 35664 641407
rect 35806 641064 35862 641073
rect 35806 640999 35862 641008
rect 39302 641064 39358 641073
rect 39302 640999 39358 641008
rect 35820 640830 35848 640999
rect 35808 640824 35860 640830
rect 35808 640766 35860 640772
rect 39316 640762 39344 640999
rect 39304 640756 39356 640762
rect 39304 640698 39356 640704
rect 35806 640656 35862 640665
rect 35806 640591 35862 640600
rect 35820 640490 35848 640591
rect 35808 640484 35860 640490
rect 35808 640426 35860 640432
rect 35624 640348 35676 640354
rect 35624 640290 35676 640296
rect 40236 640257 40264 643486
rect 41708 643346 42104 643362
rect 41696 643340 42116 643346
rect 41748 643334 42064 643340
rect 41696 643282 41748 643288
rect 42064 643282 42116 643288
rect 41696 643136 41748 643142
rect 42064 643136 42116 643142
rect 41748 643084 42064 643090
rect 41696 643078 42116 643084
rect 41708 643062 42104 643078
rect 41696 642524 41748 642530
rect 41748 642484 42104 642512
rect 41696 642466 41748 642472
rect 42076 642394 42104 642484
rect 42064 642388 42116 642394
rect 42064 642330 42116 642336
rect 40774 642288 40830 642297
rect 40774 642223 40830 642232
rect 40788 642054 40816 642223
rect 40776 642048 40828 642054
rect 40776 641990 40828 641996
rect 41696 641776 41748 641782
rect 42064 641776 42116 641782
rect 41748 641724 42064 641730
rect 41696 641718 42116 641724
rect 41708 641702 42104 641718
rect 40408 640552 40460 640558
rect 40408 640494 40460 640500
rect 40222 640248 40278 640257
rect 40222 640183 40278 640192
rect 34426 639840 34482 639849
rect 34426 639775 34482 639784
rect 34440 638246 34468 639775
rect 40420 639441 40448 640494
rect 40868 640348 40920 640354
rect 40868 640290 40920 640296
rect 35530 639432 35586 639441
rect 35530 639367 35586 639376
rect 35806 639432 35862 639441
rect 35806 639367 35862 639376
rect 40406 639432 40462 639441
rect 40406 639367 40462 639376
rect 35544 638994 35572 639367
rect 35820 639266 35848 639367
rect 35808 639260 35860 639266
rect 35808 639202 35860 639208
rect 40880 639033 40908 640290
rect 41696 639260 41748 639266
rect 41696 639202 41748 639208
rect 41708 639146 41736 639202
rect 41708 639118 42380 639146
rect 40866 639024 40922 639033
rect 35532 638988 35584 638994
rect 35532 638930 35584 638936
rect 39304 638988 39356 638994
rect 40866 638959 40922 638968
rect 39304 638930 39356 638936
rect 35622 638616 35678 638625
rect 35622 638551 35678 638560
rect 34428 638240 34480 638246
rect 34428 638182 34480 638188
rect 32402 637800 32458 637809
rect 32402 637735 32458 637744
rect 32416 629921 32444 637735
rect 35162 637392 35218 637401
rect 35162 637327 35218 637336
rect 32402 629912 32458 629921
rect 32402 629847 32458 629856
rect 35176 628590 35204 637327
rect 35636 636954 35664 638551
rect 35806 638208 35862 638217
rect 35806 638143 35862 638152
rect 35820 637906 35848 638143
rect 35808 637900 35860 637906
rect 35808 637842 35860 637848
rect 36544 637900 36596 637906
rect 36544 637842 36596 637848
rect 35806 636984 35862 636993
rect 35624 636948 35676 636954
rect 35806 636919 35862 636928
rect 35624 636890 35676 636896
rect 35820 636750 35848 636919
rect 35808 636744 35860 636750
rect 35808 636686 35860 636692
rect 35530 636576 35586 636585
rect 35530 636511 35586 636520
rect 35806 636576 35862 636585
rect 35806 636511 35862 636520
rect 35544 636274 35572 636511
rect 35820 636410 35848 636511
rect 35808 636404 35860 636410
rect 35808 636346 35860 636352
rect 35532 636268 35584 636274
rect 35532 636210 35584 636216
rect 35806 635760 35862 635769
rect 35806 635695 35862 635704
rect 35820 634846 35848 635695
rect 35808 634840 35860 634846
rect 35808 634782 35860 634788
rect 35806 634536 35862 634545
rect 35806 634471 35862 634480
rect 35820 633894 35848 634471
rect 35808 633888 35860 633894
rect 35808 633830 35860 633836
rect 35806 633720 35862 633729
rect 35806 633655 35862 633664
rect 35820 633486 35848 633655
rect 35808 633480 35860 633486
rect 35808 633422 35860 633428
rect 36556 630630 36584 637842
rect 36544 630624 36596 630630
rect 36544 630566 36596 630572
rect 39316 629241 39344 638930
rect 41696 638240 41748 638246
rect 41696 638182 41748 638188
rect 40592 636948 40644 636954
rect 40592 636890 40644 636896
rect 40132 636676 40184 636682
rect 40132 636618 40184 636624
rect 39948 634840 40000 634846
rect 39948 634782 40000 634788
rect 39960 632913 39988 634782
rect 39946 632904 40002 632913
rect 39946 632839 40002 632848
rect 40144 632505 40172 636618
rect 40604 636585 40632 636890
rect 40590 636576 40646 636585
rect 40590 636511 40646 636520
rect 40776 636472 40828 636478
rect 40776 636414 40828 636420
rect 40592 636268 40644 636274
rect 40592 636210 40644 636216
rect 40604 634545 40632 636210
rect 40590 634536 40646 634545
rect 40590 634471 40646 634480
rect 40500 633752 40552 633758
rect 40500 633694 40552 633700
rect 40130 632496 40186 632505
rect 40130 632431 40186 632440
rect 40512 630601 40540 633694
rect 40788 632233 40816 636414
rect 41512 633480 41564 633486
rect 41512 633422 41564 633428
rect 41524 633321 41552 633422
rect 41510 633312 41566 633321
rect 41510 633247 41566 633256
rect 40774 632224 40830 632233
rect 40774 632159 40830 632168
rect 41708 630674 41736 638182
rect 42156 633480 42208 633486
rect 42156 633422 42208 633428
rect 42168 633321 42196 633422
rect 42154 633312 42210 633321
rect 42154 633247 42210 633256
rect 41708 630646 42288 630674
rect 40498 630592 40554 630601
rect 40498 630527 40554 630536
rect 41604 630556 41656 630562
rect 41604 630498 41656 630504
rect 41616 630442 41644 630498
rect 41616 630414 41828 630442
rect 39302 629232 39358 629241
rect 39302 629167 39358 629176
rect 35164 628584 35216 628590
rect 35164 628526 35216 628532
rect 39672 628584 39724 628590
rect 39672 628526 39724 628532
rect 39684 628289 39712 628526
rect 39670 628280 39726 628289
rect 39670 628215 39726 628224
rect 41800 627473 41828 630414
rect 41786 627464 41842 627473
rect 41786 627399 41842 627408
rect 41786 627192 41842 627201
rect 41786 627127 41842 627136
rect 41800 626620 41828 627127
rect 42260 625274 42288 630646
rect 42168 625246 42288 625274
rect 42352 625274 42380 639118
rect 42522 636576 42578 636585
rect 42522 636511 42578 636520
rect 42536 625977 42564 636511
rect 42890 632904 42946 632913
rect 42890 632839 42946 632848
rect 42706 628280 42762 628289
rect 42706 628215 42762 628224
rect 42720 627914 42748 628215
rect 42720 627886 42840 627914
rect 42522 625968 42578 625977
rect 42522 625903 42578 625912
rect 42352 625246 42564 625274
rect 42168 624784 42196 625246
rect 42340 625184 42392 625190
rect 42340 625126 42392 625132
rect 42154 624608 42210 624617
rect 42154 624543 42210 624552
rect 42168 624172 42196 624543
rect 42352 623642 42380 625126
rect 42260 623614 42380 623642
rect 42260 623506 42288 623614
rect 41800 623478 42288 623506
rect 41800 622948 41828 623478
rect 42340 623416 42392 623422
rect 41970 623384 42026 623393
rect 42340 623358 42392 623364
rect 41970 623319 42026 623328
rect 41984 623234 42012 623319
rect 41984 623206 42288 623234
rect 42076 622169 42104 622336
rect 42062 622160 42118 622169
rect 42062 622095 42118 622104
rect 42168 621738 42196 621792
rect 42260 621738 42288 623206
rect 42168 621710 42288 621738
rect 42352 621602 42380 623358
rect 42536 623234 42564 625246
rect 42168 621574 42380 621602
rect 42444 623206 42564 623234
rect 42168 621112 42196 621574
rect 42444 621518 42472 623206
rect 42432 621512 42484 621518
rect 42432 621454 42484 621460
rect 42812 621330 42840 627886
rect 42444 621302 42840 621330
rect 41786 620936 41842 620945
rect 41786 620871 41842 620880
rect 41800 620500 41828 620871
rect 41970 620256 42026 620265
rect 41970 620191 42026 620200
rect 41984 619956 42012 620191
rect 42248 619676 42300 619682
rect 42248 619618 42300 619624
rect 42260 617454 42288 619618
rect 42182 617426 42288 617454
rect 42156 617160 42208 617166
rect 42156 617102 42208 617108
rect 42168 616978 42196 617102
rect 42076 616950 42196 616978
rect 42076 616828 42104 616950
rect 42444 616570 42472 621302
rect 42616 621240 42668 621246
rect 42616 621182 42668 621188
rect 42628 620786 42656 621182
rect 42168 616542 42472 616570
rect 42536 620758 42656 620786
rect 42536 616570 42564 620758
rect 42904 619682 42932 632839
rect 42892 619676 42944 619682
rect 42892 619618 42944 619624
rect 42708 618928 42760 618934
rect 42708 618870 42760 618876
rect 42720 617166 42748 618870
rect 42708 617160 42760 617166
rect 42708 617102 42760 617108
rect 42706 616856 42762 616865
rect 42706 616791 42762 616800
rect 42536 616542 42656 616570
rect 42168 616148 42196 616542
rect 42430 616448 42486 616457
rect 42430 616383 42486 616392
rect 42062 615904 42118 615913
rect 42062 615839 42118 615848
rect 42076 615604 42104 615839
rect 42444 613782 42472 616383
rect 42628 615913 42656 616542
rect 42720 616026 42748 616791
rect 42720 615998 42840 616026
rect 42614 615904 42670 615913
rect 42614 615839 42670 615848
rect 42812 615754 42840 615998
rect 42720 615726 42840 615754
rect 42720 615618 42748 615726
rect 42182 613754 42472 613782
rect 42536 615590 42748 615618
rect 42536 613135 42564 615590
rect 42706 615496 42762 615505
rect 42706 615431 42762 615440
rect 42720 615346 42748 615431
rect 42182 613107 42564 613135
rect 42628 615318 42748 615346
rect 42628 612490 42656 615318
rect 42800 614168 42852 614174
rect 42182 612462 42656 612490
rect 42720 614116 42800 614122
rect 42720 614110 42852 614116
rect 42720 614094 42840 614110
rect 42248 612400 42300 612406
rect 42246 612368 42248 612377
rect 42300 612368 42302 612377
rect 42246 612303 42302 612312
rect 42720 612082 42748 614094
rect 43088 612882 43116 649966
rect 43076 612876 43128 612882
rect 43076 612818 43128 612824
rect 43272 612678 43300 807434
rect 43456 773537 43484 815730
rect 44732 814292 44784 814298
rect 44732 814234 44784 814240
rect 44180 812864 44232 812870
rect 44180 812806 44232 812812
rect 43628 799128 43680 799134
rect 43628 799070 43680 799076
rect 43640 797337 43668 799070
rect 43812 797700 43864 797706
rect 43812 797642 43864 797648
rect 43626 797328 43682 797337
rect 43626 797263 43682 797272
rect 43824 795666 43852 797642
rect 43812 795660 43864 795666
rect 43812 795602 43864 795608
rect 43442 773528 43498 773537
rect 43442 773463 43498 773472
rect 44192 770098 44220 812806
rect 44364 807356 44416 807362
rect 44364 807298 44416 807304
rect 44376 794918 44404 807298
rect 44364 794912 44416 794918
rect 44364 794854 44416 794860
rect 44548 773016 44600 773022
rect 44548 772958 44600 772964
rect 44364 771452 44416 771458
rect 44364 771394 44416 771400
rect 44180 770092 44232 770098
rect 44180 770034 44232 770040
rect 43442 769448 43498 769457
rect 43442 769383 43498 769392
rect 43456 727462 43484 769383
rect 44178 764552 44234 764561
rect 44178 764487 44234 764496
rect 43626 764144 43682 764153
rect 43626 764079 43682 764088
rect 43640 750961 43668 764079
rect 44192 753574 44220 764487
rect 44180 753568 44232 753574
rect 44180 753510 44232 753516
rect 43626 750952 43682 750961
rect 43626 750887 43682 750896
rect 43626 731368 43682 731377
rect 43626 731303 43682 731312
rect 43640 730386 43668 731303
rect 43628 730380 43680 730386
rect 43628 730322 43680 730328
rect 44178 729736 44234 729745
rect 44178 729671 44234 729680
rect 43444 727456 43496 727462
rect 43444 727398 43496 727404
rect 43444 727320 43496 727326
rect 43444 727262 43496 727268
rect 43456 685137 43484 727262
rect 44192 724514 44220 729671
rect 44376 728822 44404 771394
rect 44560 730153 44588 772958
rect 44744 771662 44772 814234
rect 50344 806132 50396 806138
rect 50344 806074 50396 806080
rect 46202 773120 46258 773129
rect 46202 773055 46258 773064
rect 44732 771656 44784 771662
rect 44732 771598 44784 771604
rect 44730 765776 44786 765785
rect 44730 765711 44786 765720
rect 44744 754934 44772 765711
rect 44914 763328 44970 763337
rect 44914 763263 44970 763272
rect 44732 754928 44784 754934
rect 44732 754870 44784 754876
rect 44546 730144 44602 730153
rect 44546 730079 44602 730088
rect 44364 728816 44416 728822
rect 44364 728758 44416 728764
rect 44548 728680 44600 728686
rect 44548 728622 44600 728628
rect 44192 724486 44312 724514
rect 43994 723616 44050 723625
rect 43994 723551 44050 723560
rect 43626 721168 43682 721177
rect 43626 721103 43682 721112
rect 43442 685128 43498 685137
rect 43442 685063 43498 685072
rect 43442 684312 43498 684321
rect 43442 684247 43498 684256
rect 43456 644337 43484 684247
rect 43442 644328 43498 644337
rect 43442 644263 43498 644272
rect 43640 630674 43668 721103
rect 43812 712292 43864 712298
rect 43812 712234 43864 712240
rect 43824 711142 43852 712234
rect 43812 711136 43864 711142
rect 43812 711078 43864 711084
rect 43812 711000 43864 711006
rect 43812 710942 43864 710948
rect 43824 707713 43852 710942
rect 43810 707704 43866 707713
rect 43810 707639 43866 707648
rect 44008 703497 44036 723551
rect 43994 703488 44050 703497
rect 43994 703423 44050 703432
rect 43812 686316 43864 686322
rect 43812 686258 43864 686264
rect 43824 643346 43852 686258
rect 44284 685914 44312 724486
rect 44560 686118 44588 728622
rect 44730 722800 44786 722809
rect 44730 722735 44786 722744
rect 44744 711006 44772 722735
rect 44732 711000 44784 711006
rect 44732 710942 44784 710948
rect 44730 708520 44786 708529
rect 44730 708455 44786 708464
rect 44744 703798 44772 708455
rect 44732 703792 44784 703798
rect 44732 703734 44784 703740
rect 44548 686112 44600 686118
rect 44548 686054 44600 686060
rect 44272 685908 44324 685914
rect 44272 685850 44324 685856
rect 44364 683188 44416 683194
rect 44364 683130 44416 683136
rect 43994 679416 44050 679425
rect 43994 679351 44050 679360
rect 44008 663066 44036 679351
rect 44180 679244 44232 679250
rect 44180 679186 44232 679192
rect 44192 666942 44220 679186
rect 44180 666936 44232 666942
rect 44180 666878 44232 666884
rect 43996 663060 44048 663066
rect 43996 663002 44048 663008
rect 43812 643340 43864 643346
rect 43812 643282 43864 643288
rect 44376 641073 44404 683130
rect 44640 679040 44692 679046
rect 44640 678982 44692 678988
rect 44652 666602 44680 678982
rect 44640 666596 44692 666602
rect 44640 666538 44692 666544
rect 44362 641064 44418 641073
rect 44362 640999 44418 641008
rect 44546 640248 44602 640257
rect 44546 640183 44602 640192
rect 44362 634536 44418 634545
rect 44362 634471 44418 634480
rect 43810 632496 43866 632505
rect 43810 632431 43866 632440
rect 43640 630646 43760 630674
rect 43534 630592 43590 630601
rect 43534 630527 43590 630536
rect 43260 612672 43312 612678
rect 43260 612614 43312 612620
rect 42536 612054 42748 612082
rect 42536 611946 42564 612054
rect 42182 611918 42564 611946
rect 43548 611017 43576 630527
rect 43732 616162 43760 630646
rect 43824 627914 43852 632431
rect 43994 632224 44050 632233
rect 43994 632159 44050 632168
rect 43824 627886 43944 627914
rect 43916 618934 43944 627886
rect 44008 623914 44036 632159
rect 44180 625864 44232 625870
rect 44180 625806 44232 625812
rect 44192 624617 44220 625806
rect 44376 625190 44404 634471
rect 44364 625184 44416 625190
rect 44364 625126 44416 625132
rect 44178 624608 44234 624617
rect 44178 624543 44234 624552
rect 44008 623886 44128 623914
rect 44100 623830 44128 623886
rect 44088 623824 44140 623830
rect 44088 623766 44140 623772
rect 44178 622160 44234 622169
rect 44178 622095 44234 622104
rect 43904 618928 43956 618934
rect 43904 618870 43956 618876
rect 44192 616826 44220 622095
rect 44180 616820 44232 616826
rect 44180 616762 44232 616768
rect 43732 616134 44128 616162
rect 43904 612740 43956 612746
rect 43904 612682 43956 612688
rect 43916 611354 43944 612682
rect 44100 611590 44128 616134
rect 44088 611584 44140 611590
rect 44088 611526 44140 611532
rect 43916 611326 44128 611354
rect 44100 611266 44128 611326
rect 44100 611238 44358 611266
rect 44330 611182 44358 611238
rect 44318 611176 44370 611182
rect 44318 611118 44370 611124
rect 43534 611008 43590 611017
rect 43534 610943 43590 610952
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 40314 602032 40370 602041
rect 40314 601967 40370 601976
rect 33782 601760 33838 601769
rect 33782 601695 33838 601704
rect 33046 595232 33102 595241
rect 33046 595167 33102 595176
rect 31022 594416 31078 594425
rect 31022 594351 31078 594360
rect 31036 585750 31064 594351
rect 33060 587178 33088 595167
rect 33796 589665 33824 601695
rect 39946 601352 40002 601361
rect 39946 601287 40002 601296
rect 37922 595810 37978 595819
rect 37922 595745 37978 595754
rect 35162 594824 35218 594833
rect 35162 594759 35218 594768
rect 33782 589656 33838 589665
rect 33782 589591 33838 589600
rect 33048 587172 33100 587178
rect 33048 587114 33100 587120
rect 35176 585993 35204 594759
rect 35622 591968 35678 591977
rect 35622 591903 35678 591912
rect 35636 590714 35664 591903
rect 35806 591560 35862 591569
rect 35806 591495 35862 591504
rect 35820 590986 35848 591495
rect 35808 590980 35860 590986
rect 35808 590922 35860 590928
rect 35624 590708 35676 590714
rect 35624 590650 35676 590656
rect 35162 585984 35218 585993
rect 35162 585919 35218 585928
rect 37936 585886 37964 595745
rect 39960 594726 39988 601287
rect 40130 600944 40186 600953
rect 40130 600879 40186 600888
rect 40144 595814 40172 600879
rect 40132 595808 40184 595814
rect 40132 595750 40184 595756
rect 39948 594720 40000 594726
rect 39948 594662 40000 594668
rect 40328 592034 40356 601967
rect 44560 600545 44588 640183
rect 44928 611998 44956 763263
rect 45100 755540 45152 755546
rect 45100 755482 45152 755488
rect 45112 754322 45140 755482
rect 45100 754316 45152 754322
rect 45100 754258 45152 754264
rect 45098 751768 45154 751777
rect 45098 751703 45154 751712
rect 45112 746570 45140 751703
rect 45100 746564 45152 746570
rect 45100 746506 45152 746512
rect 46216 743782 46244 773055
rect 48964 761932 49016 761938
rect 48964 761874 49016 761880
rect 46204 743776 46256 743782
rect 46204 743718 46256 743724
rect 46202 730960 46258 730969
rect 46202 730895 46258 730904
rect 45098 721576 45154 721585
rect 45098 721511 45154 721520
rect 45112 708801 45140 721511
rect 45098 708792 45154 708801
rect 45098 708727 45154 708736
rect 46216 700330 46244 730895
rect 46204 700324 46256 700330
rect 46204 700266 46256 700272
rect 45282 687576 45338 687585
rect 45282 687511 45338 687520
rect 45100 684956 45152 684962
rect 45100 684898 45152 684904
rect 45112 642297 45140 684898
rect 45296 678974 45324 687511
rect 46202 687168 46258 687177
rect 46202 687103 46258 687112
rect 45466 680640 45522 680649
rect 45466 680575 45522 680584
rect 45204 678946 45324 678974
rect 45204 669314 45232 678946
rect 45204 669286 45416 669314
rect 45388 658986 45416 669286
rect 45480 662946 45508 680575
rect 45836 669452 45888 669458
rect 45836 669394 45888 669400
rect 45652 667956 45704 667962
rect 45652 667898 45704 667904
rect 45664 667049 45692 667898
rect 45848 667729 45876 669394
rect 45834 667720 45890 667729
rect 45834 667655 45890 667664
rect 45650 667040 45706 667049
rect 45650 666975 45706 666984
rect 45480 662930 45600 662946
rect 45480 662924 45612 662930
rect 45480 662918 45560 662924
rect 45560 662866 45612 662872
rect 45376 658980 45428 658986
rect 45376 658922 45428 658928
rect 46216 656878 46244 687103
rect 46204 656872 46256 656878
rect 46204 656814 46256 656820
rect 46202 643920 46258 643929
rect 46202 643855 46258 643864
rect 45098 642288 45154 642297
rect 45098 642223 45154 642232
rect 45284 641776 45336 641782
rect 45284 641718 45336 641724
rect 45098 639432 45154 639441
rect 45098 639367 45154 639376
rect 44916 611992 44968 611998
rect 44916 611934 44968 611940
rect 44730 611008 44786 611017
rect 44730 610943 44786 610952
rect 44744 610774 44772 610943
rect 44732 610768 44784 610774
rect 44732 610710 44784 610716
rect 44546 600536 44602 600545
rect 44546 600471 44602 600480
rect 44914 600128 44970 600137
rect 44914 600063 44970 600072
rect 44638 599312 44694 599321
rect 44638 599247 44694 599256
rect 43074 597680 43130 597689
rect 43074 597615 43130 597624
rect 43088 597446 43116 597615
rect 43076 597440 43128 597446
rect 43076 597382 43128 597388
rect 43076 597032 43128 597038
rect 42890 597000 42946 597009
rect 43076 596974 43128 596980
rect 42890 596935 42946 596944
rect 42430 596864 42486 596873
rect 42430 596799 42486 596808
rect 41326 595810 41382 595819
rect 41696 595808 41748 595814
rect 41326 595745 41382 595754
rect 41694 595776 41696 595785
rect 41748 595776 41750 595785
rect 41340 594862 41368 595745
rect 41694 595711 41750 595720
rect 41328 594856 41380 594862
rect 41328 594798 41380 594804
rect 41696 594856 41748 594862
rect 41748 594804 42012 594810
rect 41696 594798 42012 594804
rect 41708 594782 42012 594798
rect 41696 594720 41748 594726
rect 41696 594662 41748 594668
rect 41708 594561 41736 594662
rect 41694 594552 41750 594561
rect 41694 594487 41750 594496
rect 41786 593600 41842 593609
rect 41432 593558 41786 593586
rect 40328 592006 40448 592034
rect 39304 591456 39356 591462
rect 39304 591398 39356 591404
rect 37924 585880 37976 585886
rect 37924 585822 37976 585828
rect 31024 585744 31076 585750
rect 31024 585686 31076 585692
rect 39316 584633 39344 591398
rect 40420 585721 40448 592006
rect 41432 591462 41460 593558
rect 41786 593535 41842 593544
rect 41786 592376 41842 592385
rect 41616 592334 41786 592362
rect 41420 591456 41472 591462
rect 41420 591398 41472 591404
rect 40776 590980 40828 590986
rect 40776 590922 40828 590928
rect 40788 589393 40816 590922
rect 41616 590866 41644 592334
rect 41786 592311 41842 592320
rect 41984 592034 42012 594782
rect 41984 592006 42380 592034
rect 41524 590838 41644 590866
rect 40774 589384 40830 589393
rect 40774 589319 40830 589328
rect 41524 589121 41552 590838
rect 41696 590776 41748 590782
rect 41748 590724 42104 590730
rect 41696 590718 42104 590724
rect 41708 590714 42104 590718
rect 41708 590708 42116 590714
rect 41708 590702 42064 590708
rect 42064 590650 42116 590656
rect 42352 589274 42380 592006
rect 42260 589246 42380 589274
rect 41510 589112 41566 589121
rect 41510 589047 41566 589056
rect 41512 587172 41564 587178
rect 41512 587114 41564 587120
rect 40406 585712 40462 585721
rect 40406 585647 40462 585656
rect 41524 585018 41552 587114
rect 41696 585880 41748 585886
rect 42064 585880 42116 585886
rect 41748 585840 42064 585868
rect 41696 585822 41748 585828
rect 42064 585822 42116 585828
rect 41696 585744 41748 585750
rect 41748 585692 42104 585698
rect 41696 585686 42104 585692
rect 41708 585682 42104 585686
rect 41708 585676 42116 585682
rect 41708 585670 42064 585676
rect 42064 585618 42116 585624
rect 41524 584990 41828 585018
rect 39302 584624 39358 584633
rect 39302 584559 39358 584568
rect 41800 584361 41828 584990
rect 41786 584352 41842 584361
rect 41786 584287 41842 584296
rect 41786 583944 41842 583953
rect 41786 583879 41842 583888
rect 41800 583440 41828 583879
rect 42260 582457 42288 589246
rect 42444 582486 42472 596799
rect 42616 585880 42668 585886
rect 42536 585828 42616 585834
rect 42536 585822 42668 585828
rect 42536 585806 42656 585822
rect 42536 585562 42564 585806
rect 42708 585676 42760 585682
rect 42708 585618 42760 585624
rect 42536 585534 42656 585562
rect 42432 582480 42484 582486
rect 42246 582448 42302 582457
rect 42432 582422 42484 582428
rect 42246 582383 42302 582392
rect 42248 582140 42300 582146
rect 42248 582082 42300 582088
rect 42260 581618 42288 582082
rect 42182 581590 42288 581618
rect 42076 580689 42104 580961
rect 42062 580680 42118 580689
rect 42062 580615 42118 580624
rect 42432 580644 42484 580650
rect 42432 580586 42484 580592
rect 41878 580272 41934 580281
rect 41878 580207 41934 580216
rect 42246 580272 42302 580281
rect 42246 580207 42302 580216
rect 41892 579768 41920 580207
rect 42260 580106 42288 580207
rect 42248 580100 42300 580106
rect 42248 580042 42300 580048
rect 42248 579964 42300 579970
rect 42248 579906 42300 579912
rect 42260 579782 42288 579906
rect 42444 579850 42472 580586
rect 42444 579822 42564 579850
rect 42260 579754 42380 579782
rect 41786 579592 41842 579601
rect 41786 579527 41842 579536
rect 41800 579121 41828 579527
rect 42062 579320 42118 579329
rect 42352 579306 42380 579754
rect 42118 579278 42380 579306
rect 42062 579255 42118 579264
rect 42536 578762 42564 579822
rect 42444 578734 42564 578762
rect 42168 578598 42288 578626
rect 42168 578544 42196 578598
rect 42260 578558 42288 578598
rect 42444 578558 42472 578734
rect 42260 578530 42472 578558
rect 42154 578368 42210 578377
rect 42154 578303 42210 578312
rect 42168 577932 42196 578303
rect 41786 577824 41842 577833
rect 41786 577759 41842 577768
rect 41800 577281 41828 577759
rect 42628 577130 42656 585534
rect 42168 577102 42656 577130
rect 42168 576708 42196 577102
rect 42154 575784 42210 575793
rect 42154 575719 42210 575728
rect 42168 575634 42196 575719
rect 42168 575606 42288 575634
rect 41786 574696 41842 574705
rect 41786 574631 41842 574640
rect 41800 574260 41828 574631
rect 42260 573866 42288 575606
rect 42168 573838 42288 573866
rect 42168 573580 42196 573838
rect 42720 573510 42748 585618
rect 42248 573504 42300 573510
rect 42248 573446 42300 573452
rect 42708 573504 42760 573510
rect 42708 573446 42760 573452
rect 42260 572982 42288 573446
rect 42182 572954 42288 572982
rect 42614 572928 42670 572937
rect 42614 572863 42670 572872
rect 42062 572656 42118 572665
rect 42062 572591 42118 572600
rect 42076 572424 42104 572591
rect 42062 571568 42118 571577
rect 42062 571503 42118 571512
rect 42076 571282 42104 571503
rect 42430 571432 42486 571441
rect 42430 571367 42486 571376
rect 42076 571254 42380 571282
rect 42064 570988 42116 570994
rect 42064 570930 42116 570936
rect 42076 570588 42104 570930
rect 41786 570208 41842 570217
rect 41786 570143 41842 570152
rect 41800 569908 41828 570143
rect 42352 569310 42380 571254
rect 42168 569242 42196 569296
rect 42260 569282 42380 569310
rect 42260 569242 42288 569282
rect 42168 569214 42288 569242
rect 42444 568766 42472 571367
rect 42628 570994 42656 572863
rect 42616 570988 42668 570994
rect 42616 570930 42668 570936
rect 42168 568698 42196 568752
rect 42260 568738 42472 568766
rect 42260 568698 42288 568738
rect 42168 568670 42288 568698
rect 42904 567194 42932 596935
rect 42812 567166 42932 567194
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 40958 558104 41014 558113
rect 40958 558039 41014 558048
rect 37922 553408 37978 553417
rect 37922 553343 37978 553352
rect 29642 551984 29698 551993
rect 29642 551919 29698 551928
rect 29656 547194 29684 551919
rect 29644 547188 29696 547194
rect 29644 547130 29696 547136
rect 37936 542337 37964 553343
rect 40972 550526 41000 558039
rect 42812 555665 42840 567166
rect 42798 555656 42854 555665
rect 42798 555591 42854 555600
rect 43088 554849 43116 596974
rect 44362 593192 44418 593201
rect 44362 593127 44418 593136
rect 43260 590708 43312 590714
rect 43260 590650 43312 590656
rect 43272 580650 43300 590650
rect 43442 589384 43498 589393
rect 43442 589319 43498 589328
rect 43260 580644 43312 580650
rect 43260 580586 43312 580592
rect 43456 563054 43484 589319
rect 43626 581224 43682 581233
rect 43626 581159 43682 581168
rect 43640 579873 43668 581159
rect 43626 579864 43682 579873
rect 43626 579799 43682 579808
rect 44376 578377 44404 593127
rect 44362 578368 44418 578377
rect 44362 578303 44418 578312
rect 43456 563026 43576 563054
rect 43074 554840 43130 554849
rect 43074 554775 43130 554784
rect 41326 553408 41382 553417
rect 41156 553366 41326 553394
rect 40960 550520 41012 550526
rect 40960 550462 41012 550468
rect 41156 550474 41184 553366
rect 41326 553343 41382 553352
rect 43074 550760 43130 550769
rect 43074 550695 43130 550704
rect 41696 550520 41748 550526
rect 41156 550446 41460 550474
rect 42062 550488 42118 550497
rect 41748 550468 42062 550474
rect 41696 550462 42062 550468
rect 41708 550446 42062 550462
rect 41432 550338 41460 550446
rect 42062 550423 42118 550432
rect 41432 550310 42380 550338
rect 40682 549944 40738 549953
rect 40682 549879 40738 549888
rect 39578 547496 39634 547505
rect 39578 547431 39634 547440
rect 39592 542609 39620 547431
rect 40696 545601 40724 549879
rect 41326 548312 41382 548321
rect 41326 548247 41382 548256
rect 41340 548010 41368 548247
rect 41328 548004 41380 548010
rect 41328 547946 41380 547952
rect 41696 547936 41748 547942
rect 42064 547936 42116 547942
rect 41748 547884 42064 547890
rect 41696 547878 42116 547884
rect 41708 547862 42104 547878
rect 41696 547188 41748 547194
rect 41696 547130 41748 547136
rect 40682 545592 40738 545601
rect 40682 545527 40738 545536
rect 41708 543734 41736 547130
rect 42352 543734 42380 550310
rect 42798 549128 42854 549137
rect 42798 549063 42854 549072
rect 41708 543706 42288 543734
rect 42352 543706 42472 543734
rect 39578 542600 39634 542609
rect 39578 542535 39634 542544
rect 37922 542328 37978 542337
rect 37922 542263 37978 542272
rect 42260 540274 42288 543706
rect 42182 540246 42288 540274
rect 42444 538438 42472 543706
rect 42614 539608 42670 539617
rect 42614 539543 42670 539552
rect 42168 538370 42196 538424
rect 42260 538410 42472 538438
rect 42260 538370 42288 538410
rect 42168 538342 42288 538370
rect 42430 538248 42486 538257
rect 42430 538183 42486 538192
rect 42154 537976 42210 537985
rect 42154 537911 42210 537920
rect 42168 537744 42196 537911
rect 42444 536602 42472 538183
rect 42168 536466 42196 536588
rect 42260 536574 42472 536602
rect 42260 536466 42288 536574
rect 42168 536438 42288 536466
rect 42430 536480 42486 536489
rect 42430 536415 42486 536424
rect 42168 535673 42196 535908
rect 42154 535664 42210 535673
rect 42154 535599 42210 535608
rect 42444 535378 42472 536415
rect 42182 535350 42472 535378
rect 42628 534766 42656 539543
rect 42812 536874 42840 549063
rect 42168 534698 42196 534752
rect 42260 534738 42656 534766
rect 42720 536846 42840 536874
rect 42260 534698 42288 534738
rect 42168 534670 42288 534698
rect 42720 534086 42748 536846
rect 42182 534058 42748 534086
rect 42430 533896 42486 533905
rect 42430 533831 42486 533840
rect 42444 533542 42472 533831
rect 42182 533514 42472 533542
rect 42246 533352 42302 533361
rect 42246 533287 42302 533296
rect 42260 531059 42288 533287
rect 43088 532778 43116 550695
rect 43548 550634 43576 563026
rect 44362 556880 44418 556889
rect 44362 556815 44418 556824
rect 43718 554432 43774 554441
rect 43718 554367 43774 554376
rect 43732 554282 43760 554367
rect 43640 554254 43760 554282
rect 43640 550916 43668 554254
rect 43810 552392 43866 552401
rect 43810 552327 43866 552336
rect 43824 551052 43852 552327
rect 43994 551168 44050 551177
rect 43994 551103 44050 551112
rect 43824 551024 43944 551052
rect 43640 550888 43852 550916
rect 43272 550606 43576 550634
rect 43272 548026 43300 550606
rect 43272 547998 43484 548026
rect 43260 547936 43312 547942
rect 43260 547878 43312 547884
rect 42432 532772 42484 532778
rect 42432 532714 42484 532720
rect 43076 532772 43128 532778
rect 43076 532714 43128 532720
rect 42182 531031 42288 531059
rect 42444 530414 42472 532714
rect 42614 531720 42670 531729
rect 42614 531655 42670 531664
rect 42182 530386 42472 530414
rect 42430 530224 42486 530233
rect 42430 530159 42486 530168
rect 42062 529952 42118 529961
rect 42062 529887 42118 529896
rect 42076 529757 42104 529887
rect 42156 529508 42208 529514
rect 42156 529450 42208 529456
rect 42168 529205 42196 529450
rect 42444 529122 42472 530159
rect 42628 529514 42656 531655
rect 42616 529508 42668 529514
rect 42616 529450 42668 529456
rect 42260 529094 42472 529122
rect 42260 527762 42288 529094
rect 42430 529000 42486 529009
rect 42430 528935 42486 528944
rect 42614 529000 42670 529009
rect 42614 528935 42670 528944
rect 42168 527734 42288 527762
rect 42168 527340 42196 527734
rect 42064 527060 42116 527066
rect 42064 527002 42116 527008
rect 42076 526728 42104 527002
rect 42444 526091 42472 528935
rect 42628 527066 42656 528935
rect 42798 527232 42854 527241
rect 42798 527167 42854 527176
rect 42616 527060 42668 527066
rect 42616 527002 42668 527008
rect 42812 526946 42840 527167
rect 42182 526063 42472 526091
rect 42536 526918 42840 526946
rect 42168 525558 42288 525586
rect 42168 525504 42196 525558
rect 42260 525518 42288 525558
rect 42536 525518 42564 526918
rect 42260 525490 42564 525518
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 35806 430128 35862 430137
rect 35806 430063 35862 430072
rect 35820 429214 35848 430063
rect 35808 429208 35860 429214
rect 35808 429150 35860 429156
rect 41328 429208 41380 429214
rect 41328 429150 41380 429156
rect 35806 428496 35862 428505
rect 41340 428482 41368 429150
rect 41786 428496 41842 428505
rect 41340 428454 41786 428482
rect 35806 428431 35862 428440
rect 41786 428431 41842 428440
rect 35820 427990 35848 428431
rect 35808 427984 35860 427990
rect 35808 427926 35860 427932
rect 41604 427984 41656 427990
rect 41604 427926 41656 427932
rect 41616 426578 41644 427926
rect 41786 426592 41842 426601
rect 41616 426550 41786 426578
rect 41786 426527 41842 426536
rect 42890 426592 42946 426601
rect 42890 426527 42946 426536
rect 41142 426048 41198 426057
rect 41142 425983 41198 425992
rect 39302 425640 39358 425649
rect 39302 425575 39358 425584
rect 33046 424824 33102 424833
rect 33046 424759 33102 424768
rect 33060 417450 33088 424759
rect 34518 424416 34574 424425
rect 34518 424351 34574 424360
rect 33782 424008 33838 424017
rect 33782 423943 33838 423952
rect 33048 417444 33100 417450
rect 33048 417386 33100 417392
rect 33796 414633 33824 423943
rect 34532 416090 34560 424351
rect 34520 416084 34572 416090
rect 34520 416026 34572 416032
rect 39316 415313 39344 425575
rect 41156 424386 41184 425983
rect 41144 424380 41196 424386
rect 41144 424322 41196 424328
rect 41696 424380 41748 424386
rect 41696 424322 41748 424328
rect 41708 418154 41736 424322
rect 42706 422784 42762 422793
rect 42706 422719 42762 422728
rect 41878 421968 41934 421977
rect 41878 421903 41934 421912
rect 41892 418713 41920 421903
rect 41878 418704 41934 418713
rect 41878 418639 41934 418648
rect 41708 418126 42288 418154
rect 41696 417444 41748 417450
rect 41696 417386 41748 417392
rect 41708 417330 41736 417386
rect 41708 417314 42104 417330
rect 41708 417308 42116 417314
rect 41708 417302 42064 417308
rect 42064 417250 42116 417256
rect 41604 416084 41656 416090
rect 41604 416026 41656 416032
rect 41616 415970 41644 416026
rect 41616 415942 41828 415970
rect 39302 415304 39358 415313
rect 39302 415239 39358 415248
rect 33782 414624 33838 414633
rect 33782 414559 33838 414568
rect 41800 413545 41828 415942
rect 41786 413536 41842 413545
rect 41786 413471 41842 413480
rect 41786 413128 41842 413137
rect 41786 413063 41842 413072
rect 41800 412624 41828 413063
rect 42260 411346 42288 418126
rect 42524 417308 42576 417314
rect 42524 417250 42576 417256
rect 42168 411318 42288 411346
rect 42168 410788 42196 411318
rect 42182 410162 42472 410190
rect 42248 409828 42300 409834
rect 42248 409770 42300 409776
rect 42260 408966 42288 409770
rect 42182 408938 42288 408966
rect 42168 407946 42196 408340
rect 42444 407969 42472 410162
rect 42536 408494 42564 417250
rect 42720 415394 42748 422719
rect 42720 415366 42840 415394
rect 42812 409850 42840 415366
rect 42720 409834 42840 409850
rect 42708 409828 42840 409834
rect 42760 409822 42840 409828
rect 42708 409770 42760 409776
rect 42536 408466 42656 408494
rect 42430 407960 42486 407969
rect 42168 407918 42288 407946
rect 42260 407810 42288 407918
rect 42430 407895 42486 407904
rect 42076 407561 42104 407796
rect 42260 407782 42472 407810
rect 42248 407720 42300 407726
rect 42248 407662 42300 407668
rect 42062 407552 42118 407561
rect 42062 407487 42118 407496
rect 41800 407017 41828 407116
rect 41786 407008 41842 407017
rect 41786 406943 41842 406952
rect 41786 406736 41842 406745
rect 41786 406671 41842 406680
rect 41800 406504 41828 406671
rect 42260 406042 42288 407662
rect 42168 406014 42288 406042
rect 42168 405929 42196 406014
rect 42444 404977 42472 407782
rect 42628 407726 42656 408466
rect 42616 407720 42668 407726
rect 42616 407662 42668 407668
rect 42430 404968 42486 404977
rect 42430 404903 42486 404912
rect 42246 404560 42302 404569
rect 42246 404495 42302 404504
rect 42260 403458 42288 404495
rect 42182 403430 42288 403458
rect 42338 402928 42394 402937
rect 42168 402886 42338 402914
rect 42168 402801 42196 402886
rect 42338 402863 42394 402872
rect 42430 402520 42486 402529
rect 42430 402455 42486 402464
rect 42444 402166 42472 402455
rect 42182 402138 42472 402166
rect 42430 401976 42486 401985
rect 42430 401911 42486 401920
rect 42444 401622 42472 401911
rect 42182 401594 42472 401622
rect 41786 400072 41842 400081
rect 41786 400007 41842 400016
rect 41800 399772 41828 400007
rect 41970 399392 42026 399401
rect 41970 399327 42026 399336
rect 41984 399121 42012 399327
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 42168 397497 42196 397936
rect 42154 397488 42210 397497
rect 42154 397423 42210 397432
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41326 387152 41382 387161
rect 41326 387087 41382 387096
rect 41142 386744 41198 386753
rect 41142 386679 41198 386688
rect 41156 385937 41184 386679
rect 41340 386442 41368 387087
rect 41328 386436 41380 386442
rect 41328 386378 41380 386384
rect 41604 386436 41656 386442
rect 41656 386396 41828 386424
rect 41604 386378 41656 386384
rect 40866 385928 40922 385937
rect 40866 385863 40922 385872
rect 41142 385928 41198 385937
rect 41142 385863 41198 385872
rect 40880 382673 40908 385863
rect 41050 383072 41106 383081
rect 41050 383007 41106 383016
rect 41326 383072 41382 383081
rect 41326 383007 41382 383016
rect 40866 382664 40922 382673
rect 40866 382599 40922 382608
rect 40038 382256 40094 382265
rect 40038 382191 40094 382200
rect 35530 381848 35586 381857
rect 35530 381783 35586 381792
rect 33966 381032 34022 381041
rect 33966 380967 34022 380976
rect 33980 373318 34008 380967
rect 35544 374649 35572 381783
rect 39302 381440 39358 381449
rect 39302 381375 39358 381384
rect 35808 379568 35860 379574
rect 35808 379510 35860 379516
rect 35820 379409 35848 379510
rect 35806 379400 35862 379409
rect 35806 379335 35862 379344
rect 35806 377360 35862 377369
rect 35806 377295 35862 377304
rect 35820 376786 35848 377295
rect 35808 376780 35860 376786
rect 35808 376722 35860 376728
rect 35806 376544 35862 376553
rect 35806 376479 35862 376488
rect 35820 376145 35848 376479
rect 35806 376136 35862 376145
rect 35806 376071 35862 376080
rect 35530 374640 35586 374649
rect 35530 374575 35586 374584
rect 33968 373312 34020 373318
rect 33968 373254 34020 373260
rect 39316 371686 39344 381375
rect 40052 379409 40080 382191
rect 41064 381857 41092 383007
rect 41340 382566 41368 383007
rect 41328 382560 41380 382566
rect 41328 382502 41380 382508
rect 41604 382560 41656 382566
rect 41604 382502 41656 382508
rect 41050 381848 41106 381857
rect 41050 381783 41106 381792
rect 40408 379568 40460 379574
rect 40408 379510 40460 379516
rect 41616 379514 41644 382502
rect 41800 381585 41828 386396
rect 42904 385665 42932 426527
rect 42890 385656 42946 385665
rect 42890 385591 42946 385600
rect 41786 381576 41842 381585
rect 41786 381511 41842 381520
rect 42890 379944 42946 379953
rect 42890 379879 42946 379888
rect 40038 379400 40094 379409
rect 40038 379335 40094 379344
rect 40420 377369 40448 379510
rect 41616 379486 42380 379514
rect 40406 377360 40462 377369
rect 40406 377295 40462 377304
rect 41696 376780 41748 376786
rect 41696 376722 41748 376728
rect 41708 376553 41736 376722
rect 41510 376544 41566 376553
rect 41510 376479 41566 376488
rect 41694 376544 41750 376553
rect 41694 376479 41750 376488
rect 41524 376145 41552 376479
rect 41510 376136 41566 376145
rect 41510 376071 41566 376080
rect 41696 373312 41748 373318
rect 41748 373260 42288 373266
rect 41696 373254 42288 373260
rect 41708 373238 42288 373254
rect 39304 371680 39356 371686
rect 39304 371622 39356 371628
rect 41696 371680 41748 371686
rect 41748 371628 42104 371634
rect 41696 371622 42104 371628
rect 41708 371618 42104 371622
rect 41708 371612 42116 371618
rect 41708 371606 42064 371612
rect 42064 371554 42116 371560
rect 42260 369458 42288 373238
rect 42182 369430 42288 369458
rect 42352 367622 42380 379486
rect 42524 371612 42576 371618
rect 42524 371554 42576 371560
rect 42536 369854 42564 371554
rect 42182 367594 42380 367622
rect 42444 369826 42564 369854
rect 42182 366947 42288 366975
rect 42062 366208 42118 366217
rect 42062 366143 42118 366152
rect 42076 365772 42104 366143
rect 42260 365362 42288 366947
rect 42248 365356 42300 365362
rect 42248 365298 42300 365304
rect 41786 364848 41842 364857
rect 41786 364783 41842 364792
rect 41800 364548 41828 364783
rect 42168 364698 42196 365121
rect 42168 364670 42288 364698
rect 41786 364168 41842 364177
rect 41786 364103 41842 364112
rect 41800 363936 41828 364103
rect 42062 363624 42118 363633
rect 42062 363559 42118 363568
rect 42076 363256 42104 363559
rect 42260 362914 42288 364670
rect 42248 362908 42300 362914
rect 42248 362850 42300 362856
rect 42444 362794 42472 369826
rect 42614 365800 42670 365809
rect 42614 365735 42670 365744
rect 42168 362766 42288 362794
rect 42168 362712 42196 362766
rect 42260 362726 42288 362766
rect 42352 362766 42472 362794
rect 42352 362726 42380 362766
rect 42260 362698 42380 362726
rect 42248 362636 42300 362642
rect 42248 362578 42300 362584
rect 42260 362273 42288 362578
rect 42246 362264 42302 362273
rect 42246 362199 42302 362208
rect 41800 360097 41828 360264
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 42156 359984 42208 359990
rect 42156 359926 42208 359932
rect 42168 359584 42196 359926
rect 42430 359000 42486 359009
rect 42182 358958 42430 358986
rect 42430 358935 42486 358944
rect 41878 358728 41934 358737
rect 41878 358663 41934 358672
rect 41892 358428 41920 358663
rect 41786 356960 41842 356969
rect 41786 356895 41842 356904
rect 41800 356592 41828 356895
rect 42246 356144 42302 356153
rect 42246 356079 42302 356088
rect 42260 355926 42288 356079
rect 42182 355898 42288 355926
rect 42628 355314 42656 365735
rect 42904 359990 42932 379879
rect 43074 377360 43130 377369
rect 43074 377295 43130 377304
rect 43088 366217 43116 377295
rect 43074 366208 43130 366217
rect 43074 366143 43130 366152
rect 43076 365356 43128 365362
rect 43076 365298 43128 365304
rect 43088 364313 43116 365298
rect 43074 364304 43130 364313
rect 43074 364239 43130 364248
rect 42892 359984 42944 359990
rect 42892 359926 42944 359932
rect 42798 356688 42854 356697
rect 42798 356623 42854 356632
rect 42168 355178 42196 355300
rect 42260 355286 42656 355314
rect 42260 355178 42288 355286
rect 42168 355150 42288 355178
rect 42812 354770 42840 356623
rect 43272 355337 43300 547878
rect 43258 355328 43314 355337
rect 43258 355263 43314 355272
rect 42536 354742 42840 354770
rect 42536 354739 42564 354742
rect 42182 354711 42564 354739
rect 43456 354674 43484 547998
rect 43824 545986 43852 550888
rect 43640 545958 43852 545986
rect 43640 427281 43668 545958
rect 43916 540974 43944 551024
rect 43824 540946 43944 540974
rect 43824 533905 43852 540946
rect 43810 533896 43866 533905
rect 43810 533831 43866 533840
rect 44008 529961 44036 551103
rect 44178 550216 44234 550225
rect 44178 550151 44234 550160
rect 44192 538257 44220 550151
rect 44178 538248 44234 538257
rect 44178 538183 44234 538192
rect 43994 529952 44050 529961
rect 43994 529887 44050 529896
rect 44376 429729 44404 556815
rect 44652 556481 44680 599247
rect 44928 558793 44956 600063
rect 45112 598097 45140 639367
rect 45296 599729 45324 641718
rect 45466 639024 45522 639033
rect 45466 638959 45522 638968
rect 45282 599720 45338 599729
rect 45282 599655 45338 599664
rect 45480 598913 45508 638959
rect 46216 613426 46244 643855
rect 46204 613420 46256 613426
rect 46204 613362 46256 613368
rect 46204 611720 46256 611726
rect 46204 611662 46256 611668
rect 45466 598904 45522 598913
rect 45466 598839 45522 598848
rect 45098 598088 45154 598097
rect 45098 598023 45154 598032
rect 45098 580680 45154 580689
rect 45098 580615 45154 580624
rect 45112 575482 45140 580615
rect 45100 575476 45152 575482
rect 45100 575418 45152 575424
rect 44914 558784 44970 558793
rect 44914 558719 44970 558728
rect 44638 556472 44694 556481
rect 44638 556407 44694 556416
rect 44546 556064 44602 556073
rect 44546 555999 44602 556008
rect 44362 429720 44418 429729
rect 44362 429655 44418 429664
rect 44178 429312 44234 429321
rect 44178 429247 44234 429256
rect 43626 427272 43682 427281
rect 43626 427207 43682 427216
rect 43994 425232 44050 425241
rect 43994 425167 44050 425176
rect 43810 423600 43866 423609
rect 43810 423535 43866 423544
rect 43626 420744 43682 420753
rect 43626 420679 43682 420688
rect 43640 355609 43668 420679
rect 43824 402529 43852 423535
rect 43810 402520 43866 402529
rect 43810 402455 43866 402464
rect 44008 401985 44036 425167
rect 43994 401976 44050 401985
rect 43994 401911 44050 401920
rect 44192 386481 44220 429247
rect 44560 428913 44588 555999
rect 45098 555248 45154 555257
rect 45098 555183 45154 555192
rect 45112 543734 45140 555183
rect 45282 551576 45338 551585
rect 45282 551511 45338 551520
rect 45020 543706 45140 543734
rect 45296 543734 45324 551511
rect 45466 548720 45522 548729
rect 45466 548655 45522 548664
rect 45296 543706 45416 543734
rect 44730 542600 44786 542609
rect 44730 542535 44786 542544
rect 44744 534074 44772 542535
rect 45020 535514 45048 543706
rect 45190 539880 45246 539889
rect 45190 539815 45246 539824
rect 45204 537985 45232 539815
rect 45190 537976 45246 537985
rect 45190 537911 45246 537920
rect 45190 535664 45246 535673
rect 45190 535599 45246 535608
rect 45020 535486 45140 535514
rect 44744 534046 44864 534074
rect 44836 451450 44864 534046
rect 44824 451444 44876 451450
rect 44824 451386 44876 451392
rect 44822 430944 44878 430953
rect 44822 430879 44878 430888
rect 44546 428904 44602 428913
rect 44546 428839 44602 428848
rect 44362 427680 44418 427689
rect 44362 427615 44418 427624
rect 44178 386472 44234 386481
rect 44178 386407 44234 386416
rect 44376 384849 44404 427615
rect 44638 423192 44694 423201
rect 44638 423127 44694 423136
rect 44652 402937 44680 423127
rect 44638 402928 44694 402937
rect 44638 402863 44694 402872
rect 44836 400110 44864 430879
rect 45112 428097 45140 535486
rect 45204 534074 45232 535599
rect 45388 534074 45416 543706
rect 45480 536874 45508 548655
rect 45650 536888 45706 536897
rect 45480 536846 45650 536874
rect 45650 536823 45706 536832
rect 45204 534046 45324 534074
rect 45388 534046 45508 534074
rect 45296 531146 45324 534046
rect 45284 531140 45336 531146
rect 45284 531082 45336 531088
rect 45480 529009 45508 534046
rect 45466 529000 45522 529009
rect 45466 528935 45522 528944
rect 45284 528624 45336 528630
rect 45284 528566 45336 528572
rect 45296 527241 45324 528566
rect 45282 527232 45338 527241
rect 45282 527167 45338 527176
rect 45098 428088 45154 428097
rect 45098 428023 45154 428032
rect 45282 426864 45338 426873
rect 45282 426799 45338 426808
rect 45006 421152 45062 421161
rect 45006 421087 45062 421096
rect 45020 407561 45048 421087
rect 45006 407552 45062 407561
rect 45006 407487 45062 407496
rect 44824 400104 44876 400110
rect 44824 400046 44876 400052
rect 45098 385248 45154 385257
rect 45098 385183 45154 385192
rect 44362 384840 44418 384849
rect 44362 384775 44418 384784
rect 44914 384432 44970 384441
rect 44914 384367 44970 384376
rect 44546 380352 44602 380361
rect 44546 380287 44602 380296
rect 44178 378312 44234 378321
rect 44178 378247 44234 378256
rect 43810 376544 43866 376553
rect 43810 376479 43866 376488
rect 43824 355881 43852 376479
rect 44192 363633 44220 378247
rect 44178 363624 44234 363633
rect 44178 363559 44234 363568
rect 44560 359009 44588 380287
rect 44730 364304 44786 364313
rect 44730 364239 44786 364248
rect 44744 361554 44772 364239
rect 44732 361548 44784 361554
rect 44732 361490 44784 361496
rect 44546 359000 44602 359009
rect 44546 358935 44602 358944
rect 43810 355872 43866 355881
rect 43810 355807 43866 355816
rect 43626 355600 43682 355609
rect 43626 355535 43682 355544
rect 44638 355328 44694 355337
rect 44638 355263 44694 355272
rect 44652 355026 44680 355263
rect 44640 355020 44692 355026
rect 44640 354962 44692 354968
rect 44640 354884 44692 354890
rect 44640 354826 44692 354832
rect 44652 354674 44680 354826
rect 43456 354646 43852 354674
rect 44008 354657 44680 354674
rect 42706 354376 42762 354385
rect 42706 354311 42762 354320
rect 42720 351937 42748 354311
rect 43824 354226 43852 354646
rect 43994 354648 44680 354657
rect 44050 354646 44680 354648
rect 43994 354583 44050 354592
rect 44640 354544 44692 354550
rect 44284 354492 44640 354498
rect 44284 354486 44692 354492
rect 44284 354470 44680 354486
rect 43994 354376 44050 354385
rect 44284 354362 44312 354470
rect 44732 354408 44784 354414
rect 44050 354334 44312 354362
rect 44560 354356 44732 354362
rect 44560 354350 44784 354356
rect 44560 354334 44772 354350
rect 43994 354311 44050 354320
rect 44560 354226 44588 354334
rect 43824 354198 44588 354226
rect 42706 351928 42762 351937
rect 42706 351863 42762 351872
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 35530 344312 35586 344321
rect 35530 344247 35586 344256
rect 35806 344312 35862 344321
rect 35806 344247 35862 344256
rect 35544 343670 35572 344247
rect 35820 343806 35848 344247
rect 44928 343913 44956 384367
rect 45112 345014 45140 385183
rect 45296 384033 45324 426799
rect 45282 384024 45338 384033
rect 45282 383959 45338 383968
rect 45282 383616 45338 383625
rect 45282 383551 45338 383560
rect 45112 344986 45232 345014
rect 39854 343904 39910 343913
rect 39854 343839 39910 343848
rect 44914 343904 44970 343913
rect 44914 343839 44970 343848
rect 35808 343800 35860 343806
rect 35808 343742 35860 343748
rect 35532 343664 35584 343670
rect 35532 343606 35584 343612
rect 33046 343496 33102 343505
rect 33046 343431 33102 343440
rect 33060 341465 33088 343431
rect 35806 341864 35862 341873
rect 35806 341799 35862 341808
rect 33046 341456 33102 341465
rect 33046 341391 33102 341400
rect 35820 341358 35848 341799
rect 39868 341358 39896 343839
rect 40224 343800 40276 343806
rect 40224 343742 40276 343748
rect 40040 343664 40092 343670
rect 40040 343606 40092 343612
rect 40052 343505 40080 343606
rect 40038 343496 40094 343505
rect 40038 343431 40094 343440
rect 40236 342281 40264 343742
rect 45006 343496 45062 343505
rect 45006 343431 45062 343440
rect 40222 342272 40278 342281
rect 40222 342207 40278 342216
rect 45020 341873 45048 343431
rect 45204 342553 45232 344986
rect 45296 342666 45324 383551
rect 45466 382664 45522 382673
rect 45466 382599 45522 382608
rect 45480 343233 45508 382599
rect 46018 355872 46074 355881
rect 46018 355807 46074 355816
rect 45834 355600 45890 355609
rect 45834 355535 45890 355544
rect 45652 353864 45704 353870
rect 45650 353832 45652 353841
rect 45704 353832 45706 353841
rect 45650 353767 45706 353776
rect 45848 353734 45876 355535
rect 45836 353728 45888 353734
rect 45836 353670 45888 353676
rect 45652 353456 45704 353462
rect 45652 353398 45704 353404
rect 45664 352209 45692 353398
rect 46032 353258 46060 355807
rect 46020 353252 46072 353258
rect 46020 353194 46072 353200
rect 45650 352200 45706 352209
rect 45650 352135 45706 352144
rect 45466 343224 45522 343233
rect 45466 343159 45522 343168
rect 45558 342816 45614 342825
rect 45558 342751 45614 342760
rect 45296 342638 45416 342666
rect 45190 342544 45246 342553
rect 45190 342479 45246 342488
rect 44822 341864 44878 341873
rect 44822 341799 44878 341808
rect 45006 341864 45062 341873
rect 45006 341799 45062 341808
rect 35808 341352 35860 341358
rect 35808 341294 35860 341300
rect 39856 341352 39908 341358
rect 39856 341294 39908 341300
rect 35808 341216 35860 341222
rect 35808 341158 35860 341164
rect 40224 341216 40276 341222
rect 40224 341158 40276 341164
rect 35532 341080 35584 341086
rect 35530 341048 35532 341057
rect 35820 341057 35848 341158
rect 40040 341080 40092 341086
rect 35584 341048 35586 341057
rect 35530 340983 35586 340992
rect 35806 341048 35862 341057
rect 40040 341022 40092 341028
rect 35806 340983 35862 340992
rect 40052 340649 40080 341022
rect 40038 340640 40094 340649
rect 40038 340575 40094 340584
rect 40236 340241 40264 341158
rect 44836 341057 44864 341799
rect 44822 341048 44878 341057
rect 44822 340983 44878 340992
rect 45388 340649 45416 342638
rect 45374 340640 45430 340649
rect 45374 340575 45430 340584
rect 39854 340232 39910 340241
rect 39854 340167 39910 340176
rect 40222 340232 40278 340241
rect 40222 340167 40278 340176
rect 39868 339833 39896 340167
rect 35530 339824 35586 339833
rect 35530 339759 35586 339768
rect 35806 339824 35862 339833
rect 35806 339759 35862 339768
rect 39854 339824 39910 339833
rect 39854 339759 39910 339768
rect 35544 339522 35572 339759
rect 35820 339658 35848 339759
rect 35808 339652 35860 339658
rect 35808 339594 35860 339600
rect 37924 339652 37976 339658
rect 37924 339594 37976 339600
rect 35532 339516 35584 339522
rect 35532 339458 35584 339464
rect 35162 338600 35218 338609
rect 35162 338535 35218 338544
rect 35176 331809 35204 338535
rect 35806 335744 35862 335753
rect 35806 335679 35862 335688
rect 35820 335374 35848 335679
rect 35808 335368 35860 335374
rect 35808 335310 35860 335316
rect 35806 334928 35862 334937
rect 35806 334863 35862 334872
rect 35820 334150 35848 334863
rect 35808 334144 35860 334150
rect 35808 334086 35860 334092
rect 37936 332897 37964 339594
rect 38936 339516 38988 339522
rect 38936 339458 38988 339464
rect 38948 335753 38976 339458
rect 45374 338056 45430 338065
rect 45374 337991 45430 338000
rect 45388 337906 45416 337991
rect 45388 337878 45508 337906
rect 38934 335744 38990 335753
rect 38934 335679 38990 335688
rect 40224 335368 40276 335374
rect 40224 335310 40276 335316
rect 39764 334144 39816 334150
rect 40236 334121 40264 335310
rect 42062 334656 42118 334665
rect 42062 334591 42118 334600
rect 43810 334656 43866 334665
rect 43810 334591 43866 334600
rect 45098 334656 45154 334665
rect 45098 334591 45154 334600
rect 39764 334086 39816 334092
rect 40222 334112 40278 334121
rect 37922 332888 37978 332897
rect 37922 332823 37978 332832
rect 39776 332489 39804 334086
rect 40222 334047 40278 334056
rect 39762 332480 39818 332489
rect 39762 332415 39818 332424
rect 35162 331800 35218 331809
rect 35162 331735 35218 331744
rect 42076 327729 42104 334591
rect 42982 334112 43038 334121
rect 42982 334047 43038 334056
rect 42798 332480 42854 332489
rect 42798 332415 42854 332424
rect 42062 327720 42118 327729
rect 42062 327655 42118 327664
rect 42430 327040 42486 327049
rect 42430 326975 42486 326984
rect 42444 326278 42472 326975
rect 42168 326210 42196 326264
rect 42260 326250 42472 326278
rect 42260 326210 42288 326250
rect 42168 326182 42288 326210
rect 41786 324864 41842 324873
rect 41786 324799 41842 324808
rect 41800 324428 41828 324799
rect 42182 323734 42472 323762
rect 41786 322824 41842 322833
rect 41786 322759 41842 322768
rect 41800 322592 41828 322759
rect 42182 321898 42288 321926
rect 42062 321600 42118 321609
rect 42062 321535 42118 321544
rect 42076 321368 42104 321535
rect 42062 321192 42118 321201
rect 42062 321127 42118 321136
rect 42076 320725 42104 321127
rect 42260 320278 42288 321898
rect 42444 320793 42472 323734
rect 42430 320784 42486 320793
rect 42430 320719 42486 320728
rect 42248 320272 42300 320278
rect 42248 320214 42300 320220
rect 42812 320090 42840 332415
rect 42996 321201 43024 334047
rect 42982 321192 43038 321201
rect 42982 321127 43038 321136
rect 42182 320062 42840 320090
rect 42616 320000 42668 320006
rect 42616 319942 42668 319948
rect 42182 319518 42472 319546
rect 42444 319025 42472 319518
rect 42628 319433 42656 319942
rect 42614 319424 42670 319433
rect 42614 319359 42670 319368
rect 42430 319016 42486 319025
rect 42430 318951 42486 318960
rect 42246 317520 42302 317529
rect 42246 317455 42302 317464
rect 42062 317248 42118 317257
rect 42062 317183 42118 317192
rect 42076 317045 42104 317183
rect 42260 316418 42288 317455
rect 42182 316390 42288 316418
rect 41786 316024 41842 316033
rect 41786 315959 41842 315968
rect 41800 315757 41828 315959
rect 41786 315616 41842 315625
rect 41786 315551 41842 315560
rect 41800 315180 41828 315551
rect 42154 313712 42210 313721
rect 42154 313647 42210 313656
rect 42168 313344 42196 313647
rect 42430 313168 42486 313177
rect 42430 313103 42486 313112
rect 42444 312746 42472 313103
rect 42182 312718 42472 312746
rect 42246 312488 42302 312497
rect 42246 312423 42302 312432
rect 42076 311953 42104 312052
rect 42062 311944 42118 311953
rect 42062 311879 42118 311888
rect 42260 311658 42288 312423
rect 42168 311630 42288 311658
rect 42168 311508 42196 311630
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41142 300928 41198 300937
rect 41142 300863 41198 300872
rect 41156 299130 41184 300863
rect 41144 299124 41196 299130
rect 41144 299066 41196 299072
rect 41696 299124 41748 299130
rect 41696 299066 41748 299072
rect 41708 298738 41736 299066
rect 42798 299024 42854 299033
rect 42798 298959 42854 298968
rect 41970 298752 42026 298761
rect 41708 298710 41970 298738
rect 41970 298687 42026 298696
rect 41326 296440 41382 296449
rect 41326 296375 41382 296384
rect 39302 296032 39358 296041
rect 39302 295967 39358 295976
rect 33046 294808 33102 294817
rect 33046 294743 33102 294752
rect 33060 287706 33088 294743
rect 33782 294400 33838 294409
rect 33782 294335 33838 294344
rect 33048 287700 33100 287706
rect 33048 287642 33100 287648
rect 33796 284889 33824 294335
rect 35806 291952 35862 291961
rect 35806 291887 35862 291896
rect 35820 291378 35848 291887
rect 35808 291372 35860 291378
rect 35808 291314 35860 291320
rect 35162 290320 35218 290329
rect 35162 290255 35218 290264
rect 35176 286346 35204 290255
rect 35164 286340 35216 286346
rect 35164 286282 35216 286288
rect 33782 284880 33838 284889
rect 33782 284815 33838 284824
rect 39316 284345 39344 295967
rect 41340 294642 41368 296375
rect 42338 295216 42394 295225
rect 42338 295151 42394 295160
rect 41328 294636 41380 294642
rect 41328 294578 41380 294584
rect 41696 294636 41748 294642
rect 41696 294578 41748 294584
rect 41708 294522 41736 294578
rect 41708 294506 42104 294522
rect 41708 294500 42116 294506
rect 41708 294494 42064 294500
rect 42064 294442 42116 294448
rect 41786 293992 41842 294001
rect 41616 293950 41786 293978
rect 41616 292602 41644 293950
rect 41786 293927 41842 293936
rect 40592 292597 40644 292602
rect 40590 292596 40646 292597
rect 40590 292588 40592 292596
rect 40644 292588 40646 292596
rect 41604 292596 41656 292602
rect 41604 292538 41656 292544
rect 40590 292523 40646 292532
rect 41604 291372 41656 291378
rect 41604 291314 41656 291320
rect 41616 290442 41644 291314
rect 41786 290456 41842 290465
rect 41616 290414 41786 290442
rect 41786 290391 41842 290400
rect 42352 289814 42380 295151
rect 42524 294500 42576 294506
rect 42524 294442 42576 294448
rect 42536 292574 42564 294442
rect 42260 289786 42380 289814
rect 42444 292546 42564 292574
rect 42444 289814 42472 292546
rect 42444 289786 42564 289814
rect 41512 287700 41564 287706
rect 41512 287642 41564 287648
rect 41524 285410 41552 287642
rect 42260 286346 42288 289786
rect 42536 286498 42564 289786
rect 42444 286470 42564 286498
rect 41696 286340 41748 286346
rect 41696 286282 41748 286288
rect 42248 286340 42300 286346
rect 42248 286282 42300 286288
rect 41708 286226 41736 286282
rect 41708 286198 42380 286226
rect 41524 285382 42288 285410
rect 39302 284336 39358 284345
rect 39302 284271 39358 284280
rect 42260 283059 42288 285382
rect 42182 283031 42288 283059
rect 42352 281874 42380 286198
rect 42182 281846 42380 281874
rect 42168 281302 42288 281330
rect 42168 281180 42196 281302
rect 42260 281194 42288 281302
rect 42444 281194 42472 286470
rect 42616 286340 42668 286346
rect 42616 286282 42668 286288
rect 42260 281166 42472 281194
rect 42182 280554 42472 280582
rect 42154 279848 42210 279857
rect 42154 279783 42210 279792
rect 42168 279344 42196 279783
rect 42444 279449 42472 280554
rect 42430 279440 42486 279449
rect 42430 279375 42486 279384
rect 42182 278718 42472 278746
rect 41970 278488 42026 278497
rect 41970 278423 42026 278432
rect 41984 278188 42012 278423
rect 42076 277273 42104 277508
rect 42248 277364 42300 277370
rect 42248 277306 42300 277312
rect 42062 277264 42118 277273
rect 42062 277199 42118 277208
rect 42260 276910 42288 277306
rect 42182 276882 42288 276910
rect 42248 276820 42300 276826
rect 42248 276762 42300 276768
rect 42260 276570 42288 276762
rect 42444 276706 42472 278718
rect 42628 276826 42656 286282
rect 42616 276820 42668 276826
rect 42616 276762 42668 276768
rect 42444 276678 42564 276706
rect 42076 276542 42288 276570
rect 42076 276352 42104 276542
rect 42536 275913 42564 276678
rect 42522 275904 42578 275913
rect 42522 275839 42578 275848
rect 41786 274272 41842 274281
rect 41786 274207 41842 274216
rect 41800 273836 41828 274207
rect 42168 273170 42196 273224
rect 42260 273222 42472 273238
rect 42260 273216 42484 273222
rect 42260 273210 42432 273216
rect 42260 273170 42288 273210
rect 42168 273142 42288 273170
rect 42432 273158 42484 273164
rect 41786 273048 41842 273057
rect 41786 272983 41842 272992
rect 41800 272544 41828 272983
rect 41786 272232 41842 272241
rect 41786 272167 41842 272176
rect 41800 272000 41828 272167
rect 42182 270150 42472 270178
rect 41786 270056 41842 270065
rect 41786 269991 41842 270000
rect 41800 269521 41828 269991
rect 41970 269104 42026 269113
rect 41970 269039 42026 269048
rect 41984 268872 42012 269039
rect 42168 266257 42196 268328
rect 42444 267753 42472 270150
rect 42430 267744 42486 267753
rect 42430 267679 42486 267688
rect 42154 266248 42210 266257
rect 42154 266183 42210 266192
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 35806 257136 35862 257145
rect 35806 257071 35862 257080
rect 39578 257136 39634 257145
rect 39578 257071 39634 257080
rect 35820 256834 35848 257071
rect 39592 256834 39620 257071
rect 35808 256828 35860 256834
rect 35808 256770 35860 256776
rect 39580 256828 39632 256834
rect 39580 256770 39632 256776
rect 35622 255912 35678 255921
rect 35622 255847 35678 255856
rect 39946 255912 40002 255921
rect 39946 255847 40002 255856
rect 35636 255338 35664 255847
rect 35806 255504 35862 255513
rect 35806 255439 35808 255448
rect 35860 255439 35862 255448
rect 35808 255410 35860 255416
rect 35624 255332 35676 255338
rect 35624 255274 35676 255280
rect 35806 254688 35862 254697
rect 35806 254623 35862 254632
rect 35820 254386 35848 254623
rect 35808 254380 35860 254386
rect 35808 254322 35860 254328
rect 35622 254280 35678 254289
rect 35622 254215 35678 254224
rect 35636 253978 35664 254215
rect 35808 254108 35860 254114
rect 35808 254050 35860 254056
rect 35624 253972 35676 253978
rect 35624 253914 35676 253920
rect 35820 253881 35848 254050
rect 39960 253978 39988 255847
rect 40500 255468 40552 255474
rect 40500 255410 40552 255416
rect 40512 254697 40540 255410
rect 41708 255338 42104 255354
rect 42812 255338 42840 298959
rect 43166 297256 43222 297265
rect 43166 297191 43222 297200
rect 42982 293584 43038 293593
rect 42982 293519 43038 293528
rect 42996 273222 43024 293519
rect 42984 273216 43036 273222
rect 42984 273158 43036 273164
rect 43180 263594 43208 297191
rect 43350 290456 43406 290465
rect 43350 290391 43406 290400
rect 43364 277370 43392 290391
rect 43824 278361 43852 334591
rect 43994 334520 44050 334529
rect 43994 334455 44050 334464
rect 44008 278769 44036 334455
rect 44362 334384 44418 334393
rect 44362 334319 44418 334328
rect 44178 334248 44234 334257
rect 44178 334183 44234 334192
rect 44192 321609 44220 334183
rect 44178 321600 44234 321609
rect 44178 321535 44234 321544
rect 44376 317257 44404 334319
rect 44362 317248 44418 317257
rect 44362 317183 44418 317192
rect 44270 311264 44326 311273
rect 44270 311199 44326 311208
rect 44284 306374 44312 311199
rect 44284 306346 44496 306374
rect 44270 298072 44326 298081
rect 44270 298007 44326 298016
rect 43994 278760 44050 278769
rect 43994 278695 44050 278704
rect 43810 278352 43866 278361
rect 43810 278287 43866 278296
rect 43352 277364 43404 277370
rect 43352 277306 43404 277312
rect 43350 273864 43406 273873
rect 43350 273799 43406 273808
rect 43364 270494 43392 273799
rect 43364 270466 43484 270494
rect 43088 263566 43208 263594
rect 43088 255921 43116 263566
rect 43258 263256 43314 263265
rect 43258 263191 43314 263200
rect 43272 257145 43300 263191
rect 43258 257136 43314 257145
rect 43258 257071 43314 257080
rect 43074 255912 43130 255921
rect 43074 255847 43130 255856
rect 41696 255332 42116 255338
rect 41748 255326 42064 255332
rect 41696 255274 41748 255280
rect 42064 255274 42116 255280
rect 42800 255332 42852 255338
rect 42800 255274 42852 255280
rect 40498 254688 40554 254697
rect 40498 254623 40554 254632
rect 40684 254380 40736 254386
rect 40684 254322 40736 254328
rect 39948 253972 40000 253978
rect 39948 253914 40000 253920
rect 35806 253872 35862 253881
rect 35806 253807 35862 253816
rect 35622 253464 35678 253473
rect 35622 253399 35678 253408
rect 35636 252618 35664 253399
rect 40696 253065 40724 254322
rect 41512 254108 41564 254114
rect 41512 254050 41564 254056
rect 41524 253881 41552 254050
rect 41510 253872 41566 253881
rect 41510 253807 41566 253816
rect 35806 253056 35862 253065
rect 35806 252991 35862 253000
rect 40682 253056 40738 253065
rect 40682 252991 40738 253000
rect 42890 253056 42946 253065
rect 42890 252991 42946 253000
rect 35820 252754 35848 252991
rect 35808 252748 35860 252754
rect 35808 252690 35860 252696
rect 41328 252748 41380 252754
rect 41328 252690 41380 252696
rect 35624 252612 35676 252618
rect 35624 252554 35676 252560
rect 35806 252240 35862 252249
rect 35806 252175 35862 252184
rect 35820 251258 35848 252175
rect 35808 251252 35860 251258
rect 35808 251194 35860 251200
rect 37924 251252 37976 251258
rect 37924 251194 37976 251200
rect 35806 250608 35862 250617
rect 35806 250543 35862 250552
rect 35820 249966 35848 250543
rect 35808 249960 35860 249966
rect 35808 249902 35860 249908
rect 37936 242894 37964 251194
rect 40316 249960 40368 249966
rect 40316 249902 40368 249908
rect 40328 245721 40356 249902
rect 41340 248414 41368 252690
rect 41708 252618 42104 252634
rect 41696 252612 42116 252618
rect 41748 252606 42064 252612
rect 41696 252554 41748 252560
rect 42064 252554 42116 252560
rect 42708 252612 42760 252618
rect 42708 252554 42760 252560
rect 41340 248386 41552 248414
rect 40314 245712 40370 245721
rect 40314 245647 40370 245656
rect 37924 242888 37976 242894
rect 37924 242830 37976 242836
rect 41524 242706 41552 248386
rect 41696 242888 41748 242894
rect 41748 242836 42564 242842
rect 41696 242830 42564 242836
rect 41708 242814 42564 242830
rect 41524 242678 42472 242706
rect 42246 240136 42302 240145
rect 42246 240071 42302 240080
rect 42260 239850 42288 240071
rect 42182 239822 42288 239850
rect 42182 238635 42288 238663
rect 42260 238513 42288 238635
rect 42246 238504 42302 238513
rect 42246 238439 42302 238448
rect 42444 238014 42472 242678
rect 42182 237986 42472 238014
rect 41786 236600 41842 236609
rect 41786 236535 41842 236544
rect 41800 236164 41828 236535
rect 42338 235920 42394 235929
rect 42338 235855 42394 235864
rect 42352 234983 42380 235855
rect 42182 234955 42380 234983
rect 41786 234696 41842 234705
rect 41786 234631 41842 234640
rect 41800 234328 41828 234631
rect 42182 233667 42380 233695
rect 42352 233306 42380 233667
rect 42340 233300 42392 233306
rect 42340 233242 42392 233248
rect 42168 233158 42380 233186
rect 42168 233104 42196 233158
rect 42352 231985 42380 233158
rect 42338 231976 42394 231985
rect 42338 231911 42394 231920
rect 42338 231296 42394 231305
rect 42338 231231 42394 231240
rect 42352 230670 42380 231231
rect 42182 230642 42380 230670
rect 42340 230444 42392 230450
rect 42340 230386 42392 230392
rect 42154 230344 42210 230353
rect 42154 230279 42210 230288
rect 42168 229976 42196 230279
rect 42352 229378 42380 230386
rect 42182 229350 42380 229378
rect 42536 228834 42564 242814
rect 42720 237425 42748 252554
rect 42706 237416 42762 237425
rect 42706 237351 42762 237360
rect 42708 233300 42760 233306
rect 42708 233242 42760 233248
rect 42720 232257 42748 233242
rect 42706 232248 42762 232257
rect 42706 232183 42762 232192
rect 42182 228806 42564 228834
rect 41970 227352 42026 227361
rect 41970 227287 42026 227296
rect 41984 226984 42012 227287
rect 42154 226672 42210 226681
rect 42154 226607 42210 226616
rect 42168 226304 42196 226607
rect 42182 225678 42472 225706
rect 42168 223281 42196 225148
rect 42444 223553 42472 225678
rect 42430 223544 42486 223553
rect 42430 223479 42486 223488
rect 42154 223272 42210 223281
rect 42154 223207 42210 223216
rect 35806 217968 35862 217977
rect 35806 217903 35862 217912
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 35820 214713 35848 217903
rect 35806 214704 35862 214713
rect 35806 214639 35862 214648
rect 35806 214296 35862 214305
rect 35806 214231 35862 214240
rect 39762 214296 39818 214305
rect 39762 214231 39818 214240
rect 35820 214130 35848 214231
rect 39776 214130 39804 214231
rect 35808 214124 35860 214130
rect 35808 214066 35860 214072
rect 39764 214124 39816 214130
rect 39764 214066 39816 214072
rect 39854 213072 39910 213081
rect 39854 213007 39910 213016
rect 39868 212702 39896 213007
rect 35808 212696 35860 212702
rect 35806 212664 35808 212673
rect 39856 212696 39908 212702
rect 35860 212664 35862 212673
rect 39856 212638 39908 212644
rect 35806 212599 35862 212608
rect 42904 212265 42932 252991
rect 43074 245712 43130 245721
rect 43074 245647 43130 245656
rect 43088 230450 43116 245647
rect 43076 230444 43128 230450
rect 43076 230386 43128 230392
rect 43456 214305 43484 270466
rect 43626 269784 43682 269793
rect 43626 269719 43682 269728
rect 43640 263265 43668 269719
rect 43626 263256 43682 263265
rect 43626 263191 43682 263200
rect 44284 255241 44312 298007
rect 44468 297673 44496 306346
rect 44638 299704 44694 299713
rect 44638 299639 44694 299648
rect 44454 297664 44510 297673
rect 44454 297599 44510 297608
rect 44454 293176 44510 293185
rect 44454 293111 44510 293120
rect 44468 279857 44496 293111
rect 44454 279848 44510 279857
rect 44454 279783 44510 279792
rect 44652 263594 44680 299639
rect 44822 284336 44878 284345
rect 44822 284271 44878 284280
rect 44836 273254 44864 284271
rect 44560 263566 44680 263594
rect 44744 273226 44864 273254
rect 44560 256873 44588 263566
rect 44744 257689 44772 273226
rect 44730 257680 44786 257689
rect 44730 257615 44786 257624
rect 44546 256864 44602 256873
rect 44546 256799 44602 256808
rect 44914 256456 44970 256465
rect 44914 256391 44970 256400
rect 44270 255232 44326 255241
rect 44270 255167 44326 255176
rect 43810 254688 43866 254697
rect 43810 254623 43866 254632
rect 43626 253872 43682 253881
rect 43626 253807 43682 253816
rect 43640 222194 43668 253807
rect 43824 229094 43852 254623
rect 44928 253934 44956 256391
rect 44928 253906 45048 253934
rect 44454 251560 44510 251569
rect 44454 251495 44510 251504
rect 44178 250336 44234 250345
rect 44178 250271 44234 250280
rect 44192 230353 44220 250271
rect 44468 240145 44496 251495
rect 44638 251152 44694 251161
rect 44638 251087 44694 251096
rect 44454 240136 44510 240145
rect 44454 240071 44510 240080
rect 44178 230344 44234 230353
rect 44178 230279 44234 230288
rect 43548 222166 43668 222194
rect 43732 229066 43852 229094
rect 43732 222194 43760 229066
rect 44652 226681 44680 251087
rect 44638 226672 44694 226681
rect 44638 226607 44694 226616
rect 43732 222166 43852 222194
rect 43548 217410 43576 222166
rect 43548 217382 43668 217410
rect 43442 214296 43498 214305
rect 43442 214231 43498 214240
rect 40774 212256 40830 212265
rect 40774 212191 40830 212200
rect 42890 212256 42946 212265
rect 42890 212191 42946 212200
rect 35622 211848 35678 211857
rect 35622 211783 35678 211792
rect 40130 211848 40186 211857
rect 40130 211783 40186 211792
rect 35636 211206 35664 211783
rect 40144 211478 40172 211783
rect 35808 211472 35860 211478
rect 35806 211440 35808 211449
rect 40132 211472 40184 211478
rect 35860 211440 35862 211449
rect 40132 211414 40184 211420
rect 35806 211375 35862 211384
rect 40788 211206 40816 212191
rect 43640 211857 43668 217382
rect 43824 213081 43852 222166
rect 45020 215294 45048 253906
rect 44928 215266 45048 215294
rect 44928 213761 44956 215266
rect 44914 213752 44970 213761
rect 44914 213687 44970 213696
rect 43810 213072 43866 213081
rect 43810 213007 43866 213016
rect 43626 211848 43682 211857
rect 43626 211783 43682 211792
rect 35624 211200 35676 211206
rect 35624 211142 35676 211148
rect 40776 211200 40828 211206
rect 40776 211142 40828 211148
rect 35806 210216 35862 210225
rect 35806 210151 35862 210160
rect 35820 209846 35848 210151
rect 35808 209840 35860 209846
rect 35808 209782 35860 209788
rect 39212 209840 39264 209846
rect 39212 209782 39264 209788
rect 35622 209400 35678 209409
rect 35622 209335 35678 209344
rect 35636 208418 35664 209335
rect 35808 208684 35860 208690
rect 35808 208626 35860 208632
rect 35624 208412 35676 208418
rect 35624 208354 35676 208360
rect 35820 208185 35848 208626
rect 35806 208176 35862 208185
rect 35806 208111 35862 208120
rect 35806 207360 35862 207369
rect 35806 207295 35862 207304
rect 35820 207194 35848 207295
rect 35808 207188 35860 207194
rect 35808 207130 35860 207136
rect 39224 206961 39252 209782
rect 39948 208684 40000 208690
rect 39948 208626 40000 208632
rect 39210 206952 39266 206961
rect 39210 206887 39266 206896
rect 35806 206136 35862 206145
rect 35806 206071 35862 206080
rect 35820 205834 35848 206071
rect 35808 205828 35860 205834
rect 35808 205770 35860 205776
rect 39960 205329 39988 208626
rect 44454 208584 44510 208593
rect 44454 208519 44510 208528
rect 40960 208412 41012 208418
rect 40960 208354 41012 208360
rect 40972 207777 41000 208354
rect 44178 208040 44234 208049
rect 44178 207975 44234 207984
rect 40958 207768 41014 207777
rect 40958 207703 41014 207712
rect 43258 207768 43314 207777
rect 43258 207703 43314 207712
rect 40958 207360 41014 207369
rect 40958 207295 41014 207304
rect 43074 207360 43130 207369
rect 43074 207295 43130 207304
rect 40972 207194 41000 207295
rect 40960 207188 41012 207194
rect 40960 207130 41012 207136
rect 42890 206952 42946 206961
rect 42890 206887 42946 206896
rect 41696 205828 41748 205834
rect 41696 205770 41748 205776
rect 41708 205714 41736 205770
rect 41708 205686 42104 205714
rect 42076 205562 42104 205686
rect 42064 205556 42116 205562
rect 42064 205498 42116 205504
rect 39946 205320 40002 205329
rect 39946 205255 40002 205264
rect 35806 204912 35862 204921
rect 35806 204847 35862 204856
rect 41510 204912 41566 204921
rect 41510 204847 41566 204856
rect 35820 204678 35848 204847
rect 35808 204672 35860 204678
rect 35808 204614 35860 204620
rect 41524 204513 41552 204847
rect 41696 204536 41748 204542
rect 35806 204504 35862 204513
rect 35806 204439 35862 204448
rect 41510 204504 41566 204513
rect 41510 204439 41566 204448
rect 41694 204504 41696 204513
rect 41748 204504 41750 204513
rect 41694 204439 41750 204448
rect 35820 204338 35848 204439
rect 35808 204332 35860 204338
rect 35808 204274 35860 204280
rect 39396 204332 39448 204338
rect 39396 204274 39448 204280
rect 39408 204105 39436 204274
rect 39394 204096 39450 204105
rect 39394 204031 39450 204040
rect 42706 204096 42762 204105
rect 42706 204031 42762 204040
rect 35806 203688 35862 203697
rect 35806 203623 35862 203632
rect 35820 202910 35848 203623
rect 35808 202904 35860 202910
rect 35808 202846 35860 202852
rect 39304 202904 39356 202910
rect 39304 202846 39356 202852
rect 42720 202874 42748 204031
rect 42720 202846 42840 202874
rect 39316 197849 39344 202846
rect 42430 201376 42486 201385
rect 42430 201311 42486 201320
rect 39302 197840 39358 197849
rect 39302 197775 39358 197784
rect 42444 196670 42472 201311
rect 42812 197146 42840 202846
rect 42720 197130 42840 197146
rect 42708 197124 42840 197130
rect 42760 197118 42840 197124
rect 42708 197066 42760 197072
rect 42182 196642 42472 196670
rect 41878 195800 41934 195809
rect 41878 195735 41934 195744
rect 41892 195432 41920 195735
rect 42338 195528 42394 195537
rect 42338 195463 42394 195472
rect 41786 195256 41842 195265
rect 41786 195191 41842 195200
rect 41800 194820 41828 195191
rect 41786 193488 41842 193497
rect 41786 193423 41842 193432
rect 41800 192984 41828 193423
rect 42352 193225 42380 195463
rect 42338 193216 42394 193225
rect 42338 193151 42394 193160
rect 42246 192808 42302 192817
rect 42246 192743 42302 192752
rect 42076 191593 42104 191760
rect 42062 191584 42118 191593
rect 42062 191519 42118 191528
rect 42168 191026 42196 191148
rect 42260 191026 42288 192743
rect 42168 190998 42288 191026
rect 42430 190496 42486 190505
rect 42182 190454 42430 190482
rect 42430 190431 42486 190440
rect 42430 189952 42486 189961
rect 42182 189910 42430 189938
rect 42430 189887 42486 189896
rect 42430 187640 42486 187649
rect 42430 187575 42486 187584
rect 42444 187459 42472 187575
rect 42182 187431 42472 187459
rect 42432 187332 42484 187338
rect 42432 187274 42484 187280
rect 42444 186810 42472 187274
rect 42182 186782 42472 186810
rect 42338 186280 42394 186289
rect 42338 186215 42394 186224
rect 42168 186017 42196 186184
rect 42154 186008 42210 186017
rect 42154 185943 42210 185952
rect 42352 185619 42380 186215
rect 42182 185591 42380 185619
rect 42904 183779 42932 206887
rect 43088 187338 43116 207295
rect 43272 205714 43300 207703
rect 43180 205686 43300 205714
rect 43180 195974 43208 205686
rect 43352 205556 43404 205562
rect 43352 205498 43404 205504
rect 43364 205442 43392 205498
rect 43272 205414 43392 205442
rect 43272 198098 43300 205414
rect 43442 205320 43498 205329
rect 43442 205255 43498 205264
rect 43456 201385 43484 205255
rect 43810 204504 43866 204513
rect 43810 204439 43866 204448
rect 43442 201376 43498 201385
rect 43442 201311 43498 201320
rect 43272 198070 43576 198098
rect 43352 197124 43404 197130
rect 43352 197066 43404 197072
rect 43364 195974 43392 197066
rect 43180 195946 43300 195974
rect 43364 195946 43484 195974
rect 43076 187332 43128 187338
rect 43076 187274 43128 187280
rect 42182 183751 42932 183779
rect 42430 183152 42486 183161
rect 42182 183110 42430 183138
rect 42430 183087 42486 183096
rect 42182 182463 42472 182491
rect 42444 182170 42472 182463
rect 43272 182170 43300 195946
rect 42432 182164 42484 182170
rect 42432 182106 42484 182112
rect 43260 182164 43312 182170
rect 43260 182106 43312 182112
rect 42076 179353 42104 181900
rect 42062 179344 42118 179353
rect 42062 179279 42118 179288
rect 43456 44198 43484 195946
rect 43548 193214 43576 198070
rect 43548 193186 43668 193214
rect 43640 187649 43668 193186
rect 43824 191593 43852 204439
rect 43810 191584 43866 191593
rect 43810 191519 43866 191528
rect 43626 187640 43682 187649
rect 43626 187575 43682 187584
rect 44192 183161 44220 207975
rect 44468 189961 44496 208519
rect 44638 205592 44694 205601
rect 44638 205527 44694 205536
rect 44652 190505 44680 205527
rect 44638 190496 44694 190505
rect 44638 190431 44694 190440
rect 44454 189952 44510 189961
rect 44454 189887 44510 189896
rect 44178 183152 44234 183161
rect 44178 183087 44234 183096
rect 45112 74534 45140 334591
rect 45282 327040 45338 327049
rect 45480 327026 45508 337878
rect 45338 326998 45508 327026
rect 45282 326975 45338 326984
rect 45572 300121 45600 342751
rect 45742 341048 45798 341057
rect 45742 340983 45798 340992
rect 45558 300112 45614 300121
rect 45558 300047 45614 300056
rect 45756 299305 45784 340983
rect 46018 340232 46074 340241
rect 46018 340167 46074 340176
rect 45742 299296 45798 299305
rect 45742 299231 45798 299240
rect 46032 298489 46060 340167
rect 46018 298480 46074 298489
rect 46018 298415 46074 298424
rect 45282 292768 45338 292777
rect 45282 292703 45338 292712
rect 45296 282914 45324 292703
rect 45466 291544 45522 291553
rect 45466 291479 45522 291488
rect 45480 291394 45508 291479
rect 45204 282886 45324 282914
rect 45388 291366 45508 291394
rect 45204 277250 45232 282886
rect 45388 279041 45416 291366
rect 45560 284368 45612 284374
rect 45558 284336 45560 284345
rect 45612 284336 45614 284345
rect 45558 284271 45614 284280
rect 45374 279032 45430 279041
rect 45374 278967 45430 278976
rect 45466 278760 45522 278769
rect 45466 278695 45522 278704
rect 45480 277438 45508 278695
rect 45468 277432 45520 277438
rect 45468 277374 45520 277380
rect 45374 277264 45430 277273
rect 45204 277222 45374 277250
rect 45374 277199 45430 277208
rect 46216 264246 46244 611662
rect 47768 451444 47820 451450
rect 47768 451386 47820 451392
rect 46938 380760 46994 380769
rect 46938 380695 46994 380704
rect 46952 356153 46980 380695
rect 47582 376136 47638 376145
rect 47582 376071 47638 376080
rect 46938 356144 46994 356153
rect 46938 356079 46994 356088
rect 46570 338464 46626 338473
rect 46570 338399 46626 338408
rect 46386 337648 46442 337657
rect 46386 337583 46442 337592
rect 46400 313177 46428 337583
rect 46584 319025 46612 338399
rect 46570 319016 46626 319025
rect 46570 318951 46626 318960
rect 46386 313168 46442 313177
rect 46386 313103 46442 313112
rect 46938 296848 46994 296857
rect 46938 296783 46994 296792
rect 46388 285728 46440 285734
rect 46388 285670 46440 285676
rect 46204 264240 46256 264246
rect 46204 264182 46256 264188
rect 46400 258097 46428 285670
rect 46952 267753 46980 296783
rect 47596 293962 47624 376071
rect 47584 293956 47636 293962
rect 47584 293898 47636 293904
rect 47582 290728 47638 290737
rect 47582 290663 47638 290672
rect 46938 267744 46994 267753
rect 46938 267679 46994 267688
rect 46386 258088 46442 258097
rect 46386 258023 46442 258032
rect 46938 252784 46994 252793
rect 46938 252719 46994 252728
rect 45558 249112 45614 249121
rect 45558 249047 45614 249056
rect 45572 231305 45600 249047
rect 45926 248704 45982 248713
rect 45926 248639 45982 248648
rect 45742 248296 45798 248305
rect 45742 248231 45798 248240
rect 45756 235929 45784 248231
rect 45742 235920 45798 235929
rect 45742 235855 45798 235864
rect 45940 232257 45968 248639
rect 46110 247072 46166 247081
rect 46110 247007 46166 247016
rect 46124 238513 46152 247007
rect 46110 238504 46166 238513
rect 46110 238439 46166 238448
rect 45926 232248 45982 232257
rect 45926 232183 45982 232192
rect 45558 231296 45614 231305
rect 45558 231231 45614 231240
rect 46952 223553 46980 252719
rect 47122 251968 47178 251977
rect 47122 251903 47178 251912
rect 47136 231985 47164 251903
rect 47122 231976 47178 231985
rect 47122 231911 47178 231920
rect 46938 223544 46994 223553
rect 46938 223479 46994 223488
rect 46202 204912 46258 204921
rect 46202 204847 46258 204856
rect 45112 74506 45508 74534
rect 45480 53106 45508 74506
rect 45468 53100 45520 53106
rect 45468 53042 45520 53048
rect 46216 49026 46244 204847
rect 47596 52018 47624 290663
rect 47780 284986 47808 451386
rect 47768 284980 47820 284986
rect 47768 284922 47820 284928
rect 47766 247480 47822 247489
rect 47766 247415 47822 247424
rect 47584 52012 47636 52018
rect 47584 51954 47636 51960
rect 47780 50386 47808 247415
rect 48976 53242 49004 761874
rect 50160 611312 50212 611318
rect 50160 611254 50212 611260
rect 50172 610162 50200 611254
rect 50160 610156 50212 610162
rect 50160 610098 50212 610104
rect 49146 291136 49202 291145
rect 49146 291071 49202 291080
rect 48964 53236 49016 53242
rect 48964 53178 49016 53184
rect 47768 50380 47820 50386
rect 47768 50322 47820 50328
rect 49160 49162 49188 291071
rect 50356 51882 50384 806074
rect 53104 799128 53156 799134
rect 53104 799070 53156 799076
rect 53116 790770 53144 799070
rect 53104 790764 53156 790770
rect 53104 790706 53156 790712
rect 58636 786554 58664 816954
rect 61384 815652 61436 815658
rect 61384 815594 61436 815600
rect 61396 788662 61424 815594
rect 62764 814904 62816 814910
rect 62764 814846 62816 814852
rect 62212 790764 62264 790770
rect 62212 790706 62264 790712
rect 62224 790537 62252 790706
rect 62210 790528 62266 790537
rect 62210 790463 62266 790472
rect 61384 788656 61436 788662
rect 61384 788598 61436 788604
rect 62118 787400 62174 787409
rect 62118 787335 62174 787344
rect 62132 786690 62160 787335
rect 62120 786684 62172 786690
rect 62120 786626 62172 786632
rect 58624 786548 58676 786554
rect 58624 786490 58676 786496
rect 62120 786548 62172 786554
rect 62120 786490 62172 786496
rect 62132 786185 62160 786490
rect 62118 786176 62174 786185
rect 62118 786111 62174 786120
rect 62776 784961 62804 814846
rect 64144 805996 64196 806002
rect 64144 805938 64196 805944
rect 62948 797700 63000 797706
rect 62948 797642 63000 797648
rect 62960 789177 62988 797642
rect 62946 789168 63002 789177
rect 62946 789103 63002 789112
rect 62948 788656 63000 788662
rect 62948 788598 63000 788604
rect 62960 787137 62988 788598
rect 62946 787128 63002 787137
rect 62946 787063 63002 787072
rect 62762 784952 62818 784961
rect 62762 784887 62818 784896
rect 58624 774240 58676 774246
rect 58624 774182 58676 774188
rect 57244 763224 57296 763230
rect 57244 763166 57296 763172
rect 51724 712292 51776 712298
rect 51724 712234 51776 712240
rect 51736 705158 51764 712234
rect 51724 705152 51776 705158
rect 51724 705094 51776 705100
rect 55864 676252 55916 676258
rect 55864 676194 55916 676200
rect 53104 669384 53156 669390
rect 53104 669326 53156 669332
rect 53116 660958 53144 669326
rect 53104 660952 53156 660958
rect 53104 660894 53156 660900
rect 53104 612604 53156 612610
rect 53104 612546 53156 612552
rect 51722 581224 51778 581233
rect 51722 581159 51778 581168
rect 51736 574054 51764 581159
rect 51724 574048 51776 574054
rect 51724 573990 51776 573996
rect 51722 539880 51778 539889
rect 51722 539815 51778 539824
rect 51736 531282 51764 539815
rect 51724 531276 51776 531282
rect 51724 531218 51776 531224
rect 50526 419928 50582 419937
rect 50526 419863 50582 419872
rect 50540 305658 50568 419863
rect 51078 407960 51134 407969
rect 51078 407895 51134 407904
rect 51092 404326 51120 407895
rect 51446 404968 51502 404977
rect 51446 404903 51502 404912
rect 51080 404320 51132 404326
rect 51080 404262 51132 404268
rect 51460 402966 51488 404903
rect 51448 402960 51500 402966
rect 51448 402902 51500 402908
rect 51080 400240 51132 400246
rect 51080 400182 51132 400188
rect 51092 397497 51120 400182
rect 51078 397488 51134 397497
rect 51078 397423 51134 397432
rect 51078 362264 51134 362273
rect 51078 362199 51134 362208
rect 51092 360194 51120 362199
rect 51080 360188 51132 360194
rect 51080 360130 51132 360136
rect 50528 305652 50580 305658
rect 50528 305594 50580 305600
rect 51722 301336 51778 301345
rect 51722 301271 51778 301280
rect 50528 293956 50580 293962
rect 50528 293898 50580 293904
rect 50540 278322 50568 293898
rect 51736 291174 51764 301271
rect 51724 291168 51776 291174
rect 51724 291110 51776 291116
rect 51724 288516 51776 288522
rect 51724 288458 51776 288464
rect 50528 278316 50580 278322
rect 50528 278258 50580 278264
rect 50526 247888 50582 247897
rect 50526 247823 50582 247832
rect 50344 51876 50396 51882
rect 50344 51818 50396 51824
rect 49148 49156 49200 49162
rect 49148 49098 49200 49104
rect 46204 49020 46256 49026
rect 46204 48962 46256 48968
rect 50540 44334 50568 247823
rect 51736 223553 51764 288458
rect 53116 264382 53144 612546
rect 54482 558512 54538 558521
rect 54482 558447 54538 558456
rect 54496 527134 54524 558447
rect 54484 527128 54536 527134
rect 54484 527070 54536 527076
rect 54482 430536 54538 430545
rect 54482 430471 54538 430480
rect 54496 398818 54524 430471
rect 54484 398812 54536 398818
rect 54484 398754 54536 398760
rect 54482 387560 54538 387569
rect 54482 387495 54538 387504
rect 54496 356726 54524 387495
rect 54484 356720 54536 356726
rect 54484 356662 54536 356668
rect 53838 320784 53894 320793
rect 53838 320719 53894 320728
rect 53852 317422 53880 320719
rect 53840 317416 53892 317422
rect 53840 317358 53892 317364
rect 53840 314764 53892 314770
rect 53840 314706 53892 314712
rect 53852 312497 53880 314706
rect 53838 312488 53894 312497
rect 53838 312423 53894 312432
rect 54482 300520 54538 300529
rect 54482 300455 54538 300464
rect 54496 292466 54524 300455
rect 54484 292460 54536 292466
rect 54484 292402 54536 292408
rect 54484 280424 54536 280430
rect 54484 280366 54536 280372
rect 53288 280220 53340 280226
rect 53288 280162 53340 280168
rect 53104 264376 53156 264382
rect 53104 264318 53156 264324
rect 51722 223544 51778 223553
rect 51722 223479 51778 223488
rect 51908 223032 51960 223038
rect 51908 222974 51960 222980
rect 51920 179353 51948 222974
rect 53300 215121 53328 280162
rect 54496 217977 54524 280366
rect 55876 277545 55904 676194
rect 56048 292596 56100 292602
rect 56048 292538 56100 292544
rect 55862 277536 55918 277545
rect 55862 277471 55918 277480
rect 56060 266257 56088 292538
rect 56046 266248 56102 266257
rect 56046 266183 56102 266192
rect 57256 231130 57284 763166
rect 58636 742422 58664 774182
rect 61384 772880 61436 772886
rect 61384 772822 61436 772828
rect 61396 747182 61424 772822
rect 62764 755540 62816 755546
rect 62764 755482 62816 755488
rect 62776 747697 62804 755482
rect 62762 747688 62818 747697
rect 62762 747623 62818 747632
rect 61384 747176 61436 747182
rect 61384 747118 61436 747124
rect 63040 747176 63092 747182
rect 63040 747118 63092 747124
rect 62120 746564 62172 746570
rect 62120 746506 62172 746512
rect 62132 746201 62160 746506
rect 62118 746192 62174 746201
rect 62118 746127 62174 746136
rect 62118 744152 62174 744161
rect 62118 744087 62174 744096
rect 62132 743918 62160 744087
rect 62120 743912 62172 743918
rect 62120 743854 62172 743860
rect 62120 743776 62172 743782
rect 62118 743744 62120 743753
rect 62172 743744 62174 743753
rect 62118 743679 62174 743688
rect 58624 742416 58676 742422
rect 62120 742416 62172 742422
rect 58624 742358 58676 742364
rect 62118 742384 62120 742393
rect 62172 742384 62174 742393
rect 62118 742319 62174 742328
rect 63052 741849 63080 747118
rect 63038 741840 63094 741849
rect 63038 741775 63094 741784
rect 58624 730380 58676 730386
rect 58624 730322 58676 730328
rect 58636 699582 58664 730322
rect 62764 729360 62816 729366
rect 62764 729302 62816 729308
rect 61384 719024 61436 719030
rect 61384 718966 61436 718972
rect 58624 699576 58676 699582
rect 58624 699518 58676 699524
rect 58624 667956 58676 667962
rect 58624 667898 58676 667904
rect 58636 659598 58664 667898
rect 58624 659592 58676 659598
rect 58624 659534 58676 659540
rect 58624 643136 58676 643142
rect 58624 643078 58676 643084
rect 58636 614038 58664 643078
rect 58624 614032 58676 614038
rect 58624 613974 58676 613980
rect 58624 610156 58676 610162
rect 58624 610098 58676 610104
rect 57428 294092 57480 294098
rect 57428 294034 57480 294040
rect 57440 275913 57468 294034
rect 57426 275904 57482 275913
rect 57426 275839 57482 275848
rect 58636 264518 58664 610098
rect 58808 305652 58860 305658
rect 58808 305594 58860 305600
rect 58820 278458 58848 305594
rect 60004 284980 60056 284986
rect 60004 284922 60056 284928
rect 58808 278452 58860 278458
rect 58808 278394 58860 278400
rect 60016 278186 60044 284922
rect 60004 278180 60056 278186
rect 60004 278122 60056 278128
rect 58624 264512 58676 264518
rect 58624 264454 58676 264460
rect 61396 264217 61424 718966
rect 62120 705152 62172 705158
rect 62120 705094 62172 705100
rect 62132 704449 62160 705094
rect 62118 704440 62174 704449
rect 62118 704375 62174 704384
rect 62120 703792 62172 703798
rect 62120 703734 62172 703740
rect 62132 703361 62160 703734
rect 62118 703352 62174 703361
rect 62118 703287 62174 703296
rect 62210 701312 62266 701321
rect 62210 701247 62266 701256
rect 62224 701078 62252 701247
rect 62212 701072 62264 701078
rect 62212 701014 62264 701020
rect 62776 700913 62804 729302
rect 62762 700904 62818 700913
rect 62762 700839 62818 700848
rect 62120 700324 62172 700330
rect 62120 700266 62172 700272
rect 62132 698193 62160 700266
rect 62304 699576 62356 699582
rect 62302 699544 62304 699553
rect 62356 699544 62358 699553
rect 62302 699479 62358 699488
rect 62118 698184 62174 698193
rect 62118 698119 62174 698128
rect 63408 686520 63460 686526
rect 63408 686462 63460 686468
rect 62120 660952 62172 660958
rect 62118 660920 62120 660929
rect 62172 660920 62174 660929
rect 62118 660855 62174 660864
rect 62120 659592 62172 659598
rect 62118 659560 62120 659569
rect 62172 659560 62174 659569
rect 62118 659495 62174 659504
rect 62304 658980 62356 658986
rect 62304 658922 62356 658928
rect 62118 658336 62174 658345
rect 62118 658271 62174 658280
rect 62132 657558 62160 658271
rect 62120 657552 62172 657558
rect 62120 657494 62172 657500
rect 62120 656872 62172 656878
rect 62120 656814 62172 656820
rect 62132 656577 62160 656814
rect 62118 656568 62174 656577
rect 62118 656503 62174 656512
rect 62316 655353 62344 658922
rect 63420 657665 63448 686462
rect 63406 657656 63462 657665
rect 63406 657591 63462 657600
rect 62302 655344 62358 655353
rect 62302 655279 62358 655288
rect 62948 642388 63000 642394
rect 62948 642330 63000 642336
rect 62120 616820 62172 616826
rect 62120 616762 62172 616768
rect 62132 616593 62160 616762
rect 62118 616584 62174 616593
rect 62118 616519 62174 616528
rect 62118 614680 62174 614689
rect 62118 614615 62174 614624
rect 62132 614174 62160 614615
rect 62120 614168 62172 614174
rect 62120 614110 62172 614116
rect 62120 614032 62172 614038
rect 62120 613974 62172 613980
rect 62132 613873 62160 613974
rect 62118 613864 62174 613873
rect 62118 613799 62174 613808
rect 62120 613420 62172 613426
rect 62120 613362 62172 613368
rect 62132 612649 62160 613362
rect 62118 612640 62174 612649
rect 62118 612575 62174 612584
rect 62960 612105 62988 642330
rect 63408 633480 63460 633486
rect 63408 633422 63460 633428
rect 63132 625864 63184 625870
rect 63132 625806 63184 625812
rect 63144 618089 63172 625806
rect 63130 618080 63186 618089
rect 63130 618015 63186 618024
rect 62946 612096 63002 612105
rect 62946 612031 63002 612040
rect 62762 595776 62818 595785
rect 62762 595711 62818 595720
rect 62578 590064 62634 590073
rect 62578 589999 62634 590008
rect 62120 575476 62172 575482
rect 62120 575418 62172 575424
rect 62132 574841 62160 575418
rect 62118 574832 62174 574841
rect 62118 574767 62174 574776
rect 62120 574048 62172 574054
rect 62120 573990 62172 573996
rect 62132 573617 62160 573990
rect 62118 573608 62174 573617
rect 62118 573543 62174 573552
rect 62592 569945 62620 589999
rect 62776 571169 62804 595711
rect 63130 594144 63186 594153
rect 63130 594079 63186 594088
rect 62946 590744 63002 590753
rect 62946 590679 63002 590688
rect 62762 571160 62818 571169
rect 62762 571095 62818 571104
rect 62578 569936 62634 569945
rect 62578 569871 62634 569880
rect 62210 556744 62266 556753
rect 62210 556679 62266 556688
rect 62224 538214 62252 556679
rect 62762 550216 62818 550225
rect 62762 550151 62818 550160
rect 62224 538186 62344 538214
rect 62118 531312 62174 531321
rect 62118 531247 62120 531256
rect 62172 531247 62174 531256
rect 62120 531218 62172 531224
rect 62120 531140 62172 531146
rect 62120 531082 62172 531088
rect 62132 530641 62160 531082
rect 62118 530632 62174 530641
rect 62118 530567 62174 530576
rect 62120 528624 62172 528630
rect 62118 528592 62120 528601
rect 62172 528592 62174 528601
rect 62118 528527 62174 528536
rect 62316 528057 62344 538186
rect 62302 528048 62358 528057
rect 62302 527983 62358 527992
rect 62120 527128 62172 527134
rect 62118 527096 62120 527105
rect 62172 527096 62174 527105
rect 62118 527031 62174 527040
rect 62776 525745 62804 550151
rect 62762 525736 62818 525745
rect 62762 525671 62818 525680
rect 62394 428496 62450 428505
rect 62394 428431 62450 428440
rect 62120 404320 62172 404326
rect 62120 404262 62172 404268
rect 62132 404161 62160 404262
rect 62118 404152 62174 404161
rect 62118 404087 62174 404096
rect 62120 402960 62172 402966
rect 62120 402902 62172 402908
rect 62132 402665 62160 402902
rect 62118 402656 62174 402665
rect 62118 402591 62174 402600
rect 62118 400616 62174 400625
rect 62118 400551 62174 400560
rect 62132 400246 62160 400551
rect 62120 400240 62172 400246
rect 62408 400217 62436 428431
rect 62120 400182 62172 400188
rect 62394 400208 62450 400217
rect 62394 400143 62450 400152
rect 62120 400104 62172 400110
rect 62120 400046 62172 400052
rect 62132 399401 62160 400046
rect 62118 399392 62174 399401
rect 62118 399327 62174 399336
rect 62120 398812 62172 398818
rect 62120 398754 62172 398760
rect 62132 398313 62160 398754
rect 62118 398304 62174 398313
rect 62118 398239 62174 398248
rect 62762 381576 62818 381585
rect 62762 381511 62818 381520
rect 62120 361548 62172 361554
rect 62120 361490 62172 361496
rect 62132 360913 62160 361490
rect 62118 360904 62174 360913
rect 62118 360839 62174 360848
rect 62120 360188 62172 360194
rect 62120 360130 62172 360136
rect 62132 359825 62160 360130
rect 62118 359816 62174 359825
rect 62118 359751 62174 359760
rect 62302 357504 62358 357513
rect 62302 357439 62358 357448
rect 62120 356720 62172 356726
rect 62316 356697 62344 357439
rect 62120 356662 62172 356668
rect 62302 356688 62358 356697
rect 62132 356017 62160 356662
rect 62302 356623 62358 356632
rect 62118 356008 62174 356017
rect 62118 355943 62174 355952
rect 62776 354521 62804 381511
rect 62762 354512 62818 354521
rect 62762 354447 62818 354456
rect 62670 341728 62726 341737
rect 62670 341663 62726 341672
rect 62302 341456 62358 341465
rect 62302 341391 62358 341400
rect 62316 330562 62344 341391
rect 62486 332616 62542 332625
rect 62486 332551 62542 332560
rect 62316 330534 62436 330562
rect 61566 319424 61622 319433
rect 61566 319359 61622 319368
rect 61580 316033 61608 319359
rect 62120 317416 62172 317422
rect 62118 317384 62120 317393
rect 62172 317384 62174 317393
rect 62118 317319 62174 317328
rect 61566 316024 61622 316033
rect 61566 315959 61622 315968
rect 62118 314800 62174 314809
rect 62118 314735 62120 314744
rect 62172 314735 62174 314744
rect 62120 314706 62172 314712
rect 62408 314129 62436 330534
rect 62500 325694 62528 332551
rect 62684 325694 62712 341663
rect 62500 325666 62620 325694
rect 62684 325666 62804 325694
rect 62394 314120 62450 314129
rect 62394 314055 62450 314064
rect 62302 295352 62358 295361
rect 62302 295287 62358 295296
rect 62118 294128 62174 294137
rect 62118 294063 62120 294072
rect 62172 294063 62174 294072
rect 62120 294034 62172 294040
rect 62118 292496 62174 292505
rect 62118 292431 62120 292440
rect 62172 292431 62174 292440
rect 62120 292402 62172 292408
rect 62120 291168 62172 291174
rect 62120 291110 62172 291116
rect 62132 291009 62160 291110
rect 62118 291000 62174 291009
rect 62118 290935 62174 290944
rect 62118 288552 62174 288561
rect 62118 288487 62120 288496
rect 62172 288487 62174 288496
rect 62120 288458 62172 288464
rect 62118 285968 62174 285977
rect 62118 285903 62174 285912
rect 62132 285734 62160 285903
rect 62120 285728 62172 285734
rect 62120 285670 62172 285676
rect 62316 281738 62344 295287
rect 62592 287054 62620 325666
rect 62776 311817 62804 325666
rect 62762 311808 62818 311817
rect 62762 311743 62818 311752
rect 62762 292768 62818 292777
rect 62762 292703 62818 292712
rect 62776 292602 62804 292703
rect 62764 292596 62816 292602
rect 62764 292538 62816 292544
rect 62762 287192 62818 287201
rect 62762 287127 62818 287136
rect 62592 287026 62712 287054
rect 62486 282160 62542 282169
rect 62486 282095 62542 282104
rect 62132 281710 62344 281738
rect 62132 280514 62160 281710
rect 62302 280936 62358 280945
rect 62302 280871 62358 280880
rect 61948 280486 62160 280514
rect 61948 279449 61976 280486
rect 62120 280424 62172 280430
rect 62118 280392 62120 280401
rect 62172 280392 62174 280401
rect 62118 280327 62174 280336
rect 62316 280226 62344 280871
rect 62304 280220 62356 280226
rect 62304 280162 62356 280168
rect 62500 280106 62528 282095
rect 62684 280332 62712 287026
rect 62316 280078 62528 280106
rect 62592 280304 62712 280332
rect 61934 279440 61990 279449
rect 61934 279375 61990 279384
rect 62316 273873 62344 280078
rect 62592 278730 62620 280304
rect 62580 278724 62632 278730
rect 62580 278666 62632 278672
rect 62776 277394 62804 287127
rect 62960 287054 62988 590679
rect 63144 568585 63172 594079
rect 63130 568576 63186 568585
rect 63130 568511 63186 568520
rect 63130 385928 63186 385937
rect 63130 385863 63186 385872
rect 63144 357241 63172 385863
rect 63130 357232 63186 357241
rect 63130 357167 63186 357176
rect 63222 342000 63278 342009
rect 63222 341935 63278 341944
rect 63236 313041 63264 341935
rect 63222 313032 63278 313041
rect 63222 312967 63278 312976
rect 63130 298752 63186 298761
rect 63130 298687 63186 298696
rect 63144 289785 63172 298687
rect 63130 289776 63186 289785
rect 63130 289711 63186 289720
rect 62960 287026 63356 287054
rect 62946 284608 63002 284617
rect 62946 284543 63002 284552
rect 62960 284374 62988 284543
rect 62948 284368 63000 284374
rect 62948 284310 63000 284316
rect 63130 283248 63186 283257
rect 63130 283183 63186 283192
rect 62946 280120 63002 280129
rect 62946 280055 63002 280064
rect 62960 277394 62988 280055
rect 62500 277366 62804 277394
rect 62868 277366 62988 277394
rect 62302 273864 62358 273873
rect 62302 273799 62358 273808
rect 62500 269793 62528 277366
rect 62486 269784 62542 269793
rect 62486 269719 62542 269728
rect 62868 265577 62896 277366
rect 62854 265568 62910 265577
rect 62854 265503 62910 265512
rect 61382 264208 61438 264217
rect 61382 264143 61438 264152
rect 57244 231124 57296 231130
rect 57244 231066 57296 231072
rect 61384 228540 61436 228546
rect 61384 228482 61436 228488
rect 57244 228404 57296 228410
rect 57244 228346 57296 228352
rect 56508 227044 56560 227050
rect 56508 226986 56560 226992
rect 56520 218210 56548 226986
rect 55680 218204 55732 218210
rect 55680 218146 55732 218152
rect 56508 218204 56560 218210
rect 56508 218146 56560 218152
rect 54482 217968 54538 217977
rect 54482 217903 54538 217912
rect 55692 217138 55720 218146
rect 57256 218074 57284 228346
rect 60648 227452 60700 227458
rect 60648 227394 60700 227400
rect 58992 226296 59044 226302
rect 58992 226238 59044 226244
rect 57428 218204 57480 218210
rect 57428 218146 57480 218152
rect 56508 218068 56560 218074
rect 56508 218010 56560 218016
rect 57244 218068 57296 218074
rect 57244 218010 57296 218016
rect 56520 217138 56548 218010
rect 57440 217274 57468 218146
rect 58164 218068 58216 218074
rect 58164 218010 58216 218016
rect 55646 217110 55720 217138
rect 56474 217110 56548 217138
rect 57302 217246 57468 217274
rect 55646 216988 55674 217110
rect 56474 216988 56502 217110
rect 57302 216988 57330 217246
rect 58176 217138 58204 218010
rect 59004 217274 59032 226238
rect 59360 221604 59412 221610
rect 59360 221546 59412 221552
rect 59372 218074 59400 221546
rect 59820 218748 59872 218754
rect 59820 218690 59872 218696
rect 59360 218068 59412 218074
rect 59360 218010 59412 218016
rect 58130 217110 58204 217138
rect 58958 217246 59032 217274
rect 58130 216988 58158 217110
rect 58958 216988 58986 217246
rect 59832 217138 59860 218690
rect 60660 217274 60688 227394
rect 61396 218210 61424 228482
rect 63144 223038 63172 283183
rect 63328 283098 63356 287026
rect 63236 283070 63356 283098
rect 63236 278610 63264 283070
rect 63420 278769 63448 633422
rect 63406 278760 63462 278769
rect 63406 278695 63462 278704
rect 63236 278594 63356 278610
rect 63236 278588 63368 278594
rect 63236 278582 63316 278588
rect 63316 278530 63368 278536
rect 63406 278080 63462 278089
rect 63406 278015 63462 278024
rect 63590 278080 63646 278089
rect 63590 278015 63646 278024
rect 63420 223553 63448 278015
rect 63604 277545 63632 278015
rect 63590 277536 63646 277545
rect 63590 277471 63646 277480
rect 64156 231169 64184 805938
rect 653404 790832 653456 790838
rect 653404 790774 653456 790780
rect 651470 778424 651526 778433
rect 651470 778359 651526 778368
rect 651484 777646 651512 778359
rect 651472 777640 651524 777646
rect 651472 777582 651524 777588
rect 652022 777064 652078 777073
rect 652022 776999 652078 777008
rect 651470 776112 651526 776121
rect 651470 776047 651526 776056
rect 651484 775606 651512 776047
rect 651472 775600 651524 775606
rect 651472 775542 651524 775548
rect 651380 775328 651432 775334
rect 651378 775296 651380 775305
rect 651432 775296 651434 775305
rect 651378 775231 651434 775240
rect 651470 774208 651526 774217
rect 651470 774143 651472 774152
rect 651524 774143 651526 774152
rect 651472 774114 651524 774120
rect 651472 773832 651524 773838
rect 651472 773774 651524 773780
rect 651484 773401 651512 773774
rect 651470 773392 651526 773401
rect 651470 773327 651526 773336
rect 652036 768942 652064 776999
rect 653416 775334 653444 790774
rect 670608 784304 670660 784310
rect 670608 784246 670660 784252
rect 669228 784168 669280 784174
rect 669228 784110 669280 784116
rect 669044 782536 669096 782542
rect 669044 782478 669096 782484
rect 655520 781108 655572 781114
rect 655520 781050 655572 781056
rect 655060 778388 655112 778394
rect 655060 778330 655112 778336
rect 653404 775328 653456 775334
rect 653404 775270 653456 775276
rect 655072 773838 655100 778330
rect 655532 774178 655560 781050
rect 660304 777640 660356 777646
rect 660304 777582 660356 777588
rect 655520 774172 655572 774178
rect 655520 774114 655572 774120
rect 655060 773832 655112 773838
rect 655060 773774 655112 773780
rect 652024 768936 652076 768942
rect 652024 768878 652076 768884
rect 656164 768936 656216 768942
rect 656164 768878 656216 768884
rect 653404 746632 653456 746638
rect 653404 746574 653456 746580
rect 651470 734224 651526 734233
rect 651470 734159 651526 734168
rect 651484 733446 651512 734159
rect 651472 733440 651524 733446
rect 651472 733382 651524 733388
rect 652666 732864 652722 732873
rect 652666 732799 652722 732808
rect 651470 731776 651526 731785
rect 651470 731711 651526 731720
rect 651484 731474 651512 731711
rect 651472 731468 651524 731474
rect 651472 731410 651524 731416
rect 651380 731128 651432 731134
rect 651378 731096 651380 731105
rect 651432 731096 651434 731105
rect 651378 731031 651434 731040
rect 652680 730726 652708 732799
rect 653416 731134 653444 746574
rect 654784 734188 654836 734194
rect 654784 734130 654836 734136
rect 653404 731128 653456 731134
rect 653404 731070 653456 731076
rect 652668 730720 652720 730726
rect 652668 730662 652720 730668
rect 651472 730040 651524 730046
rect 651472 729982 651524 729988
rect 651484 729881 651512 729982
rect 651470 729872 651526 729881
rect 651470 729807 651526 729816
rect 654796 728550 654824 734130
rect 651472 728544 651524 728550
rect 651470 728512 651472 728521
rect 654784 728544 654836 728550
rect 651524 728512 651526 728521
rect 654784 728486 654836 728492
rect 651470 728447 651526 728456
rect 656176 716310 656204 768878
rect 657544 735616 657596 735622
rect 657544 735558 657596 735564
rect 657556 730046 657584 735558
rect 658924 731468 658976 731474
rect 658924 731410 658976 731416
rect 657544 730040 657596 730046
rect 657544 729982 657596 729988
rect 656164 716304 656216 716310
rect 656164 716246 656216 716252
rect 654784 701208 654836 701214
rect 654784 701150 654836 701156
rect 651470 689480 651526 689489
rect 651470 689415 651526 689424
rect 651484 688702 651512 689415
rect 652760 688832 652812 688838
rect 651654 688800 651710 688809
rect 652760 688774 652812 688780
rect 651654 688735 651710 688744
rect 651472 688696 651524 688702
rect 651472 688638 651524 688644
rect 651470 687440 651526 687449
rect 651470 687375 651526 687384
rect 651484 687274 651512 687375
rect 651472 687268 651524 687274
rect 651472 687210 651524 687216
rect 651472 687064 651524 687070
rect 651472 687006 651524 687012
rect 651484 686769 651512 687006
rect 651470 686760 651526 686769
rect 651470 686695 651526 686704
rect 651668 686526 651696 688735
rect 651656 686520 651708 686526
rect 651656 686462 651708 686468
rect 651472 685568 651524 685574
rect 651472 685510 651524 685516
rect 651484 685273 651512 685510
rect 651470 685264 651526 685273
rect 651470 685199 651526 685208
rect 652574 684448 652630 684457
rect 652772 684434 652800 688774
rect 654796 687070 654824 701150
rect 656440 690124 656492 690130
rect 656440 690066 656492 690072
rect 654784 687064 654836 687070
rect 654784 687006 654836 687012
rect 656452 685574 656480 690066
rect 657544 688696 657596 688702
rect 657544 688638 657596 688644
rect 656440 685568 656492 685574
rect 656440 685510 656492 685516
rect 652630 684406 652800 684434
rect 652574 684383 652630 684392
rect 653404 655580 653456 655586
rect 653404 655522 653456 655528
rect 651470 643240 651526 643249
rect 651470 643175 651526 643184
rect 651484 642394 651512 643175
rect 651472 642388 651524 642394
rect 651472 642330 651524 642336
rect 651838 641880 651894 641889
rect 651838 641815 651894 641824
rect 651470 640792 651526 640801
rect 651470 640727 651526 640736
rect 651484 640354 651512 640727
rect 651472 640348 651524 640354
rect 651472 640290 651524 640296
rect 651380 640144 651432 640150
rect 651378 640112 651380 640121
rect 651432 640112 651434 640121
rect 651378 640047 651434 640056
rect 651656 638920 651708 638926
rect 651656 638862 651708 638868
rect 651472 638784 651524 638790
rect 651472 638726 651524 638732
rect 651484 638625 651512 638726
rect 651470 638616 651526 638625
rect 651470 638551 651526 638560
rect 651668 638217 651696 638862
rect 651654 638208 651710 638217
rect 651654 638143 651710 638152
rect 651852 635526 651880 641815
rect 653416 640150 653444 655522
rect 655520 645924 655572 645930
rect 655520 645866 655572 645872
rect 655336 643136 655388 643142
rect 655336 643078 655388 643084
rect 653404 640144 653456 640150
rect 653404 640086 653456 640092
rect 655348 638926 655376 643078
rect 655336 638920 655388 638926
rect 655336 638862 655388 638868
rect 655532 638790 655560 645866
rect 655520 638784 655572 638790
rect 655520 638726 655572 638732
rect 651840 635520 651892 635526
rect 651840 635462 651892 635468
rect 657556 625190 657584 688638
rect 658936 669526 658964 731410
rect 660316 714882 660344 777582
rect 668584 733440 668636 733446
rect 668584 733382 668636 733388
rect 661684 730720 661736 730726
rect 661684 730662 661736 730668
rect 660304 714876 660356 714882
rect 660304 714818 660356 714824
rect 661696 670750 661724 730662
rect 667848 703860 667900 703866
rect 667848 703802 667900 703808
rect 666468 701072 666520 701078
rect 666468 701014 666520 701020
rect 666284 696992 666336 696998
rect 666284 696934 666336 696940
rect 661684 670744 661736 670750
rect 661684 670686 661736 670692
rect 658924 669520 658976 669526
rect 658924 669462 658976 669468
rect 660304 642388 660356 642394
rect 660304 642330 660356 642336
rect 657544 625184 657596 625190
rect 657544 625126 657596 625132
rect 653404 611380 653456 611386
rect 653404 611322 653456 611328
rect 64328 610020 64380 610026
rect 64328 609962 64380 609968
rect 64340 231266 64368 609962
rect 651470 597952 651526 597961
rect 651470 597887 651526 597896
rect 651484 597582 651512 597887
rect 651472 597576 651524 597582
rect 651472 597518 651524 597524
rect 651470 596728 651526 596737
rect 651470 596663 651526 596672
rect 651484 596222 651512 596663
rect 651472 596216 651524 596222
rect 651472 596158 651524 596164
rect 653416 595542 653444 611322
rect 657544 600364 657596 600370
rect 657544 600306 657596 600312
rect 654784 599004 654836 599010
rect 654784 598946 654836 598952
rect 651656 595536 651708 595542
rect 651656 595478 651708 595484
rect 653404 595536 653456 595542
rect 653404 595478 653456 595484
rect 651470 595368 651526 595377
rect 651470 595303 651526 595312
rect 651484 594862 651512 595303
rect 651668 595105 651696 595478
rect 651654 595096 651710 595105
rect 651654 595031 651710 595040
rect 651472 594856 651524 594862
rect 651472 594798 651524 594804
rect 651472 594720 651524 594726
rect 651472 594662 651524 594668
rect 651484 594153 651512 594662
rect 651470 594144 651526 594153
rect 651470 594079 651526 594088
rect 654796 593298 654824 598946
rect 657556 594726 657584 600306
rect 658924 594856 658976 594862
rect 658924 594798 658976 594804
rect 657544 594720 657596 594726
rect 657544 594662 657596 594668
rect 651472 593292 651524 593298
rect 651472 593234 651524 593240
rect 654784 593292 654836 593298
rect 654784 593234 654836 593240
rect 651484 592929 651512 593234
rect 651470 592920 651526 592929
rect 651470 592855 651526 592864
rect 653404 565888 653456 565894
rect 653404 565830 653456 565836
rect 651470 553480 651526 553489
rect 651470 553415 651526 553424
rect 651484 552702 651512 553415
rect 651472 552696 651524 552702
rect 651472 552638 651524 552644
rect 651470 552120 651526 552129
rect 651470 552055 651526 552064
rect 651484 549914 651512 552055
rect 652022 551032 652078 551041
rect 652022 550967 652078 550976
rect 651656 550384 651708 550390
rect 651654 550352 651656 550361
rect 651708 550352 651710 550361
rect 651654 550287 651710 550296
rect 651472 549908 651524 549914
rect 651472 549850 651524 549856
rect 651470 549264 651526 549273
rect 651470 549199 651472 549208
rect 651524 549199 651526 549208
rect 651472 549170 651524 549176
rect 651472 548888 651524 548894
rect 651472 548830 651524 548836
rect 651484 548457 651512 548830
rect 651470 548448 651526 548457
rect 651470 548383 651526 548392
rect 652036 500274 652064 550967
rect 653416 550390 653444 565830
rect 655152 553444 655204 553450
rect 655152 553386 655204 553392
rect 653404 550384 653456 550390
rect 653404 550326 653456 550332
rect 655164 548894 655192 553386
rect 655152 548888 655204 548894
rect 655152 548830 655204 548836
rect 658936 534274 658964 594798
rect 660316 579698 660344 642330
rect 661684 635520 661736 635526
rect 661684 635462 661736 635468
rect 661696 581058 661724 635462
rect 666296 619750 666324 696934
rect 666480 621110 666508 701014
rect 667204 686520 667256 686526
rect 667204 686462 667256 686468
rect 667216 626142 667244 686462
rect 667204 626136 667256 626142
rect 667204 626078 667256 626084
rect 666468 621104 666520 621110
rect 666468 621046 666520 621052
rect 666284 619744 666336 619750
rect 666284 619686 666336 619692
rect 667386 600944 667442 600953
rect 667386 600879 667442 600888
rect 667204 596216 667256 596222
rect 667204 596158 667256 596164
rect 661684 581052 661736 581058
rect 661684 580994 661736 581000
rect 660304 579692 660356 579698
rect 660304 579634 660356 579640
rect 665088 564596 665140 564602
rect 665088 564538 665140 564544
rect 661040 554804 661092 554810
rect 661040 554746 661092 554752
rect 661052 549234 661080 554746
rect 664444 549908 664496 549914
rect 664444 549850 664496 549856
rect 661040 549228 661092 549234
rect 661040 549170 661092 549176
rect 658924 534268 658976 534274
rect 658924 534210 658976 534216
rect 663800 521620 663852 521626
rect 663800 521562 663852 521568
rect 663812 514078 663840 521562
rect 656348 514072 656400 514078
rect 656348 514014 656400 514020
rect 663800 514072 663852 514078
rect 663800 514014 663852 514020
rect 656360 510678 656388 514014
rect 653404 510672 653456 510678
rect 653404 510614 653456 510620
rect 656348 510672 656400 510678
rect 656348 510614 656400 510620
rect 652024 500268 652076 500274
rect 652024 500210 652076 500216
rect 653416 494766 653444 510614
rect 650644 494760 650696 494766
rect 650644 494702 650696 494708
rect 653404 494760 653456 494766
rect 653404 494702 653456 494708
rect 649264 290828 649316 290834
rect 649264 290770 649316 290776
rect 636198 278352 636254 278361
rect 69204 278316 69256 278322
rect 649276 278322 649304 290770
rect 636198 278287 636254 278296
rect 649264 278316 649316 278322
rect 69204 278258 69256 278264
rect 65904 272542 65932 278052
rect 67100 274242 67128 278052
rect 67088 274236 67140 274242
rect 67088 274178 67140 274184
rect 65892 272536 65944 272542
rect 65892 272478 65944 272484
rect 68204 271182 68232 278052
rect 69216 278050 69244 278258
rect 69204 278044 69256 278050
rect 69204 277986 69256 277992
rect 69400 273970 69428 278052
rect 69388 273964 69440 273970
rect 69388 273906 69440 273912
rect 68192 271176 68244 271182
rect 68192 271118 68244 271124
rect 70596 269822 70624 278052
rect 71792 275330 71820 278052
rect 71780 275324 71832 275330
rect 71780 275266 71832 275272
rect 72988 272678 73016 278052
rect 74184 274718 74212 278052
rect 74172 274712 74224 274718
rect 74172 274654 74224 274660
rect 72976 272672 73028 272678
rect 72976 272614 73028 272620
rect 75380 271454 75408 278052
rect 76484 275602 76512 278052
rect 76472 275596 76524 275602
rect 76472 275538 76524 275544
rect 76840 274712 76892 274718
rect 76840 274654 76892 274660
rect 75368 271448 75420 271454
rect 75368 271390 75420 271396
rect 76852 271318 76880 274654
rect 77680 274106 77708 278052
rect 77668 274100 77720 274106
rect 77668 274042 77720 274048
rect 76840 271312 76892 271318
rect 76840 271254 76892 271260
rect 78876 270366 78904 278052
rect 78864 270360 78916 270366
rect 78864 270302 78916 270308
rect 80072 269822 80100 278052
rect 81268 274990 81296 278052
rect 81256 274984 81308 274990
rect 81256 274926 81308 274932
rect 82464 272814 82492 278052
rect 83674 278038 84148 278066
rect 84778 278038 85528 278066
rect 82452 272808 82504 272814
rect 82452 272750 82504 272756
rect 84120 270502 84148 278038
rect 84108 270496 84160 270502
rect 84108 270438 84160 270444
rect 85500 269958 85528 278038
rect 85960 274718 85988 278052
rect 86224 275596 86276 275602
rect 86224 275538 86276 275544
rect 85948 274712 86000 274718
rect 85948 274654 86000 274660
rect 85488 269952 85540 269958
rect 85488 269894 85540 269900
rect 70584 269816 70636 269822
rect 70584 269758 70636 269764
rect 79324 269816 79376 269822
rect 79324 269758 79376 269764
rect 80060 269816 80112 269822
rect 80060 269758 80112 269764
rect 79336 267034 79364 269758
rect 86236 267442 86264 275538
rect 87156 271590 87184 278052
rect 88352 273834 88380 278052
rect 89562 278038 89668 278066
rect 88340 273828 88392 273834
rect 88340 273770 88392 273776
rect 87144 271584 87196 271590
rect 87144 271526 87196 271532
rect 89640 270094 89668 278038
rect 90744 275602 90772 278052
rect 91862 278038 92428 278066
rect 90732 275596 90784 275602
rect 90732 275538 90784 275544
rect 90364 274712 90416 274718
rect 90364 274654 90416 274660
rect 89628 270088 89680 270094
rect 89628 270030 89680 270036
rect 86224 267436 86276 267442
rect 86224 267378 86276 267384
rect 90376 267170 90404 274654
rect 92400 268394 92428 278038
rect 93044 275738 93072 278052
rect 93032 275732 93084 275738
rect 93032 275674 93084 275680
rect 94240 272950 94268 278052
rect 95436 274378 95464 278052
rect 96632 275194 96660 278052
rect 96620 275188 96672 275194
rect 96620 275130 96672 275136
rect 95424 274372 95476 274378
rect 95424 274314 95476 274320
rect 94228 272944 94280 272950
rect 94228 272886 94280 272892
rect 97828 271726 97856 278052
rect 99038 278038 99328 278066
rect 97816 271720 97868 271726
rect 97816 271662 97868 271668
rect 99300 268530 99328 278038
rect 100128 275466 100156 278052
rect 100116 275460 100168 275466
rect 100116 275402 100168 275408
rect 101324 274514 101352 278052
rect 101312 274508 101364 274514
rect 101312 274450 101364 274456
rect 102520 273086 102548 278052
rect 103716 274718 103744 278052
rect 104912 277394 104940 278052
rect 104912 277366 105032 277394
rect 103704 274712 103756 274718
rect 103704 274654 103756 274660
rect 104808 274712 104860 274718
rect 104808 274654 104860 274660
rect 102508 273080 102560 273086
rect 102508 273022 102560 273028
rect 99288 268524 99340 268530
rect 99288 268466 99340 268472
rect 92388 268388 92440 268394
rect 92388 268330 92440 268336
rect 104820 267306 104848 274654
rect 105004 268666 105032 277366
rect 106016 271862 106044 278052
rect 107212 276010 107240 278052
rect 107200 276004 107252 276010
rect 107200 275946 107252 275952
rect 108408 273222 108436 278052
rect 109618 278038 110368 278066
rect 108396 273216 108448 273222
rect 108396 273158 108448 273164
rect 106004 271856 106056 271862
rect 106004 271798 106056 271804
rect 110340 268802 110368 278038
rect 110800 274718 110828 278052
rect 110788 274712 110840 274718
rect 110788 274654 110840 274660
rect 111708 274712 111760 274718
rect 111708 274654 111760 274660
rect 110328 268796 110380 268802
rect 110328 268738 110380 268744
rect 104992 268660 105044 268666
rect 104992 268602 105044 268608
rect 111720 267578 111748 274654
rect 111996 270230 112024 278052
rect 113206 278038 113496 278066
rect 113468 271046 113496 278038
rect 114388 274650 114416 278052
rect 115506 278038 115888 278066
rect 114376 274644 114428 274650
rect 114376 274586 114428 274592
rect 113456 271040 113508 271046
rect 113456 270982 113508 270988
rect 111984 270224 112036 270230
rect 111984 270166 112036 270172
rect 115860 268938 115888 278038
rect 116688 272406 116716 278052
rect 117898 278038 118648 278066
rect 116676 272400 116728 272406
rect 116676 272342 116728 272348
rect 118620 269074 118648 278038
rect 119080 273698 119108 278052
rect 120276 273834 120304 278052
rect 119344 273828 119396 273834
rect 119344 273770 119396 273776
rect 120264 273828 120316 273834
rect 120264 273770 120316 273776
rect 119068 273692 119120 273698
rect 119068 273634 119120 273640
rect 118608 269068 118660 269074
rect 118608 269010 118660 269016
rect 115848 268932 115900 268938
rect 115848 268874 115900 268880
rect 119356 267714 119384 273770
rect 121472 270638 121500 278052
rect 122590 278038 122788 278066
rect 121460 270632 121512 270638
rect 121460 270574 121512 270580
rect 122760 269686 122788 278038
rect 123772 270910 123800 278052
rect 124968 271998 124996 278052
rect 126178 278038 126928 278066
rect 124956 271992 125008 271998
rect 124956 271934 125008 271940
rect 123760 270904 123812 270910
rect 123760 270846 123812 270852
rect 122748 269680 122800 269686
rect 122748 269622 122800 269628
rect 126900 269414 126928 278038
rect 127360 272270 127388 278052
rect 128556 274786 128584 278052
rect 128544 274780 128596 274786
rect 128544 274722 128596 274728
rect 127348 272264 127400 272270
rect 127348 272206 127400 272212
rect 129660 269550 129688 278052
rect 130856 274242 130884 278052
rect 130384 274236 130436 274242
rect 130384 274178 130436 274184
rect 130844 274236 130896 274242
rect 130844 274178 130896 274184
rect 129648 269544 129700 269550
rect 129648 269486 129700 269492
rect 126888 269408 126940 269414
rect 126888 269350 126940 269356
rect 119344 267708 119396 267714
rect 119344 267650 119396 267656
rect 111708 267572 111760 267578
rect 111708 267514 111760 267520
rect 104808 267300 104860 267306
rect 104808 267242 104860 267248
rect 90364 267164 90416 267170
rect 90364 267106 90416 267112
rect 79324 267028 79376 267034
rect 79324 266970 79376 266976
rect 130396 266626 130424 274178
rect 132052 273562 132080 278052
rect 133262 278038 133828 278066
rect 132040 273556 132092 273562
rect 132040 273498 132092 273504
rect 133800 270366 133828 278038
rect 134444 270774 134472 278052
rect 134432 270768 134484 270774
rect 134432 270710 134484 270716
rect 132500 270360 132552 270366
rect 132500 270302 132552 270308
rect 133788 270360 133840 270366
rect 133788 270302 133840 270308
rect 132512 266898 132540 270302
rect 135640 268258 135668 278052
rect 136836 275058 136864 278052
rect 136824 275052 136876 275058
rect 136824 274994 136876 275000
rect 137652 275052 137704 275058
rect 137652 274994 137704 275000
rect 136824 272536 136876 272542
rect 136824 272478 136876 272484
rect 135628 268252 135680 268258
rect 135628 268194 135680 268200
rect 132500 266892 132552 266898
rect 132500 266834 132552 266840
rect 130384 266620 130436 266626
rect 130384 266562 130436 266568
rect 136836 264330 136864 272478
rect 137664 270502 137692 274994
rect 137940 272542 137968 278052
rect 139136 275874 139164 278052
rect 140346 278038 140728 278066
rect 139124 275868 139176 275874
rect 139124 275810 139176 275816
rect 139400 273964 139452 273970
rect 139400 273906 139452 273912
rect 137928 272536 137980 272542
rect 137928 272478 137980 272484
rect 138480 271176 138532 271182
rect 138480 271118 138532 271124
rect 137468 270496 137520 270502
rect 137468 270438 137520 270444
rect 137652 270496 137704 270502
rect 137652 270438 137704 270444
rect 137480 266762 137508 270438
rect 137468 266756 137520 266762
rect 137468 266698 137520 266704
rect 138112 266620 138164 266626
rect 138112 266562 138164 266568
rect 136836 264302 137310 264330
rect 138124 264316 138152 266562
rect 138492 264330 138520 271118
rect 139412 264330 139440 273906
rect 140700 268410 140728 278038
rect 141056 275324 141108 275330
rect 141056 275266 141108 275272
rect 140700 268382 140912 268410
rect 140884 268258 140912 268382
rect 140688 268252 140740 268258
rect 140688 268194 140740 268200
rect 140872 268252 140924 268258
rect 140872 268194 140924 268200
rect 140700 267034 140728 268194
rect 140228 267028 140280 267034
rect 140228 266970 140280 266976
rect 140688 267028 140740 267034
rect 140688 266970 140740 266976
rect 140240 264330 140268 266970
rect 141068 264330 141096 275266
rect 141528 271182 141556 278052
rect 142724 272678 142752 278052
rect 142160 272672 142212 272678
rect 142160 272614 142212 272620
rect 142712 272672 142764 272678
rect 142712 272614 142764 272620
rect 141516 271176 141568 271182
rect 141516 271118 141568 271124
rect 142172 264330 142200 272614
rect 142712 271448 142764 271454
rect 142712 271390 142764 271396
rect 142724 264330 142752 271390
rect 143540 271312 143592 271318
rect 143540 271254 143592 271260
rect 143552 264330 143580 271254
rect 143920 269278 143948 278052
rect 144920 274100 144972 274106
rect 144920 274042 144972 274048
rect 143908 269272 143960 269278
rect 143908 269214 143960 269220
rect 144932 267734 144960 274042
rect 145116 272134 145144 278052
rect 146220 275058 146248 278052
rect 146208 275052 146260 275058
rect 146208 274994 146260 275000
rect 145288 274916 145340 274922
rect 145288 274858 145340 274864
rect 145300 273426 145328 274858
rect 145288 273420 145340 273426
rect 145288 273362 145340 273368
rect 147416 272678 147444 278052
rect 148612 273970 148640 278052
rect 149612 275188 149664 275194
rect 149612 275130 149664 275136
rect 148600 273964 148652 273970
rect 148600 273906 148652 273912
rect 147864 273420 147916 273426
rect 147864 273362 147916 273368
rect 145564 272672 145616 272678
rect 145564 272614 145616 272620
rect 147404 272672 147456 272678
rect 147404 272614 147456 272620
rect 145104 272128 145156 272134
rect 145104 272070 145156 272076
rect 144932 267706 145144 267734
rect 144736 267436 144788 267442
rect 144736 267378 144788 267384
rect 138492 264302 138966 264330
rect 139412 264302 139794 264330
rect 140240 264302 140622 264330
rect 141068 264302 141450 264330
rect 142172 264302 142278 264330
rect 142724 264302 143106 264330
rect 143552 264302 143934 264330
rect 144748 264316 144776 267378
rect 145116 264330 145144 267706
rect 145576 267442 145604 272614
rect 146392 269816 146444 269822
rect 146392 269758 146444 269764
rect 145564 267436 145616 267442
rect 145564 267378 145616 267384
rect 145116 264302 145590 264330
rect 146404 264316 146432 269758
rect 147220 266892 147272 266898
rect 147220 266834 147272 266840
rect 147232 264316 147260 266834
rect 147876 264330 147904 273362
rect 148416 272808 148468 272814
rect 148416 272750 148468 272756
rect 148428 264330 148456 272750
rect 149428 269952 149480 269958
rect 149428 269894 149480 269900
rect 149440 264330 149468 269894
rect 149624 266626 149652 275130
rect 149808 274922 149836 278052
rect 151018 278038 151768 278066
rect 149796 274916 149848 274922
rect 149796 274858 149848 274864
rect 151084 271992 151136 271998
rect 151084 271934 151136 271940
rect 151096 266762 151124 271934
rect 151740 268122 151768 278038
rect 152004 271584 152056 271590
rect 152004 271526 152056 271532
rect 151728 268116 151780 268122
rect 151728 268058 151780 268064
rect 151360 267164 151412 267170
rect 151360 267106 151412 267112
rect 150532 266756 150584 266762
rect 150532 266698 150584 266704
rect 151084 266756 151136 266762
rect 151084 266698 151136 266704
rect 149612 266620 149664 266626
rect 149612 266562 149664 266568
rect 147876 264302 148074 264330
rect 148428 264302 148902 264330
rect 149440 264302 149730 264330
rect 150544 264316 150572 266698
rect 151372 264316 151400 267106
rect 152016 264330 152044 271526
rect 152200 271318 152228 278052
rect 152832 275732 152884 275738
rect 152832 275674 152884 275680
rect 152188 271312 152240 271318
rect 152188 271254 152240 271260
rect 152844 269958 152872 275674
rect 153396 275194 153424 278052
rect 153384 275188 153436 275194
rect 153384 275130 153436 275136
rect 154500 274106 154528 278052
rect 154764 275596 154816 275602
rect 154764 275538 154816 275544
rect 154488 274100 154540 274106
rect 154488 274042 154540 274048
rect 153844 273556 153896 273562
rect 153844 273498 153896 273504
rect 153016 270088 153068 270094
rect 153016 270030 153068 270036
rect 152832 269952 152884 269958
rect 152832 269894 152884 269900
rect 152016 264302 152214 264330
rect 153028 264316 153056 270030
rect 153476 267708 153528 267714
rect 153476 267650 153528 267656
rect 153488 264330 153516 267650
rect 153856 266898 153884 273498
rect 154776 267734 154804 275538
rect 155696 272814 155724 278052
rect 156892 275466 156920 278052
rect 158102 278038 158668 278066
rect 156880 275460 156932 275466
rect 156880 275402 156932 275408
rect 157616 274372 157668 274378
rect 157616 274314 157668 274320
rect 155960 272944 156012 272950
rect 155960 272886 156012 272892
rect 155684 272808 155736 272814
rect 155684 272750 155736 272756
rect 155500 268388 155552 268394
rect 155500 268330 155552 268336
rect 154684 267706 154804 267734
rect 153844 266892 153896 266898
rect 153844 266834 153896 266840
rect 153488 264302 153870 264330
rect 154684 264316 154712 267706
rect 155512 264316 155540 268330
rect 155972 264330 156000 272886
rect 157156 269952 157208 269958
rect 157156 269894 157208 269900
rect 155972 264302 156354 264330
rect 157168 264316 157196 269894
rect 157628 264330 157656 274314
rect 158640 269822 158668 278038
rect 159284 274378 159312 278052
rect 160480 275738 160508 278052
rect 160468 275732 160520 275738
rect 160468 275674 160520 275680
rect 159456 275324 159508 275330
rect 159456 275266 159508 275272
rect 159272 274372 159324 274378
rect 159272 274314 159324 274320
rect 158812 271720 158864 271726
rect 158812 271662 158864 271668
rect 158628 269816 158680 269822
rect 158628 269758 158680 269764
rect 157628 264302 158010 264330
rect 158824 264316 158852 271662
rect 159468 267170 159496 275266
rect 160928 274508 160980 274514
rect 160928 274450 160980 274456
rect 160468 268524 160520 268530
rect 160468 268466 160520 268472
rect 159456 267164 159508 267170
rect 159456 267106 159508 267112
rect 159640 266620 159692 266626
rect 159640 266562 159692 266568
rect 159652 264316 159680 266562
rect 160480 264316 160508 268466
rect 160940 264330 160968 274450
rect 161584 268394 161612 278052
rect 162780 277394 162808 278052
rect 162688 277366 162808 277394
rect 162688 271454 162716 277366
rect 163504 276004 163556 276010
rect 163504 275946 163556 275952
rect 162860 273080 162912 273086
rect 162860 273022 162912 273028
rect 162676 271448 162728 271454
rect 162676 271390 162728 271396
rect 161572 268388 161624 268394
rect 161572 268330 161624 268336
rect 162124 267164 162176 267170
rect 162124 267106 162176 267112
rect 160940 264302 161322 264330
rect 162136 264316 162164 267106
rect 162872 264330 162900 273022
rect 163516 266422 163544 275946
rect 163976 275466 164004 278052
rect 163964 275460 164016 275466
rect 163964 275402 164016 275408
rect 164976 271856 165028 271862
rect 164976 271798 165028 271804
rect 163780 268660 163832 268666
rect 163780 268602 163832 268608
rect 163504 266416 163556 266422
rect 163504 266358 163556 266364
rect 162872 264302 162978 264330
rect 163792 264316 163820 268602
rect 164608 267300 164660 267306
rect 164608 267242 164660 267248
rect 164620 264316 164648 267242
rect 164988 264330 165016 271798
rect 165172 271590 165200 278052
rect 165896 273216 165948 273222
rect 165896 273158 165948 273164
rect 165160 271584 165212 271590
rect 165160 271526 165212 271532
rect 165908 264330 165936 273158
rect 166368 272950 166396 278052
rect 167564 276010 167592 278052
rect 167552 276004 167604 276010
rect 167552 275946 167604 275952
rect 168288 274780 168340 274786
rect 168288 274722 168340 274728
rect 166356 272944 166408 272950
rect 166356 272886 166408 272892
rect 168104 270632 168156 270638
rect 168104 270574 168156 270580
rect 167920 268796 167972 268802
rect 167920 268738 167972 268744
rect 167092 266416 167144 266422
rect 167092 266358 167144 266364
rect 164988 264302 165462 264330
rect 165908 264302 166290 264330
rect 167104 264316 167132 266358
rect 167932 264316 167960 268738
rect 168116 267170 168144 270574
rect 168300 268802 168328 274722
rect 168760 274514 168788 278052
rect 169024 275188 169076 275194
rect 169024 275130 169076 275136
rect 168748 274508 168800 274514
rect 168748 274450 168800 274456
rect 168748 270224 168800 270230
rect 168748 270166 168800 270172
rect 168288 268796 168340 268802
rect 168288 268738 168340 268744
rect 168104 267164 168156 267170
rect 168104 267106 168156 267112
rect 168760 264316 168788 270166
rect 169036 267578 169064 275130
rect 169864 271726 169892 278052
rect 171060 275602 171088 278052
rect 171048 275596 171100 275602
rect 171048 275538 171100 275544
rect 171600 274644 171652 274650
rect 171600 274586 171652 274592
rect 169852 271720 169904 271726
rect 169852 271662 169904 271668
rect 169944 271040 169996 271046
rect 169944 270982 169996 270988
rect 169576 267708 169628 267714
rect 169576 267650 169628 267656
rect 169024 267572 169076 267578
rect 169024 267514 169076 267520
rect 169588 264316 169616 267650
rect 169956 264330 169984 270982
rect 171232 268932 171284 268938
rect 171232 268874 171284 268880
rect 169956 264302 170430 264330
rect 171244 264316 171272 268874
rect 171612 264330 171640 274586
rect 172256 273086 172284 278052
rect 173466 278038 173848 278066
rect 174662 278038 175136 278066
rect 175858 278038 176608 278066
rect 173256 273692 173308 273698
rect 173256 273634 173308 273640
rect 172244 273080 172296 273086
rect 172244 273022 172296 273028
rect 172520 272400 172572 272406
rect 172520 272342 172572 272348
rect 172532 264330 172560 272342
rect 173268 264330 173296 273634
rect 173820 269958 173848 278038
rect 174268 275868 174320 275874
rect 174268 275810 174320 275816
rect 174280 271862 174308 275810
rect 174268 271856 174320 271862
rect 174268 271798 174320 271804
rect 173808 269952 173860 269958
rect 173808 269894 173860 269900
rect 175108 269074 175136 278038
rect 175280 273828 175332 273834
rect 175280 273770 175332 273776
rect 174544 269068 174596 269074
rect 174544 269010 174596 269016
rect 175096 269068 175148 269074
rect 175096 269010 175148 269016
rect 171612 264302 172086 264330
rect 172532 264302 172914 264330
rect 173268 264302 173742 264330
rect 174556 264316 174584 269010
rect 175292 264330 175320 273770
rect 176580 270094 176608 278038
rect 176568 270088 176620 270094
rect 176568 270030 176620 270036
rect 176200 269680 176252 269686
rect 176200 269622 176252 269628
rect 175292 264302 175398 264330
rect 176212 264316 176240 269622
rect 176948 268666 176976 278052
rect 178144 275874 178172 278052
rect 178684 276004 178736 276010
rect 178684 275946 178736 275952
rect 178132 275868 178184 275874
rect 178132 275810 178184 275816
rect 177488 270904 177540 270910
rect 177488 270846 177540 270852
rect 176936 268660 176988 268666
rect 176936 268602 176988 268608
rect 177028 267164 177080 267170
rect 177028 267106 177080 267112
rect 177040 264316 177068 267106
rect 177500 264330 177528 270846
rect 178316 269408 178368 269414
rect 178316 269350 178368 269356
rect 177672 269068 177724 269074
rect 177672 269010 177724 269016
rect 177684 267170 177712 269010
rect 177672 267164 177724 267170
rect 177672 267106 177724 267112
rect 178328 264330 178356 269350
rect 178696 267714 178724 275946
rect 179340 274650 179368 278052
rect 180550 278038 180748 278066
rect 179328 274644 179380 274650
rect 179328 274586 179380 274592
rect 179880 272264 179932 272270
rect 179880 272206 179932 272212
rect 178684 267708 178736 267714
rect 178684 267650 178736 267656
rect 179512 266756 179564 266762
rect 179512 266698 179564 266704
rect 177500 264302 177882 264330
rect 178328 264302 178710 264330
rect 179524 264316 179552 266698
rect 179892 264330 179920 272206
rect 180720 268530 180748 278038
rect 181732 272542 181760 278052
rect 182942 278038 183508 278066
rect 184138 278038 184888 278066
rect 182456 274236 182508 274242
rect 182456 274178 182508 274184
rect 181720 272536 181772 272542
rect 181720 272478 181772 272484
rect 181168 269544 181220 269550
rect 181168 269486 181220 269492
rect 180708 268524 180760 268530
rect 180708 268466 180760 268472
rect 179892 264302 180366 264330
rect 181180 264316 181208 269486
rect 181996 268796 182048 268802
rect 181996 268738 182048 268744
rect 182008 264316 182036 268738
rect 182468 264330 182496 274178
rect 183480 269686 183508 278038
rect 183652 270360 183704 270366
rect 183652 270302 183704 270308
rect 183468 269680 183520 269686
rect 183468 269622 183520 269628
rect 182468 264302 182850 264330
rect 183664 264316 183692 270302
rect 184860 270230 184888 278038
rect 185228 276010 185256 278052
rect 185216 276004 185268 276010
rect 185216 275946 185268 275952
rect 185308 275052 185360 275058
rect 185308 274994 185360 275000
rect 185124 270768 185176 270774
rect 185124 270710 185176 270716
rect 184848 270224 184900 270230
rect 184848 270166 184900 270172
rect 184480 266892 184532 266898
rect 184480 266834 184532 266840
rect 184492 264316 184520 266834
rect 185136 264330 185164 270710
rect 185320 270366 185348 274994
rect 186424 273222 186452 278052
rect 187436 278038 187634 278066
rect 186412 273216 186464 273222
rect 186412 273158 186464 273164
rect 186964 272536 187016 272542
rect 186964 272478 187016 272484
rect 186136 270496 186188 270502
rect 186136 270438 186188 270444
rect 185308 270360 185360 270366
rect 185308 270302 185360 270308
rect 185136 264302 185334 264330
rect 186148 264316 186176 270438
rect 186976 267306 187004 272478
rect 187436 271046 187464 278038
rect 188816 277394 188844 278052
rect 188816 277366 188936 277394
rect 187700 272400 187752 272406
rect 187700 272342 187752 272348
rect 187424 271040 187476 271046
rect 187424 270982 187476 270988
rect 186964 267300 187016 267306
rect 186964 267242 187016 267248
rect 186964 267028 187016 267034
rect 186964 266970 187016 266976
rect 186976 264316 187004 266970
rect 187712 264330 187740 272342
rect 188908 268802 188936 277366
rect 190012 275194 190040 278052
rect 190000 275188 190052 275194
rect 190000 275130 190052 275136
rect 189080 274916 189132 274922
rect 189080 274858 189132 274864
rect 189092 272270 189120 274858
rect 189080 272264 189132 272270
rect 189080 272206 189132 272212
rect 189172 271856 189224 271862
rect 189172 271798 189224 271804
rect 188896 268796 188948 268802
rect 188896 268738 188948 268744
rect 188620 268252 188672 268258
rect 188620 268194 188672 268200
rect 187712 264302 187818 264330
rect 188632 264316 188660 268194
rect 189184 264330 189212 271798
rect 191208 271182 191236 278052
rect 192404 274242 192432 278052
rect 192392 274236 192444 274242
rect 192392 274178 192444 274184
rect 193508 273834 193536 278052
rect 194718 278038 195008 278066
rect 194784 273964 194836 273970
rect 194784 273906 194836 273912
rect 193496 273828 193548 273834
rect 193496 273770 193548 273776
rect 193220 272672 193272 272678
rect 193220 272614 193272 272620
rect 192392 272128 192444 272134
rect 192392 272070 192444 272076
rect 189816 271176 189868 271182
rect 189816 271118 189868 271124
rect 191196 271176 191248 271182
rect 191196 271118 191248 271124
rect 189828 264330 189856 271118
rect 191104 269272 191156 269278
rect 191104 269214 191156 269220
rect 190460 268796 190512 268802
rect 190460 268738 190512 268744
rect 190472 267034 190500 268738
rect 190460 267028 190512 267034
rect 190460 266970 190512 266976
rect 189184 264302 189474 264330
rect 189828 264302 190302 264330
rect 191116 264316 191144 269214
rect 191932 267436 191984 267442
rect 191932 267378 191984 267384
rect 191944 264316 191972 267378
rect 192404 264330 192432 272070
rect 193232 264330 193260 272614
rect 194416 270360 194468 270366
rect 194416 270302 194468 270308
rect 192404 264302 192786 264330
rect 193232 264302 193614 264330
rect 194428 264316 194456 270302
rect 194796 264330 194824 273906
rect 194980 272406 195008 278038
rect 195900 272542 195928 278052
rect 197096 272678 197124 278052
rect 198096 274100 198148 274106
rect 198096 274042 198148 274048
rect 197084 272672 197136 272678
rect 197084 272614 197136 272620
rect 195888 272536 195940 272542
rect 195888 272478 195940 272484
rect 194968 272400 195020 272406
rect 194968 272342 195020 272348
rect 196440 272264 196492 272270
rect 196440 272206 196492 272212
rect 196072 268116 196124 268122
rect 196072 268058 196124 268064
rect 194796 264302 195270 264330
rect 196084 264316 196112 268058
rect 196452 264330 196480 272206
rect 197360 271312 197412 271318
rect 197360 271254 197412 271260
rect 197372 264330 197400 271254
rect 198108 264330 198136 274042
rect 198292 271318 198320 278052
rect 199502 278038 199976 278066
rect 199568 275732 199620 275738
rect 199568 275674 199620 275680
rect 198280 271312 198332 271318
rect 198280 271254 198332 271260
rect 199384 267572 199436 267578
rect 199384 267514 199436 267520
rect 196452 264302 196926 264330
rect 197372 264302 197754 264330
rect 198108 264302 198582 264330
rect 199396 264316 199424 267514
rect 199580 267442 199608 275674
rect 199948 270366 199976 278038
rect 200120 272808 200172 272814
rect 200120 272750 200172 272756
rect 199936 270360 199988 270366
rect 199936 270302 199988 270308
rect 199568 267436 199620 267442
rect 199568 267378 199620 267384
rect 200132 264330 200160 272750
rect 200592 268802 200620 278052
rect 201788 277394 201816 278052
rect 201696 277366 201816 277394
rect 201040 275324 201092 275330
rect 201040 275266 201092 275272
rect 201052 270502 201080 275266
rect 201040 270496 201092 270502
rect 201040 270438 201092 270444
rect 201696 269822 201724 277366
rect 202328 274372 202380 274378
rect 202328 274314 202380 274320
rect 201868 270496 201920 270502
rect 201868 270438 201920 270444
rect 201040 269816 201092 269822
rect 201040 269758 201092 269764
rect 201684 269816 201736 269822
rect 201684 269758 201736 269764
rect 200580 268796 200632 268802
rect 200580 268738 200632 268744
rect 200132 264302 200238 264330
rect 201052 264316 201080 269758
rect 201880 264316 201908 270438
rect 202340 264330 202368 274314
rect 202984 271862 203012 278052
rect 202972 271856 203024 271862
rect 202972 271798 203024 271804
rect 204180 269550 204208 278052
rect 205376 272814 205404 278052
rect 206586 278038 206876 278066
rect 206376 275460 206428 275466
rect 206376 275402 206428 275408
rect 205364 272808 205416 272814
rect 205364 272750 205416 272756
rect 205640 271584 205692 271590
rect 205640 271526 205692 271532
rect 204720 271448 204772 271454
rect 204720 271390 204772 271396
rect 204168 269544 204220 269550
rect 204168 269486 204220 269492
rect 203524 268388 203576 268394
rect 203524 268330 203576 268336
rect 202340 264302 202722 264330
rect 203536 264316 203564 268330
rect 204352 267436 204404 267442
rect 204352 267378 204404 267384
rect 204364 264316 204392 267378
rect 204732 264330 204760 271390
rect 205456 269680 205508 269686
rect 205456 269622 205508 269628
rect 205468 267442 205496 269622
rect 205456 267436 205508 267442
rect 205456 267378 205508 267384
rect 205652 264330 205680 271526
rect 206388 264330 206416 275402
rect 206848 270502 206876 278038
rect 207768 274786 207796 278052
rect 207756 274780 207808 274786
rect 207756 274722 207808 274728
rect 208400 274508 208452 274514
rect 208400 274450 208452 274456
rect 207296 272944 207348 272950
rect 207296 272886 207348 272892
rect 206836 270496 206888 270502
rect 206836 270438 206888 270444
rect 207308 264330 207336 272886
rect 208412 264330 208440 274450
rect 208872 273970 208900 278052
rect 210068 274106 210096 278052
rect 210700 274780 210752 274786
rect 210700 274722 210752 274728
rect 210056 274100 210108 274106
rect 210056 274042 210108 274048
rect 208860 273964 208912 273970
rect 208860 273906 208912 273912
rect 209780 273080 209832 273086
rect 209780 273022 209832 273028
rect 209320 267708 209372 267714
rect 209320 267650 209372 267656
rect 204732 264302 205206 264330
rect 205652 264302 206034 264330
rect 206388 264302 206862 264330
rect 207308 264302 207690 264330
rect 208412 264302 208518 264330
rect 209332 264316 209360 267650
rect 209792 265674 209820 273022
rect 209964 271720 210016 271726
rect 209964 271662 210016 271668
rect 209780 265668 209832 265674
rect 209780 265610 209832 265616
rect 209976 264330 210004 271662
rect 210712 268394 210740 274722
rect 211264 272950 211292 278052
rect 211436 275596 211488 275602
rect 211436 275538 211488 275544
rect 211252 272944 211304 272950
rect 211252 272886 211304 272892
rect 211160 270088 211212 270094
rect 211160 270030 211212 270036
rect 210700 268388 210752 268394
rect 210700 268330 210752 268336
rect 211172 266422 211200 270030
rect 211160 266416 211212 266422
rect 211160 266358 211212 266364
rect 210700 265668 210752 265674
rect 210700 265610 210752 265616
rect 210712 264330 210740 265610
rect 211448 264330 211476 275538
rect 212460 270094 212488 278052
rect 213656 271454 213684 278052
rect 214852 275330 214880 278052
rect 214840 275324 214892 275330
rect 214840 275266 214892 275272
rect 214564 274644 214616 274650
rect 214564 274586 214616 274592
rect 213644 271448 213696 271454
rect 213644 271390 213696 271396
rect 212448 270088 212500 270094
rect 212448 270030 212500 270036
rect 212632 269952 212684 269958
rect 212632 269894 212684 269900
rect 209976 264302 210174 264330
rect 210712 264302 211002 264330
rect 211448 264302 211830 264330
rect 212644 264316 212672 269894
rect 214288 267164 214340 267170
rect 214288 267106 214340 267112
rect 213460 266416 213512 266422
rect 213460 266358 213512 266364
rect 213472 264316 213500 266358
rect 214300 264316 214328 267106
rect 214576 266422 214604 274586
rect 215956 271590 215984 278052
rect 216680 275868 216732 275874
rect 216680 275810 216732 275816
rect 215944 271584 215996 271590
rect 215944 271526 215996 271532
rect 215944 271040 215996 271046
rect 215944 270982 215996 270988
rect 215116 268660 215168 268666
rect 215116 268602 215168 268608
rect 214564 266416 214616 266422
rect 214564 266358 214616 266364
rect 215128 264316 215156 268602
rect 215956 267578 215984 270982
rect 215944 267572 215996 267578
rect 215944 267514 215996 267520
rect 215944 266416 215996 266422
rect 215944 266358 215996 266364
rect 215956 264316 215984 266358
rect 216692 264330 216720 275810
rect 217152 275738 217180 278052
rect 217140 275732 217192 275738
rect 217140 275674 217192 275680
rect 218348 275602 218376 278052
rect 218336 275596 218388 275602
rect 218336 275538 218388 275544
rect 218704 273216 218756 273222
rect 218704 273158 218756 273164
rect 217600 268524 217652 268530
rect 217600 268466 217652 268472
rect 216692 264302 216798 264330
rect 217612 264316 217640 268466
rect 218428 267436 218480 267442
rect 218428 267378 218480 267384
rect 218440 264316 218468 267378
rect 218716 266898 218744 273158
rect 219544 273086 219572 278052
rect 219532 273080 219584 273086
rect 219532 273022 219584 273028
rect 220740 272950 220768 278052
rect 221280 276004 221332 276010
rect 221280 275946 221332 275952
rect 220084 272944 220136 272950
rect 220084 272886 220136 272892
rect 220728 272944 220780 272950
rect 220728 272886 220780 272892
rect 219348 270224 219400 270230
rect 219348 270166 219400 270172
rect 219360 267458 219388 270166
rect 219360 267430 219664 267458
rect 219256 267300 219308 267306
rect 219256 267242 219308 267248
rect 218704 266892 218756 266898
rect 218704 266834 218756 266840
rect 219268 264316 219296 267242
rect 219636 264330 219664 267430
rect 220096 267170 220124 272886
rect 220084 267164 220136 267170
rect 220084 267106 220136 267112
rect 220912 266892 220964 266898
rect 220912 266834 220964 266840
rect 219636 264302 220110 264330
rect 220924 264316 220952 266834
rect 221292 264330 221320 275946
rect 221936 275466 221964 278052
rect 221924 275460 221976 275466
rect 221924 275402 221976 275408
rect 222936 275188 222988 275194
rect 222936 275130 222988 275136
rect 222568 267572 222620 267578
rect 222568 267514 222620 267520
rect 221292 264302 221766 264330
rect 222580 264316 222608 267514
rect 222948 264330 222976 275130
rect 223132 274378 223160 278052
rect 224236 275874 224264 278052
rect 224224 275868 224276 275874
rect 224224 275810 224276 275816
rect 224224 275732 224276 275738
rect 224224 275674 224276 275680
rect 223120 274372 223172 274378
rect 223120 274314 223172 274320
rect 223488 269544 223540 269550
rect 223488 269486 223540 269492
rect 223500 267306 223528 269486
rect 224236 268666 224264 275674
rect 224960 274236 225012 274242
rect 224960 274178 225012 274184
rect 224224 268660 224276 268666
rect 224224 268602 224276 268608
rect 223488 267300 223540 267306
rect 223488 267242 223540 267248
rect 224224 267028 224276 267034
rect 224224 266970 224276 266976
rect 222948 264302 223422 264330
rect 224236 264316 224264 266970
rect 224972 265674 225000 274178
rect 225432 271726 225460 278052
rect 226432 273828 226484 273834
rect 226432 273770 226484 273776
rect 225420 271720 225472 271726
rect 225420 271662 225472 271668
rect 225144 271176 225196 271182
rect 225144 271118 225196 271124
rect 224960 265668 225012 265674
rect 224960 265610 225012 265616
rect 225156 265554 225184 271118
rect 225604 265668 225656 265674
rect 225604 265610 225656 265616
rect 225064 265526 225184 265554
rect 225064 264316 225092 265526
rect 225616 264330 225644 265610
rect 226444 264330 226472 273770
rect 226628 269958 226656 278052
rect 227838 278038 228128 278066
rect 228100 272542 228128 278038
rect 229020 275738 229048 278052
rect 229008 275732 229060 275738
rect 229008 275674 229060 275680
rect 229100 272672 229152 272678
rect 229100 272614 229152 272620
rect 227904 272536 227956 272542
rect 227904 272478 227956 272484
rect 228088 272536 228140 272542
rect 228088 272478 228140 272484
rect 227168 272400 227220 272406
rect 227168 272342 227220 272348
rect 226616 269952 226668 269958
rect 226616 269894 226668 269900
rect 227180 264330 227208 272342
rect 227916 264330 227944 272478
rect 228364 271720 228416 271726
rect 228364 271662 228416 271668
rect 228376 267034 228404 271662
rect 228364 267028 228416 267034
rect 228364 266970 228416 266976
rect 229112 264330 229140 272614
rect 229560 271312 229612 271318
rect 229560 271254 229612 271260
rect 229572 264330 229600 271254
rect 230216 271182 230244 278052
rect 231334 278038 231716 278066
rect 230204 271176 230256 271182
rect 230204 271118 230256 271124
rect 230848 270360 230900 270366
rect 230848 270302 230900 270308
rect 225616 264302 225906 264330
rect 226444 264302 226734 264330
rect 227180 264302 227562 264330
rect 227916 264302 228390 264330
rect 229112 264302 229218 264330
rect 229572 264302 230046 264330
rect 230860 264316 230888 270302
rect 231308 268796 231360 268802
rect 231308 268738 231360 268744
rect 231320 264330 231348 268738
rect 231688 268530 231716 278038
rect 232516 276010 232544 278052
rect 232504 276004 232556 276010
rect 232504 275946 232556 275952
rect 232688 275868 232740 275874
rect 232688 275810 232740 275816
rect 232700 270366 232728 275810
rect 233712 272678 233740 278052
rect 234922 278038 235304 278066
rect 233884 275596 233936 275602
rect 233884 275538 233936 275544
rect 233700 272672 233752 272678
rect 233700 272614 233752 272620
rect 233240 271856 233292 271862
rect 233240 271798 233292 271804
rect 232688 270360 232740 270366
rect 232688 270302 232740 270308
rect 232504 269816 232556 269822
rect 232504 269758 232556 269764
rect 231676 268524 231728 268530
rect 231676 268466 231728 268472
rect 231320 264302 231702 264330
rect 232516 264316 232544 269758
rect 233252 264330 233280 271798
rect 233896 267442 233924 275538
rect 234804 272808 234856 272814
rect 234804 272750 234856 272756
rect 233884 267436 233936 267442
rect 233884 267378 233936 267384
rect 234160 267300 234212 267306
rect 234160 267242 234212 267248
rect 233252 264302 233358 264330
rect 234172 264316 234200 267242
rect 234816 264330 234844 272750
rect 235276 271318 235304 278038
rect 236104 275874 236132 278052
rect 236092 275868 236144 275874
rect 236092 275810 236144 275816
rect 235264 271312 235316 271318
rect 235264 271254 235316 271260
rect 235816 270496 235868 270502
rect 235816 270438 235868 270444
rect 234816 264302 235014 264330
rect 235828 264316 235856 270438
rect 237300 269822 237328 278052
rect 237840 274100 237892 274106
rect 237840 274042 237892 274048
rect 237472 273964 237524 273970
rect 237472 273906 237524 273912
rect 237288 269816 237340 269822
rect 237288 269758 237340 269764
rect 236644 268388 236696 268394
rect 236644 268330 236696 268336
rect 236656 264316 236684 268330
rect 237484 264316 237512 273906
rect 237852 264330 237880 274042
rect 238496 273970 238524 278052
rect 239600 275602 239628 278052
rect 240048 276004 240100 276010
rect 240048 275946 240100 275952
rect 239588 275596 239640 275602
rect 239588 275538 239640 275544
rect 239404 275324 239456 275330
rect 239404 275266 239456 275272
rect 238484 273964 238536 273970
rect 238484 273906 238536 273912
rect 239128 267164 239180 267170
rect 239128 267106 239180 267112
rect 237852 264302 238326 264330
rect 239140 264316 239168 267106
rect 239416 266422 239444 275266
rect 240060 274242 240088 275946
rect 240048 274236 240100 274242
rect 240048 274178 240100 274184
rect 240796 271454 240824 278052
rect 241992 277394 242020 278052
rect 241900 277366 242020 277394
rect 240416 271448 240468 271454
rect 240416 271390 240468 271396
rect 240784 271448 240836 271454
rect 240784 271390 240836 271396
rect 239956 270088 240008 270094
rect 239956 270030 240008 270036
rect 239404 266416 239456 266422
rect 239404 266358 239456 266364
rect 239968 264316 239996 270030
rect 240428 264330 240456 271390
rect 241900 270094 241928 277366
rect 243188 275330 243216 278052
rect 243728 275732 243780 275738
rect 243728 275674 243780 275680
rect 243544 275460 243596 275466
rect 243544 275402 243596 275408
rect 243176 275324 243228 275330
rect 243176 275266 243228 275272
rect 242072 271584 242124 271590
rect 242072 271526 242124 271532
rect 241888 270088 241940 270094
rect 241888 270030 241940 270036
rect 241612 266416 241664 266422
rect 241612 266358 241664 266364
rect 240428 264302 240810 264330
rect 241624 264316 241652 266358
rect 242084 264330 242112 271526
rect 243268 268660 243320 268666
rect 243268 268602 243320 268608
rect 242084 264302 242466 264330
rect 243280 264316 243308 268602
rect 243556 266422 243584 275402
rect 243740 267442 243768 275674
rect 244384 270230 244412 278052
rect 245396 278038 245502 278066
rect 246790 278038 246988 278066
rect 244556 273080 244608 273086
rect 244556 273022 244608 273028
rect 244372 270224 244424 270230
rect 244372 270166 244424 270172
rect 243728 267436 243780 267442
rect 243728 267378 243780 267384
rect 244096 267300 244148 267306
rect 244096 267242 244148 267248
rect 243544 266416 243596 266422
rect 243544 266358 243596 266364
rect 244108 264316 244136 267242
rect 244568 264330 244596 273022
rect 245396 272814 245424 278038
rect 245752 272944 245804 272950
rect 245752 272886 245804 272892
rect 245384 272808 245436 272814
rect 245384 272750 245436 272756
rect 244568 264302 244950 264330
rect 245764 264316 245792 272886
rect 246960 267170 246988 278038
rect 247224 274372 247276 274378
rect 247224 274314 247276 274320
rect 246948 267164 247000 267170
rect 246948 267106 247000 267112
rect 246580 266416 246632 266422
rect 246580 266358 246632 266364
rect 246592 264316 246620 266358
rect 247236 264330 247264 274314
rect 247880 272950 247908 278052
rect 249076 274106 249104 278052
rect 250272 275738 250300 278052
rect 250444 275868 250496 275874
rect 250444 275810 250496 275816
rect 250260 275732 250312 275738
rect 250260 275674 250312 275680
rect 249064 274100 249116 274106
rect 249064 274042 249116 274048
rect 247868 272944 247920 272950
rect 247868 272886 247920 272892
rect 249064 272536 249116 272542
rect 249064 272478 249116 272484
rect 248236 270360 248288 270366
rect 248236 270302 248288 270308
rect 247236 264302 247434 264330
rect 248248 264316 248276 270302
rect 248788 267028 248840 267034
rect 248788 266970 248840 266976
rect 248800 264330 248828 266970
rect 249076 266422 249104 272478
rect 249892 269952 249944 269958
rect 249892 269894 249944 269900
rect 249064 266416 249116 266422
rect 249064 266358 249116 266364
rect 248800 264302 249090 264330
rect 249904 264316 249932 269894
rect 250456 266558 250484 275810
rect 251468 271046 251496 278052
rect 252008 271176 252060 271182
rect 252008 271118 252060 271124
rect 251456 271040 251508 271046
rect 251456 270982 251508 270988
rect 251548 267436 251600 267442
rect 251548 267378 251600 267384
rect 250444 266552 250496 266558
rect 250444 266494 250496 266500
rect 250720 266416 250772 266422
rect 250720 266358 250772 266364
rect 250732 264316 250760 266358
rect 251560 264316 251588 267378
rect 252020 264330 252048 271118
rect 252664 268394 252692 278052
rect 253860 274718 253888 278052
rect 253848 274712 253900 274718
rect 253848 274654 253900 274660
rect 253940 274236 253992 274242
rect 253940 274178 253992 274184
rect 253204 268524 253256 268530
rect 253204 268466 253256 268472
rect 252652 268388 252704 268394
rect 252652 268330 252704 268336
rect 252020 264302 252402 264330
rect 253216 264316 253244 268466
rect 253952 264330 253980 274178
rect 254400 272672 254452 272678
rect 254400 272614 254452 272620
rect 254412 264330 254440 272614
rect 254964 272542 254992 278052
rect 255964 275596 256016 275602
rect 255964 275538 256016 275544
rect 254952 272536 255004 272542
rect 254952 272478 255004 272484
rect 255320 271312 255372 271318
rect 255320 271254 255372 271260
rect 255332 264330 255360 271254
rect 255976 267034 256004 275538
rect 256160 275466 256188 278052
rect 257356 275602 257384 278052
rect 257344 275596 257396 275602
rect 257344 275538 257396 275544
rect 256148 275460 256200 275466
rect 256148 275402 256200 275408
rect 256700 275324 256752 275330
rect 256700 275266 256752 275272
rect 256712 271318 256740 275266
rect 256884 274712 256936 274718
rect 256884 274654 256936 274660
rect 256700 271312 256752 271318
rect 256700 271254 256752 271260
rect 256896 269958 256924 274654
rect 258080 273828 258132 273834
rect 258080 273770 258132 273776
rect 256884 269952 256936 269958
rect 256884 269894 256936 269900
rect 257344 269816 257396 269822
rect 257344 269758 257396 269764
rect 255964 267028 256016 267034
rect 255964 266970 256016 266976
rect 256516 266552 256568 266558
rect 256516 266494 256568 266500
rect 253952 264302 254058 264330
rect 254412 264302 254886 264330
rect 255332 264302 255714 264330
rect 256528 264316 256556 266494
rect 257356 264316 257384 269758
rect 258092 264330 258120 273770
rect 258552 269822 258580 278052
rect 259748 277394 259776 278052
rect 259748 277366 259868 277394
rect 259368 275732 259420 275738
rect 259368 275674 259420 275680
rect 259380 273562 259408 275674
rect 259368 273556 259420 273562
rect 259368 273498 259420 273504
rect 259840 271454 259868 277366
rect 260944 275806 260972 278052
rect 260932 275800 260984 275806
rect 260932 275742 260984 275748
rect 259644 271448 259696 271454
rect 259644 271390 259696 271396
rect 259828 271448 259880 271454
rect 259828 271390 259880 271396
rect 258540 269816 258592 269822
rect 258540 269758 258592 269764
rect 259000 267028 259052 267034
rect 259000 266970 259052 266976
rect 258092 264302 258198 264330
rect 259012 264316 259040 266970
rect 259656 264330 259684 271390
rect 262048 271318 262076 278052
rect 262312 275596 262364 275602
rect 262312 275538 262364 275544
rect 262324 272814 262352 275538
rect 263244 275330 263272 278052
rect 263232 275324 263284 275330
rect 263232 275266 263284 275272
rect 264244 272944 264296 272950
rect 264244 272886 264296 272892
rect 262312 272808 262364 272814
rect 262312 272750 262364 272756
rect 262680 272672 262732 272678
rect 262680 272614 262732 272620
rect 261024 271312 261076 271318
rect 261024 271254 261076 271260
rect 262036 271312 262088 271318
rect 262036 271254 262088 271260
rect 260656 270088 260708 270094
rect 260656 270030 260708 270036
rect 259656 264302 259854 264330
rect 260668 264316 260696 270030
rect 261036 264330 261064 271254
rect 262312 270224 262364 270230
rect 262312 270166 262364 270172
rect 261036 264302 261510 264330
rect 262324 264316 262352 270166
rect 262692 264330 262720 272614
rect 264256 267734 264284 272886
rect 264440 272678 264468 278052
rect 265650 278038 266216 278066
rect 265256 274100 265308 274106
rect 265256 274042 265308 274048
rect 264428 272672 264480 272678
rect 264428 272614 264480 272620
rect 264256 267706 264376 267734
rect 263968 267164 264020 267170
rect 263968 267106 264020 267112
rect 262692 264302 263166 264330
rect 263980 264316 264008 267106
rect 264348 264330 264376 267706
rect 265268 264330 265296 274042
rect 266188 270094 266216 278038
rect 266360 275800 266412 275806
rect 266360 275742 266412 275748
rect 266372 274106 266400 275742
rect 266832 275602 266860 278052
rect 266820 275596 266872 275602
rect 266820 275538 266872 275544
rect 266360 274100 266412 274106
rect 266360 274042 266412 274048
rect 266360 273556 266412 273562
rect 266360 273498 266412 273504
rect 266176 270088 266228 270094
rect 266176 270030 266228 270036
rect 266372 264330 266400 273498
rect 268028 271182 268056 278052
rect 269224 275126 269252 278052
rect 270132 275460 270184 275466
rect 270132 275402 270184 275408
rect 269212 275120 269264 275126
rect 269212 275062 269264 275068
rect 269304 272536 269356 272542
rect 269304 272478 269356 272484
rect 268016 271176 268068 271182
rect 268016 271118 268068 271124
rect 266912 271040 266964 271046
rect 266912 270982 266964 270988
rect 266924 264330 266952 270982
rect 268936 269952 268988 269958
rect 268936 269894 268988 269900
rect 268108 268388 268160 268394
rect 268108 268330 268160 268336
rect 264348 264302 264822 264330
rect 265268 264302 265650 264330
rect 266372 264302 266478 264330
rect 266924 264302 267306 264330
rect 268120 264316 268148 268330
rect 268948 264316 268976 269894
rect 269316 264330 269344 272478
rect 270144 272354 270172 275402
rect 270328 272542 270356 278052
rect 271524 273970 271552 278052
rect 272734 278038 273116 278066
rect 271512 273964 271564 273970
rect 271512 273906 271564 273912
rect 270960 272808 271012 272814
rect 270960 272750 271012 272756
rect 270316 272536 270368 272542
rect 270316 272478 270368 272484
rect 270144 272326 270540 272354
rect 270512 264330 270540 272326
rect 270972 264330 271000 272750
rect 272616 271448 272668 271454
rect 272616 271390 272668 271396
rect 272248 269816 272300 269822
rect 272248 269758 272300 269764
rect 269316 264302 269790 264330
rect 270512 264302 270618 264330
rect 270972 264302 271446 264330
rect 272260 264316 272288 269758
rect 272628 264330 272656 271390
rect 273088 269822 273116 278038
rect 273260 275324 273312 275330
rect 273260 275266 273312 275272
rect 273076 269816 273128 269822
rect 273076 269758 273128 269764
rect 273272 269074 273300 275266
rect 273536 274100 273588 274106
rect 273536 274042 273588 274048
rect 273260 269068 273312 269074
rect 273260 269010 273312 269016
rect 273548 264330 273576 274042
rect 273916 272814 273944 278052
rect 274640 275120 274692 275126
rect 274640 275062 274692 275068
rect 273904 272808 273956 272814
rect 273904 272750 273956 272756
rect 274652 271862 274680 275062
rect 275112 274718 275140 278052
rect 276308 275330 276336 278052
rect 276480 275596 276532 275602
rect 276480 275538 276532 275544
rect 276296 275324 276348 275330
rect 276296 275266 276348 275272
rect 275100 274712 275152 274718
rect 275100 274654 275152 274660
rect 276020 272672 276072 272678
rect 276020 272614 276072 272620
rect 274640 271856 274692 271862
rect 274640 271798 274692 271804
rect 274640 271312 274692 271318
rect 274640 271254 274692 271260
rect 274652 264330 274680 271254
rect 275560 269068 275612 269074
rect 275560 269010 275612 269016
rect 272628 264302 273102 264330
rect 273548 264302 273930 264330
rect 274652 264302 274758 264330
rect 275572 264316 275600 269010
rect 276032 264330 276060 272614
rect 276492 267782 276520 275538
rect 277504 275534 277532 278052
rect 277492 275528 277544 275534
rect 277492 275470 277544 275476
rect 278044 274712 278096 274718
rect 278044 274654 278096 274660
rect 278056 270502 278084 274654
rect 278608 274106 278636 278052
rect 278596 274100 278648 274106
rect 278596 274042 278648 274048
rect 279240 271856 279292 271862
rect 279240 271798 279292 271804
rect 278780 271176 278832 271182
rect 278780 271118 278832 271124
rect 278044 270496 278096 270502
rect 278044 270438 278096 270444
rect 277216 270088 277268 270094
rect 277216 270030 277268 270036
rect 276480 267776 276532 267782
rect 276480 267718 276532 267724
rect 276032 264302 276414 264330
rect 277228 264316 277256 270030
rect 278044 267776 278096 267782
rect 278044 267718 278096 267724
rect 278056 264316 278084 267718
rect 278792 264330 278820 271118
rect 279252 264330 279280 271798
rect 279804 271182 279832 278052
rect 280344 273964 280396 273970
rect 280344 273906 280396 273912
rect 279792 271176 279844 271182
rect 279792 271118 279844 271124
rect 280356 265674 280384 273906
rect 281000 273086 281028 278052
rect 282210 278038 282776 278066
rect 280988 273080 281040 273086
rect 280988 273022 281040 273028
rect 280528 272536 280580 272542
rect 280528 272478 280580 272484
rect 280344 265668 280396 265674
rect 280344 265610 280396 265616
rect 278792 264302 278898 264330
rect 279252 264302 279726 264330
rect 280540 264316 280568 272478
rect 282184 269816 282236 269822
rect 282184 269758 282236 269764
rect 280988 265668 281040 265674
rect 280988 265610 281040 265616
rect 281000 264330 281028 265610
rect 281000 264302 281382 264330
rect 282196 264316 282224 269758
rect 282748 269278 282776 278038
rect 283104 275324 283156 275330
rect 283104 275266 283156 275272
rect 282920 272808 282972 272814
rect 282920 272750 282972 272756
rect 282736 269272 282788 269278
rect 282736 269214 282788 269220
rect 282932 264330 282960 272750
rect 283116 270366 283144 275266
rect 283392 274718 283420 278052
rect 284588 275874 284616 278052
rect 284576 275868 284628 275874
rect 284576 275810 284628 275816
rect 285128 275528 285180 275534
rect 285128 275470 285180 275476
rect 283380 274712 283432 274718
rect 283380 274654 283432 274660
rect 283840 270496 283892 270502
rect 283840 270438 283892 270444
rect 283104 270360 283156 270366
rect 283104 270302 283156 270308
rect 282932 264302 283038 264330
rect 283852 264316 283880 270438
rect 284668 270360 284720 270366
rect 284668 270302 284720 270308
rect 284680 264316 284708 270302
rect 285140 264330 285168 275470
rect 285692 275330 285720 278052
rect 286888 275738 286916 278052
rect 286876 275732 286928 275738
rect 286876 275674 286928 275680
rect 285680 275324 285732 275330
rect 285680 275266 285732 275272
rect 288084 275058 288112 278052
rect 288072 275052 288124 275058
rect 288072 274994 288124 275000
rect 289280 274922 289308 278052
rect 290096 275868 290148 275874
rect 290096 275810 290148 275816
rect 289268 274916 289320 274922
rect 289268 274858 289320 274864
rect 289176 274712 289228 274718
rect 289176 274654 289228 274660
rect 285864 274100 285916 274106
rect 285864 274042 285916 274048
rect 285876 264330 285904 274042
rect 286324 273080 286376 273086
rect 286324 273022 286376 273028
rect 286336 267034 286364 273022
rect 287060 271176 287112 271182
rect 287060 271118 287112 271124
rect 286324 267028 286376 267034
rect 286324 266970 286376 266976
rect 287072 264330 287100 271118
rect 288808 269272 288860 269278
rect 288808 269214 288860 269220
rect 287980 267028 288032 267034
rect 287980 266970 288032 266976
rect 285140 264302 285522 264330
rect 285876 264302 286350 264330
rect 287072 264302 287178 264330
rect 287992 264316 288020 266970
rect 288820 264316 288848 269214
rect 289188 264330 289216 274654
rect 290108 264330 290136 275810
rect 290476 274718 290504 278052
rect 291672 275330 291700 278052
rect 291844 275732 291896 275738
rect 291844 275674 291896 275680
rect 291292 275324 291344 275330
rect 291292 275266 291344 275272
rect 291660 275324 291712 275330
rect 291660 275266 291712 275272
rect 290464 274712 290516 274718
rect 290464 274654 290516 274660
rect 289188 264302 289662 264330
rect 290108 264302 290490 264330
rect 291304 264316 291332 275266
rect 291856 264330 291884 275674
rect 292868 275194 292896 278052
rect 292856 275188 292908 275194
rect 292856 275130 292908 275136
rect 292856 275052 292908 275058
rect 292856 274994 292908 275000
rect 292672 274916 292724 274922
rect 292672 274858 292724 274864
rect 292684 265674 292712 274858
rect 292672 265668 292724 265674
rect 292672 265610 292724 265616
rect 292868 264330 292896 274994
rect 293972 274990 294000 278052
rect 293960 274984 294012 274990
rect 293960 274926 294012 274932
rect 295168 274854 295196 278052
rect 295340 275324 295392 275330
rect 295340 275266 295392 275272
rect 295156 274848 295208 274854
rect 295156 274790 295208 274796
rect 294144 274712 294196 274718
rect 294144 274654 294196 274660
rect 293500 265668 293552 265674
rect 293500 265610 293552 265616
rect 293512 264330 293540 265610
rect 294156 264330 294184 274654
rect 295352 264330 295380 275266
rect 295800 275188 295852 275194
rect 295800 275130 295852 275136
rect 295812 264330 295840 275130
rect 296364 274718 296392 278052
rect 297560 275398 297588 278052
rect 297548 275392 297600 275398
rect 297548 275334 297600 275340
rect 298756 275262 298784 278052
rect 299952 275398 299980 278052
rect 300964 278038 301070 278066
rect 302266 278038 302464 278066
rect 299572 275392 299624 275398
rect 299572 275334 299624 275340
rect 299940 275392 299992 275398
rect 299940 275334 299992 275340
rect 298744 275256 298796 275262
rect 298744 275198 298796 275204
rect 296812 274984 296864 274990
rect 296812 274926 296864 274932
rect 296352 274712 296404 274718
rect 296352 274654 296404 274660
rect 296824 264330 296852 274926
rect 297456 274848 297508 274854
rect 297456 274790 297508 274796
rect 297468 264330 297496 274790
rect 298376 274712 298428 274718
rect 298376 274654 298428 274660
rect 298388 264330 298416 274654
rect 291856 264302 292146 264330
rect 292868 264302 292974 264330
rect 293512 264302 293802 264330
rect 294156 264302 294630 264330
rect 295352 264302 295458 264330
rect 295812 264302 296286 264330
rect 296824 264302 297114 264330
rect 297468 264302 297942 264330
rect 298388 264302 298770 264330
rect 299584 264316 299612 275334
rect 300032 275256 300084 275262
rect 300032 275198 300084 275204
rect 300044 264330 300072 275198
rect 300964 266422 300992 278038
rect 301136 275392 301188 275398
rect 301136 275334 301188 275340
rect 300952 266416 301004 266422
rect 300952 266358 301004 266364
rect 301148 264330 301176 275334
rect 302056 266416 302108 266422
rect 302056 266358 302108 266364
rect 300044 264302 300426 264330
rect 301148 264302 301254 264330
rect 302068 264316 302096 266358
rect 302436 264330 302464 278038
rect 303448 274718 303476 278052
rect 303724 278038 304658 278066
rect 305012 278038 305854 278066
rect 306392 278038 307050 278066
rect 307772 278038 308154 278066
rect 309152 278038 309350 278066
rect 303436 274712 303488 274718
rect 303436 274654 303488 274660
rect 303724 266422 303752 278038
rect 303988 274712 304040 274718
rect 303988 274654 304040 274660
rect 303712 266416 303764 266422
rect 303712 266358 303764 266364
rect 304000 264330 304028 274654
rect 304540 266416 304592 266422
rect 304540 266358 304592 266364
rect 302436 264302 302910 264330
rect 303738 264302 304028 264330
rect 304552 264316 304580 266358
rect 305012 264330 305040 278038
rect 306392 266370 306420 278038
rect 307772 267734 307800 278038
rect 306208 266342 306420 266370
rect 307496 267706 307800 267734
rect 305012 264302 305394 264330
rect 306208 264316 306236 266342
rect 307496 264330 307524 267706
rect 308680 266688 308732 266694
rect 308680 266630 308732 266636
rect 307852 266416 307904 266422
rect 307852 266358 307904 266364
rect 307050 264302 307524 264330
rect 307864 264316 307892 266358
rect 308692 264316 308720 266630
rect 309152 266422 309180 278038
rect 310532 277394 310560 278052
rect 310808 278038 311742 278066
rect 311912 278038 312938 278066
rect 313292 278038 314134 278066
rect 314672 278038 315238 278066
rect 316052 278038 316434 278066
rect 317432 278038 317630 278066
rect 318826 278038 319300 278066
rect 310532 277366 310652 277394
rect 310624 266694 310652 277366
rect 310612 266688 310664 266694
rect 310612 266630 310664 266636
rect 310336 266552 310388 266558
rect 310336 266494 310388 266500
rect 309140 266416 309192 266422
rect 309140 266358 309192 266364
rect 309508 266416 309560 266422
rect 309508 266358 309560 266364
rect 309520 264316 309548 266358
rect 310348 264316 310376 266494
rect 310808 266422 310836 278038
rect 311912 266558 311940 278038
rect 312820 266892 312872 266898
rect 312820 266834 312872 266840
rect 311900 266552 311952 266558
rect 311900 266494 311952 266500
rect 312360 266552 312412 266558
rect 312360 266494 312412 266500
rect 310796 266416 310848 266422
rect 310796 266358 310848 266364
rect 311164 266416 311216 266422
rect 311164 266358 311216 266364
rect 311176 264316 311204 266358
rect 312372 264330 312400 266494
rect 312018 264302 312400 264330
rect 312832 264316 312860 266834
rect 313292 266422 313320 278038
rect 314476 267164 314528 267170
rect 314476 267106 314528 267112
rect 313648 267028 313700 267034
rect 313648 266970 313700 266976
rect 313280 266416 313332 266422
rect 313280 266358 313332 266364
rect 313660 264316 313688 266970
rect 314488 264316 314516 267106
rect 314672 266558 314700 278038
rect 315304 267436 315356 267442
rect 315304 267378 315356 267384
rect 314660 266552 314712 266558
rect 314660 266494 314712 266500
rect 315316 264316 315344 267378
rect 316052 266898 316080 278038
rect 317432 267034 317460 278038
rect 319076 272604 319128 272610
rect 319076 272546 319128 272552
rect 318708 272468 318760 272474
rect 318708 272410 318760 272416
rect 318720 267734 318748 272410
rect 318628 267706 318748 267734
rect 317420 267028 317472 267034
rect 317420 266970 317472 266976
rect 316040 266892 316092 266898
rect 316040 266834 316092 266840
rect 317788 266824 317840 266830
rect 317788 266766 317840 266772
rect 316960 266688 317012 266694
rect 316960 266630 317012 266636
rect 316132 266552 316184 266558
rect 316132 266494 316184 266500
rect 316144 264316 316172 266494
rect 316972 264316 317000 266630
rect 317800 264316 317828 266766
rect 318628 264316 318656 267706
rect 319088 267442 319116 272546
rect 319076 267436 319128 267442
rect 319076 267378 319128 267384
rect 319272 267170 319300 278038
rect 319640 278038 320022 278066
rect 320192 278038 321218 278066
rect 321572 278038 322414 278066
rect 322952 278038 323518 278066
rect 319640 272610 319668 278038
rect 319628 272604 319680 272610
rect 319628 272546 319680 272552
rect 319444 269136 319496 269142
rect 319444 269078 319496 269084
rect 319260 267164 319312 267170
rect 319260 267106 319312 267112
rect 319456 264316 319484 269078
rect 320192 266558 320220 278038
rect 321192 274712 321244 274718
rect 321192 274654 321244 274660
rect 321204 267734 321232 274654
rect 321376 270768 321428 270774
rect 321376 270710 321428 270716
rect 321112 267706 321232 267734
rect 320180 266552 320232 266558
rect 320180 266494 320232 266500
rect 320272 266416 320324 266422
rect 320272 266358 320324 266364
rect 320284 264316 320312 266358
rect 321112 264316 321140 267706
rect 321388 266422 321416 270710
rect 321572 266694 321600 278038
rect 322756 273964 322808 273970
rect 322756 273906 322808 273912
rect 321928 267300 321980 267306
rect 321928 267242 321980 267248
rect 321560 266688 321612 266694
rect 321560 266630 321612 266636
rect 321376 266416 321428 266422
rect 321376 266358 321428 266364
rect 321940 264316 321968 267242
rect 322768 264316 322796 273906
rect 322952 266830 322980 278038
rect 324044 272672 324096 272678
rect 324044 272614 324096 272620
rect 322940 266824 322992 266830
rect 322940 266766 322992 266772
rect 324056 264330 324084 272614
rect 324700 272474 324728 278052
rect 325712 278038 325910 278066
rect 325332 272808 325384 272814
rect 325332 272750 325384 272756
rect 324688 272468 324740 272474
rect 324688 272410 324740 272416
rect 325344 266422 325372 272750
rect 325516 271448 325568 271454
rect 325516 271390 325568 271396
rect 324412 266416 324464 266422
rect 324412 266358 324464 266364
rect 325332 266416 325384 266422
rect 325332 266358 325384 266364
rect 323610 264302 324084 264330
rect 324424 264316 324452 266358
rect 325528 264330 325556 271390
rect 325712 269142 325740 278038
rect 326436 275324 326488 275330
rect 326436 275266 326488 275272
rect 325700 269136 325752 269142
rect 325700 269078 325752 269084
rect 326448 264330 326476 275266
rect 327092 270774 327120 278052
rect 328288 274718 328316 278052
rect 328276 274712 328328 274718
rect 328276 274654 328328 274660
rect 329484 273290 329512 278052
rect 330588 273970 330616 278052
rect 330576 273964 330628 273970
rect 330576 273906 330628 273912
rect 327724 273284 327776 273290
rect 327724 273226 327776 273232
rect 329472 273284 329524 273290
rect 329472 273226 329524 273232
rect 327080 270768 327132 270774
rect 327080 270710 327132 270716
rect 326896 269816 326948 269822
rect 326896 269758 326948 269764
rect 325266 264302 325556 264330
rect 326094 264302 326476 264330
rect 326908 264316 326936 269758
rect 327736 267306 327764 273226
rect 331784 272678 331812 278052
rect 331956 274304 332008 274310
rect 331956 274246 332008 274252
rect 331772 272672 331824 272678
rect 331772 272614 331824 272620
rect 329748 272536 329800 272542
rect 329748 272478 329800 272484
rect 329564 271312 329616 271318
rect 329564 271254 329616 271260
rect 327724 267300 327776 267306
rect 327724 267242 327776 267248
rect 327724 266552 327776 266558
rect 327724 266494 327776 266500
rect 327736 264316 327764 266494
rect 328552 266416 328604 266422
rect 328552 266358 328604 266364
rect 328564 264316 328592 266358
rect 329576 264330 329604 271254
rect 329760 266422 329788 272478
rect 331128 271176 331180 271182
rect 331128 271118 331180 271124
rect 330208 269952 330260 269958
rect 330208 269894 330260 269900
rect 329748 266416 329800 266422
rect 329748 266358 329800 266364
rect 329406 264302 329604 264330
rect 330220 264316 330248 269894
rect 331140 267734 331168 271118
rect 331048 267706 331168 267734
rect 331048 264316 331076 267706
rect 331968 266558 331996 274246
rect 332980 272814 333008 278052
rect 333796 272944 333848 272950
rect 333796 272886 333848 272892
rect 332968 272808 333020 272814
rect 332968 272750 333020 272756
rect 332324 272672 332376 272678
rect 332324 272614 332376 272620
rect 331956 266552 332008 266558
rect 331956 266494 332008 266500
rect 332336 264330 332364 272614
rect 332692 266892 332744 266898
rect 332692 266834 332744 266840
rect 331890 264302 332364 264330
rect 332704 264316 332732 266834
rect 333808 264330 333836 272886
rect 334176 271454 334204 278052
rect 335372 275330 335400 278052
rect 335556 278038 336582 278066
rect 335360 275324 335412 275330
rect 335360 275266 335412 275272
rect 335268 273964 335320 273970
rect 335268 273906 335320 273912
rect 334164 271448 334216 271454
rect 334164 271390 334216 271396
rect 334348 270224 334400 270230
rect 334348 270166 334400 270172
rect 333546 264302 333836 264330
rect 334360 264316 334388 270166
rect 335280 267734 335308 273906
rect 335556 269822 335584 278038
rect 337764 274310 337792 278052
rect 337752 274304 337804 274310
rect 337752 274246 337804 274252
rect 337752 274100 337804 274106
rect 337752 274042 337804 274048
rect 335544 269816 335596 269822
rect 335544 269758 335596 269764
rect 336004 269816 336056 269822
rect 336004 269758 336056 269764
rect 335188 267706 335308 267734
rect 335188 264316 335216 267706
rect 336016 264316 336044 269758
rect 337764 267734 337792 274042
rect 338868 272542 338896 278052
rect 338856 272536 338908 272542
rect 338856 272478 338908 272484
rect 339224 272536 339276 272542
rect 339224 272478 339276 272484
rect 337936 271584 337988 271590
rect 337936 271526 337988 271532
rect 337672 267706 337792 267734
rect 336832 266416 336884 266422
rect 336832 266358 336884 266364
rect 336844 264316 336872 266358
rect 337672 264316 337700 267706
rect 337948 266422 337976 271526
rect 338488 268524 338540 268530
rect 338488 268466 338540 268472
rect 337936 266416 337988 266422
rect 337936 266358 337988 266364
rect 338500 264316 338528 268466
rect 339236 264330 339264 272478
rect 340064 271318 340092 278052
rect 340892 278038 341274 278066
rect 340052 271312 340104 271318
rect 340052 271254 340104 271260
rect 340604 271312 340656 271318
rect 340604 271254 340656 271260
rect 340616 264330 340644 271254
rect 340892 269958 340920 278038
rect 342456 271182 342484 278052
rect 343652 272678 343680 278052
rect 343836 278038 344862 278066
rect 343640 272672 343692 272678
rect 343640 272614 343692 272620
rect 342444 271176 342496 271182
rect 342444 271118 342496 271124
rect 343548 271176 343600 271182
rect 343548 271118 343600 271124
rect 340880 269952 340932 269958
rect 340880 269894 340932 269900
rect 341800 269952 341852 269958
rect 341800 269894 341852 269900
rect 340972 267436 341024 267442
rect 340972 267378 341024 267384
rect 339236 264302 339342 264330
rect 340170 264302 340644 264330
rect 340984 264316 341012 267378
rect 341812 264316 341840 269894
rect 343560 267734 343588 271118
rect 343468 267706 343588 267734
rect 342628 266416 342680 266422
rect 342628 266358 342680 266364
rect 342640 264316 342668 266358
rect 343468 264316 343496 267706
rect 343836 266898 343864 278038
rect 345952 272950 345980 278052
rect 346412 278038 347162 278066
rect 345940 272944 345992 272950
rect 345940 272886 345992 272892
rect 344652 272808 344704 272814
rect 344652 272750 344704 272756
rect 343824 266892 343876 266898
rect 343824 266834 343876 266840
rect 344664 264330 344692 272750
rect 346216 272672 346268 272678
rect 346216 272614 346268 272620
rect 345296 270088 345348 270094
rect 345296 270030 345348 270036
rect 345112 266552 345164 266558
rect 345112 266494 345164 266500
rect 344310 264302 344692 264330
rect 345124 264316 345152 266494
rect 345308 266422 345336 270030
rect 345296 266416 345348 266422
rect 345296 266358 345348 266364
rect 346228 264330 346256 272614
rect 346412 270230 346440 278038
rect 348344 273970 348372 278052
rect 349172 278038 349554 278066
rect 348332 273964 348384 273970
rect 348332 273906 348384 273912
rect 348424 272944 348476 272950
rect 348424 272886 348476 272892
rect 347688 271448 347740 271454
rect 347688 271390 347740 271396
rect 346400 270224 346452 270230
rect 346400 270166 346452 270172
rect 347504 266688 347556 266694
rect 347504 266630 347556 266636
rect 346768 266416 346820 266422
rect 346768 266358 346820 266364
rect 345966 264302 346256 264330
rect 346780 264316 346808 266358
rect 347516 264330 347544 266630
rect 347700 266422 347728 271390
rect 348436 266558 348464 272886
rect 349172 269822 349200 278038
rect 350356 273964 350408 273970
rect 350356 273906 350408 273912
rect 349160 269816 349212 269822
rect 349160 269758 349212 269764
rect 348792 268388 348844 268394
rect 348792 268330 348844 268336
rect 348424 266552 348476 266558
rect 348424 266494 348476 266500
rect 347688 266416 347740 266422
rect 347688 266358 347740 266364
rect 348804 264330 348832 268330
rect 350080 266552 350132 266558
rect 350080 266494 350132 266500
rect 349252 266416 349304 266422
rect 349252 266358 349304 266364
rect 347516 264302 347622 264330
rect 348450 264302 348832 264330
rect 349264 264316 349292 266358
rect 350092 264316 350120 266494
rect 350368 266422 350396 273906
rect 350736 271590 350764 278052
rect 351932 274106 351960 278052
rect 352116 278038 353142 278066
rect 351920 274100 351972 274106
rect 351920 274042 351972 274048
rect 351184 271720 351236 271726
rect 351184 271662 351236 271668
rect 350724 271584 350776 271590
rect 350724 271526 350776 271532
rect 350908 267300 350960 267306
rect 350908 267242 350960 267248
rect 350356 266416 350408 266422
rect 350356 266358 350408 266364
rect 350920 264316 350948 267242
rect 351196 266694 351224 271662
rect 351736 269816 351788 269822
rect 351736 269758 351788 269764
rect 351184 266688 351236 266694
rect 351184 266630 351236 266636
rect 351748 264316 351776 269758
rect 352116 268530 352144 278038
rect 353944 274100 353996 274106
rect 353944 274042 353996 274048
rect 352564 268660 352616 268666
rect 352564 268602 352616 268608
rect 352104 268524 352156 268530
rect 352104 268466 352156 268472
rect 352576 264316 352604 268602
rect 353392 267028 353444 267034
rect 353392 266970 353444 266976
rect 353404 264316 353432 266970
rect 353956 266558 353984 274042
rect 354232 272542 354260 278052
rect 355152 278038 355442 278066
rect 354220 272536 354272 272542
rect 354220 272478 354272 272484
rect 354496 272536 354548 272542
rect 354496 272478 354548 272484
rect 353944 266552 353996 266558
rect 353944 266494 353996 266500
rect 354508 264330 354536 272478
rect 355152 271318 355180 278038
rect 356624 271862 356652 278052
rect 357452 278038 357834 278066
rect 358832 278038 359030 278066
rect 355324 271856 355376 271862
rect 355324 271798 355376 271804
rect 356612 271856 356664 271862
rect 356612 271798 356664 271804
rect 355140 271312 355192 271318
rect 355140 271254 355192 271260
rect 355048 270360 355100 270366
rect 355048 270302 355100 270308
rect 354246 264302 354536 264330
rect 355060 264316 355088 270302
rect 355336 267442 355364 271798
rect 357164 271312 357216 271318
rect 357164 271254 357216 271260
rect 355324 267436 355376 267442
rect 355324 267378 355376 267384
rect 355876 266552 355928 266558
rect 355876 266494 355928 266500
rect 355888 264316 355916 266494
rect 357176 264330 357204 271254
rect 357452 269958 357480 278038
rect 358636 275460 358688 275466
rect 358636 275402 358688 275408
rect 357440 269952 357492 269958
rect 357440 269894 357492 269900
rect 357532 266416 357584 266422
rect 357532 266358 357584 266364
rect 356730 264302 357204 264330
rect 357544 264316 357572 266358
rect 358648 264330 358676 275402
rect 358832 270094 358860 278038
rect 359464 274236 359516 274242
rect 359464 274178 359516 274184
rect 358820 270088 358872 270094
rect 358820 270030 358872 270036
rect 359188 269952 359240 269958
rect 359188 269894 359240 269900
rect 358386 264302 358676 264330
rect 359200 264316 359228 269894
rect 359476 266422 359504 274178
rect 360212 271182 360240 278052
rect 361212 273080 361264 273086
rect 361212 273022 361264 273028
rect 360844 271584 360896 271590
rect 360844 271526 360896 271532
rect 360200 271176 360252 271182
rect 360200 271118 360252 271124
rect 360016 267164 360068 267170
rect 360016 267106 360068 267112
rect 359464 266416 359516 266422
rect 359464 266358 359516 266364
rect 360028 264316 360056 267106
rect 360856 266558 360884 271526
rect 360844 266552 360896 266558
rect 360844 266494 360896 266500
rect 361224 264330 361252 273022
rect 361408 272814 361436 278052
rect 362512 272950 362540 278052
rect 362776 273216 362828 273222
rect 362776 273158 362828 273164
rect 362500 272944 362552 272950
rect 362500 272886 362552 272892
rect 361396 272808 361448 272814
rect 361396 272750 361448 272756
rect 362224 272808 362276 272814
rect 362224 272750 362276 272756
rect 362236 267306 362264 272750
rect 362500 267572 362552 267578
rect 362500 267514 362552 267520
rect 362224 267300 362276 267306
rect 362224 267242 362276 267248
rect 361672 266416 361724 266422
rect 361672 266358 361724 266364
rect 360870 264302 361252 264330
rect 361684 264316 361712 266358
rect 362512 264316 362540 267514
rect 362788 266422 362816 273158
rect 363708 272678 363736 278052
rect 363880 275596 363932 275602
rect 363880 275538 363932 275544
rect 363696 272672 363748 272678
rect 363696 272614 363748 272620
rect 363892 267734 363920 275538
rect 364904 271454 364932 278052
rect 365444 272944 365496 272950
rect 365444 272886 365496 272892
rect 364892 271448 364944 271454
rect 364892 271390 364944 271396
rect 364156 271176 364208 271182
rect 364156 271118 364208 271124
rect 363800 267706 363920 267734
rect 362776 266416 362828 266422
rect 362776 266358 362828 266364
rect 363800 264330 363828 267706
rect 363354 264302 363828 264330
rect 364168 264316 364196 271118
rect 365456 264330 365484 272886
rect 366100 271726 366128 278052
rect 367112 278038 367310 278066
rect 366088 271720 366140 271726
rect 366088 271662 366140 271668
rect 366364 271448 366416 271454
rect 366364 271390 366416 271396
rect 365812 267436 365864 267442
rect 365812 267378 365864 267384
rect 365010 264302 365484 264330
rect 365824 264316 365852 267378
rect 366376 267170 366404 271390
rect 366640 270088 366692 270094
rect 366640 270030 366692 270036
rect 366364 267164 366416 267170
rect 366364 267106 366416 267112
rect 366652 264316 366680 270030
rect 367112 268394 367140 278038
rect 368492 273970 368520 278052
rect 369124 274372 369176 274378
rect 369124 274314 369176 274320
rect 368480 273964 368532 273970
rect 368480 273906 368532 273912
rect 367468 268524 367520 268530
rect 367468 268466 367520 268472
rect 367100 268388 367152 268394
rect 367100 268330 367152 268336
rect 367480 264316 367508 268466
rect 369136 267578 369164 274314
rect 369596 274106 369624 278052
rect 370332 278038 370806 278066
rect 371252 278038 372002 278066
rect 372632 278038 373198 278066
rect 369584 274100 369636 274106
rect 369584 274042 369636 274048
rect 370332 272814 370360 278038
rect 371056 275324 371108 275330
rect 371056 275266 371108 275272
rect 370320 272808 370372 272814
rect 370320 272750 370372 272756
rect 370504 272808 370556 272814
rect 370504 272750 370556 272756
rect 369124 267572 369176 267578
rect 369124 267514 369176 267520
rect 368296 266756 368348 266762
rect 368296 266698 368348 266704
rect 368308 264316 368336 266698
rect 369952 266552 370004 266558
rect 369952 266494 370004 266500
rect 369124 266416 369176 266422
rect 369124 266358 369176 266364
rect 369136 264316 369164 266358
rect 369964 264316 369992 266494
rect 370516 266422 370544 272750
rect 370504 266416 370556 266422
rect 370504 266358 370556 266364
rect 371068 264330 371096 275266
rect 371252 269822 371280 278038
rect 372252 270224 372304 270230
rect 372252 270166 372304 270172
rect 371240 269816 371292 269822
rect 371240 269758 371292 269764
rect 372264 266558 372292 270166
rect 372632 268666 372660 278038
rect 374380 277394 374408 278052
rect 374380 277366 374500 277394
rect 373264 274100 373316 274106
rect 373264 274042 373316 274048
rect 372620 268660 372672 268666
rect 372620 268602 372672 268608
rect 372436 268388 372488 268394
rect 372436 268330 372488 268336
rect 372252 266552 372304 266558
rect 372252 266494 372304 266500
rect 371608 266416 371660 266422
rect 371608 266358 371660 266364
rect 370806 264302 371096 264330
rect 371620 264316 371648 266358
rect 372448 264316 372476 268330
rect 373276 266422 373304 274042
rect 374472 267306 374500 277366
rect 375576 272542 375604 278052
rect 376116 272672 376168 272678
rect 376116 272614 376168 272620
rect 375564 272536 375616 272542
rect 375564 272478 375616 272484
rect 375288 271856 375340 271862
rect 375288 271798 375340 271804
rect 374460 267300 374512 267306
rect 374460 267242 374512 267248
rect 373632 267164 373684 267170
rect 373632 267106 373684 267112
rect 373264 266416 373316 266422
rect 373264 266358 373316 266364
rect 373644 264330 373672 267106
rect 374920 266892 374972 266898
rect 374920 266834 374972 266840
rect 374092 266416 374144 266422
rect 374092 266358 374144 266364
rect 373290 264302 373672 264330
rect 374104 264316 374132 266358
rect 374932 264316 374960 266834
rect 375300 266422 375328 271798
rect 375288 266416 375340 266422
rect 375288 266358 375340 266364
rect 376128 264330 376156 272614
rect 376772 270366 376800 278052
rect 377680 273964 377732 273970
rect 377680 273906 377732 273912
rect 376760 270360 376812 270366
rect 376760 270302 376812 270308
rect 376576 269816 376628 269822
rect 376576 269758 376628 269764
rect 375774 264302 376156 264330
rect 376588 264316 376616 269758
rect 377692 264330 377720 273906
rect 377876 271590 377904 278052
rect 377864 271584 377916 271590
rect 377864 271526 377916 271532
rect 379072 271318 379100 278052
rect 380268 274242 380296 278052
rect 381464 275466 381492 278052
rect 382292 278038 382674 278066
rect 381452 275460 381504 275466
rect 381452 275402 381504 275408
rect 381544 274508 381596 274514
rect 381544 274450 381596 274456
rect 380256 274236 380308 274242
rect 380256 274178 380308 274184
rect 379428 272536 379480 272542
rect 379428 272478 379480 272484
rect 379060 271312 379112 271318
rect 379060 271254 379112 271260
rect 378784 267300 378836 267306
rect 378784 267242 378836 267248
rect 378796 266762 378824 267242
rect 378784 266756 378836 266762
rect 378784 266698 378836 266704
rect 378232 266620 378284 266626
rect 378232 266562 378284 266568
rect 377430 264302 377720 264330
rect 378244 264316 378272 266562
rect 379440 264330 379468 272478
rect 380532 270360 380584 270366
rect 380532 270302 380584 270308
rect 380544 266898 380572 270302
rect 380716 267572 380768 267578
rect 380716 267514 380768 267520
rect 380532 266892 380584 266898
rect 380532 266834 380584 266840
rect 379888 266416 379940 266422
rect 379888 266358 379940 266364
rect 379086 264302 379468 264330
rect 379900 264316 379928 266358
rect 380728 264316 380756 267514
rect 381556 267442 381584 274450
rect 382004 271720 382056 271726
rect 382004 271662 382056 271668
rect 381544 267436 381596 267442
rect 381544 267378 381596 267384
rect 382016 264330 382044 271662
rect 382292 269958 382320 278038
rect 383856 271454 383884 278052
rect 385052 274666 385080 278052
rect 384960 274638 385080 274666
rect 385880 278038 386170 278066
rect 384960 273086 384988 274638
rect 385880 273222 385908 278038
rect 386052 275460 386104 275466
rect 386052 275402 386104 275408
rect 385868 273216 385920 273222
rect 385868 273158 385920 273164
rect 384948 273080 385000 273086
rect 384948 273022 385000 273028
rect 385684 273080 385736 273086
rect 385684 273022 385736 273028
rect 384948 272128 385000 272134
rect 384948 272070 385000 272076
rect 383844 271448 383896 271454
rect 383844 271390 383896 271396
rect 384764 271448 384816 271454
rect 384764 271390 384816 271396
rect 382280 269952 382332 269958
rect 382280 269894 382332 269900
rect 383016 269952 383068 269958
rect 383016 269894 383068 269900
rect 382372 268932 382424 268938
rect 382372 268874 382424 268880
rect 381570 264302 382044 264330
rect 382384 264316 382412 268874
rect 383028 266422 383056 269894
rect 383200 267436 383252 267442
rect 383200 267378 383252 267384
rect 383016 266416 383068 266422
rect 383016 266358 383068 266364
rect 383212 264316 383240 267378
rect 384028 266416 384080 266422
rect 384028 266358 384080 266364
rect 384040 264316 384068 266358
rect 384776 264330 384804 271390
rect 384960 266422 384988 272070
rect 385696 267306 385724 273022
rect 385684 267300 385736 267306
rect 385684 267242 385736 267248
rect 384948 266416 385000 266422
rect 384948 266358 385000 266364
rect 386064 264330 386092 275402
rect 387352 274378 387380 278052
rect 388548 275602 388576 278052
rect 388536 275596 388588 275602
rect 388536 275538 388588 275544
rect 387340 274372 387392 274378
rect 387340 274314 387392 274320
rect 388996 274236 389048 274242
rect 388996 274178 389048 274184
rect 387708 271584 387760 271590
rect 387708 271526 387760 271532
rect 387340 268796 387392 268802
rect 387340 268738 387392 268744
rect 386512 266416 386564 266422
rect 386512 266358 386564 266364
rect 384776 264302 384882 264330
rect 385710 264302 386092 264330
rect 386524 264316 386552 266358
rect 387352 264316 387380 268738
rect 387720 266422 387748 271526
rect 388168 266892 388220 266898
rect 388168 266834 388220 266840
rect 387708 266416 387760 266422
rect 387708 266358 387760 266364
rect 388180 264316 388208 266834
rect 389008 264316 389036 274178
rect 389744 271182 389772 278052
rect 390940 272950 390968 278052
rect 392136 274514 392164 278052
rect 392124 274508 392176 274514
rect 392124 274450 392176 274456
rect 390928 272944 390980 272950
rect 390928 272886 390980 272892
rect 391848 272264 391900 272270
rect 391848 272206 391900 272212
rect 390284 271312 390336 271318
rect 390284 271254 390336 271260
rect 389732 271176 389784 271182
rect 389732 271118 389784 271124
rect 390296 264330 390324 271254
rect 390652 267708 390704 267714
rect 390652 267650 390704 267656
rect 389850 264302 390324 264330
rect 390664 264316 390692 267650
rect 391860 264330 391888 272206
rect 393332 270094 393360 278052
rect 393516 278038 394450 278066
rect 393320 270088 393372 270094
rect 393320 270030 393372 270036
rect 392032 269680 392084 269686
rect 392032 269622 392084 269628
rect 392044 267170 392072 269622
rect 393516 268530 393544 278038
rect 395632 273086 395660 278052
rect 395620 273080 395672 273086
rect 395620 273022 395672 273028
rect 396828 272814 396856 278052
rect 397472 278038 398038 278066
rect 397000 273828 397052 273834
rect 397000 273770 397052 273776
rect 396816 272808 396868 272814
rect 396816 272750 396868 272756
rect 395988 272400 396040 272406
rect 395988 272342 396040 272348
rect 394332 271176 394384 271182
rect 394332 271118 394384 271124
rect 393688 268660 393740 268666
rect 393688 268602 393740 268608
rect 393504 268524 393556 268530
rect 393504 268466 393556 268472
rect 392032 267164 392084 267170
rect 392032 267106 392084 267112
rect 393136 267028 393188 267034
rect 393136 266970 393188 266976
rect 392308 266416 392360 266422
rect 392308 266358 392360 266364
rect 391506 264302 391888 264330
rect 392320 264316 392348 266358
rect 393148 264316 393176 266970
rect 393700 266422 393728 268602
rect 393688 266416 393740 266422
rect 393688 266358 393740 266364
rect 394344 264330 394372 271118
rect 394700 270088 394752 270094
rect 394700 270030 394752 270036
rect 394712 266762 394740 270030
rect 394700 266756 394752 266762
rect 394700 266698 394752 266704
rect 394792 266620 394844 266626
rect 394792 266562 394844 266568
rect 393990 264302 394372 264330
rect 394804 264316 394832 266562
rect 396000 264330 396028 272342
rect 397012 267734 397040 273770
rect 397472 270230 397500 278038
rect 399220 275330 399248 278052
rect 399208 275324 399260 275330
rect 399208 275266 399260 275272
rect 400324 274106 400352 278052
rect 400508 278038 401534 278066
rect 401704 278038 402730 278066
rect 400312 274100 400364 274106
rect 400312 274042 400364 274048
rect 400036 273216 400088 273222
rect 400036 273158 400088 273164
rect 397460 270224 397512 270230
rect 397460 270166 397512 270172
rect 398748 269544 398800 269550
rect 398748 269486 398800 269492
rect 397276 268524 397328 268530
rect 397276 268466 397328 268472
rect 396920 267706 397040 267734
rect 396920 264330 396948 267706
rect 395646 264302 396028 264330
rect 396474 264302 396948 264330
rect 397288 264316 397316 268466
rect 398760 267578 398788 269486
rect 398748 267572 398800 267578
rect 398748 267514 398800 267520
rect 398104 267300 398156 267306
rect 398104 267242 398156 267248
rect 398116 264316 398144 267242
rect 399760 267164 399812 267170
rect 399760 267106 399812 267112
rect 398932 266416 398984 266422
rect 398932 266358 398984 266364
rect 398944 264316 398972 266358
rect 399772 264316 399800 267106
rect 400048 266422 400076 273158
rect 400508 268394 400536 278038
rect 401508 274100 401560 274106
rect 401508 274042 401560 274048
rect 400864 270496 400916 270502
rect 400864 270438 400916 270444
rect 400496 268388 400548 268394
rect 400496 268330 400548 268336
rect 400036 266416 400088 266422
rect 400036 266358 400088 266364
rect 400876 264330 400904 270438
rect 401520 267734 401548 274042
rect 401704 269686 401732 278038
rect 403912 271862 403940 278052
rect 404372 278038 405122 278066
rect 404176 273080 404228 273086
rect 404176 273022 404228 273028
rect 403900 271856 403952 271862
rect 403900 271798 403952 271804
rect 403624 270632 403676 270638
rect 403624 270574 403676 270580
rect 401692 269680 401744 269686
rect 401692 269622 401744 269628
rect 401692 269272 401744 269278
rect 401692 269214 401744 269220
rect 400614 264302 400904 264330
rect 401428 267706 401548 267734
rect 401428 264316 401456 267706
rect 401704 267442 401732 269214
rect 402244 268388 402296 268394
rect 402244 268330 402296 268336
rect 401692 267436 401744 267442
rect 401692 267378 401744 267384
rect 402256 264316 402284 268330
rect 403072 267436 403124 267442
rect 403072 267378 403124 267384
rect 403084 264316 403112 267378
rect 403636 266626 403664 270574
rect 403624 266620 403676 266626
rect 403624 266562 403676 266568
rect 404188 264330 404216 273022
rect 404372 270366 404400 278038
rect 405556 272944 405608 272950
rect 405556 272886 405608 272892
rect 404360 270360 404412 270366
rect 404360 270302 404412 270308
rect 404360 269680 404412 269686
rect 404360 269622 404412 269628
rect 404372 266762 404400 269622
rect 404728 267572 404780 267578
rect 404728 267514 404780 267520
rect 404360 266756 404412 266762
rect 404360 266698 404412 266704
rect 403926 264302 404216 264330
rect 404740 264316 404768 267514
rect 405568 264316 405596 272886
rect 406304 272678 406332 278052
rect 407132 278038 407514 278066
rect 406844 272808 406896 272814
rect 406844 272750 406896 272756
rect 406292 272672 406344 272678
rect 406292 272614 406344 272620
rect 406856 264330 406884 272750
rect 407132 269822 407160 278038
rect 408604 273970 408632 278052
rect 408788 278038 409814 278066
rect 408592 273964 408644 273970
rect 408592 273906 408644 273912
rect 407764 270904 407816 270910
rect 407764 270846 407816 270852
rect 407120 269816 407172 269822
rect 407120 269758 407172 269764
rect 407776 267170 407804 270846
rect 408788 270094 408816 278038
rect 410800 276004 410852 276010
rect 410800 275946 410852 275952
rect 409788 274644 409840 274650
rect 409788 274586 409840 274592
rect 409604 270224 409656 270230
rect 409604 270166 409656 270172
rect 408776 270088 408828 270094
rect 408776 270030 408828 270036
rect 408316 269408 408368 269414
rect 408316 269350 408368 269356
rect 408328 267714 408356 269350
rect 408316 267708 408368 267714
rect 408316 267650 408368 267656
rect 407764 267164 407816 267170
rect 407764 267106 407816 267112
rect 408040 266756 408092 266762
rect 408040 266698 408092 266704
rect 407212 266620 407264 266626
rect 407212 266562 407264 266568
rect 406410 264302 406884 264330
rect 407224 264316 407252 266562
rect 408052 264316 408080 266698
rect 408868 266416 408920 266422
rect 408868 266358 408920 266364
rect 408880 264316 408908 266358
rect 409616 264330 409644 270166
rect 409800 266422 409828 274586
rect 409788 266416 409840 266422
rect 409788 266358 409840 266364
rect 410812 264330 410840 275946
rect 410996 272542 411024 278052
rect 411272 278038 412206 278066
rect 412652 278038 413402 278066
rect 410984 272536 411036 272542
rect 410984 272478 411036 272484
rect 411272 269958 411300 278038
rect 412272 272672 412324 272678
rect 412272 272614 412324 272620
rect 411260 269952 411312 269958
rect 411260 269894 411312 269900
rect 412284 266422 412312 272614
rect 412456 270088 412508 270094
rect 412456 270030 412508 270036
rect 411352 266416 411404 266422
rect 411352 266358 411404 266364
rect 412272 266416 412324 266422
rect 412272 266358 412324 266364
rect 409616 264302 409722 264330
rect 410550 264302 410840 264330
rect 411364 264316 411392 266358
rect 412468 264330 412496 270030
rect 412652 269550 412680 278038
rect 413836 274508 413888 274514
rect 413836 274450 413888 274456
rect 412640 269544 412692 269550
rect 412640 269486 412692 269492
rect 413008 267164 413060 267170
rect 413008 267106 413060 267112
rect 412206 264302 412496 264330
rect 413020 264316 413048 267106
rect 413848 264316 413876 274450
rect 414584 271726 414612 278052
rect 415412 278038 415794 278066
rect 416792 278038 416898 278066
rect 414572 271720 414624 271726
rect 414572 271662 414624 271668
rect 414664 270768 414716 270774
rect 414664 270710 414716 270716
rect 414676 266626 414704 270710
rect 415032 270360 415084 270366
rect 415032 270302 415084 270308
rect 414664 266620 414716 266626
rect 414664 266562 414716 266568
rect 415044 264330 415072 270302
rect 415412 268938 415440 278038
rect 416412 275596 416464 275602
rect 416412 275538 416464 275544
rect 415400 268932 415452 268938
rect 415400 268874 415452 268880
rect 416228 268252 416280 268258
rect 416228 268194 416280 268200
rect 416240 267578 416268 268194
rect 416228 267572 416280 267578
rect 416228 267514 416280 267520
rect 416424 266422 416452 275538
rect 416596 272536 416648 272542
rect 416596 272478 416648 272484
rect 415492 266416 415544 266422
rect 415492 266358 415544 266364
rect 416412 266416 416464 266422
rect 416412 266358 416464 266364
rect 414690 264302 415072 264330
rect 415504 264316 415532 266358
rect 416608 264330 416636 272478
rect 416792 269278 416820 278038
rect 418080 272134 418108 278052
rect 418804 275324 418856 275330
rect 418804 275266 418856 275272
rect 418068 272128 418120 272134
rect 418068 272070 418120 272076
rect 417424 271040 417476 271046
rect 417424 270982 417476 270988
rect 417148 269816 417200 269822
rect 417148 269758 417200 269764
rect 416780 269272 416832 269278
rect 416780 269214 416832 269220
rect 416346 264302 416636 264330
rect 417160 264316 417188 269758
rect 417436 267306 417464 270982
rect 417424 267300 417476 267306
rect 417424 267242 417476 267248
rect 418816 266422 418844 275266
rect 419080 274372 419132 274378
rect 419080 274314 419132 274320
rect 417976 266416 418028 266422
rect 417976 266358 418028 266364
rect 418804 266416 418856 266422
rect 418804 266358 418856 266364
rect 417988 264316 418016 266358
rect 419092 264330 419120 274314
rect 419276 271454 419304 278052
rect 420472 275466 420500 278052
rect 420460 275460 420512 275466
rect 420460 275402 420512 275408
rect 420552 275052 420604 275058
rect 420552 274994 420604 275000
rect 420184 271584 420236 271590
rect 420184 271526 420236 271532
rect 419264 271448 419316 271454
rect 419264 271390 419316 271396
rect 419632 269952 419684 269958
rect 419632 269894 419684 269900
rect 418830 264302 419120 264330
rect 419644 264316 419672 269894
rect 420196 267034 420224 271526
rect 420564 267734 420592 274994
rect 421668 271726 421696 278052
rect 422312 278038 422878 278066
rect 423692 278038 423982 278066
rect 422116 273964 422168 273970
rect 422116 273906 422168 273912
rect 421656 271720 421708 271726
rect 421656 271662 421708 271668
rect 420472 267706 420592 267734
rect 420184 267028 420236 267034
rect 420184 266970 420236 266976
rect 420472 264316 420500 267706
rect 421288 267572 421340 267578
rect 421288 267514 421340 267520
rect 421300 264316 421328 267514
rect 422128 264316 422156 273906
rect 422312 268802 422340 278038
rect 423692 269686 423720 278038
rect 425164 274242 425192 278052
rect 425152 274236 425204 274242
rect 425152 274178 425204 274184
rect 425704 274236 425756 274242
rect 425704 274178 425756 274184
rect 423680 269680 423732 269686
rect 423680 269622 423732 269628
rect 423956 269680 424008 269686
rect 423956 269622 424008 269628
rect 422300 268796 422352 268802
rect 422300 268738 422352 268744
rect 422300 268116 422352 268122
rect 422300 268058 422352 268064
rect 422312 267442 422340 268058
rect 422944 267708 422996 267714
rect 422944 267650 422996 267656
rect 422300 267436 422352 267442
rect 422300 267378 422352 267384
rect 422956 264316 422984 267650
rect 423968 266762 423996 269622
rect 424600 269544 424652 269550
rect 424600 269486 424652 269492
rect 423956 266756 424008 266762
rect 423956 266698 424008 266704
rect 423772 266552 423824 266558
rect 423772 266494 423824 266500
rect 423784 264316 423812 266494
rect 424612 264316 424640 269486
rect 425716 266558 425744 274178
rect 426360 271454 426388 278052
rect 426544 278038 427570 278066
rect 426348 271448 426400 271454
rect 426348 271390 426400 271396
rect 426544 269414 426572 278038
rect 427084 275188 427136 275194
rect 427084 275130 427136 275136
rect 426532 269408 426584 269414
rect 426532 269350 426584 269356
rect 425704 266552 425756 266558
rect 425704 266494 425756 266500
rect 426256 266552 426308 266558
rect 426256 266494 426308 266500
rect 425428 266416 425480 266422
rect 425428 266358 425480 266364
rect 425440 264316 425468 266358
rect 426268 264316 426296 266494
rect 427096 266422 427124 275130
rect 428752 272270 428780 278052
rect 429212 278038 429962 278066
rect 428740 272264 428792 272270
rect 428740 272206 428792 272212
rect 428464 272128 428516 272134
rect 428464 272070 428516 272076
rect 427452 271040 427504 271046
rect 427452 270982 427504 270988
rect 427084 266416 427136 266422
rect 427084 266358 427136 266364
rect 427464 264330 427492 270982
rect 427912 266892 427964 266898
rect 427912 266834 427964 266840
rect 427110 264302 427492 264330
rect 427924 264316 427952 266834
rect 428476 266558 428504 272070
rect 429212 268666 429240 278038
rect 430212 275868 430264 275874
rect 430212 275810 430264 275816
rect 429200 268660 429252 268666
rect 429200 268602 429252 268608
rect 428740 267436 428792 267442
rect 428740 267378 428792 267384
rect 428464 266552 428516 266558
rect 428464 266494 428516 266500
rect 428752 264316 428780 267378
rect 429568 266416 429620 266422
rect 429568 266358 429620 266364
rect 429580 264316 429608 266358
rect 430224 264330 430252 275810
rect 430396 271720 430448 271726
rect 430396 271662 430448 271668
rect 430408 266422 430436 271662
rect 431144 271590 431172 278052
rect 431684 271992 431736 271998
rect 431684 271934 431736 271940
rect 431132 271584 431184 271590
rect 431132 271526 431184 271532
rect 430396 266416 430448 266422
rect 430396 266358 430448 266364
rect 431696 264330 431724 271934
rect 432248 271318 432276 278052
rect 433156 271856 433208 271862
rect 433156 271798 433208 271804
rect 432236 271312 432288 271318
rect 432236 271254 432288 271260
rect 432880 267300 432932 267306
rect 432880 267242 432932 267248
rect 432052 266416 432104 266422
rect 432052 266358 432104 266364
rect 430224 264302 430422 264330
rect 431250 264302 431724 264330
rect 432064 264316 432092 266358
rect 432892 264316 432920 267242
rect 433168 266422 433196 271798
rect 433444 270638 433472 278052
rect 434640 272406 434668 278052
rect 435640 275460 435692 275466
rect 435640 275402 435692 275408
rect 434628 272400 434680 272406
rect 434628 272342 434680 272348
rect 433432 270632 433484 270638
rect 433432 270574 433484 270580
rect 433708 268932 433760 268938
rect 433708 268874 433760 268880
rect 433156 266416 433208 266422
rect 433156 266358 433208 266364
rect 433720 264316 433748 268874
rect 434536 266756 434588 266762
rect 434536 266698 434588 266704
rect 434548 264316 434576 266698
rect 435652 264330 435680 275402
rect 435836 273834 435864 278052
rect 436112 278038 437046 278066
rect 437952 278038 438242 278066
rect 435824 273828 435876 273834
rect 435824 273770 435876 273776
rect 436112 268530 436140 278038
rect 437204 271584 437256 271590
rect 437204 271526 437256 271532
rect 436560 269068 436612 269074
rect 436560 269010 436612 269016
rect 436100 268524 436152 268530
rect 436100 268466 436152 268472
rect 436572 264330 436600 269010
rect 437216 264330 437244 271526
rect 437952 271182 437980 278038
rect 438124 273828 438176 273834
rect 438124 273770 438176 273776
rect 437940 271176 437992 271182
rect 437940 271118 437992 271124
rect 438136 267714 438164 273770
rect 439332 273222 439360 278052
rect 439320 273216 439372 273222
rect 439320 273158 439372 273164
rect 439964 271448 440016 271454
rect 439964 271390 440016 271396
rect 438676 268796 438728 268802
rect 438676 268738 438728 268744
rect 438124 267708 438176 267714
rect 438124 267650 438176 267656
rect 437848 266620 437900 266626
rect 437848 266562 437900 266568
rect 435390 264302 435680 264330
rect 436218 264302 436600 264330
rect 437046 264302 437244 264330
rect 437860 264316 437888 266562
rect 438688 264316 438716 268738
rect 439976 264330 440004 271390
rect 440528 270910 440556 278052
rect 441724 277394 441752 278052
rect 441632 277366 441752 277394
rect 440884 273556 440936 273562
rect 440884 273498 440936 273504
rect 440516 270904 440568 270910
rect 440516 270846 440568 270852
rect 440896 267578 440924 273498
rect 441344 271176 441396 271182
rect 441344 271118 441396 271124
rect 441160 268660 441212 268666
rect 441160 268602 441212 268608
rect 440884 267572 440936 267578
rect 440884 267514 440936 267520
rect 440332 266416 440384 266422
rect 440332 266358 440384 266364
rect 439530 264302 440004 264330
rect 440344 264316 440372 266358
rect 441172 264316 441200 268602
rect 441356 266422 441384 271118
rect 441632 270502 441660 277366
rect 442920 274106 442948 278052
rect 443104 278038 444130 278066
rect 444392 278038 445326 278066
rect 442908 274100 442960 274106
rect 442908 274042 442960 274048
rect 442908 271312 442960 271318
rect 442908 271254 442960 271260
rect 441620 270496 441672 270502
rect 441620 270438 441672 270444
rect 441620 269408 441672 269414
rect 441620 269350 441672 269356
rect 441632 267170 441660 269350
rect 441620 267164 441672 267170
rect 441620 267106 441672 267112
rect 442724 266892 442776 266898
rect 442724 266834 442776 266840
rect 441344 266416 441396 266422
rect 441344 266358 441396 266364
rect 441988 266416 442040 266422
rect 441988 266358 442040 266364
rect 442000 264316 442028 266358
rect 442736 264330 442764 266834
rect 442920 266422 442948 271254
rect 443104 268394 443132 278038
rect 444012 273216 444064 273222
rect 444012 273158 444064 273164
rect 443092 268388 443144 268394
rect 443092 268330 443144 268336
rect 442908 266416 442960 266422
rect 442908 266358 442960 266364
rect 444024 264330 444052 273158
rect 444392 268122 444420 278038
rect 445024 275732 445076 275738
rect 445024 275674 445076 275680
rect 445036 271182 445064 275674
rect 446508 273086 446536 278052
rect 447152 278038 447626 278066
rect 446496 273080 446548 273086
rect 446496 273022 446548 273028
rect 446864 273080 446916 273086
rect 446864 273022 446916 273028
rect 445024 271176 445076 271182
rect 445024 271118 445076 271124
rect 445668 271176 445720 271182
rect 445668 271118 445720 271124
rect 444380 268116 444432 268122
rect 444380 268058 444432 268064
rect 445300 267708 445352 267714
rect 445300 267650 445352 267656
rect 444472 266416 444524 266422
rect 444472 266358 444524 266364
rect 442736 264302 442842 264330
rect 443670 264302 444052 264330
rect 444484 264316 444512 266358
rect 445312 264316 445340 267650
rect 445680 266422 445708 271118
rect 446128 268524 446180 268530
rect 446128 268466 446180 268472
rect 445668 266416 445720 266422
rect 445668 266358 445720 266364
rect 446140 264316 446168 268466
rect 446876 264330 446904 273022
rect 447152 268258 447180 278038
rect 447784 273692 447836 273698
rect 447784 273634 447836 273640
rect 447140 268252 447192 268258
rect 447140 268194 447192 268200
rect 447796 267442 447824 273634
rect 448808 272950 448836 278052
rect 448796 272944 448848 272950
rect 448796 272886 448848 272892
rect 450004 272814 450032 278052
rect 450832 278038 451214 278066
rect 451384 278038 452410 278066
rect 449992 272808 450044 272814
rect 449992 272750 450044 272756
rect 449716 272400 449768 272406
rect 449716 272342 449768 272348
rect 449164 270904 449216 270910
rect 449164 270846 449216 270852
rect 448428 268116 448480 268122
rect 448428 268058 448480 268064
rect 447784 267436 447836 267442
rect 447784 267378 447836 267384
rect 448440 267170 448468 268058
rect 447140 267164 447192 267170
rect 447140 267106 447192 267112
rect 448428 267164 448480 267170
rect 448428 267106 448480 267112
rect 447152 266626 447180 267106
rect 449176 266762 449204 270846
rect 449164 266756 449216 266762
rect 449164 266698 449216 266704
rect 447140 266620 447192 266626
rect 447140 266562 447192 266568
rect 447784 266552 447836 266558
rect 447784 266494 447836 266500
rect 446876 264302 446982 264330
rect 447796 264316 447824 266494
rect 448612 266416 448664 266422
rect 448612 266358 448664 266364
rect 448624 264316 448652 266358
rect 449728 264330 449756 272342
rect 450544 272264 450596 272270
rect 450544 272206 450596 272212
rect 450268 267572 450320 267578
rect 450268 267514 450320 267520
rect 449466 264302 449756 264330
rect 450280 264316 450308 267514
rect 450556 266422 450584 272206
rect 450832 270774 450860 278038
rect 451188 274100 451240 274106
rect 451188 274042 451240 274048
rect 450820 270768 450872 270774
rect 450820 270710 450872 270716
rect 451200 267734 451228 274042
rect 451384 269686 451412 278038
rect 453592 274650 453620 278052
rect 454052 278038 454710 278066
rect 453580 274644 453632 274650
rect 453580 274586 453632 274592
rect 452292 272808 452344 272814
rect 452292 272750 452344 272756
rect 451372 269680 451424 269686
rect 451372 269622 451424 269628
rect 451108 267706 451228 267734
rect 450544 266416 450596 266422
rect 450544 266358 450596 266364
rect 451108 264316 451136 267706
rect 452304 264330 452332 272750
rect 453304 270632 453356 270638
rect 453304 270574 453356 270580
rect 453316 267306 453344 270574
rect 454052 270230 454080 278038
rect 455892 276010 455920 278052
rect 455880 276004 455932 276010
rect 455880 275946 455932 275952
rect 456064 276004 456116 276010
rect 456064 275946 456116 275952
rect 455328 272944 455380 272950
rect 455328 272886 455380 272892
rect 454040 270224 454092 270230
rect 454040 270166 454092 270172
rect 453580 269680 453632 269686
rect 453580 269622 453632 269628
rect 453304 267300 453356 267306
rect 453304 267242 453356 267248
rect 452752 267164 452804 267170
rect 452752 267106 452804 267112
rect 451950 264302 452332 264330
rect 452764 264316 452792 267106
rect 453592 264316 453620 269622
rect 455144 267164 455196 267170
rect 455144 267106 455196 267112
rect 454408 266416 454460 266422
rect 454408 266358 454460 266364
rect 454420 264316 454448 266358
rect 455156 264330 455184 267106
rect 455340 266422 455368 272886
rect 456076 266558 456104 275946
rect 457088 272678 457116 278052
rect 458284 277394 458312 278052
rect 458192 277366 458312 277394
rect 458468 278038 459494 278066
rect 457444 274644 457496 274650
rect 457444 274586 457496 274592
rect 457260 272944 457312 272950
rect 457260 272886 457312 272892
rect 457272 272678 457300 272886
rect 457076 272672 457128 272678
rect 457076 272614 457128 272620
rect 457260 272672 457312 272678
rect 457260 272614 457312 272620
rect 456432 270496 456484 270502
rect 456432 270438 456484 270444
rect 456064 266552 456116 266558
rect 456064 266494 456116 266500
rect 455328 266416 455380 266422
rect 455328 266358 455380 266364
rect 456444 264330 456472 270438
rect 457456 267034 457484 274586
rect 457996 272944 458048 272950
rect 457996 272886 458048 272892
rect 457444 267028 457496 267034
rect 457444 266970 457496 266976
rect 457720 266756 457772 266762
rect 457720 266698 457772 266704
rect 456892 266416 456944 266422
rect 456892 266358 456944 266364
rect 455156 264302 455262 264330
rect 456090 264302 456472 264330
rect 456904 264316 456932 266358
rect 457732 264316 457760 266698
rect 458008 266422 458036 272886
rect 458192 270094 458220 277366
rect 458180 270088 458232 270094
rect 458180 270030 458232 270036
rect 458468 269414 458496 278038
rect 460676 274514 460704 278052
rect 461228 278038 461886 278066
rect 460664 274508 460716 274514
rect 460664 274450 460716 274456
rect 460020 273352 460072 273358
rect 460020 273294 460072 273300
rect 460032 272678 460060 273294
rect 460020 272672 460072 272678
rect 460020 272614 460072 272620
rect 460204 272672 460256 272678
rect 460204 272614 460256 272620
rect 458824 270224 458876 270230
rect 458824 270166 458876 270172
rect 458456 269408 458508 269414
rect 458456 269350 458508 269356
rect 457996 266416 458048 266422
rect 457996 266358 458048 266364
rect 458836 264330 458864 270166
rect 460216 266422 460244 272614
rect 460848 272536 460900 272542
rect 460900 272484 460980 272490
rect 460848 272478 460980 272484
rect 460860 272462 460980 272478
rect 460952 272377 460980 272462
rect 460938 272368 460994 272377
rect 460938 272303 460994 272312
rect 461228 270366 461256 278038
rect 462976 275602 463004 278052
rect 463712 278038 464186 278066
rect 465092 278038 465382 278066
rect 462964 275596 463016 275602
rect 462964 275538 463016 275544
rect 463148 275596 463200 275602
rect 463148 275538 463200 275544
rect 463160 274666 463188 275538
rect 462976 274638 463188 274666
rect 461400 273352 461452 273358
rect 461400 273294 461452 273300
rect 461412 272542 461440 273294
rect 461400 272536 461452 272542
rect 461400 272478 461452 272484
rect 461216 270360 461268 270366
rect 461216 270302 461268 270308
rect 461400 270360 461452 270366
rect 461400 270302 461452 270308
rect 460480 267436 460532 267442
rect 460480 267378 460532 267384
rect 459376 266416 459428 266422
rect 459376 266358 459428 266364
rect 460204 266416 460256 266422
rect 460204 266358 460256 266364
rect 458574 264302 458864 264330
rect 459388 264316 459416 266358
rect 460492 264330 460520 267378
rect 461412 264330 461440 270302
rect 461860 268388 461912 268394
rect 461860 268330 461912 268336
rect 460230 264302 460520 264330
rect 461058 264302 461440 264330
rect 461872 264316 461900 268330
rect 462976 267306 463004 274638
rect 463240 274508 463292 274514
rect 463240 274450 463292 274456
rect 463252 267734 463280 274450
rect 463712 272377 463740 278038
rect 464802 272504 464858 272513
rect 464802 272439 464858 272448
rect 463698 272368 463754 272377
rect 463698 272303 463754 272312
rect 463516 270088 463568 270094
rect 463516 270030 463568 270036
rect 463160 267706 463280 267734
rect 462964 267300 463016 267306
rect 462964 267242 463016 267248
rect 463160 264330 463188 267706
rect 462714 264302 463188 264330
rect 463528 264316 463556 270030
rect 464816 264330 464844 272439
rect 465092 269822 465120 278038
rect 466564 275330 466592 278052
rect 466552 275324 466604 275330
rect 466552 275266 466604 275272
rect 467564 275324 467616 275330
rect 467564 275266 467616 275272
rect 465908 272944 465960 272950
rect 465908 272886 465960 272892
rect 466092 272944 466144 272950
rect 466092 272886 466144 272892
rect 465920 272678 465948 272886
rect 465908 272672 465960 272678
rect 465908 272614 465960 272620
rect 465540 272536 465592 272542
rect 466104 272490 466132 272886
rect 465592 272484 466132 272490
rect 465540 272478 466132 272484
rect 465552 272462 466132 272478
rect 465080 269816 465132 269822
rect 465080 269758 465132 269764
rect 466000 269816 466052 269822
rect 466000 269758 466052 269764
rect 465172 267300 465224 267306
rect 465172 267242 465224 267248
rect 464370 264302 464844 264330
rect 465184 264316 465212 267242
rect 466012 264316 466040 269758
rect 466828 265124 466880 265130
rect 466828 265066 466880 265072
rect 466840 264316 466868 265066
rect 467576 264330 467604 275266
rect 467760 274378 467788 278052
rect 468036 278038 468970 278066
rect 467748 274372 467800 274378
rect 467748 274314 467800 274320
rect 468036 269958 468064 278038
rect 470152 275058 470180 278052
rect 470140 275052 470192 275058
rect 470140 274994 470192 275000
rect 471256 273562 471284 278052
rect 471612 276140 471664 276146
rect 471612 276082 471664 276088
rect 471244 273556 471296 273562
rect 471244 273498 471296 273504
rect 470554 272536 470606 272542
rect 470692 272536 470744 272542
rect 470554 272478 470606 272484
rect 470690 272504 470692 272513
rect 470744 272504 470746 272513
rect 470566 272354 470594 272478
rect 470690 272439 470746 272448
rect 470566 272326 470640 272354
rect 470612 272218 470640 272326
rect 470612 272190 470824 272218
rect 470796 272134 470824 272190
rect 470554 272128 470606 272134
rect 470784 272128 470836 272134
rect 470606 272076 470640 272082
rect 470554 272070 470640 272076
rect 470784 272070 470836 272076
rect 470566 272054 470640 272070
rect 470612 271969 470640 272054
rect 470598 271960 470654 271969
rect 470598 271895 470654 271904
rect 468024 269952 468076 269958
rect 468024 269894 468076 269900
rect 468484 269952 468536 269958
rect 468484 269894 468536 269900
rect 467576 264302 467682 264330
rect 468496 264316 468524 269894
rect 470968 269408 471020 269414
rect 470968 269350 471020 269356
rect 470140 267028 470192 267034
rect 470140 266970 470192 266976
rect 469312 265260 469364 265266
rect 469312 265202 469364 265208
rect 469324 264316 469352 265202
rect 470152 264316 470180 266970
rect 470980 264316 471008 269350
rect 471624 264330 471652 276082
rect 472452 273970 472480 278052
rect 473084 274916 473136 274922
rect 473084 274858 473136 274864
rect 472440 273964 472492 273970
rect 472440 273906 472492 273912
rect 473096 264330 473124 274858
rect 473648 273834 473676 278052
rect 474844 274242 474872 278052
rect 475028 278038 476054 278066
rect 474832 274236 474884 274242
rect 474832 274178 474884 274184
rect 474648 273964 474700 273970
rect 474648 273906 474700 273912
rect 473636 273828 473688 273834
rect 473636 273770 473688 273776
rect 474280 269272 474332 269278
rect 474280 269214 474332 269220
rect 473452 266416 473504 266422
rect 473452 266358 473504 266364
rect 471624 264302 471822 264330
rect 472650 264302 473124 264330
rect 473464 264316 473492 266358
rect 474292 264316 474320 269214
rect 474660 266422 474688 273906
rect 475028 269550 475056 278038
rect 477040 276276 477092 276282
rect 477040 276218 477092 276224
rect 476764 274780 476816 274786
rect 476764 274722 476816 274728
rect 476028 273420 476080 273426
rect 476028 273362 476080 273368
rect 475016 269544 475068 269550
rect 475016 269486 475068 269492
rect 476040 267734 476068 273362
rect 475948 267706 476068 267734
rect 474648 266416 474700 266422
rect 474648 266358 474700 266364
rect 475108 266416 475160 266422
rect 475108 266358 475160 266364
rect 475120 264316 475148 266358
rect 475948 264316 475976 267706
rect 476776 266762 476804 274722
rect 476764 266756 476816 266762
rect 476764 266698 476816 266704
rect 477052 264330 477080 276218
rect 477236 275194 477264 278052
rect 478064 278038 478354 278066
rect 479168 278038 479550 278066
rect 477224 275188 477276 275194
rect 477224 275130 477276 275136
rect 478064 271969 478092 278038
rect 478696 273556 478748 273562
rect 478696 273498 478748 273504
rect 478050 271960 478106 271969
rect 478050 271895 478106 271904
rect 477592 265396 477644 265402
rect 477592 265338 477644 265344
rect 476790 264302 477080 264330
rect 477604 264316 477632 265338
rect 478708 264330 478736 273498
rect 479168 271046 479196 278038
rect 479984 276548 480036 276554
rect 479984 276490 480036 276496
rect 479522 271960 479578 271969
rect 479522 271895 479578 271904
rect 479156 271040 479208 271046
rect 479156 270982 479208 270988
rect 479536 266422 479564 271895
rect 479524 266416 479576 266422
rect 479524 266358 479576 266364
rect 479248 265532 479300 265538
rect 479248 265474 479300 265480
rect 478446 264302 478736 264330
rect 479260 264316 479288 265474
rect 479996 264330 480024 276490
rect 480732 274650 480760 278052
rect 481732 275460 481784 275466
rect 481732 275402 481784 275408
rect 481744 275194 481772 275402
rect 481732 275188 481784 275194
rect 481732 275130 481784 275136
rect 480720 274644 480772 274650
rect 480720 274586 480772 274592
rect 481364 273828 481416 273834
rect 481364 273770 481416 273776
rect 480536 271992 480588 271998
rect 480534 271960 480536 271969
rect 480588 271960 480590 271969
rect 480534 271895 480590 271904
rect 480168 271856 480220 271862
rect 480220 271804 480300 271810
rect 480168 271798 480300 271804
rect 480180 271782 480300 271798
rect 480272 270774 480300 271782
rect 480260 270768 480312 270774
rect 480260 270710 480312 270716
rect 481376 264330 481404 273770
rect 481928 273698 481956 278052
rect 483124 277394 483152 278052
rect 483124 277366 483244 277394
rect 482836 276412 482888 276418
rect 482836 276354 482888 276360
rect 481916 273692 481968 273698
rect 481916 273634 481968 273640
rect 482848 266422 482876 276354
rect 483216 271726 483244 277366
rect 484320 275874 484348 278052
rect 484688 278038 485530 278066
rect 484308 275868 484360 275874
rect 484308 275810 484360 275816
rect 483664 275460 483716 275466
rect 483664 275402 483716 275408
rect 483676 274514 483704 275402
rect 483664 274508 483716 274514
rect 483664 274450 483716 274456
rect 484216 273692 484268 273698
rect 484216 273634 484268 273640
rect 483204 271720 483256 271726
rect 483204 271662 483256 271668
rect 484228 266422 484256 273634
rect 484688 271862 484716 278038
rect 485412 272128 485464 272134
rect 485412 272070 485464 272076
rect 485044 271992 485096 271998
rect 485424 271946 485452 272070
rect 485096 271940 485452 271946
rect 485044 271934 485452 271940
rect 485056 271918 485452 271934
rect 484676 271856 484728 271862
rect 484676 271798 484728 271804
rect 485044 271040 485096 271046
rect 485044 270982 485096 270988
rect 485056 266898 485084 270982
rect 486620 270774 486648 278052
rect 486792 274644 486844 274650
rect 486792 274586 486844 274592
rect 486608 270768 486660 270774
rect 486608 270710 486660 270716
rect 485044 266892 485096 266898
rect 485044 266834 485096 266840
rect 485044 266756 485096 266762
rect 485044 266698 485096 266704
rect 481732 266416 481784 266422
rect 481732 266358 481784 266364
rect 482836 266416 482888 266422
rect 482836 266358 482888 266364
rect 483388 266416 483440 266422
rect 483388 266358 483440 266364
rect 484216 266416 484268 266422
rect 484216 266358 484268 266364
rect 479996 264302 480102 264330
rect 480930 264302 481404 264330
rect 481744 264316 481772 266358
rect 482560 266076 482612 266082
rect 482560 266018 482612 266024
rect 482572 264316 482600 266018
rect 483400 264316 483428 266358
rect 484216 266212 484268 266218
rect 484216 266154 484268 266160
rect 484228 264316 484256 266154
rect 485056 264316 485084 266698
rect 486804 266422 486832 274586
rect 486976 270768 487028 270774
rect 486976 270710 487028 270716
rect 485872 266416 485924 266422
rect 485872 266358 485924 266364
rect 486792 266416 486844 266422
rect 486792 266358 486844 266364
rect 485884 264316 485912 266358
rect 486988 264330 487016 270710
rect 487816 270638 487844 278052
rect 488552 278038 489026 278066
rect 487988 277228 488040 277234
rect 487988 277170 488040 277176
rect 487804 270632 487856 270638
rect 487804 270574 487856 270580
rect 487160 266348 487212 266354
rect 487160 266290 487212 266296
rect 487172 266082 487200 266290
rect 487160 266076 487212 266082
rect 487160 266018 487212 266024
rect 488000 264330 488028 277170
rect 488356 274508 488408 274514
rect 488356 274450 488408 274456
rect 486726 264302 487016 264330
rect 487554 264302 488028 264330
rect 488368 264316 488396 274450
rect 488552 268938 488580 278038
rect 490208 270910 490236 278052
rect 490564 275868 490616 275874
rect 490564 275810 490616 275816
rect 490196 270904 490248 270910
rect 490196 270846 490248 270852
rect 489644 270632 489696 270638
rect 489644 270574 489696 270580
rect 488540 268932 488592 268938
rect 488540 268874 488592 268880
rect 489656 264330 489684 270574
rect 490576 267714 490604 275810
rect 491404 275194 491432 278052
rect 491680 278038 492614 278066
rect 491392 275188 491444 275194
rect 491392 275130 491444 275136
rect 491680 269074 491708 278038
rect 493704 271590 493732 278052
rect 494072 278038 494914 278066
rect 495452 278038 496110 278066
rect 493692 271584 493744 271590
rect 493692 271526 493744 271532
rect 492588 270904 492640 270910
rect 492588 270846 492640 270852
rect 491668 269068 491720 269074
rect 491668 269010 491720 269016
rect 490840 267980 490892 267986
rect 490840 267922 490892 267928
rect 490564 267708 490616 267714
rect 490564 267650 490616 267656
rect 490012 266756 490064 266762
rect 490012 266698 490064 266704
rect 489210 264302 489684 264330
rect 490024 264316 490052 266698
rect 490852 264316 490880 267922
rect 492600 266490 492628 270846
rect 493324 268252 493376 268258
rect 493324 268194 493376 268200
rect 491668 266484 491720 266490
rect 491668 266426 491720 266432
rect 492588 266484 492640 266490
rect 492588 266426 492640 266432
rect 491680 264316 491708 266426
rect 492496 266076 492548 266082
rect 492496 266018 492548 266024
rect 492508 264316 492536 266018
rect 493336 264316 493364 268194
rect 494072 268122 494100 278038
rect 494704 271856 494756 271862
rect 494704 271798 494756 271804
rect 494716 271046 494744 271798
rect 494704 271040 494756 271046
rect 494704 270982 494756 270988
rect 495072 271040 495124 271046
rect 495072 270982 495124 270988
rect 494060 268116 494112 268122
rect 494060 268058 494112 268064
rect 495084 266490 495112 270982
rect 495256 269544 495308 269550
rect 495256 269486 495308 269492
rect 494152 266484 494204 266490
rect 494152 266426 494204 266432
rect 495072 266484 495124 266490
rect 495072 266426 495124 266432
rect 494164 264316 494192 266426
rect 495268 264330 495296 269486
rect 495452 268802 495480 278038
rect 497292 271590 497320 278052
rect 497924 277092 497976 277098
rect 497924 277034 497976 277040
rect 497280 271584 497332 271590
rect 497280 271526 497332 271532
rect 496544 271448 496596 271454
rect 496544 271390 496596 271396
rect 495808 269068 495860 269074
rect 495808 269010 495860 269016
rect 495440 268796 495492 268802
rect 495440 268738 495492 268744
rect 495006 264302 495296 264330
rect 495820 264316 495848 269010
rect 496556 264330 496584 271390
rect 497936 264330 497964 277034
rect 498488 275738 498516 278052
rect 499684 277394 499712 278052
rect 499592 277366 499712 277394
rect 498476 275732 498528 275738
rect 498476 275674 498528 275680
rect 498844 275732 498896 275738
rect 498844 275674 498896 275680
rect 498292 268932 498344 268938
rect 498292 268874 498344 268880
rect 496556 264302 496662 264330
rect 497490 264302 497964 264330
rect 498304 264316 498332 268874
rect 498856 267578 498884 275674
rect 499304 271720 499356 271726
rect 499304 271662 499356 271668
rect 498844 267572 498896 267578
rect 498844 267514 498896 267520
rect 499316 264330 499344 271662
rect 499592 268666 499620 277366
rect 500880 271318 500908 278052
rect 501432 278038 501998 278066
rect 501432 271862 501460 278038
rect 503180 273222 503208 278052
rect 504008 278038 504390 278066
rect 503444 275052 503496 275058
rect 503444 274994 503496 275000
rect 503168 273216 503220 273222
rect 503168 273158 503220 273164
rect 501602 271960 501658 271969
rect 501602 271895 501658 271904
rect 501420 271856 501472 271862
rect 501420 271798 501472 271804
rect 500868 271312 500920 271318
rect 500868 271254 500920 271260
rect 500776 268796 500828 268802
rect 500776 268738 500828 268744
rect 499580 268660 499632 268666
rect 499580 268602 499632 268608
rect 499948 266892 500000 266898
rect 499948 266834 500000 266840
rect 499146 264302 499344 264330
rect 499960 264316 499988 266834
rect 500788 264316 500816 268738
rect 501616 266626 501644 271895
rect 501972 271584 502024 271590
rect 501972 271526 502024 271532
rect 501604 266620 501656 266626
rect 501604 266562 501656 266568
rect 501984 264330 502012 271526
rect 503260 268660 503312 268666
rect 503260 268602 503312 268608
rect 502432 266484 502484 266490
rect 502432 266426 502484 266432
rect 501630 264302 502012 264330
rect 502444 264316 502472 266426
rect 503272 264316 503300 268602
rect 503456 266490 503484 274994
rect 504008 271182 504036 278038
rect 505572 275874 505600 278052
rect 506492 278038 506782 278066
rect 505560 275868 505612 275874
rect 505560 275810 505612 275816
rect 506204 274372 506256 274378
rect 506204 274314 506256 274320
rect 504180 273216 504232 273222
rect 504180 273158 504232 273164
rect 504192 272406 504220 273158
rect 504180 272400 504232 272406
rect 504180 272342 504232 272348
rect 504364 272400 504416 272406
rect 504364 272342 504416 272348
rect 504376 271998 504404 272342
rect 504364 271992 504416 271998
rect 504548 271992 504600 271998
rect 504364 271934 504416 271940
rect 504546 271960 504548 271969
rect 504600 271960 504602 271969
rect 504546 271895 504602 271904
rect 504364 271856 504416 271862
rect 504364 271798 504416 271804
rect 504376 271454 504404 271798
rect 504364 271448 504416 271454
rect 504364 271390 504416 271396
rect 505008 271448 505060 271454
rect 505008 271390 505060 271396
rect 503996 271176 504048 271182
rect 503996 271118 504048 271124
rect 504824 266620 504876 266626
rect 504824 266562 504876 266568
rect 503444 266484 503496 266490
rect 503444 266426 503496 266432
rect 504088 266484 504140 266490
rect 504088 266426 504140 266432
rect 504100 264316 504128 266426
rect 504836 264330 504864 266562
rect 505020 266490 505048 271390
rect 505008 266484 505060 266490
rect 505008 266426 505060 266432
rect 506216 264330 506244 274314
rect 506492 268530 506520 278038
rect 507492 275188 507544 275194
rect 507492 275130 507544 275136
rect 506480 268524 506532 268530
rect 506480 268466 506532 268472
rect 507504 267734 507532 275130
rect 507964 273086 507992 278052
rect 509068 276010 509096 278052
rect 509056 276004 509108 276010
rect 509056 275946 509108 275952
rect 507952 273080 508004 273086
rect 507952 273022 508004 273028
rect 510264 272270 510292 278052
rect 511460 273222 511488 278052
rect 511632 276956 511684 276962
rect 511632 276898 511684 276904
rect 511448 273216 511500 273222
rect 511448 273158 511500 273164
rect 510252 272264 510304 272270
rect 510252 272206 510304 272212
rect 510436 272264 510488 272270
rect 510436 272206 510488 272212
rect 507676 271312 507728 271318
rect 507676 271254 507728 271260
rect 507412 267706 507532 267734
rect 506572 266484 506624 266490
rect 506572 266426 506624 266432
rect 504836 264302 504942 264330
rect 505770 264302 506244 264330
rect 506584 264316 506612 266426
rect 507412 264316 507440 267706
rect 507688 266490 507716 271254
rect 510448 270450 510476 272206
rect 509712 270422 510476 270450
rect 509238 269920 509294 269929
rect 509238 269855 509294 269864
rect 509252 269686 509280 269855
rect 509240 269680 509292 269686
rect 509240 269622 509292 269628
rect 509146 269512 509202 269521
rect 509146 269447 509202 269456
rect 508228 268524 508280 268530
rect 508228 268466 508280 268472
rect 507860 266892 507912 266898
rect 507860 266834 507912 266840
rect 507872 266490 507900 266834
rect 507676 266484 507728 266490
rect 507676 266426 507728 266432
rect 507860 266484 507912 266490
rect 507860 266426 507912 266432
rect 508240 264316 508268 268466
rect 509160 267734 509188 269447
rect 509068 267706 509188 267734
rect 509068 264316 509096 267706
rect 509712 266762 509740 270422
rect 509884 269544 509936 269550
rect 509882 269512 509884 269521
rect 509936 269512 509938 269521
rect 509882 269447 509938 269456
rect 511644 267734 511672 276898
rect 512656 275738 512684 278052
rect 513196 276004 513248 276010
rect 513196 275946 513248 275952
rect 512644 275732 512696 275738
rect 512644 275674 512696 275680
rect 511816 274236 511868 274242
rect 511816 274178 511868 274184
rect 509884 267708 509936 267714
rect 509884 267650 509936 267656
rect 511552 267706 511672 267734
rect 509700 266756 509752 266762
rect 509700 266698 509752 266704
rect 509896 264316 509924 267650
rect 510712 266756 510764 266762
rect 510712 266698 510764 266704
rect 510724 264316 510752 266698
rect 511552 264316 511580 267706
rect 511828 266762 511856 274178
rect 513208 266762 513236 275946
rect 513852 274106 513880 278052
rect 514484 276820 514536 276826
rect 514484 276762 514536 276768
rect 513840 274100 513892 274106
rect 513840 274042 513892 274048
rect 513748 272808 513800 272814
rect 513748 272750 513800 272756
rect 513760 272406 513788 272750
rect 513748 272400 513800 272406
rect 513748 272342 513800 272348
rect 511816 266756 511868 266762
rect 511816 266698 511868 266704
rect 512368 266756 512420 266762
rect 512368 266698 512420 266704
rect 513196 266756 513248 266762
rect 513196 266698 513248 266704
rect 512380 264316 512408 266698
rect 513196 265940 513248 265946
rect 513196 265882 513248 265888
rect 513208 264316 513236 265882
rect 514496 264330 514524 276762
rect 515048 272950 515076 278052
rect 516244 275602 516272 278052
rect 516428 278038 517362 278066
rect 516232 275596 516284 275602
rect 516232 275538 516284 275544
rect 515404 273216 515456 273222
rect 515404 273158 515456 273164
rect 515036 272944 515088 272950
rect 515036 272886 515088 272892
rect 514852 267572 514904 267578
rect 514852 267514 514904 267520
rect 514050 264302 514524 264330
rect 514864 264316 514892 267514
rect 515416 267170 515444 273158
rect 516428 269929 516456 278038
rect 518348 276684 518400 276690
rect 518348 276626 518400 276632
rect 516784 275596 516836 275602
rect 516784 275538 516836 275544
rect 516414 269920 516470 269929
rect 516414 269855 516470 269864
rect 516796 267442 516824 275538
rect 517428 272400 517480 272406
rect 517428 272342 517480 272348
rect 516784 267436 516836 267442
rect 516784 267378 516836 267384
rect 515404 267164 515456 267170
rect 515404 267106 515456 267112
rect 517244 267164 517296 267170
rect 517244 267106 517296 267112
rect 516508 266756 516560 266762
rect 516508 266698 516560 266704
rect 515680 265804 515732 265810
rect 515680 265746 515732 265752
rect 515692 264316 515720 265746
rect 516520 264316 516548 266698
rect 517256 264330 517284 267106
rect 517440 266762 517468 272342
rect 517428 266756 517480 266762
rect 517428 266698 517480 266704
rect 518360 264330 518388 276626
rect 518544 273086 518572 278052
rect 519740 273222 519768 278052
rect 520292 278038 520950 278066
rect 519728 273216 519780 273222
rect 519728 273158 519780 273164
rect 518532 273080 518584 273086
rect 518532 273022 518584 273028
rect 518716 273080 518768 273086
rect 518716 273022 518768 273028
rect 518728 272270 518756 273022
rect 518716 272264 518768 272270
rect 518716 272206 518768 272212
rect 520096 272264 520148 272270
rect 520096 272206 520148 272212
rect 519820 267436 519872 267442
rect 519820 267378 519872 267384
rect 518992 266756 519044 266762
rect 518992 266698 519044 266704
rect 517256 264302 517362 264330
rect 518190 264302 518388 264330
rect 519004 264316 519032 266698
rect 519832 264316 519860 267378
rect 520108 266762 520136 272206
rect 520292 270502 520320 278038
rect 521476 273216 521528 273222
rect 521476 273158 521528 273164
rect 520280 270496 520332 270502
rect 520280 270438 520332 270444
rect 520096 266756 520148 266762
rect 520096 266698 520148 266704
rect 520648 265668 520700 265674
rect 520648 265610 520700 265616
rect 520660 264316 520688 265610
rect 521488 264316 521516 273158
rect 522132 272678 522160 278052
rect 522764 275868 522816 275874
rect 522764 275810 522816 275816
rect 522120 272672 522172 272678
rect 522120 272614 522172 272620
rect 522776 264330 522804 275810
rect 523328 274786 523356 278052
rect 524432 278038 524538 278066
rect 523316 274780 523368 274786
rect 523316 274722 523368 274728
rect 523684 274780 523736 274786
rect 523684 274722 523736 274728
rect 523132 270496 523184 270502
rect 523132 270438 523184 270444
rect 522330 264302 522804 264330
rect 523144 264316 523172 270438
rect 523696 267306 523724 274722
rect 524052 271176 524104 271182
rect 524052 271118 524104 271124
rect 524064 267734 524092 271118
rect 524432 270230 524460 278038
rect 525628 272814 525656 278052
rect 526824 275602 526852 278052
rect 527192 278038 528034 278066
rect 528572 278038 529230 278066
rect 526812 275596 526864 275602
rect 526812 275538 526864 275544
rect 525616 272808 525668 272814
rect 525616 272750 525668 272756
rect 526812 272672 526864 272678
rect 526812 272614 526864 272620
rect 525616 270360 525668 270366
rect 525616 270302 525668 270308
rect 524420 270224 524472 270230
rect 524420 270166 524472 270172
rect 523972 267706 524092 267734
rect 523684 267300 523736 267306
rect 523684 267242 523736 267248
rect 523972 264316 524000 267706
rect 524788 267300 524840 267306
rect 524788 267242 524840 267248
rect 524800 264316 524828 267242
rect 525628 264316 525656 270302
rect 526824 264330 526852 272614
rect 527192 270230 527220 278038
rect 528192 275732 528244 275738
rect 528192 275674 528244 275680
rect 527180 270224 527232 270230
rect 527180 270166 527232 270172
rect 527180 268116 527232 268122
rect 527180 268058 527232 268064
rect 527192 267170 527220 268058
rect 527180 267164 527232 267170
rect 527180 267106 527232 267112
rect 528204 266762 528232 275674
rect 528376 270224 528428 270230
rect 528376 270166 528428 270172
rect 527272 266756 527324 266762
rect 527272 266698 527324 266704
rect 528192 266756 528244 266762
rect 528192 266698 528244 266704
rect 526470 264302 526852 264330
rect 527284 264316 527312 266698
rect 528388 264330 528416 270166
rect 528572 268394 528600 278038
rect 530412 275466 530440 278052
rect 531332 278038 531622 278066
rect 530400 275460 530452 275466
rect 530400 275402 530452 275408
rect 529848 272808 529900 272814
rect 529848 272750 529900 272756
rect 528560 268388 528612 268394
rect 528560 268330 528612 268336
rect 529664 267164 529716 267170
rect 529664 267106 529716 267112
rect 528928 266756 528980 266762
rect 528928 266698 528980 266704
rect 528126 264302 528416 264330
rect 528940 264316 528968 266698
rect 529676 264330 529704 267106
rect 529860 266762 529888 272750
rect 531332 270178 531360 278038
rect 532332 275596 532384 275602
rect 532332 275538 532384 275544
rect 532344 270314 532372 275538
rect 532516 272944 532568 272950
rect 532516 272886 532568 272892
rect 532344 270286 532464 270314
rect 530780 270150 531360 270178
rect 532238 270192 532294 270201
rect 530780 270094 530808 270150
rect 532238 270127 532294 270136
rect 530768 270088 530820 270094
rect 530768 270030 530820 270036
rect 530952 270088 531004 270094
rect 530952 270030 531004 270036
rect 529848 266756 529900 266762
rect 529848 266698 529900 266704
rect 530964 264330 530992 270030
rect 532252 269822 532280 270127
rect 532240 269816 532292 269822
rect 532240 269758 532292 269764
rect 531412 266756 531464 266762
rect 531412 266698 531464 266704
rect 529676 264302 529782 264330
rect 530610 264302 530992 264330
rect 531424 264316 531452 266698
rect 532436 264330 532464 270286
rect 532528 267734 532556 272886
rect 532712 272542 532740 278052
rect 533908 274786 533936 278052
rect 534092 278038 535118 278066
rect 535748 278038 536314 278066
rect 533896 274780 533948 274786
rect 533896 274722 533948 274728
rect 532884 272808 532936 272814
rect 532884 272750 532936 272756
rect 533712 272808 533764 272814
rect 533712 272750 533764 272756
rect 532896 272542 532924 272750
rect 532700 272536 532752 272542
rect 532700 272478 532752 272484
rect 532884 272536 532936 272542
rect 532884 272478 532936 272484
rect 532988 270558 533384 270586
rect 532792 270496 532844 270502
rect 532792 270438 532844 270444
rect 532804 269686 532832 270438
rect 532988 270094 533016 270558
rect 533356 270450 533384 270558
rect 533356 270422 533568 270450
rect 533540 270366 533568 270422
rect 533528 270360 533580 270366
rect 533528 270302 533580 270308
rect 533252 270224 533304 270230
rect 533528 270224 533580 270230
rect 533304 270184 533528 270212
rect 533252 270166 533304 270172
rect 533528 270166 533580 270172
rect 532976 270088 533028 270094
rect 532976 270030 533028 270036
rect 532792 269680 532844 269686
rect 532792 269622 532844 269628
rect 532528 267706 532648 267734
rect 532620 266762 532648 267706
rect 532608 266756 532660 266762
rect 532608 266698 532660 266704
rect 533068 266756 533120 266762
rect 533068 266698 533120 266704
rect 532266 264302 532464 264330
rect 533080 264316 533108 266698
rect 533724 264330 533752 272750
rect 534092 270201 534120 278038
rect 534724 274780 534776 274786
rect 534724 274722 534776 274728
rect 534078 270192 534134 270201
rect 534078 270127 534134 270136
rect 533988 269952 534040 269958
rect 533988 269894 534040 269900
rect 534000 266762 534028 269894
rect 534736 267034 534764 274722
rect 534724 267028 534776 267034
rect 534724 266970 534776 266976
rect 535552 267028 535604 267034
rect 535552 266970 535604 266976
rect 534724 266892 534776 266898
rect 534724 266834 534776 266840
rect 533988 266756 534040 266762
rect 533988 266698 534040 266704
rect 533724 264302 533922 264330
rect 534736 264316 534764 266834
rect 535564 264316 535592 266970
rect 535748 265130 535776 278038
rect 537496 275330 537524 278052
rect 538508 278038 538706 278066
rect 537668 275460 537720 275466
rect 537668 275402 537720 275408
rect 537484 275324 537536 275330
rect 537484 275266 537536 275272
rect 536748 274100 536800 274106
rect 536748 274042 536800 274048
rect 536562 272504 536618 272513
rect 536562 272439 536618 272448
rect 535736 265124 535788 265130
rect 535736 265066 535788 265072
rect 536576 264330 536604 272439
rect 536760 267034 536788 274042
rect 536748 267028 536800 267034
rect 536748 266970 536800 266976
rect 537680 264330 537708 275402
rect 538508 273254 538536 278038
rect 539888 277394 539916 278052
rect 539888 277366 540008 277394
rect 539322 274000 539378 274009
rect 539322 273935 539378 273944
rect 538324 273226 538536 273254
rect 538324 270094 538352 273226
rect 539048 272944 539100 272950
rect 538508 272892 539048 272898
rect 538508 272886 539100 272892
rect 538508 272870 539088 272886
rect 538508 272542 538536 272870
rect 538680 272808 538732 272814
rect 538680 272750 538732 272756
rect 538692 272542 538720 272750
rect 538496 272536 538548 272542
rect 538496 272478 538548 272484
rect 538680 272536 538732 272542
rect 538680 272478 538732 272484
rect 538312 270088 538364 270094
rect 538312 270030 538364 270036
rect 539048 269952 539100 269958
rect 538692 269912 539048 269940
rect 538034 269784 538090 269793
rect 538034 269719 538090 269728
rect 536406 264302 536604 264330
rect 537234 264302 537708 264330
rect 538048 264316 538076 269719
rect 538692 269414 538720 269912
rect 539048 269894 539100 269900
rect 538864 269816 538916 269822
rect 538864 269758 538916 269764
rect 538876 269414 538904 269758
rect 538680 269408 538732 269414
rect 538680 269350 538732 269356
rect 538864 269408 538916 269414
rect 538864 269350 538916 269356
rect 539336 264330 539364 273935
rect 539692 267028 539744 267034
rect 539692 266970 539744 266976
rect 538890 264302 539364 264330
rect 539704 264316 539732 266970
rect 539980 265266 540008 277366
rect 540992 274786 541020 278052
rect 541544 278038 542202 278066
rect 540980 274780 541032 274786
rect 540980 274722 541032 274728
rect 541544 269958 541572 278038
rect 543384 276146 543412 278052
rect 543372 276140 543424 276146
rect 543372 276082 543424 276088
rect 542268 275324 542320 275330
rect 542268 275266 542320 275272
rect 542280 273254 542308 275266
rect 544580 274922 544608 278052
rect 544568 274916 544620 274922
rect 544568 274858 544620 274864
rect 545776 273970 545804 278052
rect 546512 278038 546986 278066
rect 547892 278038 548090 278066
rect 545946 274000 546002 274009
rect 545764 273964 545816 273970
rect 545946 273935 545948 273944
rect 545764 273906 545816 273912
rect 546000 273935 546002 273944
rect 545948 273906 546000 273912
rect 542188 273226 542308 273254
rect 541532 269952 541584 269958
rect 541532 269894 541584 269900
rect 540520 269816 540572 269822
rect 540520 269758 540572 269764
rect 539968 265260 540020 265266
rect 539968 265202 540020 265208
rect 540532 264316 540560 269758
rect 541348 268388 541400 268394
rect 541348 268330 541400 268336
rect 541360 264316 541388 268330
rect 542188 264316 542216 273226
rect 542452 269816 542504 269822
rect 542450 269784 542452 269793
rect 542504 269784 542506 269793
rect 542450 269719 542506 269728
rect 546512 269278 546540 278038
rect 547694 272504 547750 272513
rect 547694 272439 547750 272448
rect 547708 272134 547736 272439
rect 547512 272128 547564 272134
rect 547510 272096 547512 272105
rect 547696 272128 547748 272134
rect 547564 272096 547566 272105
rect 547892 272105 547920 278038
rect 549272 273426 549300 278052
rect 550468 276282 550496 278052
rect 550652 278038 551678 278066
rect 550456 276276 550508 276282
rect 550456 276218 550508 276224
rect 549260 273420 549312 273426
rect 549260 273362 549312 273368
rect 549904 273420 549956 273426
rect 549904 273362 549956 273368
rect 547696 272070 547748 272076
rect 547878 272096 547934 272105
rect 547510 272031 547566 272040
rect 547878 272031 547934 272040
rect 546500 269272 546552 269278
rect 546500 269214 546552 269220
rect 543004 266756 543056 266762
rect 543004 266698 543056 266704
rect 543016 264316 543044 266698
rect 549916 266490 549944 273362
rect 549904 266484 549956 266490
rect 549904 266426 549956 266432
rect 550652 265402 550680 278038
rect 552860 273562 552888 278052
rect 553412 278038 554070 278066
rect 552848 273556 552900 273562
rect 552848 273498 552900 273504
rect 553412 265538 553440 278038
rect 555252 276554 555280 278052
rect 555240 276548 555292 276554
rect 555240 276490 555292 276496
rect 556356 273834 556384 278052
rect 557552 276418 557580 278052
rect 557736 278038 558762 278066
rect 557540 276412 557592 276418
rect 557540 276354 557592 276360
rect 556344 273828 556396 273834
rect 556344 273770 556396 273776
rect 556804 273828 556856 273834
rect 556804 273770 556856 273776
rect 556816 266626 556844 273770
rect 556804 266620 556856 266626
rect 556804 266562 556856 266568
rect 557736 266354 557764 278038
rect 559944 273698 559972 278052
rect 560312 278038 561154 278066
rect 559932 273692 559984 273698
rect 559932 273634 559984 273640
rect 557724 266348 557776 266354
rect 557724 266290 557776 266296
rect 560312 266218 560340 278038
rect 562336 271998 562364 278052
rect 563440 274650 563468 278052
rect 563428 274644 563480 274650
rect 563428 274586 563480 274592
rect 562324 271992 562376 271998
rect 562324 271934 562376 271940
rect 564636 270774 564664 278052
rect 565832 277234 565860 278052
rect 565820 277228 565872 277234
rect 565820 277170 565872 277176
rect 567028 274514 567056 278052
rect 567016 274508 567068 274514
rect 567016 274450 567068 274456
rect 564624 270768 564676 270774
rect 564624 270710 564676 270716
rect 567844 270768 567896 270774
rect 567844 270710 567896 270716
rect 567856 267714 567884 270710
rect 568224 270638 568252 278052
rect 569420 273086 569448 278052
rect 569972 278038 570630 278066
rect 569408 273080 569460 273086
rect 569408 273022 569460 273028
rect 568212 270632 568264 270638
rect 568212 270574 568264 270580
rect 569972 267986 570000 278038
rect 571720 270910 571748 278052
rect 572732 278038 572930 278066
rect 571708 270904 571760 270910
rect 571708 270846 571760 270852
rect 569960 267980 570012 267986
rect 569960 267922 570012 267928
rect 567844 267708 567896 267714
rect 567844 267650 567896 267656
rect 560300 266212 560352 266218
rect 560300 266154 560352 266160
rect 572732 266082 572760 278038
rect 574112 268258 574140 278052
rect 575308 271046 575336 278052
rect 575492 278038 576518 278066
rect 576872 278038 577714 278066
rect 578528 278038 578910 278066
rect 575296 271040 575348 271046
rect 575296 270982 575348 270988
rect 575492 269414 575520 278038
rect 575480 269408 575532 269414
rect 575480 269350 575532 269356
rect 576872 269074 576900 278038
rect 578528 271862 578556 278038
rect 580000 277098 580028 278052
rect 581012 278038 581210 278066
rect 579988 277092 580040 277098
rect 579988 277034 580040 277040
rect 578516 271856 578568 271862
rect 578516 271798 578568 271804
rect 578884 271856 578936 271862
rect 578884 271798 578936 271804
rect 576860 269068 576912 269074
rect 576860 269010 576912 269016
rect 574100 268252 574152 268258
rect 574100 268194 574152 268200
rect 578896 267578 578924 271798
rect 581012 268938 581040 278038
rect 582392 271726 582420 278052
rect 583588 273426 583616 278052
rect 583772 278038 584798 278066
rect 583576 273420 583628 273426
rect 583576 273362 583628 273368
rect 582380 271720 582432 271726
rect 582380 271662 582432 271668
rect 583024 271720 583076 271726
rect 583024 271662 583076 271668
rect 581000 268932 581052 268938
rect 581000 268874 581052 268880
rect 578884 267572 578936 267578
rect 578884 267514 578936 267520
rect 583036 267442 583064 271662
rect 583772 268802 583800 278038
rect 585980 271590 586008 278052
rect 587084 275058 587112 278052
rect 587912 278038 588294 278066
rect 587072 275052 587124 275058
rect 587072 274994 587124 275000
rect 585968 271584 586020 271590
rect 585968 271526 586020 271532
rect 583760 268796 583812 268802
rect 583760 268738 583812 268744
rect 587912 268666 587940 278038
rect 589476 271454 589504 278052
rect 590672 273834 590700 278052
rect 591868 274378 591896 278052
rect 591856 274372 591908 274378
rect 591856 274314 591908 274320
rect 590660 273828 590712 273834
rect 590660 273770 590712 273776
rect 589464 271448 589516 271454
rect 589464 271390 589516 271396
rect 589924 271448 589976 271454
rect 589924 271390 589976 271396
rect 587900 268660 587952 268666
rect 587900 268602 587952 268608
rect 583024 267436 583076 267442
rect 583024 267378 583076 267384
rect 589936 266898 589964 271390
rect 593064 271318 593092 278052
rect 594260 275194 594288 278052
rect 594812 278038 595378 278066
rect 596192 278038 596574 278066
rect 594248 275188 594300 275194
rect 594248 275130 594300 275136
rect 593052 271312 593104 271318
rect 593052 271254 593104 271260
rect 594812 268530 594840 278038
rect 596192 269550 596220 278038
rect 597756 270774 597784 278052
rect 598952 274242 598980 278052
rect 600148 276962 600176 278052
rect 600136 276956 600188 276962
rect 600136 276898 600188 276904
rect 601344 276010 601372 278052
rect 601712 278038 602462 278066
rect 601332 276004 601384 276010
rect 601332 275946 601384 275952
rect 598940 274236 598992 274242
rect 598940 274178 598992 274184
rect 600780 272400 600832 272406
rect 600780 272342 600832 272348
rect 600964 272400 601016 272406
rect 600964 272342 601016 272348
rect 600792 272134 600820 272342
rect 600780 272128 600832 272134
rect 600780 272070 600832 272076
rect 600976 271998 601004 272342
rect 600964 271992 601016 271998
rect 600964 271934 601016 271940
rect 598204 271312 598256 271318
rect 598204 271254 598256 271260
rect 597744 270768 597796 270774
rect 597744 270710 597796 270716
rect 596180 269544 596232 269550
rect 596180 269486 596232 269492
rect 594800 268524 594852 268530
rect 594800 268466 594852 268472
rect 589924 266892 589976 266898
rect 589924 266834 589976 266840
rect 598216 266762 598244 271254
rect 598204 266756 598256 266762
rect 598204 266698 598256 266704
rect 572720 266076 572772 266082
rect 572720 266018 572772 266024
rect 601712 265946 601740 278038
rect 603644 276826 603672 278052
rect 603632 276820 603684 276826
rect 603632 276762 603684 276768
rect 604840 271862 604868 278052
rect 605852 278038 606050 278066
rect 604828 271856 604880 271862
rect 604828 271798 604880 271804
rect 601700 265940 601752 265946
rect 601700 265882 601752 265888
rect 605852 265810 605880 278038
rect 607232 272134 607260 278052
rect 607416 278038 608442 278066
rect 607220 272128 607272 272134
rect 607220 272070 607272 272076
rect 607416 268122 607444 278038
rect 609624 276690 609652 278052
rect 609612 276684 609664 276690
rect 609612 276626 609664 276632
rect 610728 272270 610756 278052
rect 610716 272264 610768 272270
rect 610716 272206 610768 272212
rect 611924 271726 611952 278052
rect 612752 278038 613134 278066
rect 611912 271720 611964 271726
rect 611912 271662 611964 271668
rect 612004 271584 612056 271590
rect 612004 271526 612056 271532
rect 607404 268116 607456 268122
rect 607404 268058 607456 268064
rect 612016 267306 612044 271526
rect 612004 267300 612056 267306
rect 612004 267242 612056 267248
rect 605840 265804 605892 265810
rect 605840 265746 605892 265752
rect 612752 265674 612780 278038
rect 614316 273222 614344 278052
rect 615512 275874 615540 278052
rect 616432 278038 616722 278066
rect 617352 278038 617826 278066
rect 615500 275868 615552 275874
rect 615500 275810 615552 275816
rect 614304 273216 614356 273222
rect 614304 273158 614356 273164
rect 616432 269686 616460 278038
rect 617352 271182 617380 278038
rect 619008 271590 619036 278052
rect 619652 278038 620218 278066
rect 618996 271584 619048 271590
rect 618996 271526 619048 271532
rect 617340 271176 617392 271182
rect 617340 271118 617392 271124
rect 617524 271176 617576 271182
rect 617524 271118 617576 271124
rect 616420 269680 616472 269686
rect 616420 269622 616472 269628
rect 617536 267170 617564 271118
rect 619652 270502 619680 278038
rect 621400 272678 621428 278052
rect 622596 275738 622624 278052
rect 623806 278038 624004 278066
rect 622584 275732 622636 275738
rect 622584 275674 622636 275680
rect 621388 272672 621440 272678
rect 621388 272614 621440 272620
rect 619640 270496 619692 270502
rect 619640 270438 619692 270444
rect 623976 270230 624004 278038
rect 624988 272950 625016 278052
rect 624976 272944 625028 272950
rect 624976 272886 625028 272892
rect 626092 271182 626120 278052
rect 626552 278038 627302 278066
rect 626080 271176 626132 271182
rect 626080 271118 626132 271124
rect 626552 270366 626580 278038
rect 628484 272814 628512 278052
rect 629680 275602 629708 278052
rect 630692 278038 630890 278066
rect 629668 275596 629720 275602
rect 629668 275538 629720 275544
rect 628472 272808 628524 272814
rect 628472 272750 628524 272756
rect 626540 270360 626592 270366
rect 626540 270302 626592 270308
rect 623964 270224 624016 270230
rect 623964 270166 624016 270172
rect 630692 270094 630720 278038
rect 632072 272950 632100 278052
rect 632060 272944 632112 272950
rect 632060 272886 632112 272892
rect 633268 271454 633296 278052
rect 634372 274106 634400 278052
rect 635094 277808 635150 277817
rect 635094 277743 635150 277752
rect 634360 274100 634412 274106
rect 634360 274042 634412 274048
rect 634084 272672 634136 272678
rect 634084 272614 634136 272620
rect 633256 271448 633308 271454
rect 633256 271390 633308 271396
rect 630680 270088 630732 270094
rect 630680 270030 630732 270036
rect 617524 267164 617576 267170
rect 617524 267106 617576 267112
rect 634096 267034 634124 272614
rect 634084 267028 634136 267034
rect 634084 266970 634136 266976
rect 612740 265668 612792 265674
rect 612740 265610 612792 265616
rect 553400 265532 553452 265538
rect 553400 265474 553452 265480
rect 550640 265396 550692 265402
rect 550640 265338 550692 265344
rect 554410 262168 554466 262177
rect 554410 262103 554466 262112
rect 554424 260914 554452 262103
rect 570604 261520 570656 261526
rect 570604 261462 570656 261468
rect 554412 260908 554464 260914
rect 554412 260850 554464 260856
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 554318 259992 554374 260001
rect 554318 259927 554374 259936
rect 554332 259486 554360 259927
rect 554320 259480 554372 259486
rect 554320 259422 554372 259428
rect 563704 259480 563756 259486
rect 563704 259422 563756 259428
rect 553950 257816 554006 257825
rect 553950 257751 554006 257760
rect 553964 256766 553992 257751
rect 553952 256760 554004 256766
rect 553952 256702 554004 256708
rect 560944 256760 560996 256766
rect 560944 256702 560996 256708
rect 554502 255640 554558 255649
rect 554502 255575 554504 255584
rect 554556 255575 554558 255584
rect 558184 255604 558236 255610
rect 554504 255546 554556 255552
rect 558184 255546 558236 255552
rect 554410 253464 554466 253473
rect 554410 253399 554466 253408
rect 554424 252618 554452 253399
rect 554412 252612 554464 252618
rect 554412 252554 554464 252560
rect 554134 251288 554190 251297
rect 554134 251223 554136 251232
rect 554188 251223 554190 251232
rect 556804 251252 556856 251258
rect 554136 251194 554188 251200
rect 556804 251194 556856 251200
rect 554042 249112 554098 249121
rect 554042 249047 554098 249056
rect 553858 246936 553914 246945
rect 553858 246871 553914 246880
rect 553872 245682 553900 246871
rect 553860 245676 553912 245682
rect 553860 245618 553912 245624
rect 553490 244760 553546 244769
rect 553490 244695 553546 244704
rect 553504 244322 553532 244695
rect 553492 244316 553544 244322
rect 553492 244258 553544 244264
rect 553674 242584 553730 242593
rect 553674 242519 553730 242528
rect 553688 241534 553716 242519
rect 553676 241528 553728 241534
rect 553676 241470 553728 241476
rect 553768 236836 553820 236842
rect 553768 236778 553820 236784
rect 553780 236065 553808 236778
rect 553766 236056 553822 236065
rect 553766 235991 553822 236000
rect 156984 231810 157274 231826
rect 155132 231804 155184 231810
rect 155132 231746 155184 231752
rect 156972 231804 157274 231810
rect 157024 231798 157274 231804
rect 156972 231746 157024 231752
rect 134892 231668 134944 231674
rect 134892 231610 134944 231616
rect 92388 231532 92440 231538
rect 92388 231474 92440 231480
rect 64328 231260 64380 231266
rect 64328 231202 64380 231208
rect 64142 231160 64198 231169
rect 64142 231095 64198 231104
rect 86224 230036 86276 230042
rect 86224 229978 86276 229984
rect 68284 229764 68336 229770
rect 68284 229706 68336 229712
rect 67548 228676 67600 228682
rect 67548 228618 67600 228624
rect 64788 227588 64840 227594
rect 64788 227530 64840 227536
rect 63406 223544 63462 223553
rect 63406 223479 63462 223488
rect 63132 223032 63184 223038
rect 63132 222974 63184 222980
rect 62764 222896 62816 222902
rect 62764 222838 62816 222844
rect 62304 219020 62356 219026
rect 62304 218962 62356 218968
rect 61384 218204 61436 218210
rect 61384 218146 61436 218152
rect 61476 218068 61528 218074
rect 61476 218010 61528 218016
rect 59786 217110 59860 217138
rect 60614 217246 60688 217274
rect 59786 216988 59814 217110
rect 60614 216988 60642 217246
rect 61488 217138 61516 218010
rect 62316 217274 62344 218962
rect 62776 218074 62804 222838
rect 64604 219156 64656 219162
rect 64604 219098 64656 219104
rect 63132 218884 63184 218890
rect 63132 218826 63184 218832
rect 62764 218068 62816 218074
rect 62764 218010 62816 218016
rect 61442 217110 61516 217138
rect 62270 217246 62344 217274
rect 61442 216988 61470 217110
rect 62270 216988 62298 217246
rect 63144 217138 63172 218826
rect 63960 218068 64012 218074
rect 63960 218010 64012 218016
rect 63972 217138 64000 218010
rect 64616 217274 64644 219098
rect 64800 218074 64828 227530
rect 66168 226024 66220 226030
rect 66168 225966 66220 225972
rect 66180 218074 66208 225966
rect 66904 223168 66956 223174
rect 66904 223110 66956 223116
rect 66916 219162 66944 223110
rect 66904 219156 66956 219162
rect 66904 219098 66956 219104
rect 67560 218210 67588 228618
rect 66444 218204 66496 218210
rect 66444 218146 66496 218152
rect 67548 218204 67600 218210
rect 67548 218146 67600 218152
rect 68100 218204 68152 218210
rect 68100 218146 68152 218152
rect 64788 218068 64840 218074
rect 64788 218010 64840 218016
rect 65616 218068 65668 218074
rect 65616 218010 65668 218016
rect 66168 218068 66220 218074
rect 66168 218010 66220 218016
rect 64616 217246 64782 217274
rect 63098 217110 63172 217138
rect 63926 217110 64000 217138
rect 63098 216988 63126 217110
rect 63926 216988 63954 217110
rect 64754 216988 64782 217246
rect 65628 217138 65656 218010
rect 66456 217138 66484 218146
rect 67272 218068 67324 218074
rect 67272 218010 67324 218016
rect 67284 217138 67312 218010
rect 68112 217138 68140 218146
rect 68296 218074 68324 229706
rect 82084 229628 82136 229634
rect 82084 229570 82136 229576
rect 75184 227724 75236 227730
rect 75184 227666 75236 227672
rect 72424 225616 72476 225622
rect 72424 225558 72476 225564
rect 68928 224256 68980 224262
rect 68928 224198 68980 224204
rect 68284 218068 68336 218074
rect 68284 218010 68336 218016
rect 68940 217274 68968 224198
rect 69572 223304 69624 223310
rect 69572 223246 69624 223252
rect 69584 218210 69612 223246
rect 71412 223032 71464 223038
rect 71412 222974 71464 222980
rect 69756 220516 69808 220522
rect 69756 220458 69808 220464
rect 69572 218204 69624 218210
rect 69572 218146 69624 218152
rect 69768 217274 69796 220458
rect 70584 219292 70636 219298
rect 70584 219234 70636 219240
rect 65582 217110 65656 217138
rect 66410 217110 66484 217138
rect 67238 217110 67312 217138
rect 68066 217110 68140 217138
rect 68894 217246 68968 217274
rect 69722 217246 69796 217274
rect 65582 216988 65610 217110
rect 66410 216988 66438 217110
rect 67238 216988 67266 217110
rect 68066 216988 68094 217110
rect 68894 216988 68922 217246
rect 69722 216988 69750 217246
rect 70596 217138 70624 219234
rect 71424 217274 71452 222974
rect 72436 219026 72464 225558
rect 73712 224392 73764 224398
rect 73712 224334 73764 224340
rect 73068 220380 73120 220386
rect 73068 220322 73120 220328
rect 72424 219020 72476 219026
rect 72424 218962 72476 218968
rect 72240 218068 72292 218074
rect 72240 218010 72292 218016
rect 70550 217110 70624 217138
rect 71378 217246 71452 217274
rect 70550 216988 70578 217110
rect 71378 216988 71406 217246
rect 72252 217138 72280 218010
rect 73080 217274 73108 220322
rect 73724 218074 73752 224334
rect 73896 221468 73948 221474
rect 73896 221410 73948 221416
rect 73712 218068 73764 218074
rect 73712 218010 73764 218016
rect 73908 217274 73936 221410
rect 75196 218890 75224 227666
rect 76564 225752 76616 225758
rect 76564 225694 76616 225700
rect 75828 223440 75880 223446
rect 75828 223382 75880 223388
rect 75184 218884 75236 218890
rect 75184 218826 75236 218832
rect 75552 218204 75604 218210
rect 75552 218146 75604 218152
rect 74724 218068 74776 218074
rect 74724 218010 74776 218016
rect 72206 217110 72280 217138
rect 73034 217246 73108 217274
rect 73862 217246 73936 217274
rect 72206 216988 72234 217110
rect 73034 216988 73062 217246
rect 73862 216988 73890 217246
rect 74736 217138 74764 218010
rect 75564 217138 75592 218146
rect 75840 218074 75868 223382
rect 76380 220108 76432 220114
rect 76380 220050 76432 220056
rect 75828 218068 75880 218074
rect 75828 218010 75880 218016
rect 76392 217274 76420 220050
rect 76576 218210 76604 225694
rect 79968 224664 80020 224670
rect 79968 224606 80020 224612
rect 78588 222760 78640 222766
rect 78588 222702 78640 222708
rect 77208 218884 77260 218890
rect 77208 218826 77260 218832
rect 76564 218204 76616 218210
rect 76564 218146 76616 218152
rect 74690 217110 74764 217138
rect 75518 217110 75592 217138
rect 76346 217246 76420 217274
rect 74690 216988 74718 217110
rect 75518 216988 75546 217110
rect 76346 216988 76374 217246
rect 77220 217138 77248 218826
rect 78600 218074 78628 222702
rect 79692 220244 79744 220250
rect 79692 220186 79744 220192
rect 78036 218068 78088 218074
rect 78036 218010 78088 218016
rect 78588 218068 78640 218074
rect 78588 218010 78640 218016
rect 78864 218068 78916 218074
rect 78864 218010 78916 218016
rect 78048 217138 78076 218010
rect 78876 217138 78904 218010
rect 79704 217274 79732 220186
rect 79980 218074 80008 224606
rect 81348 223576 81400 223582
rect 81348 223518 81400 223524
rect 80520 221740 80572 221746
rect 80520 221682 80572 221688
rect 79968 218068 80020 218074
rect 79968 218010 80020 218016
rect 80532 217274 80560 221682
rect 81360 217274 81388 223518
rect 82096 221474 82124 229570
rect 83464 225888 83516 225894
rect 83464 225830 83516 225836
rect 82084 221468 82136 221474
rect 82084 221410 82136 221416
rect 83004 220924 83056 220930
rect 83004 220866 83056 220872
rect 82176 218068 82228 218074
rect 82176 218010 82228 218016
rect 77174 217110 77248 217138
rect 78002 217110 78076 217138
rect 78830 217110 78904 217138
rect 79658 217246 79732 217274
rect 80486 217246 80560 217274
rect 81314 217246 81388 217274
rect 77174 216988 77202 217110
rect 78002 216988 78030 217110
rect 78830 216988 78858 217110
rect 79658 216988 79686 217246
rect 80486 216988 80514 217246
rect 81314 216988 81342 217246
rect 82188 217138 82216 218010
rect 83016 217274 83044 220866
rect 83476 218074 83504 225830
rect 85488 224528 85540 224534
rect 85488 224470 85540 224476
rect 85304 222488 85356 222494
rect 85304 222430 85356 222436
rect 83832 219020 83884 219026
rect 83832 218962 83884 218968
rect 83464 218068 83516 218074
rect 83464 218010 83516 218016
rect 82142 217110 82216 217138
rect 82970 217246 83044 217274
rect 82142 216988 82170 217110
rect 82970 216988 82998 217246
rect 83844 217138 83872 218962
rect 85316 218074 85344 222430
rect 84660 218068 84712 218074
rect 84660 218010 84712 218016
rect 85304 218068 85356 218074
rect 85304 218010 85356 218016
rect 84672 217138 84700 218010
rect 85500 217274 85528 224470
rect 86236 221746 86264 229978
rect 88248 227860 88300 227866
rect 88248 227802 88300 227808
rect 87972 222624 88024 222630
rect 87972 222566 88024 222572
rect 86224 221740 86276 221746
rect 86224 221682 86276 221688
rect 86316 221468 86368 221474
rect 86316 221410 86368 221416
rect 86328 217274 86356 221410
rect 87144 218068 87196 218074
rect 87144 218010 87196 218016
rect 83798 217110 83872 217138
rect 84626 217110 84700 217138
rect 85454 217246 85528 217274
rect 86282 217246 86356 217274
rect 83798 216988 83826 217110
rect 84626 216988 84654 217110
rect 85454 216988 85482 217246
rect 86282 216988 86310 217246
rect 87156 217138 87184 218010
rect 87984 217274 88012 222566
rect 88260 218074 88288 227802
rect 89628 227180 89680 227186
rect 89628 227122 89680 227128
rect 89444 224120 89496 224126
rect 89444 224062 89496 224068
rect 89456 218074 89484 224062
rect 88248 218068 88300 218074
rect 88248 218010 88300 218016
rect 88800 218068 88852 218074
rect 88800 218010 88852 218016
rect 89444 218068 89496 218074
rect 89444 218010 89496 218016
rect 87110 217110 87184 217138
rect 87938 217246 88012 217274
rect 87110 216988 87138 217110
rect 87938 216988 87966 217246
rect 88812 217138 88840 218010
rect 89640 217274 89668 227122
rect 91284 221332 91336 221338
rect 91284 221274 91336 221280
rect 91296 217274 91324 221274
rect 92400 219434 92428 231474
rect 128268 231396 128320 231402
rect 128268 231338 128320 231344
rect 94504 230920 94556 230926
rect 94504 230862 94556 230868
rect 93768 228812 93820 228818
rect 93768 228754 93820 228760
rect 92124 219406 92428 219434
rect 92124 217274 92152 219406
rect 93584 219156 93636 219162
rect 93584 219098 93636 219104
rect 92940 218068 92992 218074
rect 92940 218010 92992 218016
rect 88766 217110 88840 217138
rect 89594 217246 89668 217274
rect 90410 217252 90462 217258
rect 88766 216988 88794 217110
rect 89594 216988 89622 217246
rect 90410 217194 90462 217200
rect 91250 217246 91324 217274
rect 92078 217246 92152 217274
rect 90422 216988 90450 217194
rect 91250 216988 91278 217246
rect 92078 216988 92106 217246
rect 92952 217138 92980 218010
rect 93596 217274 93624 219098
rect 93780 218074 93808 228754
rect 94516 219434 94544 230862
rect 104808 230784 104860 230790
rect 104808 230726 104860 230732
rect 95240 230172 95292 230178
rect 95240 230114 95292 230120
rect 95252 227866 95280 230114
rect 102140 229492 102192 229498
rect 102140 229434 102192 229440
rect 100668 229084 100720 229090
rect 100668 229026 100720 229032
rect 95240 227860 95292 227866
rect 95240 227802 95292 227808
rect 96528 227316 96580 227322
rect 96528 227258 96580 227264
rect 96068 224936 96120 224942
rect 96068 224878 96120 224884
rect 94688 221740 94740 221746
rect 94688 221682 94740 221688
rect 94700 219434 94728 221682
rect 94424 219406 94544 219434
rect 94608 219406 94728 219434
rect 96080 219434 96108 224878
rect 96252 224256 96304 224262
rect 96252 224198 96304 224204
rect 96264 223990 96292 224198
rect 96252 223984 96304 223990
rect 96252 223926 96304 223932
rect 96540 219434 96568 227258
rect 99288 222352 99340 222358
rect 99288 222294 99340 222300
rect 97908 222012 97960 222018
rect 97908 221954 97960 221960
rect 96080 219406 96292 219434
rect 94424 219162 94452 219406
rect 94412 219156 94464 219162
rect 94412 219098 94464 219104
rect 93768 218068 93820 218074
rect 93768 218010 93820 218016
rect 94608 217274 94636 219406
rect 96264 218074 96292 219406
rect 96448 219406 96568 219434
rect 95424 218068 95476 218074
rect 95424 218010 95476 218016
rect 96252 218068 96304 218074
rect 96252 218010 96304 218016
rect 93596 217246 93762 217274
rect 92906 217110 92980 217138
rect 92906 216988 92934 217110
rect 93734 216988 93762 217246
rect 94562 217246 94636 217274
rect 94562 216988 94590 217246
rect 95436 217138 95464 218010
rect 96448 217274 96476 219406
rect 97080 218204 97132 218210
rect 97080 218146 97132 218152
rect 95390 217110 95464 217138
rect 96218 217246 96476 217274
rect 95390 216988 95418 217110
rect 96218 216988 96246 217246
rect 97092 217138 97120 218146
rect 97920 217274 97948 221954
rect 99300 218074 99328 222294
rect 100392 218612 100444 218618
rect 100392 218554 100444 218560
rect 98736 218068 98788 218074
rect 98736 218010 98788 218016
rect 99288 218068 99340 218074
rect 99288 218010 99340 218016
rect 99564 218068 99616 218074
rect 99564 218010 99616 218016
rect 97046 217110 97120 217138
rect 97874 217246 97948 217274
rect 97046 216988 97074 217110
rect 97874 216988 97902 217246
rect 98748 217138 98776 218010
rect 99576 217138 99604 218010
rect 100404 217138 100432 218554
rect 100680 218074 100708 229026
rect 102152 227458 102180 229434
rect 102140 227452 102192 227458
rect 102140 227394 102192 227400
rect 103428 227452 103480 227458
rect 103428 227394 103480 227400
rect 102048 224800 102100 224806
rect 102048 224742 102100 224748
rect 101220 220652 101272 220658
rect 101220 220594 101272 220600
rect 100668 218068 100720 218074
rect 100668 218010 100720 218016
rect 101232 217274 101260 220594
rect 102060 217274 102088 224742
rect 103440 218142 103468 227394
rect 104532 221876 104584 221882
rect 104532 221818 104584 221824
rect 102876 218136 102928 218142
rect 102876 218078 102928 218084
rect 103428 218136 103480 218142
rect 103428 218078 103480 218084
rect 103704 218136 103756 218142
rect 103704 218078 103756 218084
rect 98702 217110 98776 217138
rect 99530 217110 99604 217138
rect 100358 217110 100432 217138
rect 101186 217246 101260 217274
rect 102014 217246 102088 217274
rect 98702 216988 98730 217110
rect 99530 216988 99558 217110
rect 100358 216988 100386 217110
rect 101186 216988 101214 217246
rect 102014 216988 102042 217246
rect 102888 217138 102916 218078
rect 103716 217138 103744 218078
rect 104544 217274 104572 221818
rect 104820 218142 104848 230726
rect 118608 230648 118660 230654
rect 118608 230590 118660 230596
rect 110144 229356 110196 229362
rect 110144 229298 110196 229304
rect 106188 228948 106240 228954
rect 106188 228890 106240 228896
rect 106004 223984 106056 223990
rect 106004 223926 106056 223932
rect 106016 218142 106044 223926
rect 104808 218136 104860 218142
rect 104808 218078 104860 218084
rect 105360 218136 105412 218142
rect 105360 218078 105412 218084
rect 106004 218136 106056 218142
rect 106004 218078 106056 218084
rect 102842 217110 102916 217138
rect 103670 217110 103744 217138
rect 104498 217246 104572 217274
rect 102842 216988 102870 217110
rect 103670 216988 103698 217110
rect 104498 216988 104526 217246
rect 105372 217138 105400 218078
rect 106200 217274 106228 228890
rect 110156 227594 110184 229298
rect 112996 228268 113048 228274
rect 112996 228210 113048 228216
rect 110144 227588 110196 227594
rect 110144 227530 110196 227536
rect 110328 227588 110380 227594
rect 110328 227530 110380 227536
rect 110144 225480 110196 225486
rect 110144 225422 110196 225428
rect 108672 223848 108724 223854
rect 108672 223790 108724 223796
rect 107844 219972 107896 219978
rect 107844 219914 107896 219920
rect 107016 218476 107068 218482
rect 107016 218418 107068 218424
rect 105326 217110 105400 217138
rect 106154 217246 106228 217274
rect 105326 216988 105354 217110
rect 106154 216988 106182 217246
rect 107028 217138 107056 218418
rect 107856 217274 107884 219914
rect 108684 217274 108712 223790
rect 110156 219434 110184 225422
rect 110340 219434 110368 227530
rect 112812 223712 112864 223718
rect 112812 223654 112864 223660
rect 111156 221060 111208 221066
rect 111156 221002 111208 221008
rect 109500 219428 109552 219434
rect 110156 219406 110276 219434
rect 110340 219428 110472 219434
rect 110340 219406 110420 219428
rect 109500 219370 109552 219376
rect 106982 217110 107056 217138
rect 107810 217246 107884 217274
rect 108638 217246 108712 217274
rect 106982 216988 107010 217110
rect 107810 216988 107838 217246
rect 108638 216988 108666 217246
rect 109512 217138 109540 219370
rect 110248 217274 110276 219406
rect 110420 219370 110472 219376
rect 111168 217274 111196 221002
rect 112824 218142 112852 223654
rect 111984 218136 112036 218142
rect 111984 218078 112036 218084
rect 112812 218136 112864 218142
rect 112812 218078 112864 218084
rect 110248 217246 110322 217274
rect 109466 217110 109540 217138
rect 109466 216988 109494 217110
rect 110294 216988 110322 217246
rect 111122 217246 111196 217274
rect 111122 216988 111150 217246
rect 111996 217138 112024 218078
rect 113008 217274 113036 228210
rect 117228 226772 117280 226778
rect 117228 226714 117280 226720
rect 114284 220788 114336 220794
rect 114284 220730 114336 220736
rect 114296 219978 114324 220730
rect 114284 219972 114336 219978
rect 114284 219914 114336 219920
rect 114468 219972 114520 219978
rect 114468 219914 114520 219920
rect 113640 219428 113692 219434
rect 113640 219370 113692 219376
rect 111950 217110 112024 217138
rect 112778 217246 113036 217274
rect 111950 216988 111978 217110
rect 112778 216988 112806 217246
rect 113652 217138 113680 219370
rect 114480 217274 114508 219914
rect 117240 218142 117268 226714
rect 118424 222216 118476 222222
rect 118424 222158 118476 222164
rect 118148 221332 118200 221338
rect 118148 221274 118200 221280
rect 118160 221066 118188 221274
rect 118148 221060 118200 221066
rect 118148 221002 118200 221008
rect 118436 219434 118464 222158
rect 118436 219406 118556 219434
rect 117780 219292 117832 219298
rect 117780 219234 117832 219240
rect 117792 218346 117820 219234
rect 117964 219156 118016 219162
rect 117964 219098 118016 219104
rect 117976 218482 118004 219098
rect 117964 218476 118016 218482
rect 117964 218418 118016 218424
rect 117780 218340 117832 218346
rect 117780 218282 117832 218288
rect 117780 218204 117832 218210
rect 117780 218146 117832 218152
rect 116124 218136 116176 218142
rect 116124 218078 116176 218084
rect 117228 218136 117280 218142
rect 117228 218078 117280 218084
rect 115296 217456 115348 217462
rect 115296 217398 115348 217404
rect 113606 217110 113680 217138
rect 114434 217246 114508 217274
rect 113606 216988 113634 217110
rect 114434 216988 114462 217246
rect 115308 217138 115336 217398
rect 116136 217138 116164 218078
rect 116952 217592 117004 217598
rect 116952 217534 117004 217540
rect 116964 217138 116992 217534
rect 117792 217138 117820 218146
rect 118528 217274 118556 219406
rect 118620 218226 118648 230590
rect 126888 230444 126940 230450
rect 126888 230386 126940 230392
rect 123484 229220 123536 229226
rect 123484 229162 123536 229168
rect 119988 228132 120040 228138
rect 119988 228074 120040 228080
rect 118620 218210 118740 218226
rect 118620 218204 118752 218210
rect 118620 218198 118700 218204
rect 118700 218146 118752 218152
rect 120000 218142 120028 228074
rect 122748 226908 122800 226914
rect 122748 226850 122800 226856
rect 122564 225208 122616 225214
rect 122564 225150 122616 225156
rect 121092 219836 121144 219842
rect 121092 219778 121144 219784
rect 120264 218476 120316 218482
rect 120264 218418 120316 218424
rect 119436 218136 119488 218142
rect 119436 218078 119488 218084
rect 119988 218136 120040 218142
rect 119988 218078 120040 218084
rect 118528 217246 118602 217274
rect 115262 217110 115336 217138
rect 116090 217110 116164 217138
rect 116918 217110 116992 217138
rect 117746 217110 117820 217138
rect 115262 216988 115290 217110
rect 116090 216988 116118 217110
rect 116918 216988 116946 217110
rect 117746 216988 117774 217110
rect 118574 216988 118602 217246
rect 119448 217138 119476 218078
rect 120276 217138 120304 218418
rect 121104 217274 121132 219778
rect 122576 218142 122604 225150
rect 121920 218136 121972 218142
rect 121920 218078 121972 218084
rect 122564 218136 122616 218142
rect 122564 218078 122616 218084
rect 119402 217110 119476 217138
rect 120230 217110 120304 217138
rect 121058 217246 121132 217274
rect 119402 216988 119430 217110
rect 120230 216988 120258 217110
rect 121058 216988 121086 217246
rect 121932 217138 121960 218078
rect 122760 217274 122788 226850
rect 123496 218346 123524 229162
rect 126704 227996 126756 228002
rect 126704 227938 126756 227944
rect 125232 225072 125284 225078
rect 125232 225014 125284 225020
rect 124404 221060 124456 221066
rect 124404 221002 124456 221008
rect 123484 218340 123536 218346
rect 123484 218282 123536 218288
rect 123668 218272 123720 218278
rect 123668 218214 123720 218220
rect 123680 217274 123708 218214
rect 124416 217274 124444 221002
rect 125244 217274 125272 225014
rect 126716 218142 126744 227938
rect 126060 218136 126112 218142
rect 126060 218078 126112 218084
rect 126704 218136 126756 218142
rect 126704 218078 126756 218084
rect 121886 217110 121960 217138
rect 122714 217246 122788 217274
rect 123542 217246 123708 217274
rect 124370 217246 124444 217274
rect 125198 217246 125272 217274
rect 121886 216988 121914 217110
rect 122714 216988 122742 217246
rect 123542 216988 123570 217246
rect 124370 216988 124398 217246
rect 125198 216988 125226 217246
rect 126072 217138 126100 218078
rect 126900 217274 126928 230386
rect 127440 226160 127492 226166
rect 127440 226102 127492 226108
rect 127452 225486 127480 226102
rect 127440 225480 127492 225486
rect 127440 225422 127492 225428
rect 127440 221332 127492 221338
rect 127440 221274 127492 221280
rect 127452 221066 127480 221274
rect 127256 221060 127308 221066
rect 127256 221002 127308 221008
rect 127440 221060 127492 221066
rect 127440 221002 127492 221008
rect 127900 221060 127952 221066
rect 127900 221002 127952 221008
rect 127268 220946 127296 221002
rect 127912 220946 127940 221002
rect 127268 220918 127940 220946
rect 127624 219972 127676 219978
rect 127624 219914 127676 219920
rect 127636 219706 127664 219914
rect 127624 219700 127676 219706
rect 127624 219642 127676 219648
rect 128280 218142 128308 231338
rect 133788 230308 133840 230314
rect 133788 230250 133840 230256
rect 130384 229900 130436 229906
rect 130384 229842 130436 229848
rect 129556 226636 129608 226642
rect 129556 226578 129608 226584
rect 129372 225208 129424 225214
rect 129372 225150 129424 225156
rect 129384 218142 129412 225150
rect 127716 218136 127768 218142
rect 127716 218078 127768 218084
rect 128268 218136 128320 218142
rect 128268 218078 128320 218084
rect 128544 218136 128596 218142
rect 128544 218078 128596 218084
rect 129372 218136 129424 218142
rect 129372 218078 129424 218084
rect 126026 217110 126100 217138
rect 126854 217246 126928 217274
rect 126026 216988 126054 217110
rect 126854 216988 126882 217246
rect 127728 217138 127756 218078
rect 128556 217138 128584 218078
rect 129568 217274 129596 226578
rect 130396 226302 130424 229842
rect 133512 227860 133564 227866
rect 133512 227802 133564 227808
rect 130384 226296 130436 226302
rect 130384 226238 130436 226244
rect 132408 225072 132460 225078
rect 132408 225014 132460 225020
rect 131028 219700 131080 219706
rect 131028 219642 131080 219648
rect 130200 218340 130252 218346
rect 130200 218282 130252 218288
rect 127682 217110 127756 217138
rect 128510 217110 128584 217138
rect 129338 217246 129596 217274
rect 127682 216988 127710 217110
rect 128510 216988 128538 217110
rect 129338 216988 129366 217246
rect 130212 217138 130240 218282
rect 131040 217274 131068 219642
rect 132420 219298 132448 225014
rect 131856 219292 131908 219298
rect 131856 219234 131908 219240
rect 132408 219292 132460 219298
rect 132408 219234 132460 219240
rect 132592 219292 132644 219298
rect 132592 219234 132644 219240
rect 130166 217110 130240 217138
rect 130994 217246 131068 217274
rect 130166 216988 130194 217110
rect 130994 216988 131022 217246
rect 131868 217138 131896 219234
rect 132604 218226 132632 219234
rect 132512 218210 132632 218226
rect 132500 218204 132632 218210
rect 132552 218198 132632 218204
rect 132500 218146 132552 218152
rect 133524 218142 133552 227802
rect 133800 219434 133828 230250
rect 134904 219434 134932 231610
rect 140042 229120 140098 229129
rect 140042 229055 140098 229064
rect 137376 228540 137428 228546
rect 137376 228482 137428 228488
rect 136824 228404 136876 228410
rect 136824 228346 136876 228352
rect 136638 227896 136694 227905
rect 136836 227866 136864 228346
rect 137388 228290 137416 228482
rect 139308 228404 139360 228410
rect 139308 228346 139360 228352
rect 137204 228274 137416 228290
rect 137192 228268 137416 228274
rect 137244 228262 137416 228268
rect 137192 228210 137244 228216
rect 136638 227831 136640 227840
rect 136692 227831 136694 227840
rect 136824 227860 136876 227866
rect 136640 227802 136692 227808
rect 136824 227802 136876 227808
rect 136548 226500 136600 226506
rect 136548 226442 136600 226448
rect 135076 226296 135128 226302
rect 135076 226238 135128 226244
rect 133708 219406 133828 219434
rect 134352 219406 134932 219434
rect 132684 218136 132736 218142
rect 132684 218078 132736 218084
rect 133512 218136 133564 218142
rect 133512 218078 133564 218084
rect 132696 217138 132724 218078
rect 133708 217274 133736 219406
rect 134352 217274 134380 219406
rect 131822 217110 131896 217138
rect 132650 217110 132724 217138
rect 133478 217246 133736 217274
rect 134306 217246 134380 217274
rect 135088 217274 135116 226238
rect 136178 219328 136234 219337
rect 136178 219263 136180 219272
rect 136232 219263 136234 219272
rect 136364 219292 136416 219298
rect 136180 219234 136232 219240
rect 136364 219234 136416 219240
rect 136376 218346 136404 219234
rect 136364 218340 136416 218346
rect 136364 218282 136416 218288
rect 136560 218142 136588 226442
rect 138018 224360 138074 224369
rect 138018 224295 138074 224304
rect 138032 224210 138060 224295
rect 137986 224182 138060 224210
rect 137986 224126 138014 224182
rect 137974 224120 138026 224126
rect 137282 224088 137338 224097
rect 138112 224120 138164 224126
rect 137974 224062 138026 224068
rect 138110 224088 138112 224097
rect 138164 224088 138166 224097
rect 137282 224023 137338 224032
rect 138110 224023 138166 224032
rect 136916 220516 136968 220522
rect 136916 220458 136968 220464
rect 137100 220516 137152 220522
rect 137100 220458 137152 220464
rect 136928 219570 136956 220458
rect 137112 219842 137140 220458
rect 137100 219836 137152 219842
rect 137100 219778 137152 219784
rect 136916 219564 136968 219570
rect 136916 219506 136968 219512
rect 137296 219337 137324 224023
rect 138478 221640 138534 221649
rect 138478 221575 138534 221584
rect 137652 219564 137704 219570
rect 137652 219506 137704 219512
rect 137282 219328 137338 219337
rect 137282 219263 137338 219272
rect 136824 218340 136876 218346
rect 136824 218282 136876 218288
rect 135996 218136 136048 218142
rect 135996 218078 136048 218084
rect 136548 218136 136600 218142
rect 136548 218078 136600 218084
rect 135088 217246 135162 217274
rect 131822 216988 131850 217110
rect 132650 216988 132678 217110
rect 133478 216988 133506 217246
rect 134306 216988 134334 217246
rect 135134 216988 135162 217246
rect 136008 217138 136036 218078
rect 136836 217138 136864 218282
rect 137664 217274 137692 219506
rect 135962 217110 136036 217138
rect 136790 217110 136864 217138
rect 137618 217246 137692 217274
rect 135962 216988 135990 217110
rect 136790 216988 136818 217110
rect 137618 216988 137646 217246
rect 138492 217138 138520 221575
rect 139320 217274 139348 228346
rect 139860 223032 139912 223038
rect 139860 222974 139912 222980
rect 139872 222873 139900 222974
rect 139858 222864 139914 222873
rect 139858 222799 139914 222808
rect 140056 218754 140084 229055
rect 141160 227866 141188 231676
rect 141344 231662 141818 231690
rect 142068 231668 142120 231674
rect 141148 227860 141200 227866
rect 141148 227802 141200 227808
rect 141344 221610 141372 231662
rect 142068 231610 142120 231616
rect 142080 230602 142108 231610
rect 142080 230574 142200 230602
rect 142172 230518 142200 230574
rect 142160 230512 142212 230518
rect 142160 230454 142212 230460
rect 141976 230444 142028 230450
rect 141976 230386 142028 230392
rect 141988 229945 142016 230386
rect 142158 230208 142214 230217
rect 142158 230143 142214 230152
rect 141974 229936 142030 229945
rect 141974 229871 142030 229880
rect 142172 229770 142200 230143
rect 142160 229764 142212 229770
rect 142160 229706 142212 229712
rect 141514 227896 141570 227905
rect 141514 227831 141516 227840
rect 141568 227831 141570 227840
rect 141516 227802 141568 227808
rect 142448 227050 142476 231676
rect 142618 229936 142674 229945
rect 142618 229871 142620 229880
rect 142672 229871 142674 229880
rect 142620 229842 142672 229848
rect 143092 228274 143120 231676
rect 143552 231662 143750 231690
rect 144012 231662 144394 231690
rect 143552 229129 143580 231662
rect 143538 229120 143594 229129
rect 143538 229055 143594 229064
rect 143080 228268 143132 228274
rect 143080 228210 143132 228216
rect 143448 228268 143500 228274
rect 143448 228210 143500 228216
rect 142436 227044 142488 227050
rect 142436 226986 142488 226992
rect 143264 227044 143316 227050
rect 143264 226986 143316 226992
rect 141790 226536 141846 226545
rect 141790 226471 141792 226480
rect 141844 226471 141846 226480
rect 142250 226536 142306 226545
rect 142250 226471 142252 226480
rect 141792 226442 141844 226448
rect 142304 226471 142306 226480
rect 142252 226442 142304 226448
rect 141976 226432 142028 226438
rect 141976 226374 142028 226380
rect 142114 226432 142166 226438
rect 142166 226380 142292 226386
rect 142114 226374 142292 226380
rect 141988 224954 142016 226374
rect 142126 226358 142292 226374
rect 142264 226166 142292 226358
rect 142114 226160 142166 226166
rect 142114 226102 142166 226108
rect 142252 226160 142304 226166
rect 142252 226102 142304 226108
rect 142126 225978 142154 226102
rect 142620 226024 142672 226030
rect 142618 225992 142620 226001
rect 142804 226024 142856 226030
rect 142672 225992 142674 226001
rect 142126 225950 142292 225978
rect 142264 225622 142292 225950
rect 142804 225966 142856 225972
rect 142618 225927 142674 225936
rect 142114 225616 142166 225622
rect 142114 225558 142166 225564
rect 142252 225616 142304 225622
rect 142816 225570 142844 225966
rect 142252 225558 142304 225564
rect 142126 225434 142154 225558
rect 142448 225542 142844 225570
rect 142448 225434 142476 225542
rect 142126 225406 142476 225434
rect 141804 224926 142016 224954
rect 141514 221640 141570 221649
rect 141332 221604 141384 221610
rect 141514 221575 141516 221584
rect 141332 221546 141384 221552
rect 141568 221575 141570 221584
rect 141516 221546 141568 221552
rect 140044 218748 140096 218754
rect 140044 218690 140096 218696
rect 140964 218748 141016 218754
rect 140964 218690 141016 218696
rect 140136 218204 140188 218210
rect 140136 218146 140188 218152
rect 138446 217110 138520 217138
rect 139274 217246 139348 217274
rect 138446 216988 138474 217110
rect 139274 216988 139302 217246
rect 140148 217138 140176 218146
rect 140976 217138 141004 218690
rect 141804 217274 141832 224926
rect 142528 223168 142580 223174
rect 142526 223136 142528 223145
rect 142580 223136 142582 223145
rect 142526 223071 142582 223080
rect 142066 221640 142122 221649
rect 142066 221575 142122 221584
rect 142080 218754 142108 221575
rect 143080 219700 143132 219706
rect 143080 219642 143132 219648
rect 143092 219586 143120 219642
rect 142724 219570 143120 219586
rect 142712 219564 143120 219570
rect 142764 219558 143120 219564
rect 142712 219506 142764 219512
rect 143276 218754 143304 226986
rect 142068 218748 142120 218754
rect 142068 218690 142120 218696
rect 142620 218748 142672 218754
rect 142620 218690 142672 218696
rect 143264 218748 143316 218754
rect 143264 218690 143316 218696
rect 140102 217110 140176 217138
rect 140930 217110 141004 217138
rect 141758 217246 141832 217274
rect 140102 216988 140130 217110
rect 140930 216988 140958 217110
rect 141758 216988 141786 217246
rect 142632 217138 142660 218690
rect 143460 217274 143488 228210
rect 143816 223304 143868 223310
rect 143816 223246 143868 223252
rect 143632 223168 143684 223174
rect 143630 223136 143632 223145
rect 143684 223136 143686 223145
rect 143630 223071 143686 223080
rect 143828 222873 143856 223246
rect 144012 222902 144040 231662
rect 145024 229770 145052 231676
rect 145012 229764 145064 229770
rect 145012 229706 145064 229712
rect 145668 229498 145696 231676
rect 145656 229492 145708 229498
rect 145656 229434 145708 229440
rect 145840 229492 145892 229498
rect 145840 229434 145892 229440
rect 144642 229392 144698 229401
rect 144642 229327 144644 229336
rect 144696 229327 144698 229336
rect 144828 229356 144880 229362
rect 144644 229298 144696 229304
rect 144828 229298 144880 229304
rect 144840 224954 144868 229298
rect 145852 228274 145880 229434
rect 146024 228676 146076 228682
rect 146024 228618 146076 228624
rect 146036 228274 146064 228618
rect 145840 228268 145892 228274
rect 145840 228210 145892 228216
rect 146024 228268 146076 228274
rect 146024 228210 146076 228216
rect 145930 228032 145986 228041
rect 145930 227967 145986 227976
rect 144196 224926 144868 224954
rect 144000 222896 144052 222902
rect 143814 222864 143870 222873
rect 144000 222838 144052 222844
rect 143814 222799 143870 222808
rect 144196 219722 144224 224926
rect 145104 222896 145156 222902
rect 145104 222838 145156 222844
rect 144104 219694 144224 219722
rect 144104 219570 144132 219694
rect 144092 219564 144144 219570
rect 144092 219506 144144 219512
rect 144276 219564 144328 219570
rect 144276 219506 144328 219512
rect 142586 217110 142660 217138
rect 143414 217246 143488 217274
rect 142586 216988 142614 217110
rect 143414 216988 143442 217246
rect 144288 217138 144316 219506
rect 145116 217138 145144 222838
rect 145944 217274 145972 227967
rect 146312 227730 146340 231676
rect 146680 231662 146970 231690
rect 146680 229094 146708 231662
rect 146944 229764 146996 229770
rect 146944 229706 146996 229712
rect 146956 229226 146984 229706
rect 146944 229220 146996 229226
rect 146944 229162 146996 229168
rect 146588 229066 146708 229094
rect 146300 227724 146352 227730
rect 146300 227666 146352 227672
rect 146588 223174 146616 229066
rect 147128 228540 147180 228546
rect 147128 228482 147180 228488
rect 147140 228041 147168 228482
rect 147126 228032 147182 228041
rect 147126 227967 147182 227976
rect 147600 226030 147628 231676
rect 148244 229922 148272 231676
rect 148244 229894 148364 229922
rect 148140 229764 148192 229770
rect 148140 229706 148192 229712
rect 148152 229650 148180 229706
rect 147784 229634 148180 229650
rect 147772 229628 148180 229634
rect 147824 229622 148180 229628
rect 147772 229570 147824 229576
rect 148336 229401 148364 229894
rect 148322 229392 148378 229401
rect 148322 229327 148378 229336
rect 148324 229220 148376 229226
rect 148324 229162 148376 229168
rect 147588 226024 147640 226030
rect 147588 225966 147640 225972
rect 147772 226024 147824 226030
rect 147772 225966 147824 225972
rect 147784 225706 147812 225966
rect 147692 225678 147812 225706
rect 147692 225622 147720 225678
rect 147680 225616 147732 225622
rect 147680 225558 147732 225564
rect 146576 223168 146628 223174
rect 146576 223110 146628 223116
rect 146760 223168 146812 223174
rect 146760 223110 146812 223116
rect 146772 220946 146800 223110
rect 147586 221640 147642 221649
rect 147404 221604 147456 221610
rect 147586 221575 147588 221584
rect 147404 221546 147456 221552
rect 147640 221575 147642 221584
rect 147588 221546 147640 221552
rect 147416 221082 147444 221546
rect 147416 221066 147674 221082
rect 147416 221060 147686 221066
rect 147416 221054 147634 221060
rect 147634 221002 147686 221008
rect 146588 220918 146800 220946
rect 146588 218618 146616 220918
rect 147220 220856 147272 220862
rect 147218 220824 147220 220833
rect 147272 220824 147274 220833
rect 146760 220788 146812 220794
rect 147218 220759 147274 220768
rect 146760 220730 146812 220736
rect 146772 220538 146800 220730
rect 147036 220652 147088 220658
rect 147680 220652 147732 220658
rect 147088 220612 147680 220640
rect 147036 220594 147088 220600
rect 147680 220594 147732 220600
rect 146772 220510 147444 220538
rect 147218 220416 147274 220425
rect 147416 220386 147444 220510
rect 147588 220516 147640 220522
rect 147588 220458 147640 220464
rect 147218 220351 147220 220360
rect 147272 220351 147274 220360
rect 147404 220380 147456 220386
rect 147220 220322 147272 220328
rect 147404 220322 147456 220328
rect 146760 218748 146812 218754
rect 146760 218690 146812 218696
rect 146576 218612 146628 218618
rect 146576 218554 146628 218560
rect 144242 217110 144316 217138
rect 145070 217110 145144 217138
rect 145898 217246 145972 217274
rect 144242 216988 144270 217110
rect 145070 216988 145098 217110
rect 145898 216988 145926 217246
rect 146772 217138 146800 218690
rect 147600 217138 147628 220458
rect 148336 220425 148364 229162
rect 148888 228274 148916 231676
rect 148876 228268 148928 228274
rect 148876 228210 148928 228216
rect 148874 225448 148930 225457
rect 148874 225383 148930 225392
rect 148322 220416 148378 220425
rect 148322 220351 148378 220360
rect 148888 218618 148916 225383
rect 149532 223038 149560 231676
rect 149808 231662 150190 231690
rect 150544 231662 150834 231690
rect 149808 226001 149836 231662
rect 150544 230217 150572 231662
rect 150530 230208 150586 230217
rect 150530 230143 150586 230152
rect 151464 229362 151492 231676
rect 151452 229356 151504 229362
rect 151452 229298 151504 229304
rect 151636 229356 151688 229362
rect 151636 229298 151688 229304
rect 150346 229120 150402 229129
rect 150346 229055 150402 229064
rect 150072 227724 150124 227730
rect 150072 227666 150124 227672
rect 149794 225992 149850 226001
rect 149794 225927 149850 225936
rect 149520 223032 149572 223038
rect 149520 222974 149572 222980
rect 150084 218618 150112 227666
rect 150360 219434 150388 229055
rect 151648 227338 151676 229298
rect 151188 227310 151676 227338
rect 151188 220833 151216 227310
rect 151358 226264 151414 226273
rect 151358 226199 151414 226208
rect 151174 220824 151230 220833
rect 151174 220759 151230 220768
rect 150714 220552 150770 220561
rect 150714 220487 150716 220496
rect 150768 220487 150770 220496
rect 150900 220516 150952 220522
rect 150716 220458 150768 220464
rect 150900 220458 150952 220464
rect 150268 219406 150388 219434
rect 148416 218612 148468 218618
rect 148416 218554 148468 218560
rect 148876 218612 148928 218618
rect 148876 218554 148928 218560
rect 149244 218612 149296 218618
rect 149244 218554 149296 218560
rect 150072 218612 150124 218618
rect 150072 218554 150124 218560
rect 148428 217138 148456 218554
rect 149256 217138 149284 218554
rect 150268 217274 150296 219406
rect 150440 218884 150492 218890
rect 150440 218826 150492 218832
rect 150452 218618 150480 218826
rect 150440 218612 150492 218618
rect 150440 218554 150492 218560
rect 150912 217274 150940 220458
rect 151372 219434 151400 226199
rect 152108 223310 152136 231676
rect 152384 231662 152766 231690
rect 152384 224369 152412 231662
rect 153396 229634 153424 231676
rect 153384 229628 153436 229634
rect 153384 229570 153436 229576
rect 153844 229628 153896 229634
rect 153844 229570 153896 229576
rect 153108 228404 153160 228410
rect 153108 228346 153160 228352
rect 152370 224360 152426 224369
rect 152370 224295 152426 224304
rect 152096 223304 152148 223310
rect 152096 223246 152148 223252
rect 151910 220552 151966 220561
rect 151910 220487 151912 220496
rect 151964 220487 151966 220496
rect 151912 220458 151964 220464
rect 151556 220386 151952 220402
rect 151544 220380 151952 220386
rect 151596 220374 151952 220380
rect 151544 220322 151596 220328
rect 151726 220280 151782 220289
rect 151924 220250 151952 220374
rect 151726 220215 151728 220224
rect 151780 220215 151782 220224
rect 151912 220244 151964 220250
rect 151728 220186 151780 220192
rect 151912 220186 151964 220192
rect 151372 219406 151676 219434
rect 146726 217110 146800 217138
rect 147554 217110 147628 217138
rect 148382 217110 148456 217138
rect 149210 217110 149284 217138
rect 150038 217246 150296 217274
rect 150866 217246 150940 217274
rect 151648 217274 151676 219406
rect 152372 218884 152424 218890
rect 152372 218826 152424 218832
rect 152384 218618 152412 218826
rect 153120 218618 153148 228346
rect 153856 218890 153884 229570
rect 154040 229226 154068 231676
rect 154396 229356 154448 229362
rect 154396 229298 154448 229304
rect 154028 229220 154080 229226
rect 154028 229162 154080 229168
rect 154408 224954 154436 229298
rect 154040 224926 154436 224954
rect 154040 220250 154068 224926
rect 154684 223446 154712 231676
rect 154672 223440 154724 223446
rect 154672 223382 154724 223388
rect 154212 222896 154264 222902
rect 154212 222838 154264 222844
rect 154028 220244 154080 220250
rect 154028 220186 154080 220192
rect 153844 218884 153896 218890
rect 153844 218826 153896 218832
rect 152372 218612 152424 218618
rect 152372 218554 152424 218560
rect 152556 218612 152608 218618
rect 152556 218554 152608 218560
rect 153108 218612 153160 218618
rect 153108 218554 153160 218560
rect 153384 218612 153436 218618
rect 153384 218554 153436 218560
rect 151648 217246 151722 217274
rect 146726 216988 146754 217110
rect 147554 216988 147582 217110
rect 148382 216988 148410 217110
rect 149210 216988 149238 217110
rect 150038 216988 150066 217246
rect 150866 216988 150894 217246
rect 151694 216988 151722 217246
rect 152568 217138 152596 218554
rect 153396 217138 153424 218554
rect 154224 217274 154252 222838
rect 155144 222766 155172 231746
rect 155328 224398 155356 231676
rect 155500 231668 155552 231674
rect 155500 231610 155552 231616
rect 155512 225894 155540 231610
rect 155972 229770 156000 231676
rect 156156 231662 156630 231690
rect 157628 231662 157918 231690
rect 155960 229764 156012 229770
rect 155960 229706 156012 229712
rect 155866 227080 155922 227089
rect 155866 227015 155922 227024
rect 155500 225888 155552 225894
rect 155500 225830 155552 225836
rect 155316 224392 155368 224398
rect 155316 224334 155368 224340
rect 155132 222760 155184 222766
rect 155132 222702 155184 222708
rect 155684 222760 155736 222766
rect 155684 222702 155736 222708
rect 154394 220280 154450 220289
rect 154394 220215 154396 220224
rect 154448 220215 154450 220224
rect 154396 220186 154448 220192
rect 154672 219156 154724 219162
rect 154672 219098 154724 219104
rect 154684 218890 154712 219098
rect 154672 218884 154724 218890
rect 154672 218826 154724 218832
rect 154486 218648 154542 218657
rect 155696 218618 155724 222702
rect 154486 218583 154488 218592
rect 154540 218583 154542 218592
rect 155040 218612 155092 218618
rect 154488 218554 154540 218560
rect 155040 218554 155092 218560
rect 155684 218612 155736 218618
rect 155684 218554 155736 218560
rect 152522 217110 152596 217138
rect 153350 217110 153424 217138
rect 154178 217246 154252 217274
rect 152522 216988 152550 217110
rect 153350 216988 153378 217110
rect 154178 216988 154206 217246
rect 155052 217138 155080 218554
rect 155880 217274 155908 227015
rect 156156 220114 156184 231662
rect 157430 230208 157486 230217
rect 157430 230143 157432 230152
rect 157484 230143 157486 230152
rect 157432 230114 157484 230120
rect 157154 230072 157210 230081
rect 157154 230007 157156 230016
rect 157208 230007 157210 230016
rect 157156 229978 157208 229984
rect 157168 229894 157472 229922
rect 156328 229764 156380 229770
rect 156328 229706 156380 229712
rect 156340 229226 156368 229706
rect 157168 229362 157196 229894
rect 157444 229770 157472 229894
rect 157628 229786 157656 231662
rect 157798 230208 157854 230217
rect 157798 230143 157854 230152
rect 157812 230042 157840 230143
rect 157800 230036 157852 230042
rect 157800 229978 157852 229984
rect 157984 230036 158036 230042
rect 157984 229978 158036 229984
rect 157294 229764 157346 229770
rect 157294 229706 157346 229712
rect 157432 229764 157484 229770
rect 157628 229758 157840 229786
rect 157432 229706 157484 229712
rect 157306 229650 157334 229706
rect 157614 229664 157670 229673
rect 157306 229622 157614 229650
rect 157614 229599 157670 229608
rect 157156 229356 157208 229362
rect 157156 229298 157208 229304
rect 157340 229356 157392 229362
rect 157340 229298 157392 229304
rect 157352 229242 157380 229298
rect 156328 229220 156380 229226
rect 156328 229162 156380 229168
rect 157168 229214 157380 229242
rect 157168 229129 157196 229214
rect 157154 229120 157210 229129
rect 157154 229055 157210 229064
rect 157338 227488 157394 227497
rect 157338 227423 157394 227432
rect 157352 227338 157380 227423
rect 157306 227310 157380 227338
rect 157306 227186 157334 227310
rect 157430 227216 157486 227225
rect 157294 227180 157346 227186
rect 157430 227151 157432 227160
rect 157294 227122 157346 227128
rect 157484 227151 157486 227160
rect 157432 227122 157484 227128
rect 157154 226264 157210 226273
rect 157154 226199 157210 226208
rect 157168 226012 157196 226199
rect 157340 226024 157392 226030
rect 157168 225984 157340 226012
rect 157340 225966 157392 225972
rect 157812 225865 157840 229758
rect 156602 225856 156658 225865
rect 156602 225791 156658 225800
rect 157798 225856 157854 225865
rect 157798 225791 157854 225800
rect 156616 225690 156644 225791
rect 156604 225684 156656 225690
rect 156604 225626 156656 225632
rect 157340 225616 157392 225622
rect 157168 225564 157340 225570
rect 157168 225558 157392 225564
rect 157168 225542 157380 225558
rect 157168 225457 157196 225542
rect 157154 225448 157210 225457
rect 157154 225383 157210 225392
rect 157248 224392 157300 224398
rect 157248 224334 157300 224340
rect 156420 223304 156472 223310
rect 156420 223246 156472 223252
rect 156432 222494 156460 223246
rect 156420 222488 156472 222494
rect 156420 222430 156472 222436
rect 156604 222488 156656 222494
rect 156604 222430 156656 222436
rect 156616 222222 156644 222430
rect 156604 222216 156656 222222
rect 156604 222158 156656 222164
rect 156144 220108 156196 220114
rect 156144 220050 156196 220056
rect 156512 219428 156564 219434
rect 156512 219370 156564 219376
rect 156524 219026 156552 219370
rect 156512 219020 156564 219026
rect 156512 218962 156564 218968
rect 157260 218618 157288 224334
rect 157524 220108 157576 220114
rect 157524 220050 157576 220056
rect 156696 218612 156748 218618
rect 156696 218554 156748 218560
rect 157248 218612 157300 218618
rect 157248 218554 157300 218560
rect 155006 217110 155080 217138
rect 155834 217246 155908 217274
rect 155006 216988 155034 217110
rect 155834 216988 155862 217246
rect 156708 217138 156736 218554
rect 157536 217274 157564 220050
rect 157996 219162 158024 229978
rect 158548 229634 158576 231676
rect 158916 231662 159206 231690
rect 158718 229664 158774 229673
rect 158536 229628 158588 229634
rect 158718 229599 158720 229608
rect 158536 229570 158588 229576
rect 158772 229599 158774 229608
rect 158720 229570 158772 229576
rect 158350 220960 158406 220969
rect 158350 220895 158406 220904
rect 157984 219156 158036 219162
rect 157984 219098 158036 219104
rect 158364 217274 158392 220895
rect 158916 220250 158944 231662
rect 159836 223582 159864 231676
rect 160006 228576 160062 228585
rect 160006 228511 160062 228520
rect 159824 223576 159876 223582
rect 159824 223518 159876 223524
rect 159364 223440 159416 223446
rect 159364 223382 159416 223388
rect 158904 220244 158956 220250
rect 158904 220186 158956 220192
rect 159376 218890 159404 223382
rect 159364 218884 159416 218890
rect 159364 218826 159416 218832
rect 159824 218884 159876 218890
rect 159824 218826 159876 218832
rect 159180 218612 159232 218618
rect 159180 218554 159232 218560
rect 156662 217110 156736 217138
rect 157490 217246 157564 217274
rect 158318 217246 158392 217274
rect 156662 216988 156690 217110
rect 157490 216988 157518 217246
rect 158318 216988 158346 217246
rect 159192 217138 159220 218554
rect 159836 217274 159864 218826
rect 160020 218618 160048 228511
rect 160480 224670 160508 231676
rect 161124 230178 161152 231676
rect 161294 230208 161350 230217
rect 161112 230172 161164 230178
rect 161294 230143 161296 230152
rect 161112 230114 161164 230120
rect 161348 230143 161350 230152
rect 161296 230114 161348 230120
rect 161768 229634 161796 231676
rect 161756 229628 161808 229634
rect 161756 229570 161808 229576
rect 161940 229628 161992 229634
rect 161940 229570 161992 229576
rect 160468 224664 160520 224670
rect 160468 224606 160520 224612
rect 161952 224398 161980 229570
rect 161940 224392 161992 224398
rect 161940 224334 161992 224340
rect 162124 223576 162176 223582
rect 162124 223518 162176 223524
rect 160836 222148 160888 222154
rect 160836 222090 160888 222096
rect 160190 218648 160246 218657
rect 160008 218612 160060 218618
rect 160190 218583 160192 218592
rect 160008 218554 160060 218560
rect 160244 218583 160246 218592
rect 160192 218554 160244 218560
rect 160848 217274 160876 222090
rect 161432 221776 161488 221785
rect 161432 221711 161434 221720
rect 161486 221711 161488 221720
rect 161572 221740 161624 221746
rect 161434 221682 161486 221688
rect 161572 221682 161624 221688
rect 161584 221626 161612 221682
rect 161446 221598 161612 221626
rect 161446 221338 161474 221598
rect 161756 221468 161808 221474
rect 161756 221410 161808 221416
rect 161434 221332 161486 221338
rect 161434 221274 161486 221280
rect 161768 221082 161796 221410
rect 161446 221054 161796 221082
rect 161446 220930 161474 221054
rect 161570 220960 161626 220969
rect 161434 220924 161486 220930
rect 161570 220895 161572 220904
rect 161434 220866 161486 220872
rect 161624 220895 161626 220904
rect 161572 220866 161624 220872
rect 162136 219026 162164 223518
rect 162412 223310 162440 231676
rect 162688 231674 163070 231690
rect 162676 231668 163070 231674
rect 162728 231662 163070 231668
rect 162676 231610 162728 231616
rect 163700 230042 163728 231676
rect 163688 230036 163740 230042
rect 163688 229978 163740 229984
rect 162584 229764 162636 229770
rect 162584 229706 162636 229712
rect 164056 229764 164108 229770
rect 164056 229706 164108 229712
rect 162596 229226 162624 229706
rect 162584 229220 162636 229226
rect 162584 229162 162636 229168
rect 162768 224664 162820 224670
rect 162768 224606 162820 224612
rect 162400 223304 162452 223310
rect 162400 223246 162452 223252
rect 162124 219020 162176 219026
rect 162124 218962 162176 218968
rect 162492 219020 162544 219026
rect 162492 218962 162544 218968
rect 161664 218068 161716 218074
rect 161664 218010 161716 218016
rect 159836 217246 160002 217274
rect 159146 217110 159220 217138
rect 159146 216988 159174 217110
rect 159974 216988 160002 217246
rect 160802 217246 160876 217274
rect 160802 216988 160830 217246
rect 161676 217138 161704 218010
rect 162504 217274 162532 218962
rect 162780 218074 162808 224606
rect 164068 219434 164096 229706
rect 164344 221338 164372 231676
rect 164988 222630 165016 231676
rect 165632 224534 165660 231676
rect 166276 230178 166304 231676
rect 166552 231662 166934 231690
rect 167196 231662 167578 231690
rect 167840 231662 168222 231690
rect 168576 231662 168866 231690
rect 166264 230172 166316 230178
rect 166264 230114 166316 230120
rect 166354 228848 166410 228857
rect 166354 228783 166356 228792
rect 166408 228783 166410 228792
rect 166356 228754 166408 228760
rect 166552 227497 166580 231662
rect 166828 228682 166994 228698
rect 166828 228676 167006 228682
rect 166828 228670 166954 228676
rect 166828 228585 166856 228670
rect 166954 228618 167006 228624
rect 166814 228576 166870 228585
rect 166814 228511 166870 228520
rect 166538 227488 166594 227497
rect 166538 227423 166594 227432
rect 165620 224528 165672 224534
rect 165620 224470 165672 224476
rect 165528 224392 165580 224398
rect 165528 224334 165580 224340
rect 164976 222624 165028 222630
rect 164976 222566 165028 222572
rect 164332 221332 164384 221338
rect 164332 221274 164384 221280
rect 164240 220244 164292 220250
rect 164240 220186 164292 220192
rect 164252 220130 164280 220186
rect 163976 219406 164096 219434
rect 164160 220102 164280 220130
rect 163976 218074 164004 219406
rect 162768 218068 162820 218074
rect 162768 218010 162820 218016
rect 163320 218068 163372 218074
rect 163320 218010 163372 218016
rect 163964 218068 164016 218074
rect 163964 218010 164016 218016
rect 161630 217110 161704 217138
rect 162458 217246 162532 217274
rect 161630 216988 161658 217110
rect 162458 216988 162486 217246
rect 163332 217138 163360 218010
rect 164160 217274 164188 220102
rect 165540 218074 165568 224334
rect 166264 223032 166316 223038
rect 166264 222974 166316 222980
rect 166448 223032 166500 223038
rect 166448 222974 166500 222980
rect 166276 222766 166304 222974
rect 166264 222760 166316 222766
rect 166264 222702 166316 222708
rect 166460 222630 166488 222974
rect 166448 222624 166500 222630
rect 166448 222566 166500 222572
rect 166632 222624 166684 222630
rect 166632 222566 166684 222572
rect 166080 222148 166132 222154
rect 166080 222090 166132 222096
rect 166092 221202 166120 222090
rect 166080 221196 166132 221202
rect 166080 221138 166132 221144
rect 166644 219434 166672 222566
rect 167196 221746 167224 231662
rect 167366 229256 167422 229265
rect 167366 229191 167422 229200
rect 167380 229090 167408 229191
rect 167368 229084 167420 229090
rect 167368 229026 167420 229032
rect 167552 229084 167604 229090
rect 167552 229026 167604 229032
rect 167564 228857 167592 229026
rect 167550 228848 167606 228857
rect 167550 228783 167606 228792
rect 167840 224262 167868 231662
rect 167828 224256 167880 224262
rect 167828 224198 167880 224204
rect 168288 224256 168340 224262
rect 168288 224198 168340 224204
rect 167460 222012 167512 222018
rect 167460 221954 167512 221960
rect 167184 221740 167236 221746
rect 167184 221682 167236 221688
rect 165804 219428 165856 219434
rect 165804 219370 165856 219376
rect 166276 219406 166672 219434
rect 164976 218068 165028 218074
rect 164976 218010 165028 218016
rect 165528 218068 165580 218074
rect 165528 218010 165580 218016
rect 163286 217110 163360 217138
rect 164114 217246 164188 217274
rect 163286 216988 163314 217110
rect 164114 216988 164142 217246
rect 164988 217138 165016 218010
rect 165816 217138 165844 219370
rect 166276 218482 166304 219406
rect 166632 219156 166684 219162
rect 166632 219098 166684 219104
rect 166264 218476 166316 218482
rect 166264 218418 166316 218424
rect 166644 217138 166672 219098
rect 167472 217274 167500 221954
rect 167642 221776 167698 221785
rect 167642 221711 167644 221720
rect 167696 221711 167698 221720
rect 167644 221682 167696 221688
rect 168300 217274 168328 224198
rect 168576 217326 168604 231662
rect 169496 229090 169524 231676
rect 169772 231662 170154 231690
rect 169484 229084 169536 229090
rect 169484 229026 169536 229032
rect 169390 227352 169446 227361
rect 169390 227287 169392 227296
rect 169444 227287 169446 227296
rect 169576 227316 169628 227322
rect 169392 227258 169444 227264
rect 169576 227258 169628 227264
rect 169588 218074 169616 227258
rect 169772 221746 169800 231662
rect 170784 231538 170812 231676
rect 170772 231532 170824 231538
rect 170772 231474 170824 231480
rect 171428 230926 171456 231676
rect 171704 231662 172086 231690
rect 171416 230920 171468 230926
rect 171416 230862 171468 230868
rect 170956 230036 171008 230042
rect 170956 229978 171008 229984
rect 169760 221740 169812 221746
rect 169760 221682 169812 221688
rect 170968 219434 170996 229978
rect 171704 227361 171732 231662
rect 171690 227352 171746 227361
rect 171690 227287 171746 227296
rect 172060 227316 172112 227322
rect 172060 227258 172112 227264
rect 172072 227202 172100 227258
rect 171520 227186 172100 227202
rect 171508 227180 172100 227186
rect 171560 227174 172100 227180
rect 171508 227122 171560 227128
rect 171784 223304 171836 223310
rect 171784 223246 171836 223252
rect 171600 221740 171652 221746
rect 171600 221682 171652 221688
rect 170784 219406 170996 219434
rect 170784 218074 170812 219406
rect 170954 219328 171010 219337
rect 170954 219263 170956 219272
rect 171008 219263 171010 219272
rect 170956 219234 171008 219240
rect 170956 218476 171008 218482
rect 170956 218418 171008 218424
rect 169116 218068 169168 218074
rect 169116 218010 169168 218016
rect 169576 218068 169628 218074
rect 169576 218010 169628 218016
rect 169944 218068 169996 218074
rect 169944 218010 169996 218016
rect 170772 218068 170824 218074
rect 170772 218010 170824 218016
rect 164942 217110 165016 217138
rect 165770 217110 165844 217138
rect 166598 217110 166672 217138
rect 167426 217246 167500 217274
rect 168254 217246 168328 217274
rect 168564 217320 168616 217326
rect 168564 217262 168616 217268
rect 164942 216988 164970 217110
rect 165770 216988 165798 217110
rect 166598 216988 166626 217110
rect 167426 216988 167454 217246
rect 168254 216988 168282 217246
rect 169128 217138 169156 218010
rect 169956 217138 169984 218010
rect 170968 217274 170996 218418
rect 171612 217274 171640 221682
rect 171796 219337 171824 223246
rect 172716 222154 172744 231676
rect 172992 231662 173374 231690
rect 174018 231662 174216 231690
rect 172992 224942 173020 231662
rect 173164 228812 173216 228818
rect 173164 228754 173216 228760
rect 172980 224936 173032 224942
rect 172980 224878 173032 224884
rect 172704 222148 172756 222154
rect 172704 222090 172756 222096
rect 171782 219328 171838 219337
rect 171782 219263 171838 219272
rect 173176 218074 173204 228754
rect 173348 223168 173400 223174
rect 173348 223110 173400 223116
rect 173532 223168 173584 223174
rect 173532 223110 173584 223116
rect 173360 222358 173388 223110
rect 173544 222766 173572 223110
rect 173532 222760 173584 222766
rect 173532 222702 173584 222708
rect 173900 222624 173952 222630
rect 173900 222566 173952 222572
rect 173348 222352 173400 222358
rect 173348 222294 173400 222300
rect 173912 222222 173940 222566
rect 173900 222216 173952 222222
rect 173900 222158 173952 222164
rect 173346 221912 173402 221921
rect 173346 221847 173348 221856
rect 173400 221847 173402 221856
rect 173532 221876 173584 221882
rect 173348 221818 173400 221824
rect 173532 221818 173584 221824
rect 173544 221338 173572 221818
rect 173532 221332 173584 221338
rect 173532 221274 173584 221280
rect 174188 219434 174216 231662
rect 174372 231662 174662 231690
rect 174372 229265 174400 231662
rect 174358 229256 174414 229265
rect 174358 229191 174414 229200
rect 174912 224936 174964 224942
rect 174912 224878 174964 224884
rect 174360 222148 174412 222154
rect 174360 222090 174412 222096
rect 174372 219434 174400 222090
rect 174096 219406 174216 219434
rect 174280 219406 174400 219434
rect 172428 218068 172480 218074
rect 172428 218010 172480 218016
rect 173164 218068 173216 218074
rect 173164 218010 173216 218016
rect 173348 218068 173400 218074
rect 173348 218010 173400 218016
rect 169082 217110 169156 217138
rect 169910 217110 169984 217138
rect 170738 217246 170996 217274
rect 171566 217246 171640 217274
rect 169082 216988 169110 217110
rect 169910 216988 169938 217110
rect 170738 216988 170766 217246
rect 171566 216988 171594 217246
rect 172440 217138 172468 218010
rect 173360 217274 173388 218010
rect 174096 217938 174124 219406
rect 174084 217932 174136 217938
rect 174084 217874 174136 217880
rect 174280 217274 174308 219406
rect 174728 218340 174780 218346
rect 174728 218282 174780 218288
rect 174740 218074 174768 218282
rect 174728 218068 174780 218074
rect 174728 218010 174780 218016
rect 174924 217274 174952 224878
rect 175292 220658 175320 231676
rect 175568 231662 175950 231690
rect 176212 231662 176594 231690
rect 175568 222630 175596 231662
rect 176212 224954 176240 231662
rect 176476 230172 176528 230178
rect 176476 230114 176528 230120
rect 175752 224926 176240 224954
rect 175556 222624 175608 222630
rect 175556 222566 175608 222572
rect 175752 222358 175780 224926
rect 175924 223440 175976 223446
rect 175924 223382 175976 223388
rect 175936 222630 175964 223382
rect 175924 222624 175976 222630
rect 175924 222566 175976 222572
rect 176108 222488 176160 222494
rect 176108 222430 176160 222436
rect 175740 222352 175792 222358
rect 175740 222294 175792 222300
rect 175924 222012 175976 222018
rect 175924 221954 175976 221960
rect 175936 221474 175964 221954
rect 175924 221468 175976 221474
rect 175924 221410 175976 221416
rect 175280 220652 175332 220658
rect 175280 220594 175332 220600
rect 176120 219434 176148 222430
rect 176290 220688 176346 220697
rect 176290 220623 176346 220632
rect 175740 219428 175792 219434
rect 175740 219370 175792 219376
rect 175936 219406 176148 219434
rect 175752 219026 175780 219370
rect 175740 219020 175792 219026
rect 175740 218962 175792 218968
rect 175740 218340 175792 218346
rect 175740 218282 175792 218288
rect 172394 217110 172468 217138
rect 173222 217246 173388 217274
rect 174050 217246 174308 217274
rect 174878 217246 174952 217274
rect 172394 216988 172422 217110
rect 173222 216988 173250 217246
rect 174050 216988 174078 217246
rect 174878 216988 174906 217246
rect 175752 217138 175780 218282
rect 175936 218210 175964 219406
rect 176304 218482 176332 220623
rect 176292 218476 176344 218482
rect 176292 218418 176344 218424
rect 175924 218204 175976 218210
rect 175924 218146 175976 218152
rect 176488 217274 176516 230114
rect 177224 227458 177252 231676
rect 177408 231662 177882 231690
rect 177212 227452 177264 227458
rect 177212 227394 177264 227400
rect 177408 221921 177436 231662
rect 178512 224806 178540 231676
rect 179156 230790 179184 231676
rect 179144 230784 179196 230790
rect 179144 230726 179196 230732
rect 179800 229090 179828 231676
rect 180444 229226 180472 231676
rect 180432 229220 180484 229226
rect 180432 229162 180484 229168
rect 179788 229084 179840 229090
rect 179788 229026 179840 229032
rect 180064 229084 180116 229090
rect 180064 229026 180116 229032
rect 178500 224800 178552 224806
rect 178500 224742 178552 224748
rect 178684 224800 178736 224806
rect 178684 224742 178736 224748
rect 177394 221912 177450 221921
rect 177394 221847 177450 221856
rect 177396 220652 177448 220658
rect 177396 220594 177448 220600
rect 176660 219020 176712 219026
rect 176660 218962 176712 218968
rect 176672 218074 176700 218962
rect 176660 218068 176712 218074
rect 176660 218010 176712 218016
rect 177408 217274 177436 220594
rect 178696 218210 178724 224742
rect 179328 224528 179380 224534
rect 179328 224470 179380 224476
rect 178684 218204 178736 218210
rect 178684 218146 178736 218152
rect 179052 218204 179104 218210
rect 179052 218146 179104 218152
rect 178224 218068 178276 218074
rect 178224 218010 178276 218016
rect 176488 217246 176562 217274
rect 175706 217110 175780 217138
rect 175706 216988 175734 217110
rect 176534 216988 176562 217246
rect 177362 217246 177436 217274
rect 177362 216988 177390 217246
rect 178236 217138 178264 218010
rect 179064 217138 179092 218146
rect 179340 218074 179368 224470
rect 180076 219298 180104 229026
rect 181088 223990 181116 231676
rect 181732 229094 181760 231676
rect 181732 229066 181852 229094
rect 181444 228676 181496 228682
rect 181444 228618 181496 228624
rect 181628 228676 181680 228682
rect 181628 228618 181680 228624
rect 181456 228138 181484 228618
rect 181260 228132 181312 228138
rect 181260 228074 181312 228080
rect 181444 228132 181496 228138
rect 181444 228074 181496 228080
rect 181272 228018 181300 228074
rect 181640 228018 181668 228618
rect 181272 227990 181668 228018
rect 181260 227452 181312 227458
rect 181260 227394 181312 227400
rect 181076 223984 181128 223990
rect 181076 223926 181128 223932
rect 180798 220960 180854 220969
rect 180798 220895 180854 220904
rect 180812 220810 180840 220895
rect 180766 220794 180840 220810
rect 180754 220788 180840 220794
rect 180806 220782 180840 220788
rect 181076 220788 181128 220794
rect 180754 220730 180806 220736
rect 181076 220730 181128 220736
rect 180890 220688 180946 220697
rect 180754 220652 180806 220658
rect 180890 220623 180892 220632
rect 180754 220594 180806 220600
rect 180944 220623 180946 220632
rect 180892 220594 180944 220600
rect 180766 220538 180794 220594
rect 180766 220510 180932 220538
rect 180904 219978 180932 220510
rect 180754 219972 180806 219978
rect 180754 219914 180806 219920
rect 180892 219972 180944 219978
rect 180892 219914 180944 219920
rect 180766 219858 180794 219914
rect 181088 219858 181116 220730
rect 180766 219830 181116 219858
rect 181272 219434 181300 227394
rect 181824 222630 181852 229066
rect 182376 227594 182404 231676
rect 182652 231662 183034 231690
rect 183678 231662 183876 231690
rect 182364 227588 182416 227594
rect 182364 227530 182416 227536
rect 181812 222624 181864 222630
rect 181812 222566 181864 222572
rect 182652 222154 182680 231662
rect 183376 229220 183428 229226
rect 183376 229162 183428 229168
rect 181444 222148 181496 222154
rect 181444 222090 181496 222096
rect 182640 222148 182692 222154
rect 182640 222090 182692 222096
rect 181456 221882 181484 222090
rect 181444 221876 181496 221882
rect 181444 221818 181496 221824
rect 181628 221876 181680 221882
rect 181628 221818 181680 221824
rect 181272 219428 181496 219434
rect 181272 219406 181444 219428
rect 181444 219370 181496 219376
rect 180064 219292 180116 219298
rect 180064 219234 180116 219240
rect 180248 219292 180300 219298
rect 180248 219234 180300 219240
rect 180260 219026 180288 219234
rect 180248 219020 180300 219026
rect 180248 218962 180300 218968
rect 179880 218476 179932 218482
rect 179880 218418 179932 218424
rect 179512 218340 179564 218346
rect 179512 218282 179564 218288
rect 179524 218074 179552 218282
rect 179328 218068 179380 218074
rect 179328 218010 179380 218016
rect 179512 218068 179564 218074
rect 179512 218010 179564 218016
rect 179892 217138 179920 218418
rect 180708 218340 180760 218346
rect 180708 218282 180760 218288
rect 180720 217138 180748 218282
rect 181640 217274 181668 221818
rect 183388 219434 183416 229162
rect 183848 223854 183876 231662
rect 184032 231662 184322 231690
rect 184032 225758 184060 231662
rect 184952 228954 184980 231676
rect 185136 231662 185610 231690
rect 185872 231662 186254 231690
rect 186608 231662 186898 231690
rect 184940 228948 184992 228954
rect 184940 228890 184992 228896
rect 184020 225752 184072 225758
rect 184020 225694 184072 225700
rect 184204 225752 184256 225758
rect 184204 225694 184256 225700
rect 183836 223848 183888 223854
rect 183836 223790 183888 223796
rect 183204 219406 183416 219434
rect 183836 219428 183888 219434
rect 182364 219020 182416 219026
rect 182364 218962 182416 218968
rect 178190 217110 178264 217138
rect 179018 217110 179092 217138
rect 179846 217110 179920 217138
rect 180674 217110 180748 217138
rect 181502 217246 181668 217274
rect 178190 216988 178218 217110
rect 179018 216988 179046 217110
rect 179846 216988 179874 217110
rect 180674 216988 180702 217110
rect 181502 216988 181530 217246
rect 182376 217138 182404 218962
rect 183204 217274 183232 219406
rect 183836 219370 183888 219376
rect 183848 218074 183876 219370
rect 184216 218754 184244 225694
rect 184848 223712 184900 223718
rect 184848 223654 184900 223660
rect 184664 223440 184716 223446
rect 184664 223382 184716 223388
rect 184204 218748 184256 218754
rect 184204 218690 184256 218696
rect 184676 218074 184704 223382
rect 183836 218068 183888 218074
rect 183836 218010 183888 218016
rect 184020 218068 184072 218074
rect 184020 218010 184072 218016
rect 184664 218068 184716 218074
rect 184664 218010 184716 218016
rect 182330 217110 182404 217138
rect 183158 217246 183232 217274
rect 182330 216988 182358 217110
rect 183158 216988 183186 217246
rect 184032 217138 184060 218010
rect 184860 217274 184888 223654
rect 185136 220969 185164 231662
rect 185872 229094 185900 231662
rect 185584 229084 185636 229090
rect 185872 229066 185992 229094
rect 185584 229026 185636 229032
rect 185400 228948 185452 228954
rect 185400 228890 185452 228896
rect 185412 228682 185440 228890
rect 185596 228682 185624 229026
rect 185400 228676 185452 228682
rect 185400 228618 185452 228624
rect 185584 228676 185636 228682
rect 185584 228618 185636 228624
rect 185400 227588 185452 227594
rect 185400 227530 185452 227536
rect 185412 226914 185440 227530
rect 185584 227316 185636 227322
rect 185584 227258 185636 227264
rect 185596 226914 185624 227258
rect 185400 226908 185452 226914
rect 185400 226850 185452 226856
rect 185584 226908 185636 226914
rect 185584 226850 185636 226856
rect 185412 224998 185808 225026
rect 185412 224534 185440 224998
rect 185780 224942 185808 224998
rect 185584 224936 185636 224942
rect 185584 224878 185636 224884
rect 185768 224936 185820 224942
rect 185768 224878 185820 224884
rect 185596 224534 185624 224878
rect 185400 224528 185452 224534
rect 185400 224470 185452 224476
rect 185584 224528 185636 224534
rect 185584 224470 185636 224476
rect 185964 223854 185992 229066
rect 186136 227452 186188 227458
rect 186136 227394 186188 227400
rect 185952 223848 186004 223854
rect 185952 223790 186004 223796
rect 185768 223168 185820 223174
rect 185768 223110 185820 223116
rect 185780 222766 185808 223110
rect 185768 222760 185820 222766
rect 185768 222702 185820 222708
rect 185122 220960 185178 220969
rect 185122 220895 185178 220904
rect 185950 220824 186006 220833
rect 185950 220759 186006 220768
rect 185964 218346 185992 220759
rect 185952 218340 186004 218346
rect 185952 218282 186004 218288
rect 186148 218074 186176 227394
rect 186608 223582 186636 231662
rect 187528 226778 187556 231676
rect 188172 230654 188200 231676
rect 188448 231662 188830 231690
rect 189092 231662 189474 231690
rect 188160 230648 188212 230654
rect 188160 230590 188212 230596
rect 187516 226772 187568 226778
rect 187516 226714 187568 226720
rect 186964 223848 187016 223854
rect 186964 223790 187016 223796
rect 186596 223576 186648 223582
rect 186596 223518 186648 223524
rect 186504 218748 186556 218754
rect 186504 218690 186556 218696
rect 185676 218068 185728 218074
rect 185676 218010 185728 218016
rect 186136 218068 186188 218074
rect 186136 218010 186188 218016
rect 183986 217110 184060 217138
rect 184814 217246 184888 217274
rect 183986 216988 184014 217110
rect 184814 216988 184842 217246
rect 185688 217138 185716 218010
rect 186516 217138 186544 218690
rect 186976 218618 187004 223790
rect 187332 223576 187384 223582
rect 187332 223518 187384 223524
rect 186964 218612 187016 218618
rect 186964 218554 187016 218560
rect 187344 217274 187372 223518
rect 188448 219434 188476 231662
rect 189092 229094 189120 231662
rect 189092 229066 189212 229094
rect 188896 222352 188948 222358
rect 188896 222294 188948 222300
rect 187988 219406 188476 219434
rect 187988 217462 188016 219406
rect 188712 218612 188764 218618
rect 188712 218554 188764 218560
rect 188160 218068 188212 218074
rect 188160 218010 188212 218016
rect 187976 217456 188028 217462
rect 187976 217398 188028 217404
rect 185642 217110 185716 217138
rect 186470 217110 186544 217138
rect 187298 217246 187372 217274
rect 185642 216988 185670 217110
rect 186470 216988 186498 217110
rect 187298 216988 187326 217246
rect 188172 217138 188200 218010
rect 188724 217274 188752 218554
rect 188908 218074 188936 222294
rect 188896 218068 188948 218074
rect 188896 218010 188948 218016
rect 189184 217598 189212 229066
rect 189724 229084 189776 229090
rect 189724 229026 189776 229032
rect 189736 219026 189764 229026
rect 190104 228954 190132 231676
rect 190656 231662 190762 231690
rect 191024 231662 191406 231690
rect 190656 229094 190684 231662
rect 190472 229066 190684 229094
rect 190092 228948 190144 228954
rect 190092 228890 190144 228896
rect 190000 226772 190052 226778
rect 190000 226714 190052 226720
rect 190012 219434 190040 226714
rect 190472 220946 190500 229066
rect 191024 222222 191052 231662
rect 192036 222630 192064 231676
rect 192484 229084 192536 229090
rect 192484 229026 192536 229032
rect 192496 227866 192524 229026
rect 192484 227860 192536 227866
rect 192484 227802 192536 227808
rect 192680 227594 192708 231676
rect 193324 230194 193352 231676
rect 193600 231662 193982 231690
rect 193324 230166 193444 230194
rect 193034 228984 193090 228993
rect 193034 228919 193090 228928
rect 192668 227588 192720 227594
rect 192668 227530 192720 227536
rect 192024 222624 192076 222630
rect 192024 222566 192076 222572
rect 191012 222216 191064 222222
rect 191012 222158 191064 222164
rect 191472 222148 191524 222154
rect 191472 222090 191524 222096
rect 190380 220918 190500 220946
rect 190380 220794 190408 220918
rect 190550 220824 190606 220833
rect 190368 220788 190420 220794
rect 190550 220759 190552 220768
rect 190368 220730 190420 220736
rect 190604 220759 190606 220768
rect 190552 220730 190604 220736
rect 190000 219428 190052 219434
rect 190000 219370 190052 219376
rect 189724 219020 189776 219026
rect 189724 218962 189776 218968
rect 190644 219020 190696 219026
rect 190644 218962 190696 218968
rect 189816 218340 189868 218346
rect 189816 218282 189868 218288
rect 189172 217592 189224 217598
rect 189172 217534 189224 217540
rect 188724 217246 188982 217274
rect 188126 217110 188200 217138
rect 188126 216988 188154 217110
rect 188954 216988 188982 217246
rect 189828 217138 189856 218282
rect 190656 217138 190684 218962
rect 191484 217274 191512 222090
rect 192300 219428 192352 219434
rect 192300 219370 192352 219376
rect 192312 218754 192340 219370
rect 192300 218748 192352 218754
rect 192300 218690 192352 218696
rect 192852 218748 192904 218754
rect 192852 218690 192904 218696
rect 192300 218068 192352 218074
rect 192300 218010 192352 218016
rect 189782 217110 189856 217138
rect 190610 217110 190684 217138
rect 191438 217246 191512 217274
rect 189782 216988 189810 217110
rect 190610 216988 190638 217110
rect 191438 216988 191466 217246
rect 192312 217138 192340 218010
rect 192864 217274 192892 218690
rect 193048 218074 193076 228919
rect 193416 221338 193444 230166
rect 193600 225486 193628 231662
rect 193588 225480 193640 225486
rect 193588 225422 193640 225428
rect 193772 225480 193824 225486
rect 193772 225422 193824 225428
rect 193404 221332 193456 221338
rect 193404 221274 193456 221280
rect 193784 219434 193812 225422
rect 194612 224126 194640 231676
rect 195058 229936 195114 229945
rect 195058 229871 195060 229880
rect 195112 229871 195114 229880
rect 195060 229842 195112 229848
rect 195256 229094 195284 231676
rect 195900 231402 195928 231676
rect 196176 231662 196558 231690
rect 196912 231662 197202 231690
rect 197372 231662 197846 231690
rect 198016 231662 198490 231690
rect 195888 231396 195940 231402
rect 195888 231338 195940 231344
rect 195428 229900 195480 229906
rect 195428 229842 195480 229848
rect 195072 229066 195284 229094
rect 195072 227866 195100 229066
rect 195244 228948 195296 228954
rect 195244 228890 195296 228896
rect 195256 228138 195284 228890
rect 195244 228132 195296 228138
rect 195244 228074 195296 228080
rect 195060 227860 195112 227866
rect 195060 227802 195112 227808
rect 195244 224936 195296 224942
rect 195244 224878 195296 224884
rect 195256 224126 195284 224878
rect 194600 224120 194652 224126
rect 194600 224062 194652 224068
rect 195244 224120 195296 224126
rect 195244 224062 195296 224068
rect 194508 223168 194560 223174
rect 194508 223110 194560 223116
rect 193600 219406 193812 219434
rect 193600 218618 193628 219406
rect 193588 218612 193640 218618
rect 193588 218554 193640 218560
rect 194520 218074 194548 223110
rect 195440 219434 195468 229842
rect 195610 228984 195666 228993
rect 195610 228919 195612 228928
rect 195664 228919 195666 228928
rect 195612 228890 195664 228896
rect 196176 225350 196204 231662
rect 196912 229945 196940 231662
rect 196898 229936 196954 229945
rect 196898 229871 196954 229880
rect 197372 226642 197400 231662
rect 198016 229094 198044 231662
rect 197648 229066 198044 229094
rect 197360 226636 197412 226642
rect 197360 226578 197412 226584
rect 196164 225344 196216 225350
rect 196164 225286 196216 225292
rect 196624 225344 196676 225350
rect 196624 225286 196676 225292
rect 195612 224936 195664 224942
rect 195612 224878 195664 224884
rect 195624 223718 195652 224878
rect 195612 223712 195664 223718
rect 195612 223654 195664 223660
rect 195888 223712 195940 223718
rect 195888 223654 195940 223660
rect 195256 219406 195468 219434
rect 195256 218346 195284 219406
rect 195612 218612 195664 218618
rect 195612 218554 195664 218560
rect 195244 218340 195296 218346
rect 195244 218282 195296 218288
rect 193036 218068 193088 218074
rect 193036 218010 193088 218016
rect 193956 218068 194008 218074
rect 193956 218010 194008 218016
rect 194508 218068 194560 218074
rect 194508 218010 194560 218016
rect 194784 218068 194836 218074
rect 194784 218010 194836 218016
rect 192864 217246 193122 217274
rect 192266 217110 192340 217138
rect 192266 216988 192294 217110
rect 193094 216988 193122 217246
rect 193968 217138 193996 218010
rect 194796 217138 194824 218010
rect 195624 217138 195652 218554
rect 195900 218074 195928 223654
rect 196636 218210 196664 225286
rect 197176 222624 197228 222630
rect 197176 222566 197228 222572
rect 196624 218204 196676 218210
rect 196624 218146 196676 218152
rect 195888 218068 195940 218074
rect 195888 218010 195940 218016
rect 196440 218068 196492 218074
rect 196440 218010 196492 218016
rect 196452 217138 196480 218010
rect 197188 217274 197216 222566
rect 197648 219842 197676 229066
rect 198004 225888 198056 225894
rect 198004 225830 198056 225836
rect 197636 219836 197688 219842
rect 197636 219778 197688 219784
rect 197820 219836 197872 219842
rect 197820 219778 197872 219784
rect 197832 219026 197860 219778
rect 197820 219020 197872 219026
rect 197820 218962 197872 218968
rect 198016 218618 198044 225830
rect 199120 225214 199148 231676
rect 199108 225208 199160 225214
rect 199108 225150 199160 225156
rect 199764 223310 199792 231676
rect 200408 229090 200436 231676
rect 201052 230518 201080 231676
rect 201040 230512 201092 230518
rect 201040 230454 201092 230460
rect 200396 229084 200448 229090
rect 200396 229026 200448 229032
rect 201408 229084 201460 229090
rect 201408 229026 201460 229032
rect 200120 228540 200172 228546
rect 200120 228482 200172 228488
rect 200304 228540 200356 228546
rect 200304 228482 200356 228488
rect 200132 227866 200160 228482
rect 200316 228002 200344 228482
rect 200304 227996 200356 228002
rect 200304 227938 200356 227944
rect 200120 227860 200172 227866
rect 200120 227802 200172 227808
rect 200028 227588 200080 227594
rect 200028 227530 200080 227536
rect 199752 223304 199804 223310
rect 199752 223246 199804 223252
rect 200040 218618 200068 227530
rect 201224 223984 201276 223990
rect 201224 223926 201276 223932
rect 201236 219434 201264 223926
rect 201236 219406 201356 219434
rect 200212 219020 200264 219026
rect 200212 218962 200264 218968
rect 198004 218612 198056 218618
rect 198004 218554 198056 218560
rect 198924 218612 198976 218618
rect 198924 218554 198976 218560
rect 200028 218612 200080 218618
rect 200028 218554 200080 218560
rect 198096 218340 198148 218346
rect 198096 218282 198148 218288
rect 197188 217246 197262 217274
rect 193922 217110 193996 217138
rect 194750 217110 194824 217138
rect 195578 217110 195652 217138
rect 196406 217110 196480 217138
rect 193922 216988 193950 217110
rect 194750 216988 194778 217110
rect 195578 216988 195606 217110
rect 196406 216988 196434 217110
rect 197234 216988 197262 217246
rect 198108 217138 198136 218282
rect 198936 217138 198964 218554
rect 200224 218210 200252 218962
rect 200672 218340 200724 218346
rect 200672 218282 200724 218288
rect 200684 218226 200712 218282
rect 199752 218204 199804 218210
rect 199752 218146 199804 218152
rect 200212 218204 200264 218210
rect 200212 218146 200264 218152
rect 200408 218198 200712 218226
rect 199764 217138 199792 218146
rect 200408 218074 200436 218198
rect 200396 218068 200448 218074
rect 200396 218010 200448 218016
rect 200580 218068 200632 218074
rect 200580 218010 200632 218016
rect 200592 217138 200620 218010
rect 201328 217274 201356 219406
rect 201420 218090 201448 229026
rect 201696 225078 201724 231676
rect 202340 230314 202368 231676
rect 202328 230308 202380 230314
rect 202328 230250 202380 230256
rect 202984 226506 203012 231676
rect 203168 231662 203642 231690
rect 202972 226500 203024 226506
rect 202972 226442 203024 226448
rect 201684 225072 201736 225078
rect 201684 225014 201736 225020
rect 202236 225072 202288 225078
rect 202236 225014 202288 225020
rect 201420 218074 201540 218090
rect 201420 218068 201552 218074
rect 201420 218062 201500 218068
rect 201500 218010 201552 218016
rect 202248 217274 202276 225014
rect 203168 219706 203196 231662
rect 203524 226636 203576 226642
rect 203524 226578 203576 226584
rect 203156 219700 203208 219706
rect 203156 219642 203208 219648
rect 203536 218890 203564 226578
rect 204272 226302 204300 231676
rect 204640 231662 204930 231690
rect 204640 229094 204668 231662
rect 204548 229066 204668 229094
rect 204260 226296 204312 226302
rect 204260 226238 204312 226244
rect 204548 224806 204576 229066
rect 205560 228274 205588 231676
rect 205928 231662 206218 231690
rect 206480 231662 206862 231690
rect 205548 228268 205600 228274
rect 205548 228210 205600 228216
rect 205732 228268 205784 228274
rect 205732 228210 205784 228216
rect 205744 228154 205772 228210
rect 205468 228126 205772 228154
rect 204810 227624 204866 227633
rect 204810 227559 204866 227568
rect 204824 227458 204852 227559
rect 204812 227452 204864 227458
rect 204812 227394 204864 227400
rect 204536 224800 204588 224806
rect 204536 224742 204588 224748
rect 204720 224800 204772 224806
rect 204720 224742 204772 224748
rect 204732 224126 204760 224742
rect 204720 224120 204772 224126
rect 204720 224062 204772 224068
rect 204904 224120 204956 224126
rect 204904 224062 204956 224068
rect 204916 223718 204944 224062
rect 204904 223712 204956 223718
rect 204904 223654 204956 223660
rect 204720 223304 204772 223310
rect 204720 223246 204772 223252
rect 204732 222766 204760 223246
rect 204904 223168 204956 223174
rect 204904 223110 204956 223116
rect 204916 222766 204944 223110
rect 204720 222760 204772 222766
rect 204720 222702 204772 222708
rect 204904 222760 204956 222766
rect 204904 222702 204956 222708
rect 204168 221332 204220 221338
rect 204168 221274 204220 221280
rect 203892 219564 203944 219570
rect 203892 219506 203944 219512
rect 203524 218884 203576 218890
rect 203524 218826 203576 218832
rect 203064 218068 203116 218074
rect 203064 218010 203116 218016
rect 201328 217246 201402 217274
rect 198062 217110 198136 217138
rect 198890 217110 198964 217138
rect 199718 217110 199792 217138
rect 200546 217110 200620 217138
rect 198062 216988 198090 217110
rect 198890 216988 198918 217110
rect 199718 216988 199746 217110
rect 200546 216988 200574 217110
rect 201374 216988 201402 217246
rect 202202 217246 202276 217274
rect 202202 216988 202230 217246
rect 203076 217138 203104 218010
rect 203904 217274 203932 219506
rect 204180 218210 204208 221274
rect 204720 218612 204772 218618
rect 204720 218554 204772 218560
rect 204168 218204 204220 218210
rect 204168 218146 204220 218152
rect 203030 217110 203104 217138
rect 203858 217246 203932 217274
rect 203030 216988 203058 217110
rect 203858 216988 203886 217246
rect 204732 217138 204760 218554
rect 204904 218476 204956 218482
rect 204904 218418 204956 218424
rect 204916 218210 204944 218418
rect 204904 218204 204956 218210
rect 204904 218146 204956 218152
rect 205468 217274 205496 228126
rect 205638 227624 205694 227633
rect 205638 227559 205640 227568
rect 205692 227559 205694 227568
rect 205640 227530 205692 227536
rect 205928 221610 205956 231662
rect 206284 230308 206336 230314
rect 206284 230250 206336 230256
rect 205916 221604 205968 221610
rect 205916 221546 205968 221552
rect 206296 218074 206324 230250
rect 206480 221066 206508 231662
rect 207492 222494 207520 231676
rect 208136 227050 208164 231676
rect 208596 231662 208794 231690
rect 208124 227044 208176 227050
rect 208124 226986 208176 226992
rect 208124 226296 208176 226302
rect 208124 226238 208176 226244
rect 207480 222488 207532 222494
rect 207480 222430 207532 222436
rect 207664 222488 207716 222494
rect 207664 222430 207716 222436
rect 206468 221060 206520 221066
rect 206468 221002 206520 221008
rect 206468 218884 206520 218890
rect 206468 218826 206520 218832
rect 206284 218068 206336 218074
rect 206284 218010 206336 218016
rect 206480 217274 206508 218826
rect 207676 218618 207704 222430
rect 207664 218612 207716 218618
rect 207664 218554 207716 218560
rect 208136 218074 208164 226238
rect 208400 221604 208452 221610
rect 208400 221546 208452 221552
rect 208412 219434 208440 221546
rect 208596 219706 208624 231662
rect 209424 226166 209452 231676
rect 210068 229498 210096 231676
rect 210252 231662 210726 231690
rect 210056 229492 210108 229498
rect 210056 229434 210108 229440
rect 210252 227866 210280 231662
rect 211356 229094 211384 231676
rect 211264 229066 211384 229094
rect 211632 231662 212014 231690
rect 210424 227996 210476 228002
rect 210424 227938 210476 227944
rect 210240 227860 210292 227866
rect 210240 227802 210292 227808
rect 209412 226160 209464 226166
rect 209412 226102 209464 226108
rect 209688 226160 209740 226166
rect 209688 226102 209740 226108
rect 208584 219700 208636 219706
rect 208584 219642 208636 219648
rect 208320 219406 208440 219434
rect 207204 218068 207256 218074
rect 207204 218010 207256 218016
rect 208124 218068 208176 218074
rect 208124 218010 208176 218016
rect 205468 217246 205542 217274
rect 204686 217110 204760 217138
rect 204686 216988 204714 217110
rect 205514 216988 205542 217246
rect 206342 217246 206508 217274
rect 206342 216988 206370 217246
rect 207216 217138 207244 218010
rect 208320 217274 208348 219406
rect 209700 219162 209728 226102
rect 210436 219858 210464 227938
rect 211264 220522 211292 229066
rect 211436 223304 211488 223310
rect 211436 223246 211488 223252
rect 211448 222902 211476 223246
rect 211632 223174 211660 231662
rect 212172 226500 212224 226506
rect 212172 226442 212224 226448
rect 211620 223168 211672 223174
rect 211620 223110 211672 223116
rect 211436 222896 211488 222902
rect 211436 222838 211488 222844
rect 211804 222896 211856 222902
rect 211804 222838 211856 222844
rect 211252 220516 211304 220522
rect 211252 220458 211304 220464
rect 210344 219830 210464 219858
rect 208492 219156 208544 219162
rect 208492 219098 208544 219104
rect 208860 219156 208912 219162
rect 208860 219098 208912 219104
rect 209688 219156 209740 219162
rect 209688 219098 209740 219104
rect 208504 218482 208532 219098
rect 208492 218476 208544 218482
rect 208492 218418 208544 218424
rect 207170 217110 207244 217138
rect 207998 217246 208348 217274
rect 207170 216988 207198 217110
rect 207998 216988 208026 217246
rect 208872 217138 208900 219098
rect 209688 218340 209740 218346
rect 209688 218282 209740 218288
rect 209700 217138 209728 218282
rect 210344 218210 210372 219830
rect 210516 219700 210568 219706
rect 210516 219642 210568 219648
rect 210332 218204 210384 218210
rect 210332 218146 210384 218152
rect 210528 217274 210556 219642
rect 211816 218482 211844 222838
rect 211804 218476 211856 218482
rect 211804 218418 211856 218424
rect 211344 218204 211396 218210
rect 211344 218146 211396 218152
rect 208826 217110 208900 217138
rect 209654 217110 209728 217138
rect 210482 217246 210556 217274
rect 208826 216988 208854 217110
rect 209654 216988 209682 217110
rect 210482 216988 210510 217246
rect 211356 217138 211384 218146
rect 212184 217274 212212 226442
rect 212644 225758 212672 231676
rect 213092 230444 213144 230450
rect 213092 230386 213144 230392
rect 213104 229094 213132 230386
rect 213288 229094 213316 231676
rect 213946 231662 214144 231690
rect 213104 229066 213224 229094
rect 213288 229066 213408 229094
rect 212632 225752 212684 225758
rect 212632 225694 212684 225700
rect 213000 218476 213052 218482
rect 213000 218418 213052 218424
rect 211310 217110 211384 217138
rect 212138 217246 212212 217274
rect 211310 216988 211338 217110
rect 212138 216988 212166 217246
rect 213012 217138 213040 218418
rect 213196 218346 213224 229066
rect 213380 227730 213408 229066
rect 213368 227724 213420 227730
rect 213368 227666 213420 227672
rect 213828 227724 213880 227730
rect 213828 227666 213880 227672
rect 213644 220380 213696 220386
rect 213644 220322 213696 220328
rect 213656 219978 213684 220322
rect 213644 219972 213696 219978
rect 213644 219914 213696 219920
rect 213184 218340 213236 218346
rect 213184 218282 213236 218288
rect 213840 217274 213868 227666
rect 214116 220522 214144 231662
rect 214576 229094 214604 231676
rect 215220 229362 215248 231676
rect 215208 229356 215260 229362
rect 215208 229298 215260 229304
rect 214392 229066 214604 229094
rect 214392 225622 214420 229066
rect 215864 228410 215892 231676
rect 216232 231662 216522 231690
rect 215852 228404 215904 228410
rect 215852 228346 215904 228352
rect 214564 227588 214616 227594
rect 214564 227530 214616 227536
rect 214748 227588 214800 227594
rect 214748 227530 214800 227536
rect 214576 227050 214604 227530
rect 214564 227044 214616 227050
rect 214564 226986 214616 226992
rect 214760 226506 214788 227530
rect 214748 226500 214800 226506
rect 214748 226442 214800 226448
rect 214380 225616 214432 225622
rect 214380 225558 214432 225564
rect 215208 225616 215260 225622
rect 215208 225558 215260 225564
rect 214380 223304 214432 223310
rect 214380 223246 214432 223252
rect 214392 223122 214420 223246
rect 214392 223094 214880 223122
rect 214852 223038 214880 223094
rect 214840 223032 214892 223038
rect 214840 222974 214892 222980
rect 214104 220516 214156 220522
rect 214104 220458 214156 220464
rect 214288 220516 214340 220522
rect 214288 220458 214340 220464
rect 214300 220114 214328 220458
rect 214288 220108 214340 220114
rect 214288 220050 214340 220056
rect 214748 219972 214800 219978
rect 214748 219914 214800 219920
rect 214760 219570 214788 219914
rect 214748 219564 214800 219570
rect 214748 219506 214800 219512
rect 214288 218612 214340 218618
rect 214748 218612 214800 218618
rect 214288 218554 214340 218560
rect 214484 218572 214748 218600
rect 214300 218346 214328 218554
rect 214288 218340 214340 218346
rect 214288 218282 214340 218288
rect 214484 218210 214512 218572
rect 214748 218554 214800 218560
rect 214472 218204 214524 218210
rect 214472 218146 214524 218152
rect 215220 218074 215248 225558
rect 216232 223038 216260 231662
rect 216496 228404 216548 228410
rect 216496 228346 216548 228352
rect 216220 223032 216272 223038
rect 216220 222974 216272 222980
rect 215944 222896 215996 222902
rect 215944 222838 215996 222844
rect 215956 219298 215984 222838
rect 215944 219292 215996 219298
rect 215944 219234 215996 219240
rect 216312 218340 216364 218346
rect 216312 218282 216364 218288
rect 214656 218068 214708 218074
rect 214656 218010 214708 218016
rect 215208 218068 215260 218074
rect 215208 218010 215260 218016
rect 215484 218068 215536 218074
rect 215484 218010 215536 218016
rect 212966 217110 213040 217138
rect 213794 217246 213868 217274
rect 212966 216988 212994 217110
rect 213794 216988 213822 217246
rect 214668 217138 214696 218010
rect 215496 217138 215524 218010
rect 216324 217138 216352 218282
rect 216508 218074 216536 228346
rect 217152 226030 217180 231676
rect 217140 226024 217192 226030
rect 217140 225966 217192 225972
rect 217796 223854 217824 231676
rect 218440 226914 218468 231676
rect 218716 231662 219098 231690
rect 219544 231662 219742 231690
rect 218428 226908 218480 226914
rect 218428 226850 218480 226856
rect 217784 223848 217836 223854
rect 217784 223790 217836 223796
rect 218716 220522 218744 231662
rect 219164 227316 219216 227322
rect 219164 227258 219216 227264
rect 219176 226642 219204 227258
rect 219348 226908 219400 226914
rect 219348 226850 219400 226856
rect 219164 226636 219216 226642
rect 219164 226578 219216 226584
rect 218704 220516 218756 220522
rect 218704 220458 218756 220464
rect 217140 219700 217192 219706
rect 217140 219642 217192 219648
rect 216496 218068 216548 218074
rect 216496 218010 216548 218016
rect 217152 217274 217180 219642
rect 219360 219162 219388 226850
rect 219544 223310 219572 231662
rect 220372 229634 220400 231676
rect 220360 229628 220412 229634
rect 220360 229570 220412 229576
rect 220268 229492 220320 229498
rect 220268 229434 220320 229440
rect 220084 227316 220136 227322
rect 220084 227258 220136 227264
rect 220096 227050 220124 227258
rect 220084 227044 220136 227050
rect 220084 226986 220136 226992
rect 220280 224954 220308 229434
rect 221016 228546 221044 231676
rect 221292 231662 221674 231690
rect 221004 228540 221056 228546
rect 221004 228482 221056 228488
rect 220452 227044 220504 227050
rect 220452 226986 220504 226992
rect 220464 226506 220492 226986
rect 220452 226500 220504 226506
rect 220452 226442 220504 226448
rect 220096 224926 220308 224954
rect 219532 223304 219584 223310
rect 219532 223246 219584 223252
rect 219808 221060 219860 221066
rect 219808 221002 219860 221008
rect 219624 219292 219676 219298
rect 219624 219234 219676 219240
rect 218796 219156 218848 219162
rect 218796 219098 218848 219104
rect 219348 219156 219400 219162
rect 219348 219098 219400 219104
rect 217968 218204 218020 218210
rect 217968 218146 218020 218152
rect 214622 217110 214696 217138
rect 215450 217110 215524 217138
rect 216278 217110 216352 217138
rect 217106 217246 217180 217274
rect 214622 216988 214650 217110
rect 215450 216988 215478 217110
rect 216278 216988 216306 217110
rect 217106 216988 217134 217246
rect 217980 217138 218008 218146
rect 218808 217138 218836 219098
rect 219636 217138 219664 219234
rect 219820 218618 219848 221002
rect 219808 218612 219860 218618
rect 219808 218554 219860 218560
rect 220096 218074 220124 224926
rect 221292 221202 221320 231662
rect 221832 226500 221884 226506
rect 221832 226442 221884 226448
rect 221280 221196 221332 221202
rect 221280 221138 221332 221144
rect 220452 220516 220504 220522
rect 220452 220458 220504 220464
rect 220084 218068 220136 218074
rect 220084 218010 220136 218016
rect 220464 217274 220492 220458
rect 221844 218074 221872 226442
rect 222016 226024 222068 226030
rect 222016 225966 222068 225972
rect 221280 218068 221332 218074
rect 221280 218010 221332 218016
rect 221832 218068 221884 218074
rect 221832 218010 221884 218016
rect 217934 217110 218008 217138
rect 218762 217110 218836 217138
rect 219590 217110 219664 217138
rect 220418 217246 220492 217274
rect 217934 216988 217962 217110
rect 218762 216988 218790 217110
rect 219590 216988 219618 217110
rect 220418 216988 220446 217246
rect 221292 217138 221320 218010
rect 222028 217274 222056 225966
rect 222304 220930 222332 231676
rect 222948 227050 222976 231676
rect 222936 227044 222988 227050
rect 222936 226986 222988 226992
rect 223592 226642 223620 231676
rect 223776 231662 224250 231690
rect 224512 231662 224894 231690
rect 223580 226636 223632 226642
rect 223580 226578 223632 226584
rect 222752 221196 222804 221202
rect 222752 221138 222804 221144
rect 222292 220924 222344 220930
rect 222292 220866 222344 220872
rect 222764 218210 222792 221138
rect 223776 220250 223804 231662
rect 224512 224954 224540 231662
rect 225524 229770 225552 231676
rect 225512 229764 225564 229770
rect 225512 229706 225564 229712
rect 225604 229492 225656 229498
rect 225604 229434 225656 229440
rect 224776 228404 224828 228410
rect 224776 228346 224828 228352
rect 224052 224926 224540 224954
rect 224052 224670 224080 224926
rect 224592 224800 224644 224806
rect 224592 224742 224644 224748
rect 224040 224664 224092 224670
rect 224040 224606 224092 224612
rect 224224 220652 224276 220658
rect 224224 220594 224276 220600
rect 223764 220244 223816 220250
rect 223764 220186 223816 220192
rect 224236 219570 224264 220594
rect 224408 220380 224460 220386
rect 224408 220322 224460 220328
rect 224420 219706 224448 220322
rect 224408 219700 224460 219706
rect 224408 219642 224460 219648
rect 224224 219564 224276 219570
rect 224224 219506 224276 219512
rect 224408 219428 224460 219434
rect 224408 219370 224460 219376
rect 224224 219156 224276 219162
rect 224224 219098 224276 219104
rect 224236 218482 224264 219098
rect 224420 218482 224448 219370
rect 224224 218476 224276 218482
rect 224224 218418 224276 218424
rect 224408 218476 224460 218482
rect 224408 218418 224460 218424
rect 222752 218204 222804 218210
rect 222752 218146 222804 218152
rect 222936 218204 222988 218210
rect 222936 218146 222988 218152
rect 222028 217246 222102 217274
rect 221246 217110 221320 217138
rect 221246 216988 221274 217110
rect 222074 216988 222102 217246
rect 222948 217138 222976 218146
rect 224604 218074 224632 224742
rect 223764 218068 223816 218074
rect 223764 218010 223816 218016
rect 224592 218068 224644 218074
rect 224592 218010 224644 218016
rect 223776 217138 223804 218010
rect 224788 217274 224816 228346
rect 225616 218210 225644 229434
rect 226168 228682 226196 231676
rect 226536 231662 226826 231690
rect 226156 228676 226208 228682
rect 226156 228618 226208 228624
rect 226340 228676 226392 228682
rect 226340 228618 226392 228624
rect 226352 228562 226380 228618
rect 226168 228534 226380 228562
rect 225972 218612 226024 218618
rect 225972 218554 226024 218560
rect 225604 218204 225656 218210
rect 225604 218146 225656 218152
rect 225420 218068 225472 218074
rect 225420 218010 225472 218016
rect 222902 217110 222976 217138
rect 223730 217110 223804 217138
rect 224558 217246 224816 217274
rect 222902 216988 222930 217110
rect 223730 216988 223758 217110
rect 224558 216988 224586 217246
rect 225432 217138 225460 218010
rect 225984 217274 226012 218554
rect 226168 218074 226196 228534
rect 226536 221474 226564 231662
rect 227456 224398 227484 231676
rect 227444 224392 227496 224398
rect 227444 224334 227496 224340
rect 228100 223174 228128 231676
rect 228744 227050 228772 231676
rect 229296 231662 229402 231690
rect 228732 227044 228784 227050
rect 228732 226986 228784 226992
rect 228916 227044 228968 227050
rect 228916 226986 228968 226992
rect 228928 226506 228956 226986
rect 228916 226500 228968 226506
rect 228916 226442 228968 226448
rect 228732 224392 228784 224398
rect 228732 224334 228784 224340
rect 228088 223168 228140 223174
rect 228088 223110 228140 223116
rect 226524 221468 226576 221474
rect 226524 221410 226576 221416
rect 227904 221468 227956 221474
rect 227904 221410 227956 221416
rect 227076 219700 227128 219706
rect 227076 219642 227128 219648
rect 226156 218068 226208 218074
rect 226156 218010 226208 218016
rect 227088 217274 227116 219642
rect 227916 217274 227944 221410
rect 228744 217274 228772 224334
rect 229296 219570 229324 231662
rect 230032 224262 230060 231676
rect 230676 230042 230704 231676
rect 230664 230036 230716 230042
rect 230664 229978 230716 229984
rect 230480 229900 230532 229906
rect 230480 229842 230532 229848
rect 230020 224256 230072 224262
rect 230020 224198 230072 224204
rect 230492 223666 230520 229842
rect 231320 228818 231348 231676
rect 231978 231662 232176 231690
rect 231308 228812 231360 228818
rect 231308 228754 231360 228760
rect 231032 226636 231084 226642
rect 231032 226578 231084 226584
rect 230400 223638 230520 223666
rect 230204 223032 230256 223038
rect 230204 222974 230256 222980
rect 229284 219564 229336 219570
rect 229284 219506 229336 219512
rect 230216 219434 230244 222974
rect 230400 219434 230428 223638
rect 229560 219428 229612 219434
rect 230216 219406 230336 219434
rect 230400 219428 230532 219434
rect 230400 219406 230480 219428
rect 229560 219370 229612 219376
rect 225984 217246 226242 217274
rect 225386 217110 225460 217138
rect 225386 216988 225414 217110
rect 226214 216988 226242 217246
rect 227042 217246 227116 217274
rect 227870 217246 227944 217274
rect 228698 217246 228772 217274
rect 227042 216988 227070 217246
rect 227870 216988 227898 217246
rect 228698 216988 228726 217246
rect 229572 217138 229600 219370
rect 230308 217274 230336 219406
rect 230480 219370 230532 219376
rect 231044 218482 231072 226578
rect 231676 224256 231728 224262
rect 231676 224198 231728 224204
rect 231032 218476 231084 218482
rect 231032 218418 231084 218424
rect 231688 218074 231716 224198
rect 232148 222018 232176 231662
rect 232332 231662 232622 231690
rect 232136 222012 232188 222018
rect 232136 221954 232188 221960
rect 232332 221746 232360 231662
rect 233252 229094 233280 231676
rect 233700 229900 233752 229906
rect 233700 229842 233752 229848
rect 233712 229498 233740 229842
rect 233700 229492 233752 229498
rect 233700 229434 233752 229440
rect 233252 229066 233372 229094
rect 233148 223848 233200 223854
rect 233148 223790 233200 223796
rect 232320 221740 232372 221746
rect 232320 221682 232372 221688
rect 232872 218340 232924 218346
rect 232872 218282 232924 218288
rect 231216 218068 231268 218074
rect 231216 218010 231268 218016
rect 231676 218068 231728 218074
rect 231676 218010 231728 218016
rect 232044 218068 232096 218074
rect 232044 218010 232096 218016
rect 230308 217246 230382 217274
rect 229526 217110 229600 217138
rect 229526 216988 229554 217110
rect 230354 216988 230382 217246
rect 231228 217138 231256 218010
rect 232056 217138 232084 218010
rect 232884 217274 232912 218282
rect 233160 218074 233188 223790
rect 233344 222902 233372 229066
rect 233896 226778 233924 231676
rect 234172 231662 234554 231690
rect 233884 226772 233936 226778
rect 233884 226714 233936 226720
rect 233332 222896 233384 222902
rect 233332 222838 233384 222844
rect 233700 222012 233752 222018
rect 233700 221954 233752 221960
rect 233148 218068 233200 218074
rect 233148 218010 233200 218016
rect 233712 217274 233740 221954
rect 234172 220250 234200 231662
rect 235184 224534 235212 231676
rect 235828 230178 235856 231676
rect 235816 230172 235868 230178
rect 235816 230114 235868 230120
rect 235816 227180 235868 227186
rect 235816 227122 235868 227128
rect 235172 224528 235224 224534
rect 235172 224470 235224 224476
rect 234528 222896 234580 222902
rect 234528 222838 234580 222844
rect 234160 220244 234212 220250
rect 234160 220186 234212 220192
rect 234540 217274 234568 222838
rect 235828 218074 235856 227122
rect 236472 225350 236500 231676
rect 236656 231662 237130 231690
rect 236460 225344 236512 225350
rect 236460 225286 236512 225292
rect 236656 220794 236684 231662
rect 237288 225752 237340 225758
rect 237288 225694 237340 225700
rect 236644 220788 236696 220794
rect 236644 220730 236696 220736
rect 237012 220244 237064 220250
rect 237012 220186 237064 220192
rect 235356 218068 235408 218074
rect 235356 218010 235408 218016
rect 235816 218068 235868 218074
rect 235816 218010 235868 218016
rect 236184 218068 236236 218074
rect 236184 218010 236236 218016
rect 231182 217110 231256 217138
rect 232010 217110 232084 217138
rect 232838 217246 232912 217274
rect 233666 217246 233740 217274
rect 234494 217246 234568 217274
rect 231182 216988 231210 217110
rect 232010 216988 232038 217110
rect 232838 216988 232866 217246
rect 233666 216988 233694 217246
rect 234494 216988 234522 217246
rect 235368 217138 235396 218010
rect 236196 217138 236224 218010
rect 237024 217274 237052 220186
rect 237300 218074 237328 225694
rect 237760 224670 237788 231676
rect 238404 228002 238432 231676
rect 238576 228812 238628 228818
rect 238576 228754 238628 228760
rect 238392 227996 238444 228002
rect 238392 227938 238444 227944
rect 237748 224664 237800 224670
rect 237748 224606 237800 224612
rect 238024 223712 238076 223718
rect 238024 223654 238076 223660
rect 237840 219428 237892 219434
rect 237840 219370 237892 219376
rect 237288 218068 237340 218074
rect 237288 218010 237340 218016
rect 235322 217110 235396 217138
rect 236150 217110 236224 217138
rect 236978 217246 237052 217274
rect 235322 216988 235350 217110
rect 236150 216988 236178 217110
rect 236978 216988 237006 217246
rect 237852 217138 237880 219370
rect 238036 218482 238064 223654
rect 238024 218476 238076 218482
rect 238024 218418 238076 218424
rect 238588 217274 238616 228754
rect 239048 228138 239076 231676
rect 239036 228132 239088 228138
rect 239036 228074 239088 228080
rect 239692 223446 239720 231676
rect 240152 231662 240350 231690
rect 239680 223440 239732 223446
rect 239680 223382 239732 223388
rect 240152 221882 240180 231662
rect 240324 230172 240376 230178
rect 240324 230114 240376 230120
rect 240336 225758 240364 230114
rect 240980 229226 241008 231676
rect 240968 229220 241020 229226
rect 240968 229162 241020 229168
rect 241624 227322 241652 231676
rect 241612 227316 241664 227322
rect 241612 227258 241664 227264
rect 240324 225752 240376 225758
rect 240324 225694 240376 225700
rect 241152 225344 241204 225350
rect 241152 225286 241204 225292
rect 240140 221876 240192 221882
rect 240140 221818 240192 221824
rect 239312 221740 239364 221746
rect 239312 221682 239364 221688
rect 239324 219434 239352 221682
rect 239312 219428 239364 219434
rect 239312 219370 239364 219376
rect 239496 219428 239548 219434
rect 239496 219370 239548 219376
rect 238588 217246 238662 217274
rect 237806 217110 237880 217138
rect 237806 216988 237834 217110
rect 238634 216988 238662 217246
rect 239508 217138 239536 219370
rect 240324 218068 240376 218074
rect 240324 218010 240376 218016
rect 240336 217138 240364 218010
rect 241164 217274 241192 225286
rect 242268 223582 242296 231676
rect 242716 225208 242768 225214
rect 242716 225150 242768 225156
rect 242256 223576 242308 223582
rect 242256 223518 242308 223524
rect 241336 223168 241388 223174
rect 241336 223110 241388 223116
rect 241348 218074 241376 223110
rect 242728 220946 242756 225150
rect 242912 224942 242940 231676
rect 243280 231662 243570 231690
rect 243280 226642 243308 231662
rect 243452 226704 243504 226710
rect 243452 226646 243504 226652
rect 243268 226636 243320 226642
rect 243268 226578 243320 226584
rect 242900 224936 242952 224942
rect 242900 224878 242952 224884
rect 242728 220918 242848 220946
rect 242624 220788 242676 220794
rect 242624 220730 242676 220736
rect 242636 219434 242664 220730
rect 242820 219434 242848 220918
rect 241796 219428 241848 219434
rect 241796 219370 241848 219376
rect 241980 219428 242032 219434
rect 242636 219406 242756 219434
rect 242820 219428 242952 219434
rect 242820 219406 242900 219428
rect 241980 219370 242032 219376
rect 241808 219026 241836 219370
rect 241612 219020 241664 219026
rect 241612 218962 241664 218968
rect 241796 219020 241848 219026
rect 241796 218962 241848 218968
rect 241624 218346 241652 218962
rect 241612 218340 241664 218346
rect 241612 218282 241664 218288
rect 241336 218068 241388 218074
rect 241336 218010 241388 218016
rect 239462 217110 239536 217138
rect 240290 217110 240364 217138
rect 241118 217246 241192 217274
rect 239462 216988 239490 217110
rect 240290 216988 240318 217110
rect 241118 216988 241146 217246
rect 241992 217138 242020 219370
rect 242728 217274 242756 219406
rect 242900 219370 242952 219376
rect 243464 218754 243492 226646
rect 244200 225486 244228 231676
rect 244476 231662 244858 231690
rect 245120 231662 245502 231690
rect 244476 229094 244504 231662
rect 244384 229066 244504 229094
rect 244188 225480 244240 225486
rect 244188 225422 244240 225428
rect 244096 223440 244148 223446
rect 244096 223382 244148 223388
rect 243452 218748 243504 218754
rect 243452 218690 243504 218696
rect 244108 218074 244136 223382
rect 244384 220266 244412 229066
rect 245120 222358 245148 231662
rect 246132 229770 246160 231676
rect 246120 229764 246172 229770
rect 246120 229706 246172 229712
rect 246488 229764 246540 229770
rect 246488 229706 246540 229712
rect 246304 228132 246356 228138
rect 246304 228074 246356 228080
rect 245292 224800 245344 224806
rect 245292 224742 245344 224748
rect 245108 222352 245160 222358
rect 245108 222294 245160 222300
rect 244292 220238 244412 220266
rect 244292 220114 244320 220238
rect 244280 220108 244332 220114
rect 244280 220050 244332 220056
rect 244464 220108 244516 220114
rect 244464 220050 244516 220056
rect 243636 218068 243688 218074
rect 243636 218010 243688 218016
rect 244096 218068 244148 218074
rect 244096 218010 244148 218016
rect 242728 217246 242802 217274
rect 241946 217110 242020 217138
rect 241946 216988 241974 217110
rect 242774 216988 242802 217246
rect 243648 217138 243676 218010
rect 244476 217274 244504 220050
rect 244924 219428 244976 219434
rect 244924 219370 244976 219376
rect 244936 219026 244964 219370
rect 244924 219020 244976 219026
rect 244924 218962 244976 218968
rect 245304 217274 245332 224742
rect 246316 218346 246344 228074
rect 246500 220794 246528 229706
rect 246776 228954 246804 231676
rect 246764 228948 246816 228954
rect 246764 228890 246816 228896
rect 246856 223304 246908 223310
rect 246856 223246 246908 223252
rect 246488 220788 246540 220794
rect 246488 220730 246540 220736
rect 246304 218340 246356 218346
rect 246304 218282 246356 218288
rect 246120 218204 246172 218210
rect 246120 218146 246172 218152
rect 243602 217110 243676 217138
rect 244430 217246 244504 217274
rect 245258 217246 245332 217274
rect 243602 216988 243630 217110
rect 244430 216988 244458 217246
rect 245258 216988 245286 217246
rect 246132 217138 246160 218146
rect 246868 217274 246896 223246
rect 247420 222766 247448 231676
rect 247604 231662 248078 231690
rect 247408 222760 247460 222766
rect 247408 222702 247460 222708
rect 247604 222154 247632 231662
rect 248236 228948 248288 228954
rect 248236 228890 248288 228896
rect 247592 222148 247644 222154
rect 247592 222090 247644 222096
rect 248248 218074 248276 228890
rect 248708 226710 248736 231676
rect 248696 226704 248748 226710
rect 248696 226646 248748 226652
rect 249352 225894 249380 231676
rect 249616 226772 249668 226778
rect 249616 226714 249668 226720
rect 249340 225888 249392 225894
rect 249340 225830 249392 225836
rect 249432 218340 249484 218346
rect 249432 218282 249484 218288
rect 247776 218068 247828 218074
rect 247776 218010 247828 218016
rect 248236 218068 248288 218074
rect 248236 218010 248288 218016
rect 248604 218068 248656 218074
rect 248604 218010 248656 218016
rect 246868 217246 246942 217274
rect 246086 217110 246160 217138
rect 246086 216988 246114 217110
rect 246914 216988 246942 217246
rect 247788 217138 247816 218010
rect 248616 217138 248644 218010
rect 249444 217138 249472 218282
rect 249628 218074 249656 226714
rect 249996 222630 250024 231676
rect 250640 224126 250668 231676
rect 251284 229634 251312 231676
rect 251272 229628 251324 229634
rect 251272 229570 251324 229576
rect 251732 229628 251784 229634
rect 251732 229570 251784 229576
rect 251088 224528 251140 224534
rect 251088 224470 251140 224476
rect 250628 224120 250680 224126
rect 250628 224062 250680 224068
rect 250904 223576 250956 223582
rect 250904 223518 250956 223524
rect 249984 222624 250036 222630
rect 249984 222566 250036 222572
rect 250916 218074 250944 223518
rect 249616 218068 249668 218074
rect 249616 218010 249668 218016
rect 250260 218068 250312 218074
rect 250260 218010 250312 218016
rect 250904 218068 250956 218074
rect 250904 218010 250956 218016
rect 250272 217138 250300 218010
rect 251100 217274 251128 224470
rect 251744 218346 251772 229570
rect 251928 227458 251956 231676
rect 252572 229090 252600 231676
rect 252756 231662 253230 231690
rect 252560 229084 252612 229090
rect 252560 229026 252612 229032
rect 251916 227452 251968 227458
rect 251916 227394 251968 227400
rect 252468 225888 252520 225894
rect 252468 225830 252520 225836
rect 251732 218340 251784 218346
rect 251732 218282 251784 218288
rect 252480 218074 252508 225830
rect 252756 221338 252784 231662
rect 253860 228138 253888 231676
rect 253848 228132 253900 228138
rect 253848 228074 253900 228080
rect 254504 225078 254532 231676
rect 254780 231662 255162 231690
rect 254492 225072 254544 225078
rect 254492 225014 254544 225020
rect 252744 221332 252796 221338
rect 252744 221274 252796 221280
rect 253848 220856 253900 220862
rect 253848 220798 253900 220804
rect 253572 220652 253624 220658
rect 253572 220594 253624 220600
rect 253020 219156 253072 219162
rect 253020 219098 253072 219104
rect 252744 219020 252796 219026
rect 252744 218962 252796 218968
rect 251916 218068 251968 218074
rect 251916 218010 251968 218016
rect 252468 218068 252520 218074
rect 252468 218010 252520 218016
rect 247742 217110 247816 217138
rect 248570 217110 248644 217138
rect 249398 217110 249472 217138
rect 250226 217110 250300 217138
rect 251054 217246 251128 217274
rect 247742 216988 247770 217110
rect 248570 216988 248598 217110
rect 249398 216988 249426 217110
rect 250226 216988 250254 217110
rect 251054 216988 251082 217246
rect 251928 217138 251956 218010
rect 252756 217138 252784 218962
rect 253032 218346 253060 219098
rect 253204 218748 253256 218754
rect 253204 218690 253256 218696
rect 253020 218340 253072 218346
rect 253020 218282 253072 218288
rect 253216 218210 253244 218690
rect 253204 218204 253256 218210
rect 253204 218146 253256 218152
rect 253584 217274 253612 220594
rect 253860 218890 253888 220798
rect 254780 219978 254808 231662
rect 255228 229084 255280 229090
rect 255228 229026 255280 229032
rect 255044 225752 255096 225758
rect 255044 225694 255096 225700
rect 254768 219972 254820 219978
rect 254768 219914 254820 219920
rect 253848 218884 253900 218890
rect 253848 218826 253900 218832
rect 255056 218074 255084 225694
rect 254400 218068 254452 218074
rect 254400 218010 254452 218016
rect 255044 218068 255096 218074
rect 255044 218010 255096 218016
rect 251882 217110 251956 217138
rect 252710 217110 252784 217138
rect 253538 217246 253612 217274
rect 251882 216988 251910 217110
rect 252710 216988 252738 217110
rect 253538 216988 253566 217246
rect 254412 217138 254440 218010
rect 255240 217274 255268 229026
rect 255792 223990 255820 231676
rect 256436 230314 256464 231676
rect 256424 230308 256476 230314
rect 256424 230250 256476 230256
rect 256608 230308 256660 230314
rect 256608 230250 256660 230256
rect 255780 223984 255832 223990
rect 255780 223926 255832 223932
rect 256620 219434 256648 230250
rect 257080 228274 257108 231676
rect 257448 231662 257738 231690
rect 257068 228268 257120 228274
rect 257068 228210 257120 228216
rect 257448 226302 257476 231662
rect 257620 228268 257672 228274
rect 257620 228210 257672 228216
rect 257436 226296 257488 226302
rect 257436 226238 257488 226244
rect 257632 219434 257660 228210
rect 257804 227316 257856 227322
rect 257804 227258 257856 227264
rect 257816 219434 257844 227258
rect 258368 222494 258396 231676
rect 258644 231662 259026 231690
rect 258356 222488 258408 222494
rect 258356 222430 258408 222436
rect 258080 222148 258132 222154
rect 258080 222090 258132 222096
rect 256528 219406 256648 219434
rect 257540 219406 257660 219434
rect 257724 219406 257844 219434
rect 256528 218074 256556 219406
rect 257540 218074 257568 219406
rect 256056 218068 256108 218074
rect 256056 218010 256108 218016
rect 256516 218068 256568 218074
rect 256516 218010 256568 218016
rect 256884 218068 256936 218074
rect 256884 218010 256936 218016
rect 257528 218068 257580 218074
rect 257528 218010 257580 218016
rect 254366 217110 254440 217138
rect 255194 217246 255268 217274
rect 254366 216988 254394 217110
rect 255194 216988 255222 217246
rect 256068 217138 256096 218010
rect 256896 217138 256924 218010
rect 257724 217274 257752 219406
rect 258092 218346 258120 222090
rect 258644 220862 258672 231662
rect 259276 227452 259328 227458
rect 259276 227394 259328 227400
rect 258632 220856 258684 220862
rect 258632 220798 258684 220804
rect 259092 218884 259144 218890
rect 259092 218826 259144 218832
rect 258080 218340 258132 218346
rect 258080 218282 258132 218288
rect 258540 218068 258592 218074
rect 258540 218010 258592 218016
rect 256022 217110 256096 217138
rect 256850 217110 256924 217138
rect 257678 217246 257752 217274
rect 256022 216988 256050 217110
rect 256850 216988 256878 217110
rect 257678 216988 257706 217246
rect 258552 217138 258580 218010
rect 259104 217274 259132 218826
rect 259288 218074 259316 227394
rect 259656 226166 259684 231676
rect 259932 231662 260314 231690
rect 260852 231662 260958 231690
rect 259644 226160 259696 226166
rect 259644 226102 259696 226108
rect 259932 219842 259960 231662
rect 260852 221610 260880 231662
rect 261588 230450 261616 231676
rect 261576 230444 261628 230450
rect 261576 230386 261628 230392
rect 262232 227594 262260 231676
rect 262876 227730 262904 231676
rect 263060 231662 263534 231690
rect 263704 231662 264178 231690
rect 262864 227724 262916 227730
rect 262864 227666 262916 227672
rect 262220 227588 262272 227594
rect 262220 227530 262272 227536
rect 261852 226160 261904 226166
rect 261852 226102 261904 226108
rect 260840 221604 260892 221610
rect 260840 221546 260892 221552
rect 261024 221604 261076 221610
rect 261024 221546 261076 221552
rect 260196 220788 260248 220794
rect 260196 220730 260248 220736
rect 259920 219836 259972 219842
rect 259920 219778 259972 219784
rect 259276 218068 259328 218074
rect 259276 218010 259328 218016
rect 260208 217274 260236 220730
rect 261036 217274 261064 221546
rect 261864 217274 261892 226102
rect 263060 221066 263088 231662
rect 263508 227724 263560 227730
rect 263508 227666 263560 227672
rect 263324 221876 263376 221882
rect 263324 221818 263376 221824
rect 263048 221060 263100 221066
rect 263048 221002 263100 221008
rect 263336 219434 263364 221818
rect 263336 219406 263456 219434
rect 262680 218068 262732 218074
rect 262680 218010 262732 218016
rect 259104 217246 259362 217274
rect 258506 217110 258580 217138
rect 258506 216988 258534 217110
rect 259334 216988 259362 217246
rect 260162 217246 260236 217274
rect 260990 217246 261064 217274
rect 261818 217246 261892 217274
rect 260162 216988 260190 217246
rect 260990 216988 261018 217246
rect 261818 216988 261846 217246
rect 262692 217138 262720 218010
rect 263428 217274 263456 219406
rect 263520 218090 263548 227666
rect 263704 222154 263732 231662
rect 264808 228546 264836 231676
rect 265176 231662 265466 231690
rect 264796 228540 264848 228546
rect 264796 228482 264848 228488
rect 264152 226636 264204 226642
rect 264152 226578 264204 226584
rect 263692 222148 263744 222154
rect 263692 222090 263744 222096
rect 264164 219298 264192 226578
rect 264796 222760 264848 222766
rect 264796 222702 264848 222708
rect 264152 219292 264204 219298
rect 264152 219234 264204 219240
rect 263520 218074 263640 218090
rect 264808 218074 264836 222702
rect 265176 220386 265204 231662
rect 266096 225622 266124 231676
rect 266084 225616 266136 225622
rect 266084 225558 266136 225564
rect 266176 224936 266228 224942
rect 266176 224878 266228 224884
rect 265164 220380 265216 220386
rect 265164 220322 265216 220328
rect 265992 219156 266044 219162
rect 265992 219098 266044 219104
rect 263520 218068 263652 218074
rect 263520 218062 263600 218068
rect 263600 218010 263652 218016
rect 264336 218068 264388 218074
rect 264336 218010 264388 218016
rect 264796 218068 264848 218074
rect 264796 218010 264848 218016
rect 265164 218068 265216 218074
rect 265164 218010 265216 218016
rect 263428 217246 263502 217274
rect 262646 217110 262720 217138
rect 262646 216988 262674 217110
rect 263474 216988 263502 217246
rect 264348 217138 264376 218010
rect 265176 217138 265204 218010
rect 266004 217138 266032 219098
rect 266188 218074 266216 224878
rect 266740 223718 266768 231676
rect 267384 226914 267412 231676
rect 267936 231662 268042 231690
rect 268304 231662 268686 231690
rect 267372 226908 267424 226914
rect 267372 226850 267424 226856
rect 267004 226296 267056 226302
rect 267004 226238 267056 226244
rect 266728 223712 266780 223718
rect 266728 223654 266780 223660
rect 266820 221332 266872 221338
rect 266820 221274 266872 221280
rect 266176 218068 266228 218074
rect 266176 218010 266228 218016
rect 266832 217274 266860 221274
rect 267016 218618 267044 226238
rect 267936 220522 267964 231662
rect 268304 221202 268332 231662
rect 268936 228132 268988 228138
rect 268936 228074 268988 228080
rect 268292 221196 268344 221202
rect 268292 221138 268344 221144
rect 267924 220516 267976 220522
rect 267924 220458 267976 220464
rect 267648 220380 267700 220386
rect 267648 220322 267700 220328
rect 267004 218612 267056 218618
rect 267004 218554 267056 218560
rect 267660 217274 267688 220322
rect 268948 218074 268976 228074
rect 269316 226642 269344 231676
rect 269304 226636 269356 226642
rect 269304 226578 269356 226584
rect 269960 226030 269988 231676
rect 269948 226024 270000 226030
rect 269948 225966 270000 225972
rect 270040 225616 270092 225622
rect 270040 225558 270092 225564
rect 270052 218074 270080 225558
rect 270604 224670 270632 231676
rect 271248 227050 271276 231676
rect 271892 229906 271920 231676
rect 271880 229900 271932 229906
rect 271880 229842 271932 229848
rect 272536 228682 272564 231676
rect 272720 231662 273194 231690
rect 272524 228676 272576 228682
rect 272524 228618 272576 228624
rect 272524 228540 272576 228546
rect 272524 228482 272576 228488
rect 271236 227044 271288 227050
rect 271236 226986 271288 226992
rect 271788 227044 271840 227050
rect 271788 226986 271840 226992
rect 271144 226432 271196 226438
rect 271144 226374 271196 226380
rect 270592 224664 270644 224670
rect 270592 224606 270644 224612
rect 270224 222148 270276 222154
rect 270224 222090 270276 222096
rect 268476 218068 268528 218074
rect 268476 218010 268528 218016
rect 268936 218068 268988 218074
rect 268936 218010 268988 218016
rect 269304 218068 269356 218074
rect 269304 218010 269356 218016
rect 270040 218068 270092 218074
rect 270040 218010 270092 218016
rect 264302 217110 264376 217138
rect 265130 217110 265204 217138
rect 265958 217110 266032 217138
rect 266786 217246 266860 217274
rect 267614 217246 267688 217274
rect 264302 216988 264330 217110
rect 265130 216988 265158 217110
rect 265958 216988 265986 217110
rect 266786 216988 266814 217246
rect 267614 216988 267642 217246
rect 268488 217138 268516 218010
rect 269316 217138 269344 218010
rect 270236 217274 270264 222090
rect 271156 218482 271184 226374
rect 271144 218476 271196 218482
rect 271144 218418 271196 218424
rect 270960 218068 271012 218074
rect 270960 218010 271012 218016
rect 268442 217110 268516 217138
rect 269270 217110 269344 217138
rect 270098 217246 270264 217274
rect 268442 216988 268470 217110
rect 269270 216988 269298 217110
rect 270098 216988 270126 217246
rect 270972 217138 271000 218010
rect 271800 217274 271828 226986
rect 272340 219428 272392 219434
rect 272340 219370 272392 219376
rect 272352 218618 272380 219370
rect 272340 218612 272392 218618
rect 272340 218554 272392 218560
rect 272536 218074 272564 228482
rect 272720 219706 272748 231662
rect 273824 228410 273852 231676
rect 273812 228404 273864 228410
rect 273812 228346 273864 228352
rect 274468 226302 274496 231676
rect 275112 229094 275140 231676
rect 274928 229066 275140 229094
rect 275480 231662 275770 231690
rect 276124 231662 276414 231690
rect 274456 226296 274508 226302
rect 274456 226238 274508 226244
rect 274272 224664 274324 224670
rect 274272 224606 274324 224612
rect 273444 220516 273496 220522
rect 273444 220458 273496 220464
rect 272708 219700 272760 219706
rect 272708 219642 272760 219648
rect 272708 219428 272760 219434
rect 272708 219370 272760 219376
rect 272524 218068 272576 218074
rect 272524 218010 272576 218016
rect 272720 217274 272748 219370
rect 273456 217274 273484 220458
rect 274284 217274 274312 224606
rect 274928 224398 274956 229066
rect 274916 224392 274968 224398
rect 274916 224334 274968 224340
rect 275100 224392 275152 224398
rect 275100 224334 275152 224340
rect 275112 217274 275140 224334
rect 275480 223038 275508 231662
rect 275652 229900 275704 229906
rect 275652 229842 275704 229848
rect 275664 229094 275692 229842
rect 275664 229066 275876 229094
rect 275468 223032 275520 223038
rect 275468 222974 275520 222980
rect 270926 217110 271000 217138
rect 271754 217246 271828 217274
rect 272582 217246 272748 217274
rect 273410 217246 273484 217274
rect 274238 217246 274312 217274
rect 275066 217246 275140 217274
rect 275848 217274 275876 229066
rect 276124 221474 276152 231662
rect 277044 230042 277072 231676
rect 277032 230036 277084 230042
rect 277032 229978 277084 229984
rect 277216 230036 277268 230042
rect 277216 229978 277268 229984
rect 277228 227730 277256 229978
rect 277216 227724 277268 227730
rect 277216 227666 277268 227672
rect 277216 227588 277268 227594
rect 277216 227530 277268 227536
rect 276112 221468 276164 221474
rect 276112 221410 276164 221416
rect 277228 218074 277256 227530
rect 277688 223854 277716 231676
rect 277964 231662 278346 231690
rect 277676 223848 277728 223854
rect 277676 223790 277728 223796
rect 277964 222018 277992 231662
rect 278412 226024 278464 226030
rect 278412 225966 278464 225972
rect 277952 222012 278004 222018
rect 277952 221954 278004 221960
rect 276756 218068 276808 218074
rect 276756 218010 276808 218016
rect 277216 218068 277268 218074
rect 277216 218010 277268 218016
rect 277584 218068 277636 218074
rect 277584 218010 277636 218016
rect 275848 217246 275922 217274
rect 270926 216988 270954 217110
rect 271754 216988 271782 217246
rect 272582 216988 272610 217246
rect 273410 216988 273438 217246
rect 274238 216988 274266 217246
rect 275066 216988 275094 217246
rect 275894 216988 275922 217246
rect 276768 217138 276796 218010
rect 277596 217138 277624 218010
rect 278424 217274 278452 225966
rect 278976 224262 279004 231676
rect 279620 226438 279648 231676
rect 280264 227186 280292 231676
rect 280448 231662 280922 231690
rect 280252 227180 280304 227186
rect 280252 227122 280304 227128
rect 279608 226432 279660 226438
rect 279608 226374 279660 226380
rect 278964 224256 279016 224262
rect 278964 224198 279016 224204
rect 279424 223984 279476 223990
rect 279424 223926 279476 223932
rect 278596 223032 278648 223038
rect 278596 222974 278648 222980
rect 278608 218074 278636 222974
rect 279436 218618 279464 223926
rect 280068 222012 280120 222018
rect 280068 221954 280120 221960
rect 279424 218612 279476 218618
rect 279424 218554 279476 218560
rect 279240 218476 279292 218482
rect 279240 218418 279292 218424
rect 278596 218068 278648 218074
rect 278596 218010 278648 218016
rect 276722 217110 276796 217138
rect 277550 217110 277624 217138
rect 278378 217246 278452 217274
rect 276722 216988 276750 217110
rect 277550 216988 277578 217110
rect 278378 216988 278406 217246
rect 279252 217138 279280 218418
rect 280080 217274 280108 221954
rect 280448 220250 280476 231662
rect 281356 226908 281408 226914
rect 281356 226850 281408 226856
rect 280436 220244 280488 220250
rect 280436 220186 280488 220192
rect 281368 219434 281396 226850
rect 281552 222902 281580 231676
rect 282196 230178 282224 231676
rect 282184 230172 282236 230178
rect 282184 230114 282236 230120
rect 282644 230172 282696 230178
rect 282644 230114 282696 230120
rect 282184 227588 282236 227594
rect 282184 227530 282236 227536
rect 282196 227050 282224 227530
rect 282184 227044 282236 227050
rect 282184 226986 282236 226992
rect 282656 225622 282684 230114
rect 282840 228818 282868 231676
rect 282828 228812 282880 228818
rect 282828 228754 282880 228760
rect 282644 225616 282696 225622
rect 282644 225558 282696 225564
rect 283484 223174 283512 231676
rect 283668 231662 284142 231690
rect 283472 223168 283524 223174
rect 283472 223110 283524 223116
rect 281540 222896 281592 222902
rect 281540 222838 281592 222844
rect 282460 222896 282512 222902
rect 282460 222838 282512 222844
rect 281368 219406 281488 219434
rect 281460 218074 281488 219406
rect 282472 218074 282500 222838
rect 283668 221746 283696 231662
rect 284116 225616 284168 225622
rect 284116 225558 284168 225564
rect 283656 221740 283708 221746
rect 283656 221682 283708 221688
rect 282644 220924 282696 220930
rect 282644 220866 282696 220872
rect 280896 218068 280948 218074
rect 280896 218010 280948 218016
rect 281448 218068 281500 218074
rect 281448 218010 281500 218016
rect 281724 218068 281776 218074
rect 281724 218010 281776 218016
rect 282460 218068 282512 218074
rect 282460 218010 282512 218016
rect 279206 217110 279280 217138
rect 280034 217246 280108 217274
rect 279206 216988 279234 217110
rect 280034 216988 280062 217246
rect 280908 217138 280936 218010
rect 281736 217138 281764 218010
rect 282656 217274 282684 220866
rect 283380 220244 283432 220250
rect 283380 220186 283432 220192
rect 283392 217274 283420 220186
rect 280862 217110 280936 217138
rect 281690 217110 281764 217138
rect 282518 217246 282684 217274
rect 283346 217246 283420 217274
rect 284128 217274 284156 225558
rect 284772 223990 284800 231676
rect 285048 231662 285430 231690
rect 285048 225214 285076 231662
rect 285496 228404 285548 228410
rect 285496 228346 285548 228352
rect 285036 225208 285088 225214
rect 285036 225150 285088 225156
rect 284760 223984 284812 223990
rect 284760 223926 284812 223932
rect 285508 218074 285536 228346
rect 286060 223446 286088 231676
rect 286324 226296 286376 226302
rect 286324 226238 286376 226244
rect 286048 223440 286100 223446
rect 286048 223382 286100 223388
rect 285864 219428 285916 219434
rect 285864 219370 285916 219376
rect 285036 218068 285088 218074
rect 285036 218010 285088 218016
rect 285496 218068 285548 218074
rect 285496 218010 285548 218016
rect 284128 217246 284202 217274
rect 280862 216988 280890 217110
rect 281690 216988 281718 217110
rect 282518 216988 282546 217246
rect 283346 216988 283374 217246
rect 284174 216988 284202 217246
rect 285048 217138 285076 218010
rect 285876 217138 285904 219370
rect 286336 218754 286364 226238
rect 286704 225350 286732 231676
rect 287348 229770 287376 231676
rect 287336 229764 287388 229770
rect 287336 229706 287388 229712
rect 287704 229764 287756 229770
rect 287704 229706 287756 229712
rect 286692 225344 286744 225350
rect 286692 225286 286744 225292
rect 286692 224120 286744 224126
rect 286692 224062 286744 224068
rect 286324 218748 286376 218754
rect 286324 218690 286376 218696
rect 286704 217274 286732 224062
rect 287716 220930 287744 229706
rect 287992 224806 288020 231676
rect 287980 224800 288032 224806
rect 287980 224742 288032 224748
rect 288636 223310 288664 231676
rect 288820 231662 289294 231690
rect 288624 223304 288676 223310
rect 288624 223246 288676 223252
rect 288256 223168 288308 223174
rect 288256 223110 288308 223116
rect 287888 222352 287940 222358
rect 287888 222294 287940 222300
rect 287704 220924 287756 220930
rect 287704 220866 287756 220872
rect 287900 219026 287928 222294
rect 287888 219020 287940 219026
rect 287888 218962 287940 218968
rect 287520 218068 287572 218074
rect 287520 218010 287572 218016
rect 285002 217110 285076 217138
rect 285830 217110 285904 217138
rect 286658 217246 286732 217274
rect 285002 216988 285030 217110
rect 285830 216988 285858 217110
rect 286658 216988 286686 217246
rect 287532 217138 287560 218010
rect 288268 217274 288296 223110
rect 288820 222194 288848 231662
rect 289924 226302 289952 231676
rect 290568 226778 290596 231676
rect 290556 226772 290608 226778
rect 290556 226714 290608 226720
rect 289912 226296 289964 226302
rect 289912 226238 289964 226244
rect 291016 226296 291068 226302
rect 291016 226238 291068 226244
rect 290832 224256 290884 224262
rect 290832 224198 290884 224204
rect 289728 223304 289780 223310
rect 289728 223246 289780 223252
rect 288544 222166 288848 222194
rect 288544 220114 288572 222166
rect 288532 220108 288584 220114
rect 288532 220050 288584 220056
rect 288716 220108 288768 220114
rect 288716 220050 288768 220056
rect 288728 218074 288756 220050
rect 289740 218074 289768 223246
rect 288716 218068 288768 218074
rect 288716 218010 288768 218016
rect 289176 218068 289228 218074
rect 289176 218010 289228 218016
rect 289728 218068 289780 218074
rect 289728 218010 289780 218016
rect 290004 218068 290056 218074
rect 290004 218010 290056 218016
rect 288268 217246 288342 217274
rect 287486 217110 287560 217138
rect 287486 216988 287514 217110
rect 288314 216988 288342 217246
rect 289188 217138 289216 218010
rect 290016 217138 290044 218010
rect 290844 217274 290872 224198
rect 291028 219434 291056 226238
rect 291212 223582 291240 231676
rect 291856 228954 291884 231676
rect 292500 229634 292528 231676
rect 292488 229628 292540 229634
rect 292488 229570 292540 229576
rect 291844 228948 291896 228954
rect 291844 228890 291896 228896
rect 291844 228812 291896 228818
rect 291844 228754 291896 228760
rect 291200 223576 291252 223582
rect 291200 223518 291252 223524
rect 291028 219406 291148 219434
rect 291120 218074 291148 219406
rect 291660 218884 291712 218890
rect 291660 218826 291712 218832
rect 291108 218068 291160 218074
rect 291108 218010 291160 218016
rect 289142 217110 289216 217138
rect 289970 217110 290044 217138
rect 290798 217246 290872 217274
rect 289142 216988 289170 217110
rect 289970 216988 289998 217110
rect 290798 216988 290826 217246
rect 291672 217138 291700 218826
rect 291856 218754 291884 228754
rect 293144 225894 293172 231676
rect 293328 231662 293802 231690
rect 293132 225888 293184 225894
rect 293132 225830 293184 225836
rect 292488 221468 292540 221474
rect 292488 221410 292540 221416
rect 291844 218748 291896 218754
rect 291844 218690 291896 218696
rect 292500 217274 292528 221410
rect 293328 220658 293356 231662
rect 293776 226908 293828 226914
rect 293776 226850 293828 226856
rect 293316 220652 293368 220658
rect 293316 220594 293368 220600
rect 293788 218074 293816 226850
rect 294432 224534 294460 231676
rect 294420 224528 294472 224534
rect 294420 224470 294472 224476
rect 295076 222358 295104 231676
rect 295720 229090 295748 231676
rect 295708 229084 295760 229090
rect 295708 229026 295760 229032
rect 296364 228274 296392 231676
rect 296628 228676 296680 228682
rect 296628 228618 296680 228624
rect 296352 228268 296404 228274
rect 296352 228210 296404 228216
rect 296444 225888 296496 225894
rect 296444 225830 296496 225836
rect 295064 222352 295116 222358
rect 295064 222294 295116 222300
rect 294972 219972 295024 219978
rect 294972 219914 295024 219920
rect 294144 218476 294196 218482
rect 294144 218418 294196 218424
rect 293316 218068 293368 218074
rect 293316 218010 293368 218016
rect 293776 218068 293828 218074
rect 293776 218010 293828 218016
rect 291626 217110 291700 217138
rect 292454 217246 292528 217274
rect 291626 216988 291654 217110
rect 292454 216988 292482 217246
rect 293328 217138 293356 218010
rect 294156 217138 294184 218418
rect 294984 217274 295012 219914
rect 296456 219434 296484 225830
rect 296456 219406 296576 219434
rect 295800 219156 295852 219162
rect 295800 219098 295852 219104
rect 293282 217110 293356 217138
rect 294110 217110 294184 217138
rect 294938 217246 295012 217274
rect 293282 216988 293310 217110
rect 294110 216988 294138 217110
rect 294938 216988 294966 217246
rect 295812 217138 295840 219098
rect 296548 217274 296576 219406
rect 296640 219178 296668 228618
rect 297008 225758 297036 231676
rect 297652 230314 297680 231676
rect 297640 230308 297692 230314
rect 297640 230250 297692 230256
rect 297824 230308 297876 230314
rect 297824 230250 297876 230256
rect 297836 229094 297864 230250
rect 297744 229066 297864 229094
rect 296996 225752 297048 225758
rect 296996 225694 297048 225700
rect 297272 225004 297324 225010
rect 297272 224946 297324 224952
rect 296640 219162 296760 219178
rect 296640 219156 296772 219162
rect 296640 219150 296720 219156
rect 296720 219098 296772 219104
rect 297284 219026 297312 224946
rect 297744 223310 297772 229066
rect 298296 227458 298324 231676
rect 298572 231662 298954 231690
rect 298284 227452 298336 227458
rect 298284 227394 298336 227400
rect 297916 223576 297968 223582
rect 297916 223518 297968 223524
rect 297732 223304 297784 223310
rect 297732 223246 297784 223252
rect 297272 219020 297324 219026
rect 297272 218962 297324 218968
rect 297928 218074 297956 223518
rect 298572 220794 298600 231662
rect 299584 227322 299612 231676
rect 300228 228818 300256 231676
rect 300216 228812 300268 228818
rect 300216 228754 300268 228760
rect 300676 228812 300728 228818
rect 300676 228754 300728 228760
rect 299572 227316 299624 227322
rect 299572 227258 299624 227264
rect 299296 224528 299348 224534
rect 299296 224470 299348 224476
rect 299112 223304 299164 223310
rect 299112 223246 299164 223252
rect 298560 220788 298612 220794
rect 298560 220730 298612 220736
rect 299124 218074 299152 223246
rect 297456 218068 297508 218074
rect 297456 218010 297508 218016
rect 297916 218068 297968 218074
rect 297916 218010 297968 218016
rect 298284 218068 298336 218074
rect 298284 218010 298336 218016
rect 299112 218068 299164 218074
rect 299112 218010 299164 218016
rect 296548 217246 296622 217274
rect 295766 217110 295840 217138
rect 295766 216988 295794 217110
rect 296594 216988 296622 217246
rect 297468 217138 297496 218010
rect 298296 217138 298324 218010
rect 299308 217274 299336 224470
rect 300492 218884 300544 218890
rect 300492 218826 300544 218832
rect 299940 218068 299992 218074
rect 299940 218010 299992 218016
rect 297422 217110 297496 217138
rect 298250 217110 298324 217138
rect 299078 217246 299336 217274
rect 297422 216988 297450 217110
rect 298250 216988 298278 217110
rect 299078 216988 299106 217246
rect 299952 217138 299980 218010
rect 300504 217274 300532 218826
rect 300688 218074 300716 228754
rect 300872 226166 300900 231676
rect 301148 231662 301530 231690
rect 301792 231662 302174 231690
rect 300860 226160 300912 226166
rect 300860 226102 300912 226108
rect 301148 221882 301176 231662
rect 301136 221876 301188 221882
rect 301136 221818 301188 221824
rect 301792 221610 301820 231662
rect 302804 230042 302832 231676
rect 302792 230036 302844 230042
rect 302792 229978 302844 229984
rect 303252 230036 303304 230042
rect 303252 229978 303304 229984
rect 302148 228948 302200 228954
rect 302148 228890 302200 228896
rect 301964 221876 302016 221882
rect 301964 221818 302016 221824
rect 301780 221604 301832 221610
rect 301780 221546 301832 221552
rect 301976 219298 302004 221818
rect 301964 219292 302016 219298
rect 301964 219234 302016 219240
rect 302160 218074 302188 228890
rect 303264 223582 303292 229978
rect 303448 224874 303476 231676
rect 303816 231662 304106 231690
rect 304368 231662 304750 231690
rect 303436 224868 303488 224874
rect 303436 224810 303488 224816
rect 303252 223576 303304 223582
rect 303252 223518 303304 223524
rect 303252 221740 303304 221746
rect 303252 221682 303304 221688
rect 302424 220652 302476 220658
rect 302424 220594 302476 220600
rect 300676 218068 300728 218074
rect 300676 218010 300728 218016
rect 301596 218068 301648 218074
rect 301596 218010 301648 218016
rect 302148 218068 302200 218074
rect 302148 218010 302200 218016
rect 300504 217246 300762 217274
rect 299906 217110 299980 217138
rect 299906 216988 299934 217110
rect 300734 216988 300762 217246
rect 301608 217138 301636 218010
rect 302436 217274 302464 220594
rect 303264 217274 303292 221682
rect 303816 221338 303844 231662
rect 304368 222766 304396 231662
rect 304908 227452 304960 227458
rect 304908 227394 304960 227400
rect 304356 222760 304408 222766
rect 304356 222702 304408 222708
rect 304724 222692 304776 222698
rect 304724 222634 304776 222640
rect 303804 221332 303856 221338
rect 303804 221274 303856 221280
rect 304736 218074 304764 222634
rect 304080 218068 304132 218074
rect 304080 218010 304132 218016
rect 304724 218068 304776 218074
rect 304724 218010 304776 218016
rect 301562 217110 301636 217138
rect 302390 217246 302464 217274
rect 303218 217246 303292 217274
rect 301562 216988 301590 217110
rect 302390 216988 302418 217246
rect 303218 216988 303246 217246
rect 304092 217138 304120 218010
rect 304920 217274 304948 227394
rect 305380 225010 305408 231676
rect 305552 229084 305604 229090
rect 305552 229026 305604 229032
rect 305368 225004 305420 225010
rect 305368 224946 305420 224952
rect 305564 218618 305592 229026
rect 306024 228138 306052 231676
rect 306576 231662 306682 231690
rect 306944 231662 307326 231690
rect 306012 228132 306064 228138
rect 306012 228074 306064 228080
rect 306196 227180 306248 227186
rect 306196 227122 306248 227128
rect 305552 218612 305604 218618
rect 305552 218554 305604 218560
rect 306208 218074 306236 227122
rect 306576 222154 306604 231662
rect 306564 222148 306616 222154
rect 306564 222090 306616 222096
rect 306944 220386 306972 231662
rect 307956 230178 307984 231676
rect 307944 230172 307996 230178
rect 307944 230114 307996 230120
rect 308128 230172 308180 230178
rect 308128 230114 308180 230120
rect 307668 223576 307720 223582
rect 307668 223518 307720 223524
rect 306932 220380 306984 220386
rect 306932 220322 306984 220328
rect 307392 219020 307444 219026
rect 307392 218962 307444 218968
rect 305736 218068 305788 218074
rect 305736 218010 305788 218016
rect 306196 218068 306248 218074
rect 306196 218010 306248 218016
rect 306564 218068 306616 218074
rect 306564 218010 306616 218016
rect 304046 217110 304120 217138
rect 304874 217246 304948 217274
rect 304046 216988 304074 217110
rect 304874 216988 304902 217246
rect 305748 217138 305776 218010
rect 306576 217138 306604 218010
rect 307404 217274 307432 218962
rect 307680 218074 307708 223518
rect 308140 222698 308168 230114
rect 308600 227594 308628 231676
rect 308588 227588 308640 227594
rect 308588 227530 308640 227536
rect 309048 226160 309100 226166
rect 309048 226102 309100 226108
rect 308128 222692 308180 222698
rect 308128 222634 308180 222640
rect 308864 221604 308916 221610
rect 308864 221546 308916 221552
rect 308876 219434 308904 221546
rect 309060 219434 309088 226102
rect 309244 220522 309272 231676
rect 309888 228546 309916 231676
rect 310546 231662 310744 231690
rect 310716 229094 310744 231662
rect 310716 229066 310928 229094
rect 309876 228540 309928 228546
rect 309876 228482 309928 228488
rect 310428 227316 310480 227322
rect 310428 227258 310480 227264
rect 309232 220516 309284 220522
rect 309232 220458 309284 220464
rect 308220 219428 308272 219434
rect 308876 219406 308996 219434
rect 309060 219428 309192 219434
rect 309060 219406 309140 219428
rect 308220 219370 308272 219376
rect 307668 218068 307720 218074
rect 307668 218010 307720 218016
rect 305702 217110 305776 217138
rect 306530 217110 306604 217138
rect 307358 217246 307432 217274
rect 305702 216988 305730 217110
rect 306530 216988 306558 217110
rect 307358 216988 307386 217246
rect 308232 217138 308260 219370
rect 308968 217274 308996 219406
rect 309140 219370 309192 219376
rect 310440 218074 310468 227258
rect 310704 222148 310756 222154
rect 310704 222090 310756 222096
rect 309876 218068 309928 218074
rect 309876 218010 309928 218016
rect 310428 218068 310480 218074
rect 310428 218010 310480 218016
rect 308968 217246 309042 217274
rect 308186 217110 308260 217138
rect 308186 216988 308214 217110
rect 309014 216988 309042 217246
rect 309888 217138 309916 218010
rect 310716 217274 310744 222090
rect 310900 221882 310928 229066
rect 311176 224398 311204 231676
rect 311820 227730 311848 231676
rect 311992 230444 312044 230450
rect 311992 230386 312044 230392
rect 312004 229906 312032 230386
rect 311992 229900 312044 229906
rect 311992 229842 312044 229848
rect 311808 227724 311860 227730
rect 311808 227666 311860 227672
rect 311532 224800 311584 224806
rect 311532 224742 311584 224748
rect 311164 224392 311216 224398
rect 311164 224334 311216 224340
rect 310888 221876 310940 221882
rect 310888 221818 310940 221824
rect 311544 217274 311572 224742
rect 312464 224670 312492 231676
rect 313108 230450 313136 231676
rect 313292 231662 313766 231690
rect 313936 231662 314410 231690
rect 313096 230444 313148 230450
rect 313096 230386 313148 230392
rect 312636 229900 312688 229906
rect 312636 229842 312688 229848
rect 312452 224664 312504 224670
rect 312452 224606 312504 224612
rect 312648 222154 312676 229842
rect 313292 226030 313320 231662
rect 313936 229094 313964 231662
rect 313752 229066 313964 229094
rect 313280 226024 313332 226030
rect 313280 225966 313332 225972
rect 312912 223440 312964 223446
rect 312912 223382 312964 223388
rect 312636 222148 312688 222154
rect 312636 222090 312688 222096
rect 312924 218074 312952 223382
rect 313752 222018 313780 229066
rect 313924 228540 313976 228546
rect 313924 228482 313976 228488
rect 313740 222012 313792 222018
rect 313740 221954 313792 221960
rect 313188 221876 313240 221882
rect 313188 221818 313240 221824
rect 312360 218068 312412 218074
rect 312360 218010 312412 218016
rect 312912 218068 312964 218074
rect 312912 218010 312964 218016
rect 309842 217110 309916 217138
rect 310670 217246 310744 217274
rect 311498 217246 311572 217274
rect 309842 216988 309870 217110
rect 310670 216988 310698 217246
rect 311498 216988 311526 217246
rect 312372 217138 312400 218010
rect 313200 217274 313228 221818
rect 313936 219298 313964 228482
rect 315040 223038 315068 231676
rect 315684 229090 315712 231676
rect 315672 229084 315724 229090
rect 315672 229026 315724 229032
rect 315672 225752 315724 225758
rect 315672 225694 315724 225700
rect 315028 223032 315080 223038
rect 315028 222974 315080 222980
rect 314844 220380 314896 220386
rect 314844 220322 314896 220328
rect 313924 219292 313976 219298
rect 313924 219234 313976 219240
rect 314016 219156 314068 219162
rect 314016 219098 314068 219104
rect 312326 217110 312400 217138
rect 313154 217246 313228 217274
rect 312326 216988 312354 217110
rect 313154 216988 313182 217246
rect 314028 217138 314056 219098
rect 314856 217274 314884 220322
rect 315684 217274 315712 225694
rect 316328 222902 316356 231676
rect 316512 231662 316986 231690
rect 316316 222896 316368 222902
rect 316316 222838 316368 222844
rect 316512 221218 316540 231662
rect 317616 227050 317644 231676
rect 318260 229770 318288 231676
rect 318248 229764 318300 229770
rect 318248 229706 318300 229712
rect 318064 229628 318116 229634
rect 318064 229570 318116 229576
rect 317604 227044 317656 227050
rect 317604 226986 317656 226992
rect 316684 223032 316736 223038
rect 316684 222974 316736 222980
rect 316328 221190 316540 221218
rect 316328 220250 316356 221190
rect 316316 220244 316368 220250
rect 316316 220186 316368 220192
rect 316500 220244 316552 220250
rect 316500 220186 316552 220192
rect 316512 217274 316540 220186
rect 316696 218482 316724 222974
rect 318076 219434 318104 229570
rect 318904 228410 318932 231676
rect 318892 228404 318944 228410
rect 318892 228346 318944 228352
rect 319548 224126 319576 231676
rect 320192 225622 320220 231676
rect 320836 228546 320864 231676
rect 321112 231662 321494 231690
rect 320824 228540 320876 228546
rect 320824 228482 320876 228488
rect 320180 225616 320232 225622
rect 320180 225558 320232 225564
rect 319996 224664 320048 224670
rect 319996 224606 320048 224612
rect 319812 224392 319864 224398
rect 319812 224334 319864 224340
rect 319536 224120 319588 224126
rect 319536 224062 319588 224068
rect 318248 222012 318300 222018
rect 318248 221954 318300 221960
rect 318260 219434 318288 221954
rect 317984 219406 318104 219434
rect 318168 219406 318288 219434
rect 316684 218476 316736 218482
rect 316684 218418 316736 218424
rect 317984 218074 318012 219406
rect 317328 218068 317380 218074
rect 317328 218010 317380 218016
rect 317972 218068 318024 218074
rect 317972 218010 318024 218016
rect 313982 217110 314056 217138
rect 314810 217246 314884 217274
rect 315638 217246 315712 217274
rect 316466 217246 316540 217274
rect 313982 216988 314010 217110
rect 314810 216988 314838 217246
rect 315638 216988 315666 217246
rect 316466 216988 316494 217246
rect 317340 217138 317368 218010
rect 318168 217274 318196 219406
rect 319824 218074 319852 224334
rect 318984 218068 319036 218074
rect 318984 218010 319036 218016
rect 319812 218068 319864 218074
rect 319812 218010 319864 218016
rect 317294 217110 317368 217138
rect 318122 217246 318196 217274
rect 317294 216988 317322 217110
rect 318122 216988 318150 217246
rect 318996 217138 319024 218010
rect 320008 217274 320036 224606
rect 321112 223174 321140 231662
rect 322124 226302 322152 231676
rect 322400 231662 322782 231690
rect 322112 226296 322164 226302
rect 322112 226238 322164 226244
rect 321376 225616 321428 225622
rect 321376 225558 321428 225564
rect 321100 223168 321152 223174
rect 321100 223110 321152 223116
rect 320640 219292 320692 219298
rect 320640 219234 320692 219240
rect 318950 217110 319024 217138
rect 319778 217246 320036 217274
rect 318950 216988 318978 217110
rect 319778 216988 319806 217246
rect 320652 217138 320680 219234
rect 321388 217274 321416 225558
rect 321560 220788 321612 220794
rect 321560 220730 321612 220736
rect 321572 218754 321600 220730
rect 322400 220114 322428 231662
rect 323412 230314 323440 231676
rect 323688 231662 324070 231690
rect 324516 231662 324714 231690
rect 324976 231662 325358 231690
rect 325896 231662 326002 231690
rect 326264 231662 326646 231690
rect 323400 230308 323452 230314
rect 323400 230250 323452 230256
rect 322848 227044 322900 227050
rect 322848 226986 322900 226992
rect 322388 220108 322440 220114
rect 322388 220050 322440 220056
rect 321560 218748 321612 218754
rect 321560 218690 321612 218696
rect 322860 218074 322888 226986
rect 323688 224262 323716 231662
rect 323676 224256 323728 224262
rect 323676 224198 323728 224204
rect 323952 224256 324004 224262
rect 323952 224198 324004 224204
rect 322296 218068 322348 218074
rect 322296 218010 322348 218016
rect 322848 218068 322900 218074
rect 322848 218010 322900 218016
rect 323124 218068 323176 218074
rect 323124 218010 323176 218016
rect 321388 217246 321462 217274
rect 320606 217110 320680 217138
rect 320606 216988 320634 217110
rect 321434 216988 321462 217246
rect 322308 217138 322336 218010
rect 323136 217138 323164 218010
rect 323964 217274 323992 224198
rect 324136 222896 324188 222902
rect 324136 222838 324188 222844
rect 324148 218074 324176 222838
rect 324516 220794 324544 231662
rect 324976 226914 325004 231662
rect 325424 228540 325476 228546
rect 325424 228482 325476 228488
rect 324964 226908 325016 226914
rect 324964 226850 325016 226856
rect 324504 220788 324556 220794
rect 324504 220730 324556 220736
rect 325436 218074 325464 228482
rect 325608 220108 325660 220114
rect 325608 220050 325660 220056
rect 324136 218068 324188 218074
rect 324136 218010 324188 218016
rect 324780 218068 324832 218074
rect 324780 218010 324832 218016
rect 325424 218068 325476 218074
rect 325424 218010 325476 218016
rect 322262 217110 322336 217138
rect 323090 217110 323164 217138
rect 323918 217246 323992 217274
rect 322262 216988 322290 217110
rect 323090 216988 323118 217110
rect 323918 216988 323946 217246
rect 324792 217138 324820 218010
rect 325620 217274 325648 220050
rect 325896 219978 325924 231662
rect 326264 221474 326292 231662
rect 326896 229084 326948 229090
rect 326896 229026 326948 229032
rect 326252 221468 326304 221474
rect 326252 221410 326304 221416
rect 325884 219972 325936 219978
rect 325884 219914 325936 219920
rect 326908 218074 326936 229026
rect 327276 223038 327304 231676
rect 327552 231662 327934 231690
rect 327552 225894 327580 231662
rect 327540 225888 327592 225894
rect 327540 225830 327592 225836
rect 327724 225004 327776 225010
rect 327724 224946 327776 224952
rect 327264 223032 327316 223038
rect 327264 222974 327316 222980
rect 327736 218890 327764 224946
rect 328564 223310 328592 231676
rect 329208 228682 329236 231676
rect 329852 230042 329880 231676
rect 329840 230036 329892 230042
rect 329840 229978 329892 229984
rect 330496 228818 330524 231676
rect 330944 230036 330996 230042
rect 330944 229978 330996 229984
rect 330956 229094 330984 229978
rect 330956 229066 331076 229094
rect 330484 228812 330536 228818
rect 330484 228754 330536 228760
rect 329196 228676 329248 228682
rect 329196 228618 329248 228624
rect 330484 228404 330536 228410
rect 330484 228346 330536 228352
rect 329748 226024 329800 226030
rect 329748 225966 329800 225972
rect 328552 223304 328604 223310
rect 328552 223246 328604 223252
rect 328092 223032 328144 223038
rect 328092 222974 328144 222980
rect 327724 218884 327776 218890
rect 327724 218826 327776 218832
rect 327264 218748 327316 218754
rect 327264 218690 327316 218696
rect 326436 218068 326488 218074
rect 326436 218010 326488 218016
rect 326896 218068 326948 218074
rect 326896 218010 326948 218016
rect 324746 217110 324820 217138
rect 325574 217246 325648 217274
rect 324746 216988 324774 217110
rect 325574 216988 325602 217246
rect 326448 217138 326476 218010
rect 327276 217138 327304 218690
rect 328104 217274 328132 222974
rect 328920 218204 328972 218210
rect 328920 218146 328972 218152
rect 326402 217110 326476 217138
rect 327230 217110 327304 217138
rect 328058 217246 328132 217274
rect 326402 216988 326430 217110
rect 327230 216988 327258 217110
rect 328058 216988 328086 217246
rect 328932 217138 328960 218146
rect 329760 217274 329788 225966
rect 330496 218210 330524 228346
rect 330484 218204 330536 218210
rect 330484 218146 330536 218152
rect 331048 218074 331076 229066
rect 331140 228970 331168 231676
rect 331140 228954 331260 228970
rect 331140 228948 331272 228954
rect 331140 228942 331220 228948
rect 331220 228890 331272 228896
rect 331784 224534 331812 231676
rect 332060 231662 332442 231690
rect 332796 231662 333086 231690
rect 332060 225010 332088 231662
rect 332232 225888 332284 225894
rect 332232 225830 332284 225836
rect 332048 225004 332100 225010
rect 332048 224946 332100 224952
rect 331772 224528 331824 224534
rect 331772 224470 331824 224476
rect 331404 222148 331456 222154
rect 331404 222090 331456 222096
rect 330576 218068 330628 218074
rect 330576 218010 330628 218016
rect 331036 218068 331088 218074
rect 331036 218010 331088 218016
rect 328886 217110 328960 217138
rect 329714 217246 329788 217274
rect 328886 216988 328914 217110
rect 329714 216988 329742 217246
rect 330588 217138 330616 218010
rect 331416 217274 331444 222090
rect 332244 217274 332272 225830
rect 332796 221746 332824 231662
rect 333716 227458 333744 231676
rect 334084 231662 334374 231690
rect 333704 227452 333756 227458
rect 333704 227394 333756 227400
rect 333888 227452 333940 227458
rect 333888 227394 333940 227400
rect 332784 221740 332836 221746
rect 332784 221682 332836 221688
rect 332692 219564 332744 219570
rect 332692 219506 332744 219512
rect 332704 219026 332732 219506
rect 333704 219428 333756 219434
rect 333704 219370 333756 219376
rect 332692 219020 332744 219026
rect 332692 218962 332744 218968
rect 333060 218068 333112 218074
rect 333060 218010 333112 218016
rect 330542 217110 330616 217138
rect 331370 217246 331444 217274
rect 332198 217246 332272 217274
rect 330542 216988 330570 217110
rect 331370 216988 331398 217246
rect 332198 216988 332226 217246
rect 333072 217138 333100 218010
rect 333716 217274 333744 219370
rect 333900 218074 333928 227394
rect 334084 220658 334112 231662
rect 335004 230178 335032 231676
rect 334992 230172 335044 230178
rect 334992 230114 335044 230120
rect 335176 230172 335228 230178
rect 335176 230114 335228 230120
rect 335188 229094 335216 230114
rect 335004 229066 335216 229094
rect 335004 224262 335032 229066
rect 335176 224528 335228 224534
rect 335176 224470 335228 224476
rect 334992 224256 335044 224262
rect 334992 224198 335044 224204
rect 334072 220652 334124 220658
rect 334072 220594 334124 220600
rect 335188 218074 335216 224470
rect 335648 223582 335676 231676
rect 336292 226166 336320 231676
rect 336464 228676 336516 228682
rect 336464 228618 336516 228624
rect 336280 226160 336332 226166
rect 336280 226102 336332 226108
rect 335636 223576 335688 223582
rect 335636 223518 335688 223524
rect 336004 223372 336056 223378
rect 336004 223314 336056 223320
rect 336016 219162 336044 223314
rect 336476 219434 336504 228618
rect 336936 227186 336964 231676
rect 337212 231662 337594 231690
rect 336924 227180 336976 227186
rect 336924 227122 336976 227128
rect 337212 219570 337240 231662
rect 338224 227322 338252 231676
rect 338212 227316 338264 227322
rect 338212 227258 338264 227264
rect 338672 227180 338724 227186
rect 338672 227122 338724 227128
rect 338028 220516 338080 220522
rect 338028 220458 338080 220464
rect 337200 219564 337252 219570
rect 337200 219506 337252 219512
rect 336384 219406 336504 219434
rect 336004 219156 336056 219162
rect 336004 219098 336056 219104
rect 333888 218068 333940 218074
rect 333888 218010 333940 218016
rect 334716 218068 334768 218074
rect 334716 218010 334768 218016
rect 335176 218068 335228 218074
rect 335176 218010 335228 218016
rect 335544 218068 335596 218074
rect 335544 218010 335596 218016
rect 333716 217246 333882 217274
rect 333026 217110 333100 217138
rect 333026 216988 333054 217110
rect 333854 216988 333882 217246
rect 334728 217138 334756 218010
rect 335556 217138 335584 218010
rect 336384 217274 336412 219406
rect 337200 219020 337252 219026
rect 337200 218962 337252 218968
rect 334682 217110 334756 217138
rect 335510 217110 335584 217138
rect 336338 217246 336412 217274
rect 334682 216988 334710 217110
rect 335510 216988 335538 217110
rect 336338 216988 336366 217246
rect 337212 217138 337240 218962
rect 338040 217274 338068 220458
rect 338684 218074 338712 227122
rect 338868 224806 338896 231676
rect 339526 231662 339724 231690
rect 338856 224800 338908 224806
rect 338856 224742 338908 224748
rect 339408 224256 339460 224262
rect 339408 224198 339460 224204
rect 339420 218074 339448 224198
rect 339696 221610 339724 231662
rect 340156 229906 340184 231676
rect 340432 231662 340814 231690
rect 341076 231662 341458 231690
rect 340144 229900 340196 229906
rect 340144 229842 340196 229848
rect 340432 221882 340460 231662
rect 340696 227316 340748 227322
rect 340696 227258 340748 227264
rect 340420 221876 340472 221882
rect 340420 221818 340472 221824
rect 339684 221604 339736 221610
rect 339684 221546 339736 221552
rect 340512 218884 340564 218890
rect 340512 218826 340564 218832
rect 338672 218068 338724 218074
rect 338672 218010 338724 218016
rect 338856 218068 338908 218074
rect 338856 218010 338908 218016
rect 339408 218068 339460 218074
rect 339408 218010 339460 218016
rect 339684 218068 339736 218074
rect 339684 218010 339736 218016
rect 337166 217110 337240 217138
rect 337994 217246 338068 217274
rect 337166 216988 337194 217110
rect 337994 216988 338022 217246
rect 338868 217138 338896 218010
rect 339696 217138 339724 218010
rect 340524 217138 340552 218826
rect 340708 218074 340736 227258
rect 341076 220386 341104 231662
rect 342088 223514 342116 231676
rect 342272 231662 342746 231690
rect 342916 231662 343390 231690
rect 343836 231662 344034 231690
rect 342076 223508 342128 223514
rect 342076 223450 342128 223456
rect 342272 223378 342300 231662
rect 342916 229094 342944 231662
rect 342640 229066 342944 229094
rect 342260 223372 342312 223378
rect 342260 223314 342312 223320
rect 341340 221604 341392 221610
rect 341340 221546 341392 221552
rect 341064 220380 341116 220386
rect 341064 220322 341116 220328
rect 340696 218068 340748 218074
rect 340696 218010 340748 218016
rect 341352 217274 341380 221546
rect 342168 221468 342220 221474
rect 342168 221410 342220 221416
rect 342180 217274 342208 221410
rect 342640 220250 342668 229066
rect 342812 223440 342864 223446
rect 342812 223382 342864 223388
rect 342628 220244 342680 220250
rect 342628 220186 342680 220192
rect 342824 219298 342852 223382
rect 343836 222018 343864 231662
rect 344664 225758 344692 231676
rect 345308 229770 345336 231676
rect 345664 229900 345716 229906
rect 345664 229842 345716 229848
rect 345296 229764 345348 229770
rect 345296 229706 345348 229712
rect 344652 225752 344704 225758
rect 344652 225694 344704 225700
rect 344652 223168 344704 223174
rect 344652 223110 344704 223116
rect 343824 222012 343876 222018
rect 343824 221954 343876 221960
rect 342996 220380 343048 220386
rect 342996 220322 343048 220328
rect 342812 219292 342864 219298
rect 342812 219234 342864 219240
rect 343008 217274 343036 220322
rect 343824 219156 343876 219162
rect 343824 219098 343876 219104
rect 338822 217110 338896 217138
rect 339650 217110 339724 217138
rect 340478 217110 340552 217138
rect 341306 217246 341380 217274
rect 342134 217246 342208 217274
rect 342962 217246 343036 217274
rect 338822 216988 338850 217110
rect 339650 216988 339678 217110
rect 340478 216988 340506 217110
rect 341306 216988 341334 217246
rect 342134 216988 342162 217246
rect 342962 216988 342990 217246
rect 343836 217138 343864 219098
rect 344664 217274 344692 223110
rect 345676 219026 345704 229842
rect 345952 224670 345980 231676
rect 346596 225622 346624 231676
rect 346584 225616 346636 225622
rect 346584 225558 346636 225564
rect 347044 225616 347096 225622
rect 347044 225558 347096 225564
rect 345940 224664 345992 224670
rect 345940 224606 345992 224612
rect 346216 224664 346268 224670
rect 346216 224606 346268 224612
rect 345664 219020 345716 219026
rect 345664 218962 345716 218968
rect 345480 218068 345532 218074
rect 345480 218010 345532 218016
rect 343790 217110 343864 217138
rect 344618 217246 344692 217274
rect 343790 216988 343818 217110
rect 344618 216988 344646 217246
rect 345492 217138 345520 218010
rect 346228 217274 346256 224606
rect 347056 218074 347084 225558
rect 347240 224398 347268 231676
rect 347228 224392 347280 224398
rect 347228 224334 347280 224340
rect 347884 223446 347912 231676
rect 347872 223440 347924 223446
rect 347872 223382 347924 223388
rect 347228 223304 347280 223310
rect 347228 223246 347280 223252
rect 347240 219434 347268 223246
rect 348528 222902 348556 231676
rect 349172 228546 349200 231676
rect 349160 228540 349212 228546
rect 349160 228482 349212 228488
rect 349816 227050 349844 231676
rect 350460 230178 350488 231676
rect 350448 230172 350500 230178
rect 350448 230114 350500 230120
rect 351104 229090 351132 231676
rect 351472 231662 351762 231690
rect 352116 231662 352406 231690
rect 351092 229084 351144 229090
rect 351092 229026 351144 229032
rect 350448 228540 350500 228546
rect 350448 228482 350500 228488
rect 349804 227044 349856 227050
rect 349804 226986 349856 226992
rect 350264 226364 350316 226370
rect 350264 226306 350316 226312
rect 348516 222896 348568 222902
rect 348516 222838 348568 222844
rect 349068 222896 349120 222902
rect 349068 222838 349120 222844
rect 348792 220244 348844 220250
rect 348792 220186 348844 220192
rect 347228 219428 347280 219434
rect 347228 219370 347280 219376
rect 347228 219020 347280 219026
rect 347228 218962 347280 218968
rect 347044 218068 347096 218074
rect 347044 218010 347096 218016
rect 347240 217274 347268 218962
rect 347964 218068 348016 218074
rect 347964 218010 348016 218016
rect 346228 217246 346302 217274
rect 345446 217110 345520 217138
rect 345446 216988 345474 217110
rect 346274 216988 346302 217246
rect 347102 217246 347268 217274
rect 347102 216988 347130 217246
rect 347976 217138 348004 218010
rect 348804 217274 348832 220186
rect 349080 218074 349108 222838
rect 350276 219434 350304 226306
rect 350460 219434 350488 228482
rect 351092 226500 351144 226506
rect 351092 226442 351144 226448
rect 349620 219428 349672 219434
rect 350276 219406 350396 219434
rect 350460 219428 350592 219434
rect 350460 219406 350540 219428
rect 349620 219370 349672 219376
rect 349068 218068 349120 218074
rect 349068 218010 349120 218016
rect 347930 217110 348004 217138
rect 348758 217246 348832 217274
rect 347930 216988 347958 217110
rect 348758 216988 348786 217246
rect 349632 217138 349660 219370
rect 350368 217274 350396 219406
rect 350540 219370 350592 219376
rect 351104 218754 351132 226442
rect 351472 223038 351500 231662
rect 351736 229764 351788 229770
rect 351736 229706 351788 229712
rect 351748 226370 351776 229706
rect 351736 226364 351788 226370
rect 351736 226306 351788 226312
rect 351460 223032 351512 223038
rect 351460 222974 351512 222980
rect 351276 221876 351328 221882
rect 351276 221818 351328 221824
rect 351092 218748 351144 218754
rect 351092 218690 351144 218696
rect 351288 217274 351316 221818
rect 352116 220114 352144 231662
rect 353036 226506 353064 231676
rect 353024 226500 353076 226506
rect 353024 226442 353076 226448
rect 353680 226030 353708 231676
rect 353864 231662 354338 231690
rect 353668 226024 353720 226030
rect 353668 225966 353720 225972
rect 352932 225752 352984 225758
rect 352932 225694 352984 225700
rect 352104 220108 352156 220114
rect 352104 220050 352156 220056
rect 352104 219428 352156 219434
rect 352104 219370 352156 219376
rect 350368 217246 350442 217274
rect 349586 217110 349660 217138
rect 349586 216988 349614 217110
rect 350414 216988 350442 217246
rect 351242 217246 351316 217274
rect 351242 216988 351270 217246
rect 352116 217138 352144 219370
rect 352944 217274 352972 225694
rect 353864 223122 353892 231662
rect 354968 228410 354996 231676
rect 355612 230042 355640 231676
rect 355600 230036 355652 230042
rect 355600 229978 355652 229984
rect 354956 228404 355008 228410
rect 354956 228346 355008 228352
rect 355324 228404 355376 228410
rect 355324 228346 355376 228352
rect 354588 226024 354640 226030
rect 354588 225966 354640 225972
rect 353772 223094 353892 223122
rect 353772 222154 353800 223094
rect 353944 223032 353996 223038
rect 353944 222974 353996 222980
rect 353760 222148 353812 222154
rect 353760 222090 353812 222096
rect 353956 219162 353984 222974
rect 353944 219156 353996 219162
rect 353944 219098 353996 219104
rect 353760 218748 353812 218754
rect 353760 218690 353812 218696
rect 352070 217110 352144 217138
rect 352898 217246 352972 217274
rect 352070 216988 352098 217110
rect 352898 216988 352926 217246
rect 353772 217138 353800 218690
rect 354600 217274 354628 225966
rect 355336 219434 355364 228346
rect 356256 227458 356284 231676
rect 356244 227452 356296 227458
rect 356244 227394 356296 227400
rect 355876 227044 355928 227050
rect 355876 226986 355928 226992
rect 355324 219428 355376 219434
rect 355324 219370 355376 219376
rect 355888 218074 355916 226986
rect 356900 224534 356928 231676
rect 357072 227452 357124 227458
rect 357072 227394 357124 227400
rect 356888 224528 356940 224534
rect 356888 224470 356940 224476
rect 357084 222034 357112 227394
rect 357544 225894 357572 231676
rect 357912 231662 358202 231690
rect 357532 225888 357584 225894
rect 357532 225830 357584 225836
rect 357912 223310 357940 231662
rect 358832 228682 358860 231676
rect 359016 231662 359490 231690
rect 358820 228676 358872 228682
rect 358820 228618 358872 228624
rect 358084 224120 358136 224126
rect 358084 224062 358136 224068
rect 357900 223304 357952 223310
rect 357900 223246 357952 223252
rect 356992 222006 357112 222034
rect 356992 218074 357020 222006
rect 357164 221740 357216 221746
rect 357164 221682 357216 221688
rect 355416 218068 355468 218074
rect 355416 218010 355468 218016
rect 355876 218068 355928 218074
rect 355876 218010 355928 218016
rect 356244 218068 356296 218074
rect 356244 218010 356296 218016
rect 356980 218068 357032 218074
rect 356980 218010 357032 218016
rect 353726 217110 353800 217138
rect 354554 217246 354628 217274
rect 353726 216988 353754 217110
rect 354554 216988 354582 217246
rect 355428 217138 355456 218010
rect 356256 217138 356284 218010
rect 357176 217274 357204 221682
rect 357900 220652 357952 220658
rect 357900 220594 357952 220600
rect 357912 217274 357940 220594
rect 358096 218890 358124 224062
rect 359016 220522 359044 231662
rect 359924 228676 359976 228682
rect 359924 228618 359976 228624
rect 359004 220516 359056 220522
rect 359004 220458 359056 220464
rect 358820 220108 358872 220114
rect 358820 220050 358872 220056
rect 358832 219434 358860 220050
rect 358740 219406 358860 219434
rect 359936 219434 359964 228618
rect 360120 227186 360148 231676
rect 360764 229906 360792 231676
rect 360752 229900 360804 229906
rect 360752 229842 360804 229848
rect 361212 229900 361264 229906
rect 361212 229842 361264 229848
rect 361224 229094 361252 229842
rect 361040 229066 361252 229094
rect 360108 227180 360160 227186
rect 360108 227122 360160 227128
rect 359936 219406 360148 219434
rect 358084 218884 358136 218890
rect 358084 218826 358136 218832
rect 358740 217274 358768 219406
rect 360120 218074 360148 219406
rect 361040 218074 361068 229066
rect 361408 227322 361436 231676
rect 361776 231662 362066 231690
rect 362328 231662 362710 231690
rect 361396 227316 361448 227322
rect 361396 227258 361448 227264
rect 361212 224392 361264 224398
rect 361212 224334 361264 224340
rect 359556 218068 359608 218074
rect 359556 218010 359608 218016
rect 360108 218068 360160 218074
rect 360108 218010 360160 218016
rect 360384 218068 360436 218074
rect 360384 218010 360436 218016
rect 361028 218068 361080 218074
rect 361028 218010 361080 218016
rect 355382 217110 355456 217138
rect 356210 217110 356284 217138
rect 357038 217246 357204 217274
rect 357866 217246 357940 217274
rect 358694 217246 358768 217274
rect 355382 216988 355410 217110
rect 356210 216988 356238 217110
rect 357038 216988 357066 217246
rect 357866 216988 357894 217246
rect 358694 216988 358722 217246
rect 359568 217138 359596 218010
rect 360396 217138 360424 218010
rect 361224 217274 361252 224334
rect 361776 221610 361804 231662
rect 362328 224262 362356 231662
rect 363340 229094 363368 231676
rect 363524 231662 363998 231690
rect 363524 229094 363552 231662
rect 363248 229066 363368 229094
rect 363432 229066 363552 229094
rect 362776 227180 362828 227186
rect 362776 227122 362828 227128
rect 362316 224256 362368 224262
rect 362316 224198 362368 224204
rect 361764 221604 361816 221610
rect 361764 221546 361816 221552
rect 362040 219428 362092 219434
rect 362040 219370 362092 219376
rect 359522 217110 359596 217138
rect 360350 217110 360424 217138
rect 361178 217246 361252 217274
rect 359522 216988 359550 217110
rect 360350 216988 360378 217110
rect 361178 216988 361206 217246
rect 362052 217138 362080 219370
rect 362788 217274 362816 227122
rect 363248 224126 363276 229066
rect 363236 224120 363288 224126
rect 363236 224062 363288 224068
rect 363432 220386 363460 229066
rect 363604 224256 363656 224262
rect 363604 224198 363656 224204
rect 363420 220380 363472 220386
rect 363420 220322 363472 220328
rect 363616 219026 363644 224198
rect 364628 223174 364656 231676
rect 364812 231662 365286 231690
rect 364616 223168 364668 223174
rect 364616 223110 364668 223116
rect 364812 221474 364840 231662
rect 365536 223168 365588 223174
rect 365536 223110 365588 223116
rect 364800 221468 364852 221474
rect 364800 221410 364852 221416
rect 363604 219020 363656 219026
rect 363604 218962 363656 218968
rect 363696 218884 363748 218890
rect 363696 218826 363748 218832
rect 362788 217246 362862 217274
rect 362006 217110 362080 217138
rect 362006 216988 362034 217110
rect 362834 216988 362862 217246
rect 363708 217138 363736 218826
rect 365352 218204 365404 218210
rect 365352 218146 365404 218152
rect 364524 218068 364576 218074
rect 364524 218010 364576 218016
rect 364536 217138 364564 218010
rect 365364 217138 365392 218146
rect 365548 218074 365576 223110
rect 365916 223038 365944 231676
rect 366560 224670 366588 231676
rect 366548 224664 366600 224670
rect 366548 224606 366600 224612
rect 366732 224528 366784 224534
rect 366732 224470 366784 224476
rect 365904 223032 365956 223038
rect 365904 222974 365956 222980
rect 366744 218074 366772 224470
rect 366916 223032 366968 223038
rect 366916 222974 366968 222980
rect 365536 218068 365588 218074
rect 365536 218010 365588 218016
rect 366180 218068 366232 218074
rect 366180 218010 366232 218016
rect 366732 218068 366784 218074
rect 366732 218010 366784 218016
rect 366192 217138 366220 218010
rect 366928 217274 366956 222974
rect 367204 222902 367232 231676
rect 367848 225622 367876 231676
rect 367836 225616 367888 225622
rect 367836 225558 367888 225564
rect 368492 224262 368520 231676
rect 369136 228546 369164 231676
rect 369320 231662 369794 231690
rect 369964 231662 370438 231690
rect 369124 228540 369176 228546
rect 369124 228482 369176 228488
rect 369124 225004 369176 225010
rect 369124 224946 369176 224952
rect 368480 224256 368532 224262
rect 368480 224198 368532 224204
rect 367192 222896 367244 222902
rect 367192 222838 367244 222844
rect 368388 222896 368440 222902
rect 368388 222838 368440 222844
rect 367652 222012 367704 222018
rect 367652 221954 367704 221960
rect 367664 219434 367692 221954
rect 367652 219428 367704 219434
rect 367652 219370 367704 219376
rect 368400 218074 368428 222838
rect 368664 219020 368716 219026
rect 368664 218962 368716 218968
rect 367836 218068 367888 218074
rect 367836 218010 367888 218016
rect 368388 218068 368440 218074
rect 368388 218010 368440 218016
rect 366928 217246 367002 217274
rect 363662 217110 363736 217138
rect 364490 217110 364564 217138
rect 365318 217110 365392 217138
rect 366146 217110 366220 217138
rect 363662 216988 363690 217110
rect 364490 216988 364518 217110
rect 365318 216988 365346 217110
rect 366146 216988 366174 217110
rect 366974 216988 367002 217246
rect 367848 217138 367876 218010
rect 368676 217138 368704 218962
rect 369136 218754 369164 224946
rect 369320 221882 369348 231662
rect 369308 221876 369360 221882
rect 369308 221818 369360 221824
rect 369492 221604 369544 221610
rect 369492 221546 369544 221552
rect 369124 218748 369176 218754
rect 369124 218690 369176 218696
rect 369504 217274 369532 221546
rect 369964 220250 369992 231662
rect 371068 229770 371096 231676
rect 371056 229764 371108 229770
rect 371056 229706 371108 229712
rect 371712 229094 371740 231676
rect 371620 229066 371740 229094
rect 371056 228540 371108 228546
rect 371056 228482 371108 228488
rect 369952 220244 370004 220250
rect 369952 220186 370004 220192
rect 370504 220244 370556 220250
rect 370504 220186 370556 220192
rect 370516 218890 370544 220186
rect 370504 218884 370556 218890
rect 370504 218826 370556 218832
rect 370320 218748 370372 218754
rect 370320 218690 370372 218696
rect 370332 217274 370360 218690
rect 367802 217110 367876 217138
rect 368630 217110 368704 217138
rect 369458 217246 369532 217274
rect 370286 217246 370360 217274
rect 371068 217274 371096 228482
rect 371620 225758 371648 229066
rect 372356 226030 372384 231676
rect 373000 228410 373028 231676
rect 372988 228404 373040 228410
rect 372988 228346 373040 228352
rect 373448 228404 373500 228410
rect 373448 228346 373500 228352
rect 372344 226024 372396 226030
rect 372344 225966 372396 225972
rect 371608 225752 371660 225758
rect 371608 225694 371660 225700
rect 371792 225752 371844 225758
rect 371792 225694 371844 225700
rect 371804 218210 371832 225694
rect 372528 225616 372580 225622
rect 372528 225558 372580 225564
rect 371792 218204 371844 218210
rect 371792 218146 371844 218152
rect 372540 218074 372568 225558
rect 373460 218074 373488 228346
rect 373644 225010 373672 231676
rect 374288 227458 374316 231676
rect 374472 231662 374946 231690
rect 374276 227452 374328 227458
rect 374276 227394 374328 227400
rect 373816 225888 373868 225894
rect 373816 225830 373868 225836
rect 373632 225004 373684 225010
rect 373632 224946 373684 224952
rect 373828 219434 373856 225830
rect 374472 220658 374500 231662
rect 374644 230444 374696 230450
rect 374644 230386 374696 230392
rect 374656 221746 374684 230386
rect 375576 227050 375604 231676
rect 376220 230450 376248 231676
rect 376208 230444 376260 230450
rect 376208 230386 376260 230392
rect 376024 228812 376076 228818
rect 376024 228754 376076 228760
rect 375564 227044 375616 227050
rect 375564 226986 375616 226992
rect 374644 221740 374696 221746
rect 374644 221682 374696 221688
rect 375288 221468 375340 221474
rect 375288 221410 375340 221416
rect 374460 220652 374512 220658
rect 374460 220594 374512 220600
rect 373644 219406 373856 219434
rect 371976 218068 372028 218074
rect 371976 218010 372028 218016
rect 372528 218068 372580 218074
rect 372528 218010 372580 218016
rect 372804 218068 372856 218074
rect 372804 218010 372856 218016
rect 373448 218068 373500 218074
rect 373448 218010 373500 218016
rect 371068 217246 371142 217274
rect 367802 216988 367830 217110
rect 368630 216988 368658 217110
rect 369458 216988 369486 217246
rect 370286 216988 370314 217246
rect 371114 216988 371142 217246
rect 371988 217138 372016 218010
rect 372816 217138 372844 218010
rect 373644 217274 373672 219406
rect 374460 218204 374512 218210
rect 374460 218146 374512 218152
rect 371942 217110 372016 217138
rect 372770 217110 372844 217138
rect 373598 217246 373672 217274
rect 371942 216988 371970 217110
rect 372770 216988 372798 217110
rect 373598 216988 373626 217246
rect 374472 217138 374500 218146
rect 375300 217274 375328 221410
rect 376036 218210 376064 228754
rect 376864 228682 376892 231676
rect 376852 228676 376904 228682
rect 376852 228618 376904 228624
rect 376668 227044 376720 227050
rect 376668 226986 376720 226992
rect 376024 218204 376076 218210
rect 376024 218146 376076 218152
rect 376680 218074 376708 226986
rect 377508 224398 377536 231676
rect 378166 231662 378364 231690
rect 377680 229764 377732 229770
rect 377680 229706 377732 229712
rect 377692 225894 377720 229706
rect 377680 225888 377732 225894
rect 377680 225830 377732 225836
rect 377864 225888 377916 225894
rect 377864 225830 377916 225836
rect 377496 224392 377548 224398
rect 377496 224334 377548 224340
rect 377404 224052 377456 224058
rect 377404 223994 377456 224000
rect 377416 219026 377444 223994
rect 377876 219434 377904 225830
rect 378336 220114 378364 231662
rect 378796 229906 378824 231676
rect 378784 229900 378836 229906
rect 378784 229842 378836 229848
rect 379440 227186 379468 231676
rect 379624 231662 380098 231690
rect 380268 231662 380742 231690
rect 381096 231662 381386 231690
rect 381648 231662 382030 231690
rect 382384 231662 382674 231690
rect 382844 231662 383318 231690
rect 379428 227180 379480 227186
rect 379428 227122 379480 227128
rect 379244 224256 379296 224262
rect 379244 224198 379296 224204
rect 378324 220108 378376 220114
rect 378324 220050 378376 220056
rect 377784 219406 377904 219434
rect 377404 219020 377456 219026
rect 377404 218962 377456 218968
rect 376944 218884 376996 218890
rect 376944 218826 376996 218832
rect 376116 218068 376168 218074
rect 376116 218010 376168 218016
rect 376668 218068 376720 218074
rect 376668 218010 376720 218016
rect 374426 217110 374500 217138
rect 375254 217246 375328 217274
rect 374426 216988 374454 217110
rect 375254 216988 375282 217246
rect 376128 217138 376156 218010
rect 376956 217138 376984 218826
rect 377784 217274 377812 219406
rect 379256 218074 379284 224198
rect 379624 223174 379652 231662
rect 379612 223168 379664 223174
rect 379612 223110 379664 223116
rect 380072 223168 380124 223174
rect 380072 223110 380124 223116
rect 379428 220108 379480 220114
rect 379428 220050 379480 220056
rect 378600 218068 378652 218074
rect 378600 218010 378652 218016
rect 379244 218068 379296 218074
rect 379244 218010 379296 218016
rect 376082 217110 376156 217138
rect 376910 217110 376984 217138
rect 377738 217246 377812 217274
rect 376082 216988 376110 217110
rect 376910 216988 376938 217110
rect 377738 216988 377766 217246
rect 378612 217138 378640 218010
rect 379440 217274 379468 220050
rect 380084 218754 380112 223110
rect 380268 222018 380296 231662
rect 380256 222012 380308 222018
rect 380256 221954 380308 221960
rect 381096 220250 381124 231662
rect 381648 224534 381676 231662
rect 382096 227180 382148 227186
rect 382096 227122 382148 227128
rect 381636 224528 381688 224534
rect 381636 224470 381688 224476
rect 381084 220244 381136 220250
rect 381084 220186 381136 220192
rect 380256 219428 380308 219434
rect 380256 219370 380308 219376
rect 380072 218748 380124 218754
rect 380072 218690 380124 218696
rect 378566 217110 378640 217138
rect 379394 217246 379468 217274
rect 378566 216988 378594 217110
rect 379394 216988 379422 217246
rect 380268 217138 380296 219370
rect 381912 218204 381964 218210
rect 381912 218146 381964 218152
rect 381084 218068 381136 218074
rect 381084 218010 381136 218016
rect 381096 217138 381124 218010
rect 381924 217138 381952 218146
rect 382108 218074 382136 227122
rect 382384 222902 382412 231662
rect 382844 229094 382872 231662
rect 382752 229066 382872 229094
rect 382752 225758 382780 229066
rect 382740 225752 382792 225758
rect 382740 225694 382792 225700
rect 382924 225752 382976 225758
rect 382924 225694 382976 225700
rect 382372 222896 382424 222902
rect 382372 222838 382424 222844
rect 382740 218884 382792 218890
rect 382740 218826 382792 218832
rect 382096 218068 382148 218074
rect 382096 218010 382148 218016
rect 382752 217138 382780 218826
rect 382936 218210 382964 225694
rect 383948 223038 383976 231676
rect 384132 231662 384606 231690
rect 383936 223032 383988 223038
rect 383936 222974 383988 222980
rect 383476 222896 383528 222902
rect 383476 222838 383528 222844
rect 383488 218890 383516 222838
rect 384132 221610 384160 231662
rect 385236 228546 385264 231676
rect 385224 228540 385276 228546
rect 385224 228482 385276 228488
rect 385880 224058 385908 231676
rect 386052 228540 386104 228546
rect 386052 228482 386104 228488
rect 385868 224052 385920 224058
rect 385868 223994 385920 224000
rect 384304 223032 384356 223038
rect 384304 222974 384356 222980
rect 384120 221604 384172 221610
rect 384120 221546 384172 221552
rect 384316 219434 384344 222974
rect 384488 221604 384540 221610
rect 384488 221546 384540 221552
rect 384500 219434 384528 221546
rect 385224 220788 385276 220794
rect 385224 220730 385276 220736
rect 384212 219428 384344 219434
rect 384264 219406 384344 219428
rect 384408 219406 384528 219434
rect 384212 219370 384264 219376
rect 383476 218884 383528 218890
rect 383476 218826 383528 218832
rect 383568 218748 383620 218754
rect 383568 218690 383620 218696
rect 382924 218204 382976 218210
rect 382924 218146 382976 218152
rect 383580 217138 383608 218690
rect 384408 217274 384436 219406
rect 385236 217274 385264 220730
rect 386064 217274 386092 228482
rect 386524 223174 386552 231676
rect 387168 228410 387196 231676
rect 387432 230376 387484 230382
rect 387432 230318 387484 230324
rect 387156 228404 387208 228410
rect 387156 228346 387208 228352
rect 387444 225622 387472 230318
rect 387812 228818 387840 231676
rect 388456 230382 388484 231676
rect 388444 230376 388496 230382
rect 388444 230318 388496 230324
rect 389100 229770 389128 231676
rect 389088 229764 389140 229770
rect 389088 229706 389140 229712
rect 388628 229628 388680 229634
rect 388628 229570 388680 229576
rect 388640 229094 388668 229570
rect 388640 229066 388760 229094
rect 387800 228812 387852 228818
rect 387800 228754 387852 228760
rect 388536 226364 388588 226370
rect 388536 226306 388588 226312
rect 387432 225616 387484 225622
rect 387432 225558 387484 225564
rect 387708 224392 387760 224398
rect 387708 224334 387760 224340
rect 386512 223168 386564 223174
rect 386512 223110 386564 223116
rect 386880 219020 386932 219026
rect 386880 218962 386932 218968
rect 380222 217110 380296 217138
rect 381050 217110 381124 217138
rect 381878 217110 381952 217138
rect 382706 217110 382780 217138
rect 383534 217110 383608 217138
rect 384362 217246 384436 217274
rect 385190 217246 385264 217274
rect 386018 217246 386092 217274
rect 380222 216988 380250 217110
rect 381050 216988 381078 217110
rect 381878 216988 381906 217110
rect 382706 216988 382734 217110
rect 383534 216988 383562 217110
rect 384362 216988 384390 217246
rect 385190 216988 385218 217246
rect 386018 216988 386046 217246
rect 386892 217138 386920 218962
rect 387720 217274 387748 224334
rect 388548 218890 388576 226306
rect 388732 220794 388760 229066
rect 389744 227050 389772 231676
rect 390008 228404 390060 228410
rect 390008 228346 390060 228352
rect 389732 227044 389784 227050
rect 389732 226986 389784 226992
rect 388720 220788 388772 220794
rect 388720 220730 388772 220736
rect 388720 220244 388772 220250
rect 388720 220186 388772 220192
rect 388536 218884 388588 218890
rect 388536 218826 388588 218832
rect 388732 217274 388760 220186
rect 390020 218074 390048 228346
rect 390388 225894 390416 231676
rect 390756 231662 391046 231690
rect 390376 225888 390428 225894
rect 390376 225830 390428 225836
rect 390192 225616 390244 225622
rect 390192 225558 390244 225564
rect 389364 218068 389416 218074
rect 389364 218010 389416 218016
rect 390008 218068 390060 218074
rect 390008 218010 390060 218016
rect 386846 217110 386920 217138
rect 387674 217246 387748 217274
rect 388502 217246 388760 217274
rect 386846 216988 386874 217110
rect 387674 216988 387702 217246
rect 388502 216988 388530 217246
rect 389376 217138 389404 218010
rect 390204 217274 390232 225558
rect 390756 221474 390784 231662
rect 391676 226370 391704 231676
rect 392136 231662 392334 231690
rect 391848 227044 391900 227050
rect 391848 226986 391900 226992
rect 391664 226364 391716 226370
rect 391664 226306 391716 226312
rect 391020 221740 391072 221746
rect 391020 221682 391072 221688
rect 390744 221468 390796 221474
rect 390744 221410 390796 221416
rect 391032 217274 391060 221682
rect 391860 219434 391888 226986
rect 392136 220114 392164 231662
rect 392964 227186 392992 231676
rect 392952 227180 393004 227186
rect 392952 227122 393004 227128
rect 393136 227180 393188 227186
rect 393136 227122 393188 227128
rect 392124 220108 392176 220114
rect 392124 220050 392176 220056
rect 389330 217110 389404 217138
rect 390158 217246 390232 217274
rect 390986 217246 391060 217274
rect 391768 219406 391888 219434
rect 391768 217274 391796 219406
rect 393148 218074 393176 227122
rect 393608 224262 393636 231676
rect 393976 231662 394266 231690
rect 393596 224256 393648 224262
rect 393596 224198 393648 224204
rect 393976 223038 394004 231662
rect 394332 225888 394384 225894
rect 394332 225830 394384 225836
rect 393964 223032 394016 223038
rect 393964 222974 394016 222980
rect 392676 218068 392728 218074
rect 392676 218010 392728 218016
rect 393136 218068 393188 218074
rect 393136 218010 393188 218016
rect 393504 218068 393556 218074
rect 393504 218010 393556 218016
rect 391768 217246 391842 217274
rect 389330 216988 389358 217110
rect 390158 216988 390186 217246
rect 390986 216988 391014 217246
rect 391814 216988 391842 217246
rect 392688 217138 392716 218010
rect 393516 217138 393544 218010
rect 394344 217274 394372 225830
rect 394516 224256 394568 224262
rect 394516 224198 394568 224204
rect 394528 218074 394556 224198
rect 394896 222902 394924 231676
rect 395172 231662 395554 231690
rect 394884 222896 394936 222902
rect 394884 222838 394936 222844
rect 395172 221610 395200 231662
rect 396184 225758 396212 231676
rect 396368 231662 396842 231690
rect 396172 225752 396224 225758
rect 396172 225694 396224 225700
rect 395804 222896 395856 222902
rect 395804 222838 395856 222844
rect 395160 221604 395212 221610
rect 395160 221546 395212 221552
rect 395816 218074 395844 222838
rect 395988 220108 396040 220114
rect 395988 220050 396040 220056
rect 394516 218068 394568 218074
rect 394516 218010 394568 218016
rect 395160 218068 395212 218074
rect 395160 218010 395212 218016
rect 395804 218068 395856 218074
rect 395804 218010 395856 218016
rect 392642 217110 392716 217138
rect 393470 217110 393544 217138
rect 394298 217246 394372 217274
rect 392642 216988 392670 217110
rect 393470 216988 393498 217110
rect 394298 216988 394326 217246
rect 395172 217138 395200 218010
rect 396000 217274 396028 220050
rect 396368 219434 396396 231662
rect 397472 228546 397500 231676
rect 397840 231662 398130 231690
rect 397460 228540 397512 228546
rect 397460 228482 397512 228488
rect 397840 224398 397868 231662
rect 398104 230376 398156 230382
rect 398104 230318 398156 230324
rect 397828 224392 397880 224398
rect 397828 224334 397880 224340
rect 396816 221468 396868 221474
rect 396816 221410 396868 221416
rect 396276 219406 396396 219434
rect 396276 218754 396304 219406
rect 396264 218748 396316 218754
rect 396264 218690 396316 218696
rect 396828 217274 396856 221410
rect 398116 219026 398144 230318
rect 398760 229634 398788 231676
rect 399404 230382 399432 231676
rect 399392 230376 399444 230382
rect 399392 230318 399444 230324
rect 399852 229764 399904 229770
rect 399852 229706 399904 229712
rect 398748 229628 398800 229634
rect 398748 229570 398800 229576
rect 399864 219434 399892 229706
rect 400048 228410 400076 231676
rect 400232 231662 400706 231690
rect 400968 231662 401350 231690
rect 400232 229094 400260 231662
rect 400232 229066 400352 229094
rect 400036 228404 400088 228410
rect 400036 228346 400088 228352
rect 400128 228132 400180 228138
rect 400128 228074 400180 228080
rect 400140 219434 400168 228074
rect 400324 221746 400352 229066
rect 400312 221740 400364 221746
rect 400312 221682 400364 221688
rect 400680 221604 400732 221610
rect 400680 221546 400732 221552
rect 399300 219428 399352 219434
rect 399864 219406 400076 219434
rect 400140 219428 400272 219434
rect 400140 219406 400220 219428
rect 399300 219370 399352 219376
rect 398104 219020 398156 219026
rect 398104 218962 398156 218968
rect 398472 218612 398524 218618
rect 398472 218554 398524 218560
rect 397644 218068 397696 218074
rect 397644 218010 397696 218016
rect 395126 217110 395200 217138
rect 395954 217246 396028 217274
rect 396782 217246 396856 217274
rect 395126 216988 395154 217110
rect 395954 216988 395982 217246
rect 396782 216988 396810 217246
rect 397656 217138 397684 218010
rect 398484 217138 398512 218554
rect 399312 217138 399340 219370
rect 400048 217274 400076 219406
rect 400220 219370 400272 219376
rect 400692 218074 400720 221546
rect 400968 220250 400996 231662
rect 401980 225622 402008 231676
rect 402624 227322 402652 231676
rect 402796 228404 402848 228410
rect 402796 228346 402848 228352
rect 402612 227316 402664 227322
rect 402612 227258 402664 227264
rect 402244 227180 402296 227186
rect 402244 227122 402296 227128
rect 401968 225616 402020 225622
rect 401968 225558 402020 225564
rect 400956 220244 401008 220250
rect 400956 220186 401008 220192
rect 401784 218204 401836 218210
rect 401784 218146 401836 218152
rect 400680 218068 400732 218074
rect 400680 218010 400732 218016
rect 400956 218068 401008 218074
rect 400956 218010 401008 218016
rect 400048 217246 400122 217274
rect 397610 217110 397684 217138
rect 398438 217110 398512 217138
rect 399266 217110 399340 217138
rect 397610 216988 397638 217110
rect 398438 216988 398466 217110
rect 399266 216988 399294 217110
rect 400094 216988 400122 217246
rect 400968 217138 400996 218010
rect 401796 217138 401824 218146
rect 402256 218074 402284 227122
rect 402612 218884 402664 218890
rect 402612 218826 402664 218832
rect 402244 218068 402296 218074
rect 402244 218010 402296 218016
rect 402624 217138 402652 218826
rect 402808 218210 402836 228346
rect 403268 225894 403296 231676
rect 403544 231662 403926 231690
rect 403544 227050 403572 231662
rect 403532 227044 403584 227050
rect 403532 226986 403584 226992
rect 403992 226500 404044 226506
rect 403992 226442 404044 226448
rect 403256 225888 403308 225894
rect 403256 225830 403308 225836
rect 402796 218204 402848 218210
rect 402796 218146 402848 218152
rect 404004 218074 404032 226442
rect 404176 225004 404228 225010
rect 404176 224946 404228 224952
rect 403440 218068 403492 218074
rect 403440 218010 403492 218016
rect 403992 218068 404044 218074
rect 403992 218010 404044 218016
rect 403452 217138 403480 218010
rect 404188 217274 404216 224946
rect 404556 224262 404584 231676
rect 404832 231662 405214 231690
rect 404544 224256 404596 224262
rect 404544 224198 404596 224204
rect 404832 220114 404860 231662
rect 405556 224256 405608 224262
rect 405556 224198 405608 224204
rect 404820 220108 404872 220114
rect 404820 220050 404872 220056
rect 405568 218074 405596 224198
rect 405844 221610 405872 231676
rect 406488 222902 406516 231676
rect 407146 231662 407344 231690
rect 406752 223576 406804 223582
rect 406752 223518 406804 223524
rect 406476 222896 406528 222902
rect 406476 222838 406528 222844
rect 405832 221604 405884 221610
rect 405832 221546 405884 221552
rect 405924 219496 405976 219502
rect 405924 219438 405976 219444
rect 405096 218068 405148 218074
rect 405096 218010 405148 218016
rect 405556 218068 405608 218074
rect 405556 218010 405608 218016
rect 404188 217246 404262 217274
rect 400922 217110 400996 217138
rect 401750 217110 401824 217138
rect 402578 217110 402652 217138
rect 403406 217110 403480 217138
rect 400922 216988 400950 217110
rect 401750 216988 401778 217110
rect 402578 216988 402606 217110
rect 403406 216988 403434 217110
rect 404234 216988 404262 217246
rect 405108 217138 405136 218010
rect 405936 217274 405964 219438
rect 406764 217274 406792 223518
rect 407316 221474 407344 231662
rect 407776 228546 407804 231676
rect 407764 228540 407816 228546
rect 407764 228482 407816 228488
rect 408420 227186 408448 231676
rect 408696 231662 409078 231690
rect 408408 227180 408460 227186
rect 408408 227122 408460 227128
rect 408696 226370 408724 231662
rect 409708 229770 409736 231676
rect 409696 229764 409748 229770
rect 409696 229706 409748 229712
rect 409788 228540 409840 228546
rect 409788 228482 409840 228488
rect 409052 227792 409104 227798
rect 409052 227734 409104 227740
rect 407764 226364 407816 226370
rect 407764 226306 407816 226312
rect 408684 226364 408736 226370
rect 408684 226306 408736 226312
rect 407304 221468 407356 221474
rect 407304 221410 407356 221416
rect 407776 218618 407804 226306
rect 408408 221468 408460 221474
rect 408408 221410 408460 221416
rect 407764 218612 407816 218618
rect 407764 218554 407816 218560
rect 407580 218204 407632 218210
rect 407580 218146 407632 218152
rect 405062 217110 405136 217138
rect 405890 217246 405964 217274
rect 406718 217246 406792 217274
rect 405062 216988 405090 217110
rect 405890 216988 405918 217246
rect 406718 216988 406746 217246
rect 407592 217138 407620 218146
rect 408420 217274 408448 221410
rect 409064 218890 409092 227734
rect 409052 218884 409104 218890
rect 409052 218826 409104 218832
rect 409800 218074 409828 228482
rect 410352 227798 410380 231676
rect 410720 231662 411010 231690
rect 410720 229094 410748 231662
rect 410892 229900 410944 229906
rect 410892 229842 410944 229848
rect 410904 229094 410932 229842
rect 410628 229066 410748 229094
rect 410812 229066 410932 229094
rect 410340 227792 410392 227798
rect 410340 227734 410392 227740
rect 410628 225010 410656 229066
rect 410616 225004 410668 225010
rect 410616 224946 410668 224952
rect 410812 219434 410840 229066
rect 411640 228410 411668 231676
rect 411628 228404 411680 228410
rect 411628 228346 411680 228352
rect 411904 227792 411956 227798
rect 411904 227734 411956 227740
rect 410984 225616 411036 225622
rect 410984 225558 411036 225564
rect 410996 219434 411024 225558
rect 410720 219406 410840 219434
rect 410904 219406 411024 219434
rect 410720 218074 410748 219406
rect 409236 218068 409288 218074
rect 409236 218010 409288 218016
rect 409788 218068 409840 218074
rect 409788 218010 409840 218016
rect 410064 218068 410116 218074
rect 410064 218010 410116 218016
rect 410708 218068 410760 218074
rect 410708 218010 410760 218016
rect 407546 217110 407620 217138
rect 408374 217246 408448 217274
rect 407546 216988 407574 217110
rect 408374 216988 408402 217246
rect 409248 217138 409276 218010
rect 410076 217138 410104 218010
rect 410904 217274 410932 219406
rect 411720 218884 411772 218890
rect 411720 218826 411772 218832
rect 409202 217110 409276 217138
rect 410030 217110 410104 217138
rect 410858 217246 410932 217274
rect 409202 216988 409230 217110
rect 410030 216988 410058 217110
rect 410858 216988 410886 217246
rect 411732 217138 411760 218826
rect 411916 218210 411944 227734
rect 412284 226506 412312 231676
rect 412744 231662 412942 231690
rect 412548 227044 412600 227050
rect 412548 226986 412600 226992
rect 412272 226500 412324 226506
rect 412272 226442 412324 226448
rect 412560 218890 412588 226986
rect 412744 219502 412772 231662
rect 413572 227798 413600 231676
rect 413836 229356 413888 229362
rect 413836 229298 413888 229304
rect 413560 227792 413612 227798
rect 413560 227734 413612 227740
rect 412732 219496 412784 219502
rect 412732 219438 412784 219444
rect 412548 218884 412600 218890
rect 412548 218826 412600 218832
rect 412548 218748 412600 218754
rect 412548 218690 412600 218696
rect 411904 218204 411956 218210
rect 411904 218146 411956 218152
rect 412560 217138 412588 218690
rect 413848 218074 413876 229298
rect 414216 224262 414244 231676
rect 414204 224256 414256 224262
rect 414204 224198 414256 224204
rect 414860 223582 414888 231676
rect 415504 228546 415532 231676
rect 415492 228540 415544 228546
rect 415492 228482 415544 228488
rect 415032 228064 415084 228070
rect 415032 228006 415084 228012
rect 414848 223576 414900 223582
rect 414848 223518 414900 223524
rect 414204 220788 414256 220794
rect 414204 220730 414256 220736
rect 413376 218068 413428 218074
rect 413376 218010 413428 218016
rect 413836 218068 413888 218074
rect 413836 218010 413888 218016
rect 413388 217138 413416 218010
rect 414216 217274 414244 220730
rect 415044 217274 415072 228006
rect 416148 225622 416176 231676
rect 416792 229094 416820 231676
rect 417436 229906 417464 231676
rect 417712 231662 418094 231690
rect 418356 231662 418738 231690
rect 417424 229900 417476 229906
rect 417424 229842 417476 229848
rect 417712 229094 417740 231662
rect 416792 229066 416912 229094
rect 416688 227928 416740 227934
rect 416688 227870 416740 227876
rect 416136 225616 416188 225622
rect 416136 225558 416188 225564
rect 416504 225004 416556 225010
rect 416504 224946 416556 224952
rect 416516 219434 416544 224946
rect 416700 219434 416728 227870
rect 416884 221474 416912 229066
rect 417160 229066 417740 229094
rect 416872 221468 416924 221474
rect 416872 221410 416924 221416
rect 415860 219428 415912 219434
rect 416516 219406 416636 219434
rect 416700 219428 416832 219434
rect 416700 219406 416780 219428
rect 415860 219370 415912 219376
rect 411686 217110 411760 217138
rect 412514 217110 412588 217138
rect 413342 217110 413416 217138
rect 414170 217246 414244 217274
rect 414998 217246 415072 217274
rect 411686 216988 411714 217110
rect 412514 216988 412542 217110
rect 413342 216988 413370 217110
rect 414170 216988 414198 217246
rect 414998 216988 415026 217246
rect 415872 217138 415900 219370
rect 416608 217274 416636 219406
rect 416780 219370 416832 219376
rect 417160 218754 417188 229066
rect 418356 224954 418384 231662
rect 419368 227050 419396 231676
rect 420012 229362 420040 231676
rect 420000 229356 420052 229362
rect 420000 229298 420052 229304
rect 420656 227934 420684 231676
rect 421024 231662 421314 231690
rect 420644 227928 420696 227934
rect 420644 227870 420696 227876
rect 420644 227792 420696 227798
rect 420644 227734 420696 227740
rect 419356 227044 419408 227050
rect 419356 226986 419408 226992
rect 418172 224926 418384 224954
rect 418172 220794 418200 224926
rect 418344 220856 418396 220862
rect 418344 220798 418396 220804
rect 418160 220788 418212 220794
rect 418160 220730 418212 220736
rect 417516 219428 417568 219434
rect 417516 219370 417568 219376
rect 417148 218748 417200 218754
rect 417148 218690 417200 218696
rect 416608 217246 416682 217274
rect 415826 217110 415900 217138
rect 415826 216988 415854 217110
rect 416654 216988 416682 217246
rect 417528 217138 417556 219370
rect 418356 217274 418384 220798
rect 420656 219434 420684 227734
rect 420828 222896 420880 222902
rect 420828 222838 420880 222844
rect 420656 219406 420776 219434
rect 419172 219292 419224 219298
rect 419172 219234 419224 219240
rect 419184 217274 419212 219234
rect 420000 218068 420052 218074
rect 420000 218010 420052 218016
rect 417482 217110 417556 217138
rect 418310 217246 418384 217274
rect 419138 217246 419212 217274
rect 417482 216988 417510 217110
rect 418310 216988 418338 217246
rect 419138 216988 419166 217246
rect 420012 217138 420040 218010
rect 420748 217274 420776 219406
rect 420840 218090 420868 222838
rect 421024 219502 421052 231662
rect 421944 228070 421972 231676
rect 422312 231662 422602 231690
rect 422864 231662 423246 231690
rect 422312 229094 422340 231662
rect 422220 229066 422340 229094
rect 421932 228064 421984 228070
rect 421932 228006 421984 228012
rect 422220 225010 422248 229066
rect 422208 225004 422260 225010
rect 422208 224946 422260 224952
rect 421656 220108 421708 220114
rect 421656 220050 421708 220056
rect 421012 219496 421064 219502
rect 421012 219438 421064 219444
rect 420840 218074 420960 218090
rect 420840 218068 420972 218074
rect 420840 218062 420920 218068
rect 420920 218010 420972 218016
rect 421668 217274 421696 220050
rect 422864 219434 422892 231662
rect 423496 229152 423548 229158
rect 423496 229094 423548 229100
rect 423508 219434 423536 229094
rect 423876 227798 423904 231676
rect 424060 231662 424534 231690
rect 423864 227792 423916 227798
rect 423864 227734 423916 227740
rect 424060 220862 424088 231662
rect 425164 222902 425192 231676
rect 425440 231662 425822 231690
rect 425152 222896 425204 222902
rect 425152 222838 425204 222844
rect 424968 221944 425020 221950
rect 424968 221886 425020 221892
rect 424048 220856 424100 220862
rect 424048 220798 424100 220804
rect 422680 219406 422892 219434
rect 423324 219406 423536 219434
rect 422680 219298 422708 219406
rect 422668 219292 422720 219298
rect 422668 219234 422720 219240
rect 422484 218204 422536 218210
rect 422484 218146 422536 218152
rect 420748 217246 420822 217274
rect 419966 217110 420040 217138
rect 419966 216988 419994 217110
rect 420794 216988 420822 217246
rect 421622 217246 421696 217274
rect 421622 216988 421650 217246
rect 422496 217138 422524 218146
rect 423324 217274 423352 219406
rect 424140 218068 424192 218074
rect 424140 218010 424192 218016
rect 422450 217110 422524 217138
rect 423278 217246 423352 217274
rect 422450 216988 422478 217110
rect 423278 216988 423306 217246
rect 424152 217138 424180 218010
rect 424980 217274 425008 221886
rect 425440 218210 425468 231662
rect 426452 222562 426480 231676
rect 426728 231662 427110 231690
rect 426440 222556 426492 222562
rect 426440 222498 426492 222504
rect 426728 220114 426756 231662
rect 427740 229158 427768 231676
rect 427924 231662 428398 231690
rect 428752 231662 429042 231690
rect 429212 231662 429686 231690
rect 429856 231662 430330 231690
rect 430684 231662 430974 231690
rect 431236 231662 431618 231690
rect 432064 231662 432262 231690
rect 432708 231662 432906 231690
rect 433550 231662 433748 231690
rect 427728 229152 427780 229158
rect 427728 229094 427780 229100
rect 426992 222556 427044 222562
rect 426992 222498 427044 222504
rect 426716 220108 426768 220114
rect 426716 220050 426768 220056
rect 426624 218340 426676 218346
rect 426624 218282 426676 218288
rect 425428 218204 425480 218210
rect 425428 218146 425480 218152
rect 425796 218204 425848 218210
rect 425796 218146 425848 218152
rect 424106 217110 424180 217138
rect 424934 217246 425008 217274
rect 424106 216988 424134 217110
rect 424934 216988 424962 217246
rect 425808 217138 425836 218146
rect 426636 217138 426664 218282
rect 427004 218074 427032 222498
rect 427924 218210 427952 231662
rect 428752 219434 428780 231662
rect 429212 221950 429240 231662
rect 429200 221944 429252 221950
rect 429200 221886 429252 221892
rect 429856 219434 429884 231662
rect 430684 219434 430712 231662
rect 431236 219434 431264 231662
rect 432064 219570 432092 231662
rect 432236 220516 432288 220522
rect 432236 220458 432288 220464
rect 432052 219564 432104 219570
rect 432052 219506 432104 219512
rect 432248 219434 432276 220458
rect 428280 219428 428332 219434
rect 428280 219370 428332 219376
rect 428476 219406 428780 219434
rect 429396 219406 429884 219434
rect 430592 219406 430712 219434
rect 430776 219406 431264 219434
rect 431972 219406 432276 219434
rect 427912 218204 427964 218210
rect 427912 218146 427964 218152
rect 426992 218068 427044 218074
rect 426992 218010 427044 218016
rect 427452 218068 427504 218074
rect 427452 218010 427504 218016
rect 427464 217138 427492 218010
rect 428292 217138 428320 219370
rect 428476 218074 428504 219406
rect 429396 218346 429424 219406
rect 429936 218748 429988 218754
rect 429936 218690 429988 218696
rect 429384 218340 429436 218346
rect 429384 218282 429436 218288
rect 428464 218068 428516 218074
rect 428464 218010 428516 218016
rect 429108 218068 429160 218074
rect 429108 218010 429160 218016
rect 429120 217138 429148 218010
rect 429948 217138 429976 218690
rect 430592 218074 430620 219406
rect 430580 218068 430632 218074
rect 430580 218010 430632 218016
rect 430776 217274 430804 219406
rect 431972 218090 432000 219406
rect 432708 218754 432736 231662
rect 433524 229832 433576 229838
rect 433524 229774 433576 229780
rect 433536 229094 433564 229774
rect 433720 229094 433748 231662
rect 434180 229838 434208 231676
rect 434168 229832 434220 229838
rect 434168 229774 434220 229780
rect 433536 229066 433656 229094
rect 433720 229066 433840 229094
rect 432696 218748 432748 218754
rect 432696 218690 432748 218696
rect 433248 218204 433300 218210
rect 433248 218146 433300 218152
rect 425762 217110 425836 217138
rect 426590 217110 426664 217138
rect 427418 217110 427492 217138
rect 428246 217110 428320 217138
rect 429074 217110 429148 217138
rect 429902 217110 429976 217138
rect 430730 217246 430804 217274
rect 431604 218062 432000 218090
rect 432420 218068 432472 218074
rect 425762 216988 425790 217110
rect 426590 216988 426618 217110
rect 427418 216988 427446 217110
rect 428246 216988 428274 217110
rect 429074 216988 429102 217110
rect 429902 216988 429930 217110
rect 430730 216988 430758 217246
rect 431604 217138 431632 218062
rect 432420 218010 432472 218016
rect 432432 217138 432460 218010
rect 433260 217138 433288 218146
rect 433628 217274 433656 229066
rect 433812 218074 433840 229066
rect 434824 220522 434852 231676
rect 435192 231662 435482 231690
rect 436126 231662 436324 231690
rect 434812 220516 434864 220522
rect 434812 220458 434864 220464
rect 435192 219434 435220 231662
rect 434732 219406 435220 219434
rect 434732 218210 434760 219406
rect 434720 218204 434772 218210
rect 434720 218146 434772 218152
rect 434904 218204 434956 218210
rect 434904 218146 434956 218152
rect 433800 218068 433852 218074
rect 433800 218010 433852 218016
rect 433628 217246 434070 217274
rect 431558 217110 431632 217138
rect 432386 217110 432460 217138
rect 433214 217110 433288 217138
rect 431558 216988 431586 217110
rect 432386 216988 432414 217110
rect 433214 216988 433242 217110
rect 434042 216988 434070 217246
rect 434916 217138 434944 218146
rect 436296 218074 436324 231662
rect 436572 231662 436770 231690
rect 437032 231662 437414 231690
rect 437768 231662 438058 231690
rect 436572 229094 436600 231662
rect 436572 229066 436692 229094
rect 435732 218068 435784 218074
rect 435732 218010 435784 218016
rect 436284 218068 436336 218074
rect 436284 218010 436336 218016
rect 436468 218068 436520 218074
rect 436468 218010 436520 218016
rect 435744 217138 435772 218010
rect 434870 217110 434944 217138
rect 435698 217110 435772 217138
rect 436480 217138 436508 218010
rect 436664 217546 436692 229066
rect 437032 219434 437060 231662
rect 436848 219406 437060 219434
rect 436848 218210 436876 219406
rect 436836 218204 436888 218210
rect 436836 218146 436888 218152
rect 437768 218074 437796 231662
rect 438688 230382 438716 231676
rect 439332 230586 439360 231676
rect 439516 231662 439990 231690
rect 440344 231662 440634 231690
rect 439320 230580 439372 230586
rect 439320 230522 439372 230528
rect 439516 230466 439544 231662
rect 438964 230438 439544 230466
rect 438676 230376 438728 230382
rect 438676 230318 438728 230324
rect 438964 224954 438992 230438
rect 439320 230376 439372 230382
rect 439320 230318 439372 230324
rect 439332 224954 439360 230318
rect 438872 224926 438992 224954
rect 439056 224926 439360 224954
rect 438872 219434 438900 224926
rect 438216 219428 438268 219434
rect 438216 219370 438268 219376
rect 438860 219428 438912 219434
rect 438860 219370 438912 219376
rect 437756 218068 437808 218074
rect 437756 218010 437808 218016
rect 436664 217518 437336 217546
rect 437308 217274 437336 217518
rect 437308 217246 437382 217274
rect 436480 217110 436554 217138
rect 434870 216988 434898 217110
rect 435698 216988 435726 217110
rect 436526 216988 436554 217110
rect 437354 216988 437382 217246
rect 438228 217138 438256 219370
rect 439056 217274 439084 224926
rect 440344 219434 440372 231662
rect 440700 230444 440752 230450
rect 440700 230386 440752 230392
rect 439872 219428 439924 219434
rect 439872 219370 439924 219376
rect 440332 219428 440384 219434
rect 440332 219370 440384 219376
rect 438182 217110 438256 217138
rect 439010 217246 439084 217274
rect 438182 216988 438210 217110
rect 439010 216988 439038 217246
rect 439884 217138 439912 219370
rect 440712 217274 440740 230386
rect 441264 229158 441292 231676
rect 441908 230450 441936 231676
rect 442092 231662 442566 231690
rect 443104 231662 443210 231690
rect 441896 230444 441948 230450
rect 441896 230386 441948 230392
rect 442092 230330 442120 231662
rect 441724 230302 442120 230330
rect 441252 229152 441304 229158
rect 441252 229094 441304 229100
rect 441724 224954 441752 230302
rect 442080 229152 442132 229158
rect 442080 229094 442132 229100
rect 442092 229066 442304 229094
rect 441632 224926 441752 224954
rect 441632 218090 441660 224926
rect 441540 218062 441660 218090
rect 441540 217274 441568 218062
rect 439838 217110 439912 217138
rect 440666 217246 440740 217274
rect 441494 217246 441568 217274
rect 442276 217274 442304 229066
rect 443104 217274 443132 231662
rect 443460 230444 443512 230450
rect 443460 230386 443512 230392
rect 443472 229094 443500 230386
rect 443840 230246 443868 231676
rect 444484 230450 444512 231676
rect 444668 231662 445142 231690
rect 444472 230444 444524 230450
rect 444472 230386 444524 230392
rect 444668 230330 444696 231662
rect 444484 230302 444696 230330
rect 443828 230240 443880 230246
rect 443828 230182 443880 230188
rect 443472 229066 443960 229094
rect 443932 217274 443960 229066
rect 444484 224954 444512 230302
rect 444656 230240 444708 230246
rect 444656 230182 444708 230188
rect 444668 224954 444696 230182
rect 445772 229094 445800 231676
rect 446416 229430 446444 231676
rect 446404 229424 446456 229430
rect 446404 229366 446456 229372
rect 445772 229066 446444 229094
rect 444484 224926 444604 224954
rect 444668 224926 445616 224954
rect 444576 217274 444604 224926
rect 445588 217274 445616 224926
rect 446416 217274 446444 229066
rect 447060 227934 447088 231676
rect 447244 231662 447718 231690
rect 447048 227928 447100 227934
rect 447048 227870 447100 227876
rect 447244 219434 447272 231662
rect 447600 230444 447652 230450
rect 447600 230386 447652 230392
rect 447612 219434 447640 230386
rect 448348 229094 448376 231676
rect 448992 229566 449020 231676
rect 449636 229906 449664 231676
rect 449624 229900 449676 229906
rect 449624 229842 449676 229848
rect 448980 229560 449032 229566
rect 448980 229502 449032 229508
rect 448980 229424 449032 229430
rect 448980 229366 449032 229372
rect 448348 229066 448652 229094
rect 447152 219406 447272 219434
rect 447336 219406 447640 219434
rect 442276 217246 442350 217274
rect 443104 217246 443178 217274
rect 443932 217246 444006 217274
rect 444576 217246 444834 217274
rect 445588 217246 445662 217274
rect 446416 217246 446490 217274
rect 447152 217258 447180 219406
rect 447336 217274 447364 219406
rect 439838 216988 439866 217110
rect 440666 216988 440694 217246
rect 441494 216988 441522 217246
rect 442322 216988 442350 217246
rect 443150 216988 443178 217246
rect 443978 216988 444006 217246
rect 444806 216988 444834 217246
rect 445634 216988 445662 217246
rect 446462 216988 446490 217246
rect 447140 217252 447192 217258
rect 447140 217194 447192 217200
rect 447290 217246 447364 217274
rect 448624 217258 448652 229066
rect 448992 217274 449020 229366
rect 450280 229294 450308 231676
rect 450544 229900 450596 229906
rect 450544 229842 450596 229848
rect 450268 229288 450320 229294
rect 450268 229230 450320 229236
rect 450556 229094 450584 229842
rect 450924 229430 450952 231676
rect 451568 230450 451596 231676
rect 452226 231662 452516 231690
rect 451556 230444 451608 230450
rect 451556 230386 451608 230392
rect 451372 229560 451424 229566
rect 451372 229502 451424 229508
rect 450912 229424 450964 229430
rect 450912 229366 450964 229372
rect 450556 229066 450768 229094
rect 450544 227928 450596 227934
rect 450544 227870 450596 227876
rect 448106 217252 448158 217258
rect 447290 216988 447318 217246
rect 448106 217194 448158 217200
rect 448612 217252 448664 217258
rect 448612 217194 448664 217200
rect 448946 217246 449020 217274
rect 450556 217274 450584 227870
rect 450740 218346 450768 229066
rect 450728 218340 450780 218346
rect 450728 218282 450780 218288
rect 451384 217870 451412 229502
rect 451740 229288 451792 229294
rect 451740 229230 451792 229236
rect 451752 219434 451780 229230
rect 452488 222154 452516 231662
rect 452856 230246 452884 231676
rect 453304 230444 453356 230450
rect 453304 230386 453356 230392
rect 452844 230240 452896 230246
rect 452844 230182 452896 230188
rect 452660 229424 452712 229430
rect 452660 229366 452712 229372
rect 452672 229094 452700 229366
rect 452672 229066 453068 229094
rect 452476 222148 452528 222154
rect 452476 222090 452528 222096
rect 451568 219406 451780 219434
rect 451372 217864 451424 217870
rect 451372 217806 451424 217812
rect 451568 217274 451596 219406
rect 452200 217864 452252 217870
rect 452200 217806 452252 217812
rect 449762 217252 449814 217258
rect 448118 216988 448146 217194
rect 448946 216988 448974 217246
rect 450556 217246 450630 217274
rect 449762 217194 449814 217200
rect 449774 216988 449802 217194
rect 450602 216988 450630 217246
rect 451430 217246 451596 217274
rect 451430 216988 451458 217246
rect 452212 217138 452240 217806
rect 453040 217274 453068 229066
rect 453316 218074 453344 230386
rect 453500 229974 453528 231676
rect 454144 230110 454172 231676
rect 454316 230240 454368 230246
rect 454316 230182 454368 230188
rect 454132 230104 454184 230110
rect 454132 230046 454184 230052
rect 453488 229968 453540 229974
rect 453488 229910 453540 229916
rect 454328 229094 454356 230182
rect 454788 229094 454816 231676
rect 455432 230382 455460 231676
rect 455420 230376 455472 230382
rect 455420 230318 455472 230324
rect 455328 230104 455380 230110
rect 455328 230046 455380 230052
rect 454328 229066 454724 229094
rect 454788 229066 454908 229094
rect 453856 218340 453908 218346
rect 453856 218282 453908 218288
rect 453304 218068 453356 218074
rect 453304 218010 453356 218016
rect 453040 217246 453114 217274
rect 452212 217110 452286 217138
rect 452258 216988 452286 217110
rect 453086 216988 453114 217246
rect 453868 217138 453896 218282
rect 454696 217274 454724 229066
rect 454880 223582 454908 229066
rect 454868 223576 454920 223582
rect 454868 223518 454920 223524
rect 455340 220794 455368 230046
rect 455788 229968 455840 229974
rect 455788 229910 455840 229916
rect 455604 222148 455656 222154
rect 455604 222090 455656 222096
rect 455328 220788 455380 220794
rect 455328 220730 455380 220736
rect 455616 218074 455644 222090
rect 455800 219434 455828 229910
rect 456076 224534 456104 231676
rect 456064 224528 456116 224534
rect 456064 224470 456116 224476
rect 456720 220930 456748 231676
rect 457168 230376 457220 230382
rect 457168 230318 457220 230324
rect 456708 220924 456760 220930
rect 456708 220866 456760 220872
rect 457180 219434 457208 230318
rect 457364 229906 457392 231676
rect 457352 229900 457404 229906
rect 457352 229842 457404 229848
rect 458008 229094 458036 231676
rect 458008 229066 458128 229094
rect 455800 219406 456380 219434
rect 457180 219406 458036 219434
rect 455420 218068 455472 218074
rect 455420 218010 455472 218016
rect 455604 218068 455656 218074
rect 455604 218010 455656 218016
rect 455432 217274 455460 218010
rect 456352 217274 456380 219406
rect 457168 218068 457220 218074
rect 457168 218010 457220 218016
rect 454696 217246 454770 217274
rect 455432 217246 455598 217274
rect 456352 217246 456426 217274
rect 453868 217110 453942 217138
rect 453914 216988 453942 217110
rect 454742 216988 454770 217246
rect 455570 216988 455598 217246
rect 456398 216988 456426 217246
rect 457180 217138 457208 218010
rect 458008 217274 458036 219406
rect 458100 218498 458128 229066
rect 458652 226302 458680 231676
rect 459310 231662 459508 231690
rect 458640 226296 458692 226302
rect 458640 226238 458692 226244
rect 458824 220788 458876 220794
rect 458824 220730 458876 220736
rect 458100 218470 458220 218498
rect 458192 218414 458220 218470
rect 458180 218408 458232 218414
rect 458180 218350 458232 218356
rect 458836 217274 458864 220730
rect 459480 220250 459508 231662
rect 459744 224528 459796 224534
rect 459744 224470 459796 224476
rect 459468 220244 459520 220250
rect 459468 220186 459520 220192
rect 459756 217274 459784 224470
rect 459940 222902 459968 231676
rect 460584 223718 460612 231676
rect 461242 231662 461716 231690
rect 461886 231662 462176 231690
rect 461688 229094 461716 231662
rect 461688 229066 461992 229094
rect 460572 223712 460624 223718
rect 460572 223654 460624 223660
rect 460480 223576 460532 223582
rect 460480 223518 460532 223524
rect 459928 222896 459980 222902
rect 459928 222838 459980 222844
rect 458008 217246 458082 217274
rect 458836 217246 458910 217274
rect 457180 217110 457254 217138
rect 457226 216988 457254 217110
rect 458054 216988 458082 217246
rect 458882 216988 458910 217246
rect 459710 217246 459784 217274
rect 460492 217274 460520 223518
rect 461308 218340 461360 218346
rect 461308 218282 461360 218288
rect 460492 217246 460566 217274
rect 459710 216988 459738 217246
rect 460538 216988 460566 217246
rect 461320 217138 461348 218282
rect 461964 218210 461992 229066
rect 462148 222154 462176 231662
rect 462516 224806 462544 231676
rect 462964 226296 463016 226302
rect 462964 226238 463016 226244
rect 462504 224800 462556 224806
rect 462504 224742 462556 224748
rect 462136 222148 462188 222154
rect 462136 222090 462188 222096
rect 462136 220856 462188 220862
rect 462136 220798 462188 220804
rect 461952 218204 462004 218210
rect 461952 218146 462004 218152
rect 462148 217274 462176 220798
rect 462976 217274 463004 226238
rect 463160 225418 463188 231676
rect 463804 229634 463832 231676
rect 464462 231662 465028 231690
rect 465106 231662 465488 231690
rect 465750 231662 465948 231690
rect 464068 229900 464120 229906
rect 464068 229842 464120 229848
rect 463792 229628 463844 229634
rect 463792 229570 463844 229576
rect 463148 225412 463200 225418
rect 463148 225354 463200 225360
rect 463148 223712 463200 223718
rect 463148 223654 463200 223660
rect 463160 218074 463188 223654
rect 464080 219434 464108 229842
rect 465000 219638 465028 231662
rect 465460 229498 465488 231662
rect 465724 229628 465776 229634
rect 465724 229570 465776 229576
rect 465448 229492 465500 229498
rect 465448 229434 465500 229440
rect 465736 220726 465764 229570
rect 465920 227662 465948 231662
rect 466104 231662 466394 231690
rect 465908 227656 465960 227662
rect 465908 227598 465960 227604
rect 466104 220862 466132 231662
rect 467024 229770 467052 231676
rect 467012 229764 467064 229770
rect 467012 229706 467064 229712
rect 467472 229492 467524 229498
rect 467472 229434 467524 229440
rect 467288 225412 467340 225418
rect 467288 225354 467340 225360
rect 467104 222896 467156 222902
rect 467104 222838 467156 222844
rect 466092 220856 466144 220862
rect 466092 220798 466144 220804
rect 465724 220720 465776 220726
rect 465724 220662 465776 220668
rect 465448 220244 465500 220250
rect 465448 220186 465500 220192
rect 464988 219632 465040 219638
rect 464988 219574 465040 219580
rect 463896 219406 464108 219434
rect 463148 218068 463200 218074
rect 463148 218010 463200 218016
rect 463896 217274 463924 219406
rect 464620 218068 464672 218074
rect 464620 218010 464672 218016
rect 462148 217246 462222 217274
rect 462976 217246 463050 217274
rect 461320 217110 461394 217138
rect 461366 216988 461394 217110
rect 462194 216988 462222 217246
rect 463022 216988 463050 217246
rect 463850 217246 463924 217274
rect 463850 216988 463878 217246
rect 464632 217138 464660 218010
rect 465460 217274 465488 220186
rect 466276 218204 466328 218210
rect 466276 218146 466328 218152
rect 465460 217246 465534 217274
rect 464632 217110 464706 217138
rect 464678 216988 464706 217110
rect 465506 216988 465534 217246
rect 466288 217138 466316 218146
rect 467116 217274 467144 222838
rect 467300 218074 467328 225354
rect 467484 222902 467512 229434
rect 467668 225622 467696 231676
rect 468312 230246 468340 231676
rect 468300 230240 468352 230246
rect 468300 230182 468352 230188
rect 467656 225616 467708 225622
rect 467656 225558 467708 225564
rect 467472 222896 467524 222902
rect 467472 222838 467524 222844
rect 468760 222148 468812 222154
rect 468760 222090 468812 222096
rect 467288 218068 467340 218074
rect 467288 218010 467340 218016
rect 467932 218068 467984 218074
rect 467932 218010 467984 218016
rect 467116 217246 467190 217274
rect 466288 217110 466362 217138
rect 466334 216988 466362 217110
rect 467162 216988 467190 217246
rect 467944 217138 467972 218010
rect 468772 217274 468800 222090
rect 468956 221474 468984 231676
rect 469128 230240 469180 230246
rect 469128 230182 469180 230188
rect 468944 221468 468996 221474
rect 468944 221410 468996 221416
rect 469140 220522 469168 230182
rect 469600 229906 469628 231676
rect 469588 229900 469640 229906
rect 469588 229842 469640 229848
rect 469864 227656 469916 227662
rect 469864 227598 469916 227604
rect 469312 224800 469364 224806
rect 469312 224742 469364 224748
rect 469128 220516 469180 220522
rect 469128 220458 469180 220464
rect 468772 217246 468846 217274
rect 469324 217258 469352 224742
rect 469588 220720 469640 220726
rect 469588 220662 469640 220668
rect 469600 217274 469628 220662
rect 469876 218618 469904 227598
rect 470244 224262 470272 231676
rect 470888 230382 470916 231676
rect 470876 230376 470928 230382
rect 470876 230318 470928 230324
rect 471532 227798 471560 231676
rect 471888 230376 471940 230382
rect 471888 230318 471940 230324
rect 471520 227792 471572 227798
rect 471520 227734 471572 227740
rect 470232 224256 470284 224262
rect 470232 224198 470284 224204
rect 471900 222154 471928 230318
rect 472176 229362 472204 231676
rect 472834 231662 473216 231690
rect 472164 229356 472216 229362
rect 472164 229298 472216 229304
rect 472992 229356 473044 229362
rect 472992 229298 473044 229304
rect 471888 222148 471940 222154
rect 471888 222090 471940 222096
rect 471428 220856 471480 220862
rect 471428 220798 471480 220804
rect 469864 218612 469916 218618
rect 469864 218554 469916 218560
rect 471244 218612 471296 218618
rect 471244 218554 471296 218560
rect 467944 217110 468018 217138
rect 467990 216988 468018 217110
rect 468818 216988 468846 217246
rect 469312 217252 469364 217258
rect 469600 217246 469674 217274
rect 469312 217194 469364 217200
rect 469646 216988 469674 217246
rect 470462 217252 470514 217258
rect 470462 217194 470514 217200
rect 470474 216988 470502 217194
rect 471256 217138 471284 218554
rect 471440 218074 471468 220798
rect 473004 220386 473032 229298
rect 472992 220380 473044 220386
rect 472992 220322 473044 220328
rect 473188 220250 473216 231662
rect 473464 223582 473492 231676
rect 474122 231662 474504 231690
rect 474004 229764 474056 229770
rect 474004 229706 474056 229712
rect 473452 223576 473504 223582
rect 473452 223518 473504 223524
rect 473728 222896 473780 222902
rect 473728 222838 473780 222844
rect 473176 220244 473228 220250
rect 473176 220186 473228 220192
rect 472072 219632 472124 219638
rect 472072 219574 472124 219580
rect 471428 218068 471480 218074
rect 471428 218010 471480 218016
rect 472084 217274 472112 219574
rect 472900 218068 472952 218074
rect 472900 218010 472952 218016
rect 472084 217246 472158 217274
rect 471256 217110 471330 217138
rect 471302 216988 471330 217110
rect 472130 216988 472158 217246
rect 472912 217138 472940 218010
rect 473740 217274 473768 222838
rect 474016 220794 474044 229706
rect 474476 228410 474504 231662
rect 474464 228404 474516 228410
rect 474464 228346 474516 228352
rect 474752 226506 474780 231676
rect 475410 231662 475976 231690
rect 474740 226500 474792 226506
rect 474740 226442 474792 226448
rect 475568 223576 475620 223582
rect 475568 223518 475620 223524
rect 474004 220788 474056 220794
rect 474004 220730 474056 220736
rect 475384 220788 475436 220794
rect 475384 220730 475436 220736
rect 474556 220516 474608 220522
rect 474556 220458 474608 220464
rect 474568 217274 474596 220458
rect 475396 217274 475424 220730
rect 475580 218618 475608 223518
rect 475948 221746 475976 231662
rect 476040 230466 476068 231676
rect 476040 230450 476160 230466
rect 476040 230444 476172 230450
rect 476040 230438 476120 230444
rect 476120 230386 476172 230392
rect 476684 230042 476712 231676
rect 476672 230036 476724 230042
rect 476672 229978 476724 229984
rect 476764 229900 476816 229906
rect 476764 229842 476816 229848
rect 476580 225616 476632 225622
rect 476580 225558 476632 225564
rect 475936 221740 475988 221746
rect 475936 221682 475988 221688
rect 476212 221468 476264 221474
rect 476212 221410 476264 221416
rect 475568 218612 475620 218618
rect 475568 218554 475620 218560
rect 476224 217274 476252 221410
rect 476592 217274 476620 225558
rect 476776 220794 476804 229842
rect 477328 225622 477356 231676
rect 477986 231662 478368 231690
rect 478630 231662 478828 231690
rect 477316 225616 477368 225622
rect 477316 225558 477368 225564
rect 477868 222148 477920 222154
rect 477868 222090 477920 222096
rect 476764 220788 476816 220794
rect 476764 220730 476816 220736
rect 477880 217274 477908 222090
rect 478340 220114 478368 231662
rect 478604 230444 478656 230450
rect 478604 230386 478656 230392
rect 478616 227186 478644 230386
rect 478800 229094 478828 231662
rect 479260 229770 479288 231676
rect 479248 229764 479300 229770
rect 479248 229706 479300 229712
rect 478800 229066 478920 229094
rect 478892 228818 478920 229066
rect 478880 228812 478932 228818
rect 478880 228754 478932 228760
rect 479524 227792 479576 227798
rect 479524 227734 479576 227740
rect 478604 227180 478656 227186
rect 478604 227122 478656 227128
rect 478696 220788 478748 220794
rect 478696 220730 478748 220736
rect 478328 220108 478380 220114
rect 478328 220050 478380 220056
rect 478708 217274 478736 220730
rect 479536 217274 479564 227734
rect 479904 222902 479932 231676
rect 480548 224398 480576 231676
rect 480824 231662 481206 231690
rect 480536 224392 480588 224398
rect 480536 224334 480588 224340
rect 480444 224256 480496 224262
rect 480444 224198 480496 224204
rect 479892 222896 479944 222902
rect 479892 222838 479944 222844
rect 480456 217274 480484 224198
rect 480824 221610 480852 231662
rect 481640 230036 481692 230042
rect 481640 229978 481692 229984
rect 481652 226370 481680 229978
rect 481836 229906 481864 231676
rect 482494 231662 482968 231690
rect 481824 229900 481876 229906
rect 481824 229842 481876 229848
rect 482744 226500 482796 226506
rect 482744 226442 482796 226448
rect 481640 226364 481692 226370
rect 481640 226306 481692 226312
rect 482756 223038 482784 226442
rect 482744 223032 482796 223038
rect 482744 222974 482796 222980
rect 480812 221604 480864 221610
rect 480812 221546 480864 221552
rect 481180 220380 481232 220386
rect 481180 220322 481232 220328
rect 473740 217246 473814 217274
rect 474568 217246 474642 217274
rect 475396 217246 475470 217274
rect 476224 217246 476298 217274
rect 476592 217246 477126 217274
rect 477880 217246 477954 217274
rect 478708 217246 478782 217274
rect 479536 217246 479610 217274
rect 472912 217110 472986 217138
rect 472958 216988 472986 217110
rect 473786 216988 473814 217246
rect 474614 216988 474642 217246
rect 475442 216988 475470 217246
rect 476270 216988 476298 217246
rect 477098 216988 477126 217246
rect 477926 216988 477954 217246
rect 478754 216988 478782 217246
rect 479582 216988 479610 217246
rect 480410 217246 480484 217274
rect 481192 217274 481220 220322
rect 482008 220244 482060 220250
rect 482008 220186 482060 220192
rect 482020 217274 482048 220186
rect 482756 218754 482784 222974
rect 482940 220250 482968 231662
rect 483124 223310 483152 231676
rect 483768 225894 483796 231676
rect 484412 230042 484440 231676
rect 484400 230036 484452 230042
rect 484400 229978 484452 229984
rect 485056 228546 485084 231676
rect 485700 228682 485728 231676
rect 486358 231662 486648 231690
rect 485688 228676 485740 228682
rect 485688 228618 485740 228624
rect 485044 228540 485096 228546
rect 485044 228482 485096 228488
rect 484492 228404 484544 228410
rect 484492 228346 484544 228352
rect 483756 225888 483808 225894
rect 483756 225830 483808 225836
rect 483112 223304 483164 223310
rect 483112 223246 483164 223252
rect 484504 222358 484532 228346
rect 486620 224262 486648 231662
rect 486792 227180 486844 227186
rect 486792 227122 486844 227128
rect 486804 224954 486832 227122
rect 486988 227050 487016 231676
rect 487632 230246 487660 231676
rect 488290 231662 488488 231690
rect 488460 230330 488488 231662
rect 488460 230302 488672 230330
rect 487620 230240 487672 230246
rect 487620 230182 487672 230188
rect 488448 230240 488500 230246
rect 488448 230182 488500 230188
rect 486976 227044 487028 227050
rect 486976 226986 487028 226992
rect 487804 226364 487856 226370
rect 487804 226306 487856 226312
rect 486804 224926 487016 224954
rect 486608 224256 486660 224262
rect 486608 224198 486660 224204
rect 484492 222352 484544 222358
rect 484492 222294 484544 222300
rect 483756 221468 483808 221474
rect 483756 221410 483808 221416
rect 482928 220244 482980 220250
rect 482928 220186 482980 220192
rect 482744 218748 482796 218754
rect 482744 218690 482796 218696
rect 482836 218612 482888 218618
rect 482836 218554 482888 218560
rect 481192 217246 481266 217274
rect 482020 217246 482094 217274
rect 480410 216988 480438 217246
rect 481238 216988 481266 217246
rect 482066 216988 482094 217246
rect 482848 217138 482876 218554
rect 483768 217274 483796 221410
rect 483722 217246 483796 217274
rect 484504 217274 484532 222294
rect 486148 221740 486200 221746
rect 486148 221682 486200 221688
rect 485320 218748 485372 218754
rect 485320 218690 485372 218696
rect 484504 217246 484578 217274
rect 482848 217110 482922 217138
rect 482894 216988 482922 217110
rect 483722 216988 483750 217246
rect 484550 216988 484578 217246
rect 485332 217138 485360 218690
rect 486160 217138 486188 221682
rect 486988 220289 487016 224926
rect 486974 220280 487030 220289
rect 486974 220215 487030 220224
rect 486988 217274 487016 220215
rect 487816 218113 487844 226306
rect 488460 220522 488488 230182
rect 488644 223174 488672 230302
rect 488920 225758 488948 231676
rect 489564 227186 489592 231676
rect 489920 229764 489972 229770
rect 489920 229706 489972 229712
rect 489552 227180 489604 227186
rect 489552 227122 489604 227128
rect 488908 225752 488960 225758
rect 488908 225694 488960 225700
rect 488816 225616 488868 225622
rect 488816 225558 488868 225564
rect 488632 223168 488684 223174
rect 488632 223110 488684 223116
rect 488448 220516 488500 220522
rect 488448 220458 488500 220464
rect 487802 218104 487858 218113
rect 487802 218039 487858 218048
rect 487816 217274 487844 218039
rect 488828 217274 488856 225558
rect 489932 222494 489960 229706
rect 490208 228410 490236 231676
rect 490866 231662 491248 231690
rect 491220 229094 491248 231662
rect 491496 230110 491524 231676
rect 491484 230104 491536 230110
rect 491484 230046 491536 230052
rect 492140 229770 492168 231676
rect 492798 231662 493088 231690
rect 492496 230104 492548 230110
rect 492496 230046 492548 230052
rect 492128 229764 492180 229770
rect 492128 229706 492180 229712
rect 491220 229066 491340 229094
rect 490380 228812 490432 228818
rect 490380 228754 490432 228760
rect 490196 228404 490248 228410
rect 490196 228346 490248 228352
rect 489920 222488 489972 222494
rect 489920 222430 489972 222436
rect 489460 220108 489512 220114
rect 489460 220050 489512 220056
rect 486988 217246 487062 217274
rect 487816 217246 487890 217274
rect 485332 217110 485406 217138
rect 486160 217110 486234 217138
rect 485378 216988 485406 217110
rect 486206 216988 486234 217110
rect 487034 216988 487062 217246
rect 487862 216988 487890 217246
rect 488690 217246 488856 217274
rect 488690 216988 488718 217246
rect 488828 217161 488856 217246
rect 488814 217152 488870 217161
rect 489472 217138 489500 220050
rect 490392 218074 490420 228754
rect 491312 224534 491340 229066
rect 491300 224528 491352 224534
rect 491300 224470 491352 224476
rect 491944 222896 491996 222902
rect 491944 222838 491996 222844
rect 491116 222488 491168 222494
rect 491116 222430 491168 222436
rect 490380 218068 490432 218074
rect 490380 218010 490432 218016
rect 490392 217274 490420 218010
rect 490346 217246 490420 217274
rect 489472 217110 489546 217138
rect 488814 217087 488870 217096
rect 489518 216988 489546 217110
rect 490346 216988 490374 217246
rect 491128 217138 491156 222430
rect 491956 218210 491984 222838
rect 492508 220114 492536 230046
rect 492772 224392 492824 224398
rect 492772 224334 492824 224340
rect 492496 220108 492548 220114
rect 492496 220050 492548 220056
rect 491944 218204 491996 218210
rect 491944 218146 491996 218152
rect 491956 217138 491984 218146
rect 492784 217138 492812 224334
rect 493060 223446 493088 231662
rect 493428 230382 493456 231676
rect 493416 230376 493468 230382
rect 493416 230318 493468 230324
rect 493692 229900 493744 229906
rect 493692 229842 493744 229848
rect 493704 225010 493732 229842
rect 494072 225622 494100 231676
rect 494716 227322 494744 231676
rect 495164 230240 495216 230246
rect 495164 230182 495216 230188
rect 494704 227316 494756 227322
rect 494704 227258 494756 227264
rect 494060 225616 494112 225622
rect 494060 225558 494112 225564
rect 495176 225010 495204 230182
rect 495360 229294 495388 231676
rect 496004 229906 496032 231676
rect 496188 231662 496662 231690
rect 495992 229900 496044 229906
rect 495992 229842 496044 229848
rect 495348 229288 495400 229294
rect 495348 229230 495400 229236
rect 496188 229094 496216 231662
rect 497292 230382 497320 231676
rect 497476 231662 497950 231690
rect 496360 230376 496412 230382
rect 496360 230318 496412 230324
rect 497280 230376 497332 230382
rect 497280 230318 497332 230324
rect 496372 229094 496400 230318
rect 496188 229066 496308 229094
rect 496372 229066 496492 229094
rect 493692 225004 493744 225010
rect 493692 224946 493744 224952
rect 494704 225004 494756 225010
rect 494704 224946 494756 224952
rect 495164 225004 495216 225010
rect 495164 224946 495216 224952
rect 493048 223440 493100 223446
rect 493048 223382 493100 223388
rect 492956 221604 493008 221610
rect 492956 221546 493008 221552
rect 492968 219745 492996 221546
rect 492954 219736 493010 219745
rect 492954 219671 493010 219680
rect 493690 219736 493746 219745
rect 493690 219671 493746 219680
rect 493704 217138 493732 219671
rect 494716 218385 494744 224946
rect 495176 222086 495204 224946
rect 496084 223304 496136 223310
rect 496084 223246 496136 223252
rect 495164 222080 495216 222086
rect 495164 222022 495216 222028
rect 495256 220244 495308 220250
rect 495256 220186 495308 220192
rect 494702 218376 494758 218385
rect 494532 218334 494702 218362
rect 494532 217274 494560 218334
rect 494702 218311 494758 218320
rect 495268 217274 495296 220186
rect 496096 217274 496124 223246
rect 496280 221746 496308 229066
rect 496268 221740 496320 221746
rect 496268 221682 496320 221688
rect 496464 220386 496492 229066
rect 497280 225888 497332 225894
rect 497280 225830 497332 225836
rect 496452 220380 496504 220386
rect 496452 220322 496504 220328
rect 497292 219434 497320 225830
rect 497476 221610 497504 231662
rect 498108 230376 498160 230382
rect 498108 230318 498160 230324
rect 498120 226030 498148 230318
rect 498580 228682 498608 231676
rect 498292 228676 498344 228682
rect 498292 228618 498344 228624
rect 498568 228676 498620 228682
rect 498568 228618 498620 228624
rect 498108 226024 498160 226030
rect 498108 225966 498160 225972
rect 497740 222080 497792 222086
rect 497740 222022 497792 222028
rect 497464 221604 497516 221610
rect 497464 221546 497516 221552
rect 497292 219406 497504 219434
rect 497476 218346 497504 219406
rect 497464 218340 497516 218346
rect 497464 218282 497516 218288
rect 497476 218074 497504 218282
rect 497004 218068 497056 218074
rect 497004 218010 497056 218016
rect 497464 218068 497516 218074
rect 497464 218010 497516 218016
rect 497016 217274 497044 218010
rect 491128 217110 491202 217138
rect 491956 217110 492030 217138
rect 492784 217110 492858 217138
rect 491174 216988 491202 217110
rect 492002 216988 492030 217110
rect 492830 216988 492858 217110
rect 493658 217110 493732 217138
rect 494486 217246 494560 217274
rect 495176 217246 495342 217274
rect 496096 217246 496170 217274
rect 493658 216988 493686 217110
rect 494486 216988 494514 217246
rect 495176 217161 495204 217246
rect 495162 217152 495218 217161
rect 495162 217087 495218 217096
rect 495314 216988 495342 217246
rect 496142 216988 496170 217246
rect 496970 217246 497044 217274
rect 497752 217274 497780 222022
rect 498304 219434 498332 228618
rect 498660 228540 498712 228546
rect 498660 228482 498712 228488
rect 498212 219406 498332 219434
rect 497752 217246 497826 217274
rect 498212 217258 498240 219406
rect 498672 217274 498700 228482
rect 499224 224398 499252 231676
rect 499868 228818 499896 231676
rect 500526 231662 500816 231690
rect 500224 229288 500276 229294
rect 500224 229230 500276 229236
rect 499856 228812 499908 228818
rect 499856 228754 499908 228760
rect 499212 224392 499264 224398
rect 499212 224334 499264 224340
rect 500236 220658 500264 229230
rect 500408 224256 500460 224262
rect 500408 224198 500460 224204
rect 500224 220652 500276 220658
rect 500224 220594 500276 220600
rect 500420 218754 500448 224198
rect 500788 222902 500816 231662
rect 500960 227044 501012 227050
rect 500960 226986 501012 226992
rect 500776 222896 500828 222902
rect 500776 222838 500828 222844
rect 500972 220368 501000 226986
rect 501156 225894 501184 231676
rect 501340 231662 501814 231690
rect 501144 225888 501196 225894
rect 501144 225830 501196 225836
rect 500972 220340 501184 220368
rect 501156 219570 501184 220340
rect 501340 220250 501368 231662
rect 502444 228546 502472 231676
rect 503102 231662 503392 231690
rect 502432 228540 502484 228546
rect 502432 228482 502484 228488
rect 503364 223174 503392 231662
rect 503732 229158 503760 231676
rect 503720 229152 503772 229158
rect 503720 229094 503772 229100
rect 504180 227180 504232 227186
rect 504180 227122 504232 227128
rect 503628 225752 503680 225758
rect 503628 225694 503680 225700
rect 503168 223168 503220 223174
rect 503168 223110 503220 223116
rect 503352 223168 503404 223174
rect 503352 223110 503404 223116
rect 501880 220516 501932 220522
rect 501880 220458 501932 220464
rect 501328 220244 501380 220250
rect 501328 220186 501380 220192
rect 501144 219564 501196 219570
rect 501144 219506 501196 219512
rect 500408 218748 500460 218754
rect 500408 218690 500460 218696
rect 500420 217274 500448 218690
rect 501156 217274 501184 219506
rect 496970 216988 496998 217246
rect 497798 216988 497826 217246
rect 498200 217252 498252 217258
rect 498200 217194 498252 217200
rect 498626 217246 498700 217274
rect 499442 217252 499494 217258
rect 498626 217122 498654 217246
rect 499442 217194 499494 217200
rect 500282 217246 500448 217274
rect 501110 217246 501184 217274
rect 501892 217274 501920 220458
rect 503180 218482 503208 223110
rect 503640 219910 503668 225694
rect 503628 219904 503680 219910
rect 503628 219846 503680 219852
rect 502800 218476 502852 218482
rect 502800 218418 502852 218424
rect 503168 218476 503220 218482
rect 503168 218418 503220 218424
rect 502248 218204 502300 218210
rect 502248 218146 502300 218152
rect 502260 217297 502288 218146
rect 502246 217288 502302 217297
rect 501892 217246 501966 217274
rect 498614 217116 498666 217122
rect 498614 217058 498666 217064
rect 498626 216988 498654 217058
rect 499454 216988 499482 217194
rect 500282 216988 500310 217246
rect 501110 216988 501138 217246
rect 501938 216988 501966 217246
rect 502246 217223 502302 217232
rect 502812 217138 502840 218418
rect 503640 217274 503668 219846
rect 504192 219434 504220 227122
rect 504376 224262 504404 231676
rect 505020 227050 505048 231676
rect 505664 229294 505692 231676
rect 506216 231662 506322 231690
rect 505652 229288 505704 229294
rect 505652 229230 505704 229236
rect 505192 228404 505244 228410
rect 505192 228346 505244 228352
rect 505008 227044 505060 227050
rect 505008 226986 505060 226992
rect 505204 224670 505232 228346
rect 506216 227186 506244 231662
rect 506388 229900 506440 229906
rect 506388 229842 506440 229848
rect 506400 228954 506428 229842
rect 506388 228948 506440 228954
rect 506388 228890 506440 228896
rect 506204 227180 506256 227186
rect 506204 227122 506256 227128
rect 506952 224806 506980 231676
rect 507596 229906 507624 231676
rect 507584 229900 507636 229906
rect 507584 229842 507636 229848
rect 507124 229764 507176 229770
rect 507124 229706 507176 229712
rect 506940 224800 506992 224806
rect 506940 224742 506992 224748
rect 505192 224664 505244 224670
rect 505192 224606 505244 224612
rect 504364 224256 504416 224262
rect 504364 224198 504416 224204
rect 504364 222488 504416 222494
rect 504364 222430 504416 222436
rect 504376 222222 504404 222430
rect 504364 222216 504416 222222
rect 504364 222158 504416 222164
rect 504192 219406 504404 219434
rect 502766 217110 502840 217138
rect 503594 217246 503668 217274
rect 504376 217274 504404 219406
rect 505204 217274 505232 224606
rect 506020 224528 506072 224534
rect 506020 224470 506072 224476
rect 506032 217274 506060 224470
rect 506848 220108 506900 220114
rect 506848 220050 506900 220056
rect 506860 217274 506888 220050
rect 507136 218210 507164 229706
rect 508240 222766 508268 231676
rect 508884 225758 508912 231676
rect 509528 229702 509556 231676
rect 509516 229696 509568 229702
rect 509516 229638 509568 229644
rect 509884 229152 509936 229158
rect 509884 229094 509936 229100
rect 508872 225752 508924 225758
rect 508872 225694 508924 225700
rect 509700 225616 509752 225622
rect 509700 225558 509752 225564
rect 509712 224126 509740 225558
rect 509700 224120 509752 224126
rect 509700 224062 509752 224068
rect 508596 223440 508648 223446
rect 508596 223382 508648 223388
rect 508228 222760 508280 222766
rect 508228 222702 508280 222708
rect 508044 218748 508096 218754
rect 508044 218690 508096 218696
rect 507676 218612 507728 218618
rect 507676 218554 507728 218560
rect 507688 218210 507716 218554
rect 508056 218482 508084 218690
rect 507860 218476 507912 218482
rect 507860 218418 507912 218424
rect 508044 218476 508096 218482
rect 508044 218418 508096 218424
rect 507872 218210 507900 218418
rect 507124 218204 507176 218210
rect 507124 218146 507176 218152
rect 507676 218204 507728 218210
rect 507676 218146 507728 218152
rect 507860 218204 507912 218210
rect 507860 218146 507912 218152
rect 504376 217246 504450 217274
rect 505204 217246 505278 217274
rect 506032 217246 506106 217274
rect 506860 217246 506934 217274
rect 502766 216988 502794 217110
rect 503594 216988 503622 217246
rect 504422 216988 504450 217246
rect 505250 216988 505278 217246
rect 506078 217190 506106 217246
rect 506066 217184 506118 217190
rect 506066 217126 506118 217132
rect 506078 216988 506106 217126
rect 506906 216988 506934 217246
rect 507688 217138 507716 218146
rect 508608 217326 508636 223382
rect 509896 221882 509924 229094
rect 510172 225622 510200 231676
rect 510816 230382 510844 231676
rect 510804 230376 510856 230382
rect 510804 230318 510856 230324
rect 511460 230246 511488 231676
rect 511908 230376 511960 230382
rect 511908 230318 511960 230324
rect 511448 230240 511500 230246
rect 511448 230182 511500 230188
rect 510620 229288 510672 229294
rect 510620 229230 510672 229236
rect 510632 227322 510660 229230
rect 511920 229094 511948 230318
rect 511828 229066 511948 229094
rect 510620 227316 510672 227322
rect 510620 227258 510672 227264
rect 510988 226908 511040 226914
rect 510988 226850 511040 226856
rect 510160 225616 510212 225622
rect 510160 225558 510212 225564
rect 510160 224120 510212 224126
rect 510160 224062 510212 224068
rect 509884 221876 509936 221882
rect 509884 221818 509936 221824
rect 509332 220380 509384 220386
rect 509332 220322 509384 220328
rect 508596 217320 508648 217326
rect 508596 217262 508648 217268
rect 509344 217274 509372 220322
rect 510172 217274 510200 224062
rect 511000 217569 511028 226850
rect 511828 220794 511856 229066
rect 512104 228410 512132 231676
rect 512762 231662 513144 231690
rect 512736 228948 512788 228954
rect 512736 228890 512788 228896
rect 512092 228404 512144 228410
rect 512092 228346 512144 228352
rect 511816 220788 511868 220794
rect 511816 220730 511868 220736
rect 511816 220652 511868 220658
rect 511816 220594 511868 220600
rect 510986 217560 511042 217569
rect 510986 217495 511042 217504
rect 508608 217138 508636 217262
rect 509344 217246 509418 217274
rect 510172 217246 510246 217274
rect 507688 217110 507762 217138
rect 507734 216988 507762 217110
rect 508562 217110 508636 217138
rect 508562 216988 508590 217110
rect 509390 216988 509418 217246
rect 510218 216988 510246 217246
rect 511000 217138 511028 217495
rect 511828 217274 511856 220594
rect 512748 218890 512776 228890
rect 513116 220114 513144 231662
rect 513392 229294 513420 231676
rect 513380 229288 513432 229294
rect 513380 229230 513432 229236
rect 514036 227458 514064 231676
rect 514024 227452 514076 227458
rect 514024 227394 514076 227400
rect 514300 226024 514352 226030
rect 514300 225966 514352 225972
rect 513564 221740 513616 221746
rect 513564 221682 513616 221688
rect 513576 221513 513604 221682
rect 513562 221504 513618 221513
rect 513562 221439 513618 221448
rect 513104 220108 513156 220114
rect 513104 220050 513156 220056
rect 512736 218884 512788 218890
rect 512736 218826 512788 218832
rect 512748 217274 512776 218826
rect 513576 217274 513604 221439
rect 511828 217246 511902 217274
rect 511000 217110 511074 217138
rect 511046 216988 511074 217110
rect 511874 216988 511902 217246
rect 512702 217246 512776 217274
rect 513530 217246 513604 217274
rect 514312 217274 514340 225966
rect 514680 223310 514708 231676
rect 515324 229158 515352 231676
rect 515496 229696 515548 229702
rect 515496 229638 515548 229644
rect 515312 229152 515364 229158
rect 515312 229094 515364 229100
rect 514668 223304 514720 223310
rect 514668 223246 514720 223252
rect 515508 222086 515536 229638
rect 515772 228676 515824 228682
rect 515772 228618 515824 228624
rect 515496 222080 515548 222086
rect 515496 222022 515548 222028
rect 515128 221604 515180 221610
rect 515128 221546 515180 221552
rect 515140 220017 515168 221546
rect 515784 221241 515812 228618
rect 515968 224534 515996 231676
rect 516612 226030 516640 231676
rect 517256 230042 517284 231676
rect 517520 230240 517572 230246
rect 517520 230182 517572 230188
rect 517244 230036 517296 230042
rect 517244 229978 517296 229984
rect 516784 229900 516836 229906
rect 516784 229842 516836 229848
rect 516796 229094 516824 229842
rect 516796 229066 517008 229094
rect 516600 226024 516652 226030
rect 516600 225966 516652 225972
rect 515956 224528 516008 224534
rect 515956 224470 516008 224476
rect 516784 224392 516836 224398
rect 516784 224334 516836 224340
rect 515770 221232 515826 221241
rect 515770 221167 515826 221176
rect 515126 220008 515182 220017
rect 515126 219943 515182 219952
rect 515140 217274 515168 219943
rect 515784 219434 515812 221167
rect 515784 219406 516088 219434
rect 516060 217274 516088 219406
rect 514312 217246 514386 217274
rect 515140 217246 515214 217274
rect 512702 216988 512730 217246
rect 513530 216988 513558 217246
rect 514358 216988 514386 217246
rect 515186 216988 515214 217246
rect 516014 217246 516088 217274
rect 516796 217274 516824 224334
rect 516980 220386 517008 229066
rect 517532 223446 517560 230182
rect 517900 228682 517928 231676
rect 518544 228818 518572 231676
rect 519188 229906 519216 231676
rect 519176 229900 519228 229906
rect 519176 229842 519228 229848
rect 519084 229288 519136 229294
rect 519084 229230 519136 229236
rect 518164 228812 518216 228818
rect 518164 228754 518216 228760
rect 518532 228812 518584 228818
rect 518532 228754 518584 228760
rect 517888 228676 517940 228682
rect 517888 228618 517940 228624
rect 517520 223440 517572 223446
rect 517520 223382 517572 223388
rect 517520 222896 517572 222902
rect 517520 222838 517572 222844
rect 517532 220862 517560 222838
rect 517520 220856 517572 220862
rect 517520 220798 517572 220804
rect 516968 220380 517020 220386
rect 516968 220322 517020 220328
rect 518176 218754 518204 228754
rect 519096 223990 519124 229230
rect 519268 225888 519320 225894
rect 519268 225830 519320 225836
rect 519084 223984 519136 223990
rect 519084 223926 519136 223932
rect 518532 220856 518584 220862
rect 518532 220798 518584 220804
rect 517704 218748 517756 218754
rect 517704 218690 517756 218696
rect 518164 218748 518216 218754
rect 518164 218690 518216 218696
rect 517716 217274 517744 218690
rect 518544 217274 518572 220798
rect 516796 217246 516870 217274
rect 516014 216988 516042 217246
rect 516842 216988 516870 217246
rect 517670 217246 517744 217274
rect 518498 217246 518572 217274
rect 519280 217274 519308 225830
rect 519832 222902 519860 231676
rect 520476 223650 520504 231676
rect 521120 230382 521148 231676
rect 521108 230376 521160 230382
rect 521108 230318 521160 230324
rect 520924 229152 520976 229158
rect 520924 229094 520976 229100
rect 520464 223644 520516 223650
rect 520464 223586 520516 223592
rect 519820 222896 519872 222902
rect 519820 222838 519872 222844
rect 520936 220658 520964 229094
rect 521108 228540 521160 228546
rect 521108 228482 521160 228488
rect 521120 221270 521148 228482
rect 521764 225894 521792 231676
rect 522422 231662 522896 231690
rect 521752 225888 521804 225894
rect 521752 225830 521804 225836
rect 521752 223168 521804 223174
rect 521752 223110 521804 223116
rect 521108 221264 521160 221270
rect 521108 221206 521160 221212
rect 520924 220652 520976 220658
rect 520924 220594 520976 220600
rect 520188 220244 520240 220250
rect 520188 220186 520240 220192
rect 520200 219473 520228 220186
rect 520186 219464 520242 219473
rect 521120 219434 521148 221206
rect 520186 219399 520242 219408
rect 521028 219406 521148 219434
rect 520004 218748 520056 218754
rect 520004 218690 520056 218696
rect 520016 217569 520044 218690
rect 520002 217560 520058 217569
rect 520002 217495 520058 217504
rect 520200 217274 520228 219399
rect 521028 217274 521056 219406
rect 519280 217246 519354 217274
rect 517670 216988 517698 217246
rect 518498 216988 518526 217246
rect 519326 216988 519354 217246
rect 520154 217246 520228 217274
rect 520982 217246 521056 217274
rect 521764 217274 521792 223110
rect 522580 221876 522632 221882
rect 522580 221818 522632 221824
rect 522592 220969 522620 221818
rect 522868 221610 522896 231662
rect 523052 229770 523080 231676
rect 523040 229764 523092 229770
rect 523040 229706 523092 229712
rect 523696 227050 523724 231676
rect 524248 231662 524354 231690
rect 523040 227044 523092 227050
rect 523040 226986 523092 226992
rect 523684 227044 523736 227050
rect 523684 226986 523736 226992
rect 522856 221604 522908 221610
rect 522856 221546 522908 221552
rect 522578 220960 522634 220969
rect 522578 220895 522634 220904
rect 522592 217274 522620 220895
rect 523052 217870 523080 226986
rect 523500 224256 523552 224262
rect 523500 224198 523552 224204
rect 523512 221134 523540 224198
rect 523684 222488 523736 222494
rect 523684 222430 523736 222436
rect 523696 222222 523724 222430
rect 523684 222216 523736 222222
rect 523684 222158 523736 222164
rect 524248 221746 524276 231662
rect 524604 230036 524656 230042
rect 524604 229978 524656 229984
rect 524616 227594 524644 229978
rect 524984 229158 525012 231676
rect 524972 229152 525024 229158
rect 524972 229094 525024 229100
rect 524604 227588 524656 227594
rect 524604 227530 524656 227536
rect 524420 227316 524472 227322
rect 524420 227258 524472 227264
rect 524432 224262 524460 227258
rect 525628 224398 525656 231676
rect 526272 227322 526300 231676
rect 526444 230376 526496 230382
rect 526444 230318 526496 230324
rect 526456 228954 526484 230318
rect 526916 229634 526944 231676
rect 526904 229628 526956 229634
rect 526904 229570 526956 229576
rect 526444 228948 526496 228954
rect 526444 228890 526496 228896
rect 527560 228546 527588 231676
rect 528218 231662 528416 231690
rect 527548 228540 527600 228546
rect 527548 228482 527600 228488
rect 526260 227316 526312 227322
rect 526260 227258 526312 227264
rect 525984 227180 526036 227186
rect 525984 227122 526036 227128
rect 525616 224392 525668 224398
rect 525616 224334 525668 224340
rect 524420 224256 524472 224262
rect 524420 224198 524472 224204
rect 525064 224256 525116 224262
rect 525064 224198 525116 224204
rect 524236 221740 524288 221746
rect 524236 221682 524288 221688
rect 523500 221128 523552 221134
rect 523500 221070 523552 221076
rect 523040 217864 523092 217870
rect 523040 217806 523092 217812
rect 523512 217274 523540 221070
rect 524236 217864 524288 217870
rect 524236 217806 524288 217812
rect 521764 217246 521838 217274
rect 522592 217246 522666 217274
rect 520154 216988 520182 217246
rect 520982 216988 521010 217246
rect 521810 216988 521838 217246
rect 522638 216988 522666 217246
rect 523466 217246 523540 217274
rect 523466 216988 523494 217246
rect 524248 217138 524276 217806
rect 525076 217274 525104 224198
rect 525996 220998 526024 227122
rect 526720 224800 526772 224806
rect 526720 224742 526772 224748
rect 525984 220992 526036 220998
rect 525984 220934 526036 220940
rect 525996 217274 526024 220934
rect 525076 217246 525150 217274
rect 524248 217110 524322 217138
rect 524294 216988 524322 217110
rect 525122 216988 525150 217246
rect 525950 217246 526024 217274
rect 526732 217274 526760 224742
rect 527824 222760 527876 222766
rect 527824 222702 527876 222708
rect 527548 220380 527600 220386
rect 527548 220322 527600 220328
rect 527560 219638 527588 220322
rect 527548 219632 527600 219638
rect 527548 219574 527600 219580
rect 527560 217274 527588 219574
rect 527836 217734 527864 222702
rect 528388 220250 528416 231662
rect 528848 230042 528876 231676
rect 528836 230036 528888 230042
rect 528836 229978 528888 229984
rect 528560 229900 528612 229906
rect 528560 229842 528612 229848
rect 528572 226166 528600 229842
rect 528560 226160 528612 226166
rect 528560 226102 528612 226108
rect 529204 225752 529256 225758
rect 529204 225694 529256 225700
rect 528376 220244 528428 220250
rect 528376 220186 528428 220192
rect 527824 217728 527876 217734
rect 527824 217670 527876 217676
rect 528376 217728 528428 217734
rect 528376 217670 528428 217676
rect 526732 217246 526806 217274
rect 527560 217246 527634 217274
rect 525950 216988 525978 217246
rect 526778 216988 526806 217246
rect 527606 216988 527634 217246
rect 528388 217138 528416 217670
rect 529216 217274 529244 225694
rect 529492 222494 529520 231676
rect 530136 230382 530164 231676
rect 530124 230376 530176 230382
rect 530124 230318 530176 230324
rect 530780 230246 530808 231676
rect 531136 230376 531188 230382
rect 531136 230318 531188 230324
rect 530768 230240 530820 230246
rect 530768 230182 530820 230188
rect 529940 229152 529992 229158
rect 529940 229094 529992 229100
rect 529952 224806 529980 229094
rect 530952 225616 531004 225622
rect 530952 225558 531004 225564
rect 529940 224800 529992 224806
rect 529940 224742 529992 224748
rect 529848 222624 529900 222630
rect 529848 222566 529900 222572
rect 529480 222488 529532 222494
rect 529480 222430 529532 222436
rect 529860 222086 529888 222566
rect 529848 222080 529900 222086
rect 529848 222022 529900 222028
rect 529860 221354 529888 222022
rect 529860 221326 530072 221354
rect 530044 217274 530072 221326
rect 530964 217462 530992 225558
rect 531148 220386 531176 230318
rect 531424 225622 531452 231676
rect 531412 225616 531464 225622
rect 531412 225558 531464 225564
rect 531504 223440 531556 223446
rect 531504 223382 531556 223388
rect 531136 220380 531188 220386
rect 531136 220322 531188 220328
rect 531516 217569 531544 223382
rect 532068 223174 532096 231676
rect 532712 230178 532740 231676
rect 532700 230172 532752 230178
rect 532700 230114 532752 230120
rect 533356 227186 533384 231676
rect 533528 230308 533580 230314
rect 533528 230250 533580 230256
rect 533540 230042 533568 230250
rect 533528 230036 533580 230042
rect 533528 229978 533580 229984
rect 533528 228404 533580 228410
rect 533528 228346 533580 228352
rect 533344 227180 533396 227186
rect 533344 227122 533396 227128
rect 532056 223168 532108 223174
rect 532056 223110 532108 223116
rect 531688 220516 531740 220522
rect 531688 220458 531740 220464
rect 531502 217560 531558 217569
rect 531502 217495 531558 217504
rect 530952 217456 531004 217462
rect 530952 217398 531004 217404
rect 529216 217246 529290 217274
rect 530044 217246 530118 217274
rect 528388 217110 528462 217138
rect 528434 216988 528462 217110
rect 529262 216988 529290 217246
rect 530090 216988 530118 217246
rect 530964 217138 530992 217398
rect 531700 217274 531728 220458
rect 533540 219434 533568 228346
rect 534000 222086 534028 231676
rect 534644 230042 534672 231676
rect 534632 230036 534684 230042
rect 534632 229978 534684 229984
rect 534724 229764 534776 229770
rect 534724 229706 534776 229712
rect 534736 223446 534764 229706
rect 535288 223990 535316 231676
rect 535736 227452 535788 227458
rect 535736 227394 535788 227400
rect 535276 223984 535328 223990
rect 535276 223926 535328 223932
rect 535092 223780 535144 223786
rect 535092 223722 535144 223728
rect 534724 223440 534776 223446
rect 534724 223382 534776 223388
rect 533988 222080 534040 222086
rect 533988 222022 534040 222028
rect 534172 220108 534224 220114
rect 534172 220050 534224 220056
rect 533448 219406 533568 219434
rect 533448 217598 533476 219406
rect 533436 217592 533488 217598
rect 532514 217560 532570 217569
rect 533436 217534 533488 217540
rect 532514 217495 532570 217504
rect 531700 217246 531774 217274
rect 530918 217110 530992 217138
rect 530918 216988 530946 217110
rect 531746 216988 531774 217246
rect 532528 217138 532556 217495
rect 533448 217138 533476 217534
rect 532528 217110 532602 217138
rect 532574 216988 532602 217110
rect 533402 217110 533476 217138
rect 534184 217138 534212 220050
rect 535104 217138 535132 223722
rect 535748 222057 535776 227394
rect 535932 225758 535960 231676
rect 536576 229906 536604 231676
rect 536564 229900 536616 229906
rect 536564 229842 536616 229848
rect 536104 229628 536156 229634
rect 536104 229570 536156 229576
rect 535920 225752 535972 225758
rect 535920 225694 535972 225700
rect 536116 222086 536144 229570
rect 537220 228410 537248 231676
rect 537878 231662 538168 231690
rect 537208 228404 537260 228410
rect 537208 228346 537260 228352
rect 536656 223304 536708 223310
rect 536656 223246 536708 223252
rect 536104 222080 536156 222086
rect 535734 222048 535790 222057
rect 536104 222022 536156 222028
rect 535734 221983 535790 221992
rect 535748 217274 535776 221983
rect 536380 217864 536432 217870
rect 536380 217806 536432 217812
rect 536392 217598 536420 217806
rect 536380 217592 536432 217598
rect 536380 217534 536432 217540
rect 535748 217246 535914 217274
rect 534184 217110 534258 217138
rect 533402 216988 533430 217110
rect 534230 216988 534258 217110
rect 535058 217110 535132 217138
rect 535058 216988 535086 217110
rect 535886 216988 535914 217246
rect 536668 217138 536696 223246
rect 537484 220652 537536 220658
rect 537484 220594 537536 220600
rect 537496 218754 537524 220594
rect 538140 220114 538168 231662
rect 538312 230308 538364 230314
rect 538312 230250 538364 230256
rect 538324 227458 538352 230250
rect 538508 229770 538536 231676
rect 538784 231662 539166 231690
rect 538496 229764 538548 229770
rect 538496 229706 538548 229712
rect 538784 229094 538812 231662
rect 539600 230444 539652 230450
rect 539600 230386 539652 230392
rect 538508 229066 538812 229094
rect 538312 227452 538364 227458
rect 538312 227394 538364 227400
rect 538312 224528 538364 224534
rect 538312 224470 538364 224476
rect 538324 221354 538352 224470
rect 538508 221474 538536 229066
rect 539612 228682 539640 230386
rect 547144 230172 547196 230178
rect 547144 230114 547196 230120
rect 544016 228948 544068 228954
rect 544016 228890 544068 228896
rect 541624 228812 541676 228818
rect 541624 228754 541676 228760
rect 539416 228676 539468 228682
rect 539416 228618 539468 228624
rect 539600 228676 539652 228682
rect 539600 228618 539652 228624
rect 539428 228274 539456 228618
rect 539416 228268 539468 228274
rect 539416 228210 539468 228216
rect 540796 228268 540848 228274
rect 540796 228210 540848 228216
rect 539968 227588 540020 227594
rect 539968 227530 540020 227536
rect 538680 226024 538732 226030
rect 538680 225966 538732 225972
rect 538692 224954 538720 225966
rect 538692 224926 539180 224954
rect 538864 224528 538916 224534
rect 538864 224470 538916 224476
rect 538876 224262 538904 224470
rect 538864 224256 538916 224262
rect 538864 224198 538916 224204
rect 538496 221468 538548 221474
rect 538496 221410 538548 221416
rect 538680 221400 538732 221406
rect 538324 221348 538680 221354
rect 538324 221342 538732 221348
rect 538324 221326 538720 221342
rect 538128 220108 538180 220114
rect 538128 220050 538180 220056
rect 537484 218748 537536 218754
rect 537484 218690 537536 218696
rect 537496 217138 537524 218690
rect 538324 217138 538352 221326
rect 539152 217274 539180 224926
rect 539324 224256 539376 224262
rect 539324 224198 539376 224204
rect 539336 223990 539364 224198
rect 539324 223984 539376 223990
rect 539324 223926 539376 223932
rect 539980 223922 540008 227530
rect 539968 223916 540020 223922
rect 539968 223858 540020 223864
rect 539600 222080 539652 222086
rect 539784 222080 539836 222086
rect 539600 222022 539652 222028
rect 539782 222048 539784 222057
rect 539836 222048 539838 222057
rect 539612 221814 539640 222022
rect 539782 221983 539838 221992
rect 539324 221808 539376 221814
rect 539324 221750 539376 221756
rect 539600 221808 539652 221814
rect 539600 221750 539652 221756
rect 539336 221542 539364 221750
rect 539324 221536 539376 221542
rect 539324 221478 539376 221484
rect 539980 217274 540008 223858
rect 540808 219774 540836 228210
rect 540796 219768 540848 219774
rect 540796 219710 540848 219716
rect 540808 217274 540836 219710
rect 541636 217274 541664 228754
rect 542636 226160 542688 226166
rect 542636 226102 542688 226108
rect 542360 222896 542412 222902
rect 542360 222838 542412 222844
rect 542372 217598 542400 222838
rect 542648 219162 542676 226102
rect 544028 223650 544056 228890
rect 545764 225888 545816 225894
rect 545764 225830 545816 225836
rect 543832 223644 543884 223650
rect 543832 223586 543884 223592
rect 544016 223644 544068 223650
rect 544016 223586 544068 223592
rect 544936 223644 544988 223650
rect 544936 223586 544988 223592
rect 542636 219156 542688 219162
rect 542636 219098 542688 219104
rect 542360 217592 542412 217598
rect 542360 217534 542412 217540
rect 542648 217274 542676 219098
rect 543280 217592 543332 217598
rect 543280 217534 543332 217540
rect 539152 217246 539226 217274
rect 539980 217246 540054 217274
rect 540808 217246 540882 217274
rect 541636 217246 541710 217274
rect 536668 217110 536742 217138
rect 537496 217110 537570 217138
rect 538324 217110 538398 217138
rect 536714 216988 536742 217110
rect 537542 216988 537570 217110
rect 538370 216988 538398 217110
rect 539198 216988 539226 217246
rect 540026 216988 540054 217246
rect 540854 216988 540882 217246
rect 541682 216988 541710 217246
rect 542510 217246 542676 217274
rect 542510 216988 542538 217246
rect 543292 217138 543320 217534
rect 543844 217274 543872 223586
rect 544948 217274 544976 223586
rect 545776 220726 545804 225830
rect 547156 221678 547184 230114
rect 549260 230036 549312 230042
rect 549260 229978 549312 229984
rect 548340 227044 548392 227050
rect 548340 226986 548392 226992
rect 547420 223440 547472 223446
rect 547420 223382 547472 223388
rect 546592 221672 546644 221678
rect 546592 221614 546644 221620
rect 547144 221672 547196 221678
rect 547144 221614 547196 221620
rect 545764 220720 545816 220726
rect 545764 220662 545816 220668
rect 545776 217274 545804 220662
rect 546604 217274 546632 221614
rect 547432 219026 547460 223382
rect 547834 221808 547886 221814
rect 547832 221776 547834 221785
rect 547972 221808 548024 221814
rect 547886 221776 547888 221785
rect 547972 221750 548024 221756
rect 547832 221711 547888 221720
rect 547984 221626 548012 221750
rect 547846 221598 548012 221626
rect 547846 221542 547874 221598
rect 547834 221536 547886 221542
rect 547834 221478 547886 221484
rect 547972 221536 548024 221542
rect 547972 221478 548024 221484
rect 547984 220726 548012 221478
rect 547972 220720 548024 220726
rect 547972 220662 548024 220668
rect 548352 220522 548380 226986
rect 549272 224874 549300 229978
rect 553308 228540 553360 228546
rect 553308 228482 553360 228488
rect 551560 227316 551612 227322
rect 551560 227258 551612 227264
rect 549260 224868 549312 224874
rect 549260 224810 549312 224816
rect 549076 224800 549128 224806
rect 549128 224748 549300 224754
rect 549076 224742 549300 224748
rect 549088 224726 549300 224742
rect 549272 224505 549300 224726
rect 549258 224496 549314 224505
rect 549258 224431 549314 224440
rect 549902 224496 549958 224505
rect 549902 224431 549958 224440
rect 549076 221808 549128 221814
rect 549260 221808 549312 221814
rect 549076 221750 549128 221756
rect 549258 221776 549260 221785
rect 549312 221776 549314 221785
rect 548340 220516 548392 220522
rect 548340 220458 548392 220464
rect 548156 219292 548208 219298
rect 548156 219234 548208 219240
rect 547420 219020 547472 219026
rect 547420 218962 547472 218968
rect 547432 217274 547460 218962
rect 548168 218890 548196 219234
rect 548156 218884 548208 218890
rect 548156 218826 548208 218832
rect 548352 217274 548380 220458
rect 543844 217246 544194 217274
rect 544948 217246 545022 217274
rect 545776 217246 545850 217274
rect 546604 217246 546678 217274
rect 547432 217246 547506 217274
rect 543292 217110 543366 217138
rect 543338 216988 543366 217110
rect 544166 216988 544194 217246
rect 544994 216988 545022 217246
rect 545822 216988 545850 217246
rect 546650 216988 546678 217246
rect 547478 216988 547506 217246
rect 548306 217246 548380 217274
rect 549088 217274 549116 221750
rect 549258 221711 549314 221720
rect 549916 217274 549944 224431
rect 550824 224392 550876 224398
rect 550824 224334 550876 224340
rect 550836 220658 550864 224334
rect 550824 220652 550876 220658
rect 550824 220594 550876 220600
rect 550836 217274 550864 220594
rect 549088 217246 549162 217274
rect 549916 217246 549990 217274
rect 548306 216988 548334 217246
rect 549134 216988 549162 217246
rect 549962 216988 549990 217246
rect 550790 217246 550864 217274
rect 551572 217274 551600 227258
rect 552848 224528 552900 224534
rect 552846 224496 552848 224505
rect 552900 224496 552902 224505
rect 552846 224431 552902 224440
rect 552480 222760 552532 222766
rect 552480 222702 552532 222708
rect 552492 222494 552520 222702
rect 552480 222488 552532 222494
rect 552480 222430 552532 222436
rect 552664 222488 552716 222494
rect 552664 222430 552716 222436
rect 552676 222222 552704 222430
rect 552664 222216 552716 222222
rect 552664 222158 552716 222164
rect 552848 222216 552900 222222
rect 552848 222158 552900 222164
rect 552860 221814 552888 222158
rect 553320 221814 553348 228482
rect 554056 222902 554084 249047
rect 555424 244316 555476 244322
rect 555424 244258 555476 244264
rect 554502 240408 554558 240417
rect 554502 240343 554558 240352
rect 554516 240174 554544 240343
rect 554504 240168 554556 240174
rect 554504 240110 554556 240116
rect 554320 238740 554372 238746
rect 554320 238682 554372 238688
rect 554332 238241 554360 238682
rect 554318 238232 554374 238241
rect 554318 238167 554374 238176
rect 554412 234592 554464 234598
rect 554412 234534 554464 234540
rect 554424 233889 554452 234534
rect 554410 233880 554466 233889
rect 554410 233815 554466 233824
rect 555436 227050 555464 244258
rect 556816 228546 556844 251194
rect 557172 228676 557224 228682
rect 557172 228618 557224 228624
rect 556804 228540 556856 228546
rect 556804 228482 556856 228488
rect 556068 227452 556120 227458
rect 556068 227394 556120 227400
rect 555424 227044 555476 227050
rect 555424 226986 555476 226992
rect 556080 224954 556108 227394
rect 555804 224926 556108 224954
rect 557184 224954 557212 228618
rect 558196 225894 558224 255546
rect 559564 246356 559616 246362
rect 559564 246298 559616 246304
rect 559576 236842 559604 246298
rect 559564 236836 559616 236842
rect 559564 236778 559616 236784
rect 560956 230110 560984 256702
rect 562324 252612 562376 252618
rect 562324 252554 562376 252560
rect 560944 230104 560996 230110
rect 560944 230046 560996 230052
rect 559564 229900 559616 229906
rect 559564 229842 559616 229848
rect 558184 225888 558236 225894
rect 558184 225830 558236 225836
rect 558276 225616 558328 225622
rect 558276 225558 558328 225564
rect 558288 224954 558316 225558
rect 557184 224926 557396 224954
rect 558288 224926 558408 224954
rect 554778 224904 554834 224913
rect 554778 224839 554780 224848
rect 554832 224839 554834 224848
rect 554780 224810 554832 224816
rect 555804 224806 555832 224926
rect 556080 224890 556108 224926
rect 556080 224862 556384 224890
rect 554964 224800 555016 224806
rect 554964 224742 555016 224748
rect 555792 224800 555844 224806
rect 555792 224742 555844 224748
rect 555976 224800 556028 224806
rect 555976 224742 556028 224748
rect 554044 222896 554096 222902
rect 554044 222838 554096 222844
rect 553950 221912 554006 221921
rect 553950 221847 554006 221856
rect 552112 221808 552164 221814
rect 552112 221750 552164 221756
rect 552848 221808 552900 221814
rect 552848 221750 552900 221756
rect 553308 221808 553360 221814
rect 553308 221750 553360 221756
rect 552124 219434 552152 221750
rect 552296 221536 552348 221542
rect 552296 221478 552348 221484
rect 552308 221354 552336 221478
rect 553124 221400 553176 221406
rect 552308 221348 553124 221354
rect 552308 221342 553176 221348
rect 552308 221326 553164 221342
rect 552124 219406 552428 219434
rect 552400 217274 552428 219406
rect 553320 217274 553348 221750
rect 553964 221678 553992 221847
rect 553952 221672 554004 221678
rect 553952 221614 554004 221620
rect 554044 220244 554096 220250
rect 554044 220186 554096 220192
rect 551572 217246 551646 217274
rect 552400 217246 552474 217274
rect 550790 216988 550818 217246
rect 551618 216988 551646 217246
rect 552446 216988 552474 217246
rect 553274 217246 553348 217274
rect 553274 216988 553302 217246
rect 554056 217138 554084 220186
rect 554976 217274 555004 224742
rect 555988 224262 556016 224742
rect 556356 224398 556384 224862
rect 556344 224392 556396 224398
rect 556344 224334 556396 224340
rect 555976 224256 556028 224262
rect 555976 224198 556028 224204
rect 555700 222760 555752 222766
rect 555700 222702 555752 222708
rect 555712 220250 555740 222702
rect 556528 220380 556580 220386
rect 556528 220322 556580 220328
rect 555700 220244 555752 220250
rect 555700 220186 555752 220192
rect 554930 217246 555004 217274
rect 554056 217110 554130 217138
rect 554102 216988 554130 217110
rect 554930 216988 554958 217246
rect 555712 217138 555740 220186
rect 556540 217138 556568 220322
rect 557368 219026 557396 224926
rect 558184 222760 558236 222766
rect 558184 222702 558236 222708
rect 558196 222222 558224 222702
rect 558184 222216 558236 222222
rect 558184 222158 558236 222164
rect 557998 220552 558054 220561
rect 557998 220487 558054 220496
rect 558012 220250 558040 220487
rect 558380 220250 558408 224926
rect 559012 223168 559064 223174
rect 559012 223110 559064 223116
rect 558552 222216 558604 222222
rect 558552 222158 558604 222164
rect 558564 221921 558592 222158
rect 558550 221912 558606 221921
rect 558550 221847 558606 221856
rect 558736 220720 558788 220726
rect 558736 220662 558788 220668
rect 558552 220652 558604 220658
rect 558552 220594 558604 220600
rect 558000 220244 558052 220250
rect 558000 220186 558052 220192
rect 558368 220244 558420 220250
rect 558368 220186 558420 220192
rect 558380 220130 558408 220186
rect 558196 220102 558408 220130
rect 557356 219020 557408 219026
rect 557356 218962 557408 218968
rect 557368 217274 557396 218962
rect 558196 217274 558224 220102
rect 558368 220040 558420 220046
rect 558368 219982 558420 219988
rect 558380 219638 558408 219982
rect 558564 219638 558592 220594
rect 558748 220561 558776 220662
rect 558734 220552 558790 220561
rect 558734 220487 558790 220496
rect 558368 219632 558420 219638
rect 558368 219574 558420 219580
rect 558552 219632 558604 219638
rect 558552 219574 558604 219580
rect 557368 217246 557442 217274
rect 558196 217246 558270 217274
rect 555712 217110 555786 217138
rect 556540 217110 556614 217138
rect 555758 216988 555786 217110
rect 556586 216988 556614 217110
rect 557414 216988 557442 217246
rect 558242 216988 558270 217246
rect 559024 217138 559052 223110
rect 559576 221950 559604 229842
rect 560944 227180 560996 227186
rect 560944 227122 560996 227128
rect 560956 224954 560984 227122
rect 560772 224926 560984 224954
rect 559932 222216 559984 222222
rect 559932 222158 559984 222164
rect 559380 221944 559432 221950
rect 559378 221912 559380 221921
rect 559564 221944 559616 221950
rect 559432 221912 559434 221921
rect 559564 221886 559616 221892
rect 559378 221847 559434 221856
rect 559944 217138 559972 222158
rect 560772 217569 560800 224926
rect 561678 224904 561734 224913
rect 561678 224839 561734 224848
rect 561692 223174 561720 224839
rect 562336 224806 562364 252554
rect 563716 225010 563744 259422
rect 568120 230104 568172 230110
rect 568120 230046 568172 230052
rect 566832 229764 566884 229770
rect 566832 229706 566884 229712
rect 565636 228404 565688 228410
rect 565636 228346 565688 228352
rect 563980 225752 564032 225758
rect 563980 225694 564032 225700
rect 563704 225004 563756 225010
rect 563704 224946 563756 224952
rect 562140 224800 562192 224806
rect 562138 224768 562140 224777
rect 562324 224800 562376 224806
rect 562192 224768 562194 224777
rect 562324 224742 562376 224748
rect 563794 224768 563850 224777
rect 562138 224703 562194 224712
rect 563794 224703 563850 224712
rect 561680 223168 561732 223174
rect 561680 223110 561732 223116
rect 562416 223168 562468 223174
rect 562416 223110 562468 223116
rect 561494 221912 561550 221921
rect 561494 221847 561550 221856
rect 560758 217560 560814 217569
rect 560758 217495 560814 217504
rect 560772 217274 560800 217495
rect 559024 217110 559098 217138
rect 559070 216988 559098 217110
rect 559898 217110 559972 217138
rect 560726 217246 560800 217274
rect 559898 216988 559926 217110
rect 560726 216988 560754 217246
rect 561508 217138 561536 221847
rect 562428 217138 562456 223110
rect 563808 221785 563836 224703
rect 563794 221776 563850 221785
rect 563794 221711 563850 221720
rect 562968 220720 563020 220726
rect 563152 220720 563204 220726
rect 563020 220668 563054 220674
rect 562968 220662 563054 220668
rect 563152 220662 563204 220668
rect 562980 220646 563054 220662
rect 562874 220552 562930 220561
rect 562874 220487 562930 220496
rect 562888 220250 562916 220487
rect 563026 220266 563054 220646
rect 563164 220402 563192 220662
rect 563334 220552 563390 220561
rect 563334 220487 563390 220496
rect 563164 220386 563238 220402
rect 563348 220386 563376 220487
rect 563164 220380 563250 220386
rect 563164 220374 563198 220380
rect 563198 220322 563250 220328
rect 563336 220380 563388 220386
rect 563336 220322 563388 220328
rect 563026 220250 563100 220266
rect 562876 220244 562928 220250
rect 563026 220244 563112 220250
rect 563026 220238 563060 220244
rect 562876 220186 562928 220192
rect 563060 220186 563112 220192
rect 562704 219422 563284 219450
rect 562704 218890 562732 219422
rect 563256 219298 563284 219422
rect 563060 219292 563112 219298
rect 563060 219234 563112 219240
rect 563244 219292 563296 219298
rect 563244 219234 563296 219240
rect 562874 219192 562930 219201
rect 562874 219127 562876 219136
rect 562928 219127 562930 219136
rect 562876 219098 562928 219104
rect 562692 218884 562744 218890
rect 562692 218826 562744 218832
rect 563072 218657 563100 219234
rect 563518 219192 563574 219201
rect 563518 219127 563520 219136
rect 563572 219127 563574 219136
rect 563520 219098 563572 219104
rect 563426 218920 563482 218929
rect 563348 218864 563426 218872
rect 563348 218855 563482 218864
rect 563612 218884 563664 218890
rect 563348 218844 563468 218855
rect 563348 218754 563376 218844
rect 563612 218826 563664 218832
rect 563336 218748 563388 218754
rect 563336 218690 563388 218696
rect 563058 218648 563114 218657
rect 563058 218583 563114 218592
rect 563198 218612 563250 218618
rect 563624 218600 563652 218826
rect 563250 218572 563652 218600
rect 563198 218554 563250 218560
rect 562876 218204 562928 218210
rect 562876 218146 562928 218152
rect 562888 217841 562916 218146
rect 563612 218000 563664 218006
rect 563072 217948 563612 217954
rect 563072 217942 563664 217948
rect 563072 217926 563652 217942
rect 562874 217832 562930 217841
rect 562874 217767 562930 217776
rect 563072 217682 563100 217926
rect 563026 217654 563100 217682
rect 563026 217326 563054 217654
rect 563150 217560 563206 217569
rect 563150 217495 563206 217504
rect 563164 217326 563192 217495
rect 563014 217320 563066 217326
rect 563014 217262 563066 217268
rect 563152 217320 563204 217326
rect 563152 217262 563204 217268
rect 563808 217138 563836 221711
rect 563992 217274 564020 225694
rect 564624 223304 564676 223310
rect 564624 223246 564676 223252
rect 564636 222494 564664 223246
rect 564808 223168 564860 223174
rect 564808 223110 564860 223116
rect 564820 222494 564848 223110
rect 564624 222488 564676 222494
rect 564624 222430 564676 222436
rect 564808 222488 564860 222494
rect 564808 222430 564860 222436
rect 564808 221944 564860 221950
rect 564808 221886 564860 221892
rect 564820 218929 564848 221886
rect 565648 220697 565676 228346
rect 566844 223514 566872 229706
rect 567016 225140 567068 225146
rect 567016 225082 567068 225088
rect 567028 224806 567056 225082
rect 567016 224800 567068 224806
rect 567016 224742 567068 224748
rect 567844 224800 567896 224806
rect 567844 224742 567896 224748
rect 567856 223650 567884 224742
rect 567844 223644 567896 223650
rect 567844 223586 567896 223592
rect 566832 223508 566884 223514
rect 566832 223450 566884 223456
rect 566844 220726 566872 223450
rect 566464 220720 566516 220726
rect 565634 220688 565690 220697
rect 566464 220662 566516 220668
rect 566832 220720 566884 220726
rect 566832 220662 566884 220668
rect 567292 220720 567344 220726
rect 567292 220662 567344 220668
rect 565634 220623 565690 220632
rect 564162 218920 564218 218929
rect 564162 218855 564218 218864
rect 564806 218920 564862 218929
rect 564806 218855 564862 218864
rect 564176 218754 564204 218855
rect 564164 218748 564216 218754
rect 564164 218690 564216 218696
rect 563992 217246 564066 217274
rect 561508 217110 561582 217138
rect 561554 216988 561582 217110
rect 562382 217110 562456 217138
rect 563210 217110 563836 217138
rect 562382 216988 562410 217110
rect 563210 216988 563238 217110
rect 564038 216988 564066 217246
rect 564820 217138 564848 218855
rect 565648 217274 565676 220623
rect 565648 217246 565722 217274
rect 564820 217110 564894 217138
rect 564866 216988 564894 217110
rect 565694 216988 565722 217246
rect 566476 217138 566504 220662
rect 567304 217274 567332 220662
rect 568132 217274 568160 230046
rect 568592 220658 568620 260850
rect 570616 234598 570644 261462
rect 596824 245676 596876 245682
rect 596824 245618 596876 245624
rect 576124 242208 576176 242214
rect 576124 242150 576176 242156
rect 576136 238746 576164 242150
rect 577504 240168 577556 240174
rect 577504 240110 577556 240116
rect 576124 238740 576176 238746
rect 576124 238682 576176 238688
rect 570604 234592 570656 234598
rect 570604 234534 570656 234540
rect 570604 228540 570656 228546
rect 570604 228482 570656 228488
rect 568948 224936 569000 224942
rect 568948 224878 569000 224884
rect 568580 220652 568632 220658
rect 568580 220594 568632 220600
rect 568304 218544 568356 218550
rect 568304 218486 568356 218492
rect 568316 217841 568344 218486
rect 568302 217832 568358 217841
rect 568302 217767 568358 217776
rect 567304 217246 567378 217274
rect 568132 217246 568206 217274
rect 566476 217110 566550 217138
rect 566522 216988 566550 217110
rect 567350 216988 567378 217246
rect 568178 216988 568206 217246
rect 568960 217138 568988 224878
rect 569958 220688 570014 220697
rect 569776 220652 569828 220658
rect 569958 220623 569960 220632
rect 569776 220594 569828 220600
rect 570012 220623 570014 220632
rect 569960 220594 570012 220600
rect 569788 217138 569816 220594
rect 570616 217274 570644 228482
rect 572260 225888 572312 225894
rect 572260 225830 572312 225836
rect 571432 225140 571484 225146
rect 571432 225082 571484 225088
rect 571444 217274 571472 225082
rect 572272 220561 572300 225830
rect 572626 221776 572682 221785
rect 572626 221711 572682 221720
rect 572640 220658 572668 221711
rect 572444 220652 572496 220658
rect 572444 220594 572496 220600
rect 572628 220652 572680 220658
rect 572628 220594 572680 220600
rect 572258 220552 572314 220561
rect 572258 220487 572314 220496
rect 572456 220130 572484 220594
rect 572456 220114 572714 220130
rect 572456 220108 572726 220114
rect 572456 220102 572674 220108
rect 572674 220050 572726 220056
rect 572536 220040 572588 220046
rect 572536 219982 572588 219988
rect 572548 219450 572576 219982
rect 572548 219422 572714 219450
rect 572686 219366 572714 219422
rect 572674 219360 572726 219366
rect 572674 219302 572726 219308
rect 574376 219224 574428 219230
rect 572074 219192 572130 219201
rect 574376 219166 574428 219172
rect 574558 219192 574614 219201
rect 572074 219127 572076 219136
rect 572128 219127 572130 219136
rect 572076 219098 572128 219104
rect 572076 218884 572128 218890
rect 572076 218826 572128 218832
rect 572088 218770 572116 218826
rect 572088 218742 572852 218770
rect 572824 218618 572852 218742
rect 572812 218612 572864 218618
rect 572812 218554 572864 218560
rect 572444 218544 572496 218550
rect 572496 218492 573036 218498
rect 572444 218486 573036 218492
rect 572456 218470 573036 218486
rect 572076 218408 572128 218414
rect 572076 218350 572128 218356
rect 571892 218000 571944 218006
rect 571892 217942 571944 217948
rect 571904 217682 571932 217942
rect 572088 217841 572116 218350
rect 572812 218340 572864 218346
rect 572812 218282 572864 218288
rect 572536 218272 572588 218278
rect 572824 218226 572852 218282
rect 572588 218220 572852 218226
rect 572536 218214 572852 218220
rect 572548 218198 572852 218214
rect 573008 218210 573036 218470
rect 572996 218204 573048 218210
rect 572996 218146 573048 218152
rect 572074 217832 572130 217841
rect 572074 217767 572130 217776
rect 571904 217654 572760 217682
rect 572258 217560 572314 217569
rect 572258 217495 572314 217504
rect 570616 217246 570690 217274
rect 571444 217246 571518 217274
rect 568960 217110 569034 217138
rect 569788 217110 569862 217138
rect 569006 216988 569034 217110
rect 569834 216988 569862 217110
rect 570662 216988 570690 217246
rect 571490 216988 571518 217246
rect 572272 217138 572300 217495
rect 572732 217326 572760 217654
rect 572902 217560 572958 217569
rect 572902 217495 572958 217504
rect 574190 217560 574246 217569
rect 574190 217495 574246 217504
rect 572536 217320 572588 217326
rect 572536 217262 572588 217268
rect 572720 217320 572772 217326
rect 572720 217262 572772 217268
rect 572548 217138 572576 217262
rect 572916 217138 572944 217495
rect 572272 217110 572346 217138
rect 572548 217110 572944 217138
rect 572318 216988 572346 217110
rect 574204 217054 574232 217495
rect 574192 217048 574244 217054
rect 574192 216990 574244 216996
rect 53286 215112 53342 215121
rect 53286 215047 53342 215056
rect 574388 214606 574416 219166
rect 574558 219127 574614 219136
rect 574572 214742 574600 219127
rect 574742 218920 574798 218929
rect 574742 218855 574744 218864
rect 574796 218855 574798 218864
rect 574744 218826 574796 218832
rect 574742 218648 574798 218657
rect 574742 218583 574798 218592
rect 574756 214878 574784 218583
rect 574928 218476 574980 218482
rect 574928 218418 574980 218424
rect 574940 217841 574968 218418
rect 574926 217832 574982 217841
rect 574926 217767 574982 217776
rect 575478 216744 575534 216753
rect 575478 216679 575534 216688
rect 574744 214872 574796 214878
rect 574744 214814 574796 214820
rect 574560 214736 574612 214742
rect 574560 214678 574612 214684
rect 574376 214600 574428 214606
rect 574376 214542 574428 214548
rect 575492 213246 575520 216679
rect 575480 213240 575532 213246
rect 575480 213182 575532 213188
rect 51906 179344 51962 179353
rect 51906 179279 51962 179288
rect 577516 99142 577544 240110
rect 593972 223032 594024 223038
rect 593972 222974 594024 222980
rect 589108 219966 589504 219994
rect 589108 219502 589136 219966
rect 589476 219910 589504 219966
rect 589280 219904 589332 219910
rect 589280 219846 589332 219852
rect 589464 219904 589516 219910
rect 589464 219846 589516 219852
rect 589096 219496 589148 219502
rect 589096 219438 589148 219444
rect 589292 219230 589320 219846
rect 589280 219224 589332 219230
rect 589280 219166 589332 219172
rect 578882 214024 578938 214033
rect 578882 213959 578938 213968
rect 578514 211712 578570 211721
rect 578514 211647 578570 211656
rect 578528 211206 578556 211647
rect 578516 211200 578568 211206
rect 578516 211142 578568 211148
rect 578896 208350 578924 213959
rect 592684 212696 592736 212702
rect 592684 212638 592736 212644
rect 591304 212560 591356 212566
rect 591304 212502 591356 212508
rect 580908 211200 580960 211206
rect 580908 211142 580960 211148
rect 579528 209840 579580 209846
rect 579526 209808 579528 209817
rect 579580 209808 579582 209817
rect 579526 209743 579582 209752
rect 578884 208344 578936 208350
rect 578884 208286 578936 208292
rect 579526 207496 579582 207505
rect 579582 207454 579752 207482
rect 579526 207431 579582 207440
rect 579526 205864 579582 205873
rect 579526 205799 579528 205808
rect 579580 205799 579582 205808
rect 579528 205770 579580 205776
rect 579724 204270 579752 207454
rect 580920 206922 580948 211142
rect 582288 209840 582340 209846
rect 582288 209782 582340 209788
rect 581644 208616 581696 208622
rect 581644 208558 581696 208564
rect 580908 206916 580960 206922
rect 580908 206858 580960 206864
rect 581000 205828 581052 205834
rect 581000 205770 581052 205776
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578330 203280 578386 203289
rect 578330 203215 578386 203224
rect 578344 202910 578372 203215
rect 578332 202904 578384 202910
rect 578332 202846 578384 202852
rect 580264 202904 580316 202910
rect 580264 202846 580316 202852
rect 578790 200832 578846 200841
rect 578790 200767 578846 200776
rect 578804 200190 578832 200767
rect 578792 200184 578844 200190
rect 578792 200126 578844 200132
rect 580276 200054 580304 202846
rect 581012 202842 581040 205770
rect 581000 202836 581052 202842
rect 581000 202778 581052 202784
rect 580264 200048 580316 200054
rect 580264 199990 580316 199996
rect 579526 198928 579582 198937
rect 579526 198863 579582 198872
rect 579540 198762 579568 198863
rect 579528 198756 579580 198762
rect 579528 198698 579580 198704
rect 578514 196480 578570 196489
rect 578514 196415 578570 196424
rect 578528 196042 578556 196415
rect 578516 196036 578568 196042
rect 578516 195978 578568 195984
rect 579526 194984 579582 194993
rect 579526 194919 579582 194928
rect 579540 194614 579568 194919
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 579526 192264 579582 192273
rect 579526 192199 579582 192208
rect 579540 191894 579568 192199
rect 579528 191888 579580 191894
rect 579528 191830 579580 191836
rect 579526 190768 579582 190777
rect 579526 190703 579582 190712
rect 579540 190534 579568 190703
rect 579528 190528 579580 190534
rect 579528 190470 579580 190476
rect 579526 188048 579582 188057
rect 579526 187983 579582 187992
rect 579540 187746 579568 187983
rect 579528 187740 579580 187746
rect 579528 187682 579580 187688
rect 579528 186312 579580 186318
rect 579526 186280 579528 186289
rect 579580 186280 579582 186289
rect 579526 186215 579582 186224
rect 579528 184884 579580 184890
rect 579528 184826 579580 184832
rect 579540 184385 579568 184826
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 579528 182164 579580 182170
rect 579528 182106 579580 182112
rect 579540 181937 579568 182106
rect 579526 181928 579582 181937
rect 579526 181863 579582 181872
rect 578792 180804 578844 180810
rect 578792 180746 578844 180752
rect 578804 180169 578832 180746
rect 578790 180160 578846 180169
rect 578790 180095 578846 180104
rect 578792 178084 578844 178090
rect 578792 178026 578844 178032
rect 578804 175137 578832 178026
rect 579528 177948 579580 177954
rect 579528 177890 579580 177896
rect 579540 177721 579568 177890
rect 579526 177712 579582 177721
rect 579526 177647 579582 177656
rect 579988 175296 580040 175302
rect 579988 175238 580040 175244
rect 578790 175128 578846 175137
rect 578790 175063 578846 175072
rect 578424 174548 578476 174554
rect 578424 174490 578476 174496
rect 578436 173505 578464 174490
rect 578422 173496 578478 173505
rect 578422 173431 578478 173440
rect 580000 172922 580028 175238
rect 578240 172916 578292 172922
rect 578240 172858 578292 172864
rect 579988 172916 580040 172922
rect 579988 172858 580040 172864
rect 578252 171057 578280 172858
rect 580908 172576 580960 172582
rect 580908 172518 580960 172524
rect 580264 171148 580316 171154
rect 580264 171090 580316 171096
rect 578238 171048 578294 171057
rect 578238 170983 578294 170992
rect 578700 169788 578752 169794
rect 578700 169730 578752 169736
rect 578712 169289 578740 169730
rect 578698 169280 578754 169289
rect 578698 169215 578754 169224
rect 580276 167346 580304 171090
rect 580920 169794 580948 172518
rect 580908 169788 580960 169794
rect 580908 169730 580960 169736
rect 578240 167340 578292 167346
rect 578240 167282 578292 167288
rect 580264 167340 580316 167346
rect 580264 167282 580316 167288
rect 578252 166977 578280 167282
rect 579988 167068 580040 167074
rect 579988 167010 580040 167016
rect 578238 166968 578294 166977
rect 578238 166903 578294 166912
rect 579528 166320 579580 166326
rect 579528 166262 579580 166268
rect 579344 165232 579396 165238
rect 579344 165174 579396 165180
rect 578240 163668 578292 163674
rect 578240 163610 578292 163616
rect 578252 159905 578280 163610
rect 579356 162761 579384 165174
rect 579540 164529 579568 166262
rect 579526 164520 579582 164529
rect 579526 164455 579582 164464
rect 580000 163674 580028 167010
rect 579988 163668 580040 163674
rect 579988 163610 580040 163616
rect 580908 162920 580960 162926
rect 580908 162862 580960 162868
rect 579342 162752 579398 162761
rect 578424 162716 578476 162722
rect 579342 162687 579398 162696
rect 578424 162658 578476 162664
rect 578238 159896 578294 159905
rect 578238 159831 578294 159840
rect 578436 158409 578464 162658
rect 580540 161492 580592 161498
rect 580540 161434 580592 161440
rect 578884 158772 578936 158778
rect 578884 158714 578936 158720
rect 578422 158400 578478 158409
rect 578422 158335 578478 158344
rect 578896 155961 578924 158714
rect 578882 155952 578938 155961
rect 578882 155887 578938 155896
rect 580552 154698 580580 161434
rect 580724 160132 580776 160138
rect 580724 160074 580776 160080
rect 578332 154692 578384 154698
rect 578332 154634 578384 154640
rect 580540 154692 580592 154698
rect 580540 154634 580592 154640
rect 578344 154057 578372 154634
rect 578330 154048 578386 154057
rect 578330 153983 578386 153992
rect 580736 152794 580764 160074
rect 580920 158778 580948 162862
rect 580908 158772 580960 158778
rect 580908 158714 580960 158720
rect 578240 152788 578292 152794
rect 578240 152730 578292 152736
rect 580724 152788 580776 152794
rect 580724 152730 580776 152736
rect 578252 151745 578280 152730
rect 580264 151836 580316 151842
rect 580264 151778 580316 151784
rect 578238 151736 578294 151745
rect 578238 151671 578294 151680
rect 578884 150612 578936 150618
rect 578884 150554 578936 150560
rect 578896 149705 578924 150554
rect 578882 149696 578938 149705
rect 578882 149631 578938 149640
rect 579528 148368 579580 148374
rect 579528 148310 579580 148316
rect 579540 147529 579568 148310
rect 579526 147520 579582 147529
rect 579526 147455 579582 147464
rect 578884 146328 578936 146334
rect 578884 146270 578936 146276
rect 578608 140752 578660 140758
rect 578608 140694 578660 140700
rect 578620 140593 578648 140694
rect 578606 140584 578662 140593
rect 578606 140519 578662 140528
rect 578608 139324 578660 139330
rect 578608 139266 578660 139272
rect 578620 138825 578648 139266
rect 578606 138816 578662 138825
rect 578606 138751 578662 138760
rect 578896 136649 578924 146270
rect 579252 144696 579304 144702
rect 579250 144664 579252 144673
rect 579304 144664 579306 144673
rect 579250 144599 579306 144608
rect 579528 143472 579580 143478
rect 579528 143414 579580 143420
rect 579540 143041 579568 143414
rect 579526 143032 579582 143041
rect 579526 142967 579582 142976
rect 580276 140758 580304 151778
rect 580448 140820 580500 140826
rect 580448 140762 580500 140768
rect 580264 140752 580316 140758
rect 580264 140694 580316 140700
rect 579528 138712 579580 138718
rect 579528 138654 579580 138660
rect 579068 137352 579120 137358
rect 579068 137294 579120 137300
rect 578882 136640 578938 136649
rect 578882 136575 578938 136584
rect 579080 132297 579108 137294
rect 579540 134473 579568 138654
rect 580264 134564 580316 134570
rect 580264 134506 580316 134512
rect 579526 134464 579582 134473
rect 579526 134399 579582 134408
rect 579066 132288 579122 132297
rect 579066 132223 579122 132232
rect 578884 131164 578936 131170
rect 578884 131106 578936 131112
rect 578896 129713 578924 131106
rect 578882 129704 578938 129713
rect 578882 129639 578938 129648
rect 579528 129056 579580 129062
rect 579528 128998 579580 129004
rect 579540 127945 579568 128998
rect 579526 127936 579582 127945
rect 579526 127871 579582 127880
rect 579068 127016 579120 127022
rect 579068 126958 579120 126964
rect 578332 125656 578384 125662
rect 578332 125598 578384 125604
rect 578344 125361 578372 125598
rect 578330 125352 578386 125361
rect 578330 125287 578386 125296
rect 578424 123616 578476 123622
rect 578422 123584 578424 123593
rect 578476 123584 578478 123593
rect 578422 123519 578478 123528
rect 578884 122188 578936 122194
rect 578884 122130 578936 122136
rect 578896 121417 578924 122130
rect 578882 121408 578938 121417
rect 578882 121343 578938 121352
rect 578516 118448 578568 118454
rect 578514 118416 578516 118425
rect 578568 118416 578570 118425
rect 578514 118351 578570 118360
rect 578332 108724 578384 108730
rect 578332 108666 578384 108672
rect 578344 108361 578372 108666
rect 578330 108352 578386 108361
rect 578330 108287 578386 108296
rect 578884 107636 578936 107642
rect 578884 107578 578936 107584
rect 578608 99272 578660 99278
rect 578606 99240 578608 99249
rect 578660 99240 578662 99249
rect 578606 99175 578662 99184
rect 577504 99136 577556 99142
rect 577504 99078 577556 99084
rect 578332 97980 578384 97986
rect 578332 97922 578384 97928
rect 578344 97481 578372 97922
rect 578330 97472 578386 97481
rect 578330 97407 578386 97416
rect 578516 93492 578568 93498
rect 578516 93434 578568 93440
rect 578528 93129 578556 93434
rect 578514 93120 578570 93129
rect 578514 93055 578570 93064
rect 578896 80073 578924 107578
rect 579080 105913 579108 126958
rect 580276 118454 580304 134506
rect 580460 125662 580488 140762
rect 580448 125656 580500 125662
rect 580448 125598 580500 125604
rect 580448 124228 580500 124234
rect 580448 124170 580500 124176
rect 580264 118448 580316 118454
rect 580264 118390 580316 118396
rect 579528 116952 579580 116958
rect 579526 116920 579528 116929
rect 579580 116920 579582 116929
rect 579526 116855 579582 116864
rect 579252 114504 579304 114510
rect 579250 114472 579252 114481
rect 579304 114472 579306 114481
rect 579250 114407 579306 114416
rect 579528 112872 579580 112878
rect 579528 112814 579580 112820
rect 579540 112577 579568 112814
rect 579526 112568 579582 112577
rect 579526 112503 579582 112512
rect 579344 110152 579396 110158
rect 579342 110120 579344 110129
rect 579396 110120 579398 110129
rect 579342 110055 579398 110064
rect 579066 105904 579122 105913
rect 579066 105839 579122 105848
rect 580264 104916 580316 104922
rect 580264 104858 580316 104864
rect 579528 103488 579580 103494
rect 579528 103430 579580 103436
rect 579540 103329 579568 103430
rect 579526 103320 579582 103329
rect 579526 103255 579582 103264
rect 579528 101856 579580 101862
rect 579528 101798 579580 101804
rect 579540 101697 579568 101798
rect 579526 101688 579582 101697
rect 579526 101623 579582 101632
rect 579068 99408 579120 99414
rect 579068 99350 579120 99356
rect 579080 90953 579108 99350
rect 579528 95056 579580 95062
rect 579526 95024 579528 95033
rect 579580 95024 579582 95033
rect 579526 94959 579582 94968
rect 579344 91112 579396 91118
rect 579344 91054 579396 91060
rect 579066 90944 579122 90953
rect 579066 90879 579122 90888
rect 579356 86465 579384 91054
rect 579528 88120 579580 88126
rect 579526 88088 579528 88097
rect 579580 88088 579582 88097
rect 579526 88023 579582 88032
rect 579342 86456 579398 86465
rect 579342 86391 579398 86400
rect 579160 84176 579212 84182
rect 579160 84118 579212 84124
rect 579172 84017 579200 84118
rect 579158 84008 579214 84017
rect 579158 83943 579214 83952
rect 579068 82408 579120 82414
rect 579068 82350 579120 82356
rect 579080 82249 579108 82350
rect 579066 82240 579122 82249
rect 579066 82175 579122 82184
rect 579528 82136 579580 82142
rect 579528 82078 579580 82084
rect 578882 80064 578938 80073
rect 578882 79999 578938 80008
rect 579068 79348 579120 79354
rect 579068 79290 579120 79296
rect 578240 75880 578292 75886
rect 578240 75822 578292 75828
rect 578252 75585 578280 75822
rect 578238 75576 578294 75585
rect 578238 75511 578294 75520
rect 579080 73137 579108 79290
rect 579540 77897 579568 82078
rect 579526 77888 579582 77897
rect 579526 77823 579582 77832
rect 580276 75886 580304 104858
rect 580460 99278 580488 124170
rect 580632 122052 580684 122058
rect 580632 121994 580684 122000
rect 580644 108730 580672 121994
rect 581656 114510 581684 208558
rect 582300 205562 582328 209782
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208049 589504 208286
rect 589462 208040 589518 208049
rect 589462 207975 589518 207984
rect 589464 206916 589516 206922
rect 589464 206858 589516 206864
rect 589476 206417 589504 206858
rect 589462 206408 589518 206417
rect 589462 206343 589518 206352
rect 582288 205556 582340 205562
rect 582288 205498 582340 205504
rect 589464 205556 589516 205562
rect 589464 205498 589516 205504
rect 589476 204785 589504 205498
rect 589462 204776 589518 204785
rect 589462 204711 589518 204720
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203153 589504 204206
rect 589462 203144 589518 203153
rect 589462 203079 589518 203088
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 201521 589504 202778
rect 589462 201512 589518 201521
rect 589462 201447 589518 201456
rect 590384 200184 590436 200190
rect 590384 200126 590436 200132
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 589464 198756 589516 198762
rect 589464 198698 589516 198704
rect 589476 196625 589504 198698
rect 590396 198257 590424 200126
rect 590382 198248 590438 198257
rect 590382 198183 590438 198192
rect 589462 196616 589518 196625
rect 589462 196551 589518 196560
rect 589280 196036 589332 196042
rect 589280 195978 589332 195984
rect 589292 194993 589320 195978
rect 589278 194984 589334 194993
rect 589278 194919 589334 194928
rect 589464 194608 589516 194614
rect 589464 194550 589516 194556
rect 589476 193361 589504 194550
rect 589462 193352 589518 193361
rect 589462 193287 589518 193296
rect 589464 191888 589516 191894
rect 589464 191830 589516 191836
rect 589476 191729 589504 191830
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 590568 190528 590620 190534
rect 590568 190470 590620 190476
rect 590580 190097 590608 190470
rect 590566 190088 590622 190097
rect 590566 190023 590622 190032
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 589464 187740 589516 187746
rect 589464 187682 589516 187688
rect 589476 186833 589504 187682
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 589660 186318 589688 188391
rect 589648 186312 589700 186318
rect 589648 186254 589700 186260
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184890 589504 185127
rect 589464 184884 589516 184890
rect 589464 184826 589516 184832
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182170 589504 183495
rect 589464 182164 589516 182170
rect 589464 182106 589516 182112
rect 590566 181928 590622 181937
rect 590566 181863 590622 181872
rect 590580 180810 590608 181863
rect 590568 180804 590620 180810
rect 590568 180746 590620 180752
rect 589646 180296 589702 180305
rect 589646 180231 589702 180240
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 589660 177954 589688 180231
rect 589648 177948 589700 177954
rect 589648 177890 589700 177896
rect 589646 177032 589702 177041
rect 589646 176967 589702 176976
rect 589462 175400 589518 175409
rect 589462 175335 589464 175344
rect 589516 175335 589518 175344
rect 589464 175306 589516 175312
rect 589660 174554 589688 176967
rect 589648 174548 589700 174554
rect 589648 174490 589700 174496
rect 589462 173768 589518 173777
rect 589462 173703 589518 173712
rect 589476 172582 589504 173703
rect 589464 172576 589516 172582
rect 589464 172518 589516 172524
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 589646 170504 589702 170513
rect 589646 170439 589702 170448
rect 589462 168872 589518 168881
rect 589462 168807 589518 168816
rect 589476 168434 589504 168807
rect 582380 168428 582432 168434
rect 582380 168370 582432 168376
rect 589464 168428 589516 168434
rect 589464 168370 589516 168376
rect 582392 165238 582420 168370
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 589660 166326 589688 170439
rect 589648 166320 589700 166326
rect 589648 166262 589700 166268
rect 589462 165608 589518 165617
rect 589462 165543 589518 165552
rect 582380 165232 582432 165238
rect 582380 165174 582432 165180
rect 589476 164286 589504 165543
rect 582472 164280 582524 164286
rect 582472 164222 582524 164228
rect 589464 164280 589516 164286
rect 589464 164222 589516 164228
rect 582484 162722 582512 164222
rect 589462 163976 589518 163985
rect 589462 163911 589518 163920
rect 589476 162926 589504 163911
rect 589464 162920 589516 162926
rect 589464 162862 589516 162868
rect 582472 162716 582524 162722
rect 582472 162658 582524 162664
rect 589462 162344 589518 162353
rect 589462 162279 589518 162288
rect 589476 161498 589504 162279
rect 589464 161492 589516 161498
rect 589464 161434 589516 161440
rect 589462 160712 589518 160721
rect 589462 160647 589518 160656
rect 589476 160138 589504 160647
rect 589464 160132 589516 160138
rect 589464 160074 589516 160080
rect 589462 159080 589518 159089
rect 589462 159015 589518 159024
rect 589476 158778 589504 159015
rect 585784 158772 585836 158778
rect 585784 158714 585836 158720
rect 589464 158772 589516 158778
rect 589464 158714 589516 158720
rect 584404 154624 584456 154630
rect 584404 154566 584456 154572
rect 583024 153264 583076 153270
rect 583024 153206 583076 153212
rect 583036 143478 583064 153206
rect 584416 144702 584444 154566
rect 585796 150618 585824 158714
rect 589278 157448 589334 157457
rect 587164 157412 587216 157418
rect 589278 157383 589280 157392
rect 587164 157354 587216 157360
rect 589332 157383 589334 157392
rect 589280 157354 589332 157360
rect 585784 150612 585836 150618
rect 585784 150554 585836 150560
rect 585140 149116 585192 149122
rect 585140 149058 585192 149064
rect 585152 146334 585180 149058
rect 587176 148374 587204 157354
rect 589462 155816 589518 155825
rect 589462 155751 589518 155760
rect 589476 154630 589504 155751
rect 589464 154624 589516 154630
rect 589464 154566 589516 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589462 152552 589518 152561
rect 589462 152487 589518 152496
rect 589476 151842 589504 152487
rect 589464 151836 589516 151842
rect 589464 151778 589516 151784
rect 590014 150920 590070 150929
rect 590014 150855 590070 150864
rect 589462 149288 589518 149297
rect 589462 149223 589518 149232
rect 589476 149122 589504 149223
rect 589464 149116 589516 149122
rect 589464 149058 589516 149064
rect 587164 148368 587216 148374
rect 587164 148310 587216 148316
rect 588542 147656 588598 147665
rect 588542 147591 588598 147600
rect 585140 146328 585192 146334
rect 585140 146270 585192 146276
rect 584772 144968 584824 144974
rect 584772 144910 584824 144916
rect 584404 144696 584456 144702
rect 584404 144638 584456 144644
rect 583024 143472 583076 143478
rect 583024 143414 583076 143420
rect 583024 139460 583076 139466
rect 583024 139402 583076 139408
rect 581828 131300 581880 131306
rect 581828 131242 581880 131248
rect 581644 114504 581696 114510
rect 581644 114446 581696 114452
rect 581644 110492 581696 110498
rect 581644 110434 581696 110440
rect 580632 108724 580684 108730
rect 580632 108666 580684 108672
rect 580448 99272 580500 99278
rect 580448 99214 580500 99220
rect 581656 84182 581684 110434
rect 581840 110158 581868 131242
rect 583036 123622 583064 139402
rect 584784 137358 584812 144910
rect 585968 143608 586020 143614
rect 585968 143550 586020 143556
rect 584772 137352 584824 137358
rect 584772 137294 584824 137300
rect 584588 136672 584640 136678
rect 584588 136614 584640 136620
rect 583208 129192 583260 129198
rect 583208 129134 583260 129140
rect 583024 123616 583076 123622
rect 583024 123558 583076 123564
rect 583220 116958 583248 129134
rect 584404 122868 584456 122874
rect 584404 122810 584456 122816
rect 583208 116952 583260 116958
rect 583208 116894 583260 116900
rect 583208 115252 583260 115258
rect 583208 115194 583260 115200
rect 583024 113212 583076 113218
rect 583024 113154 583076 113160
rect 581828 110152 581880 110158
rect 581828 110094 581880 110100
rect 581644 84176 581696 84182
rect 581644 84118 581696 84124
rect 583036 82414 583064 113154
rect 583220 95062 583248 115194
rect 584416 101862 584444 122810
rect 584600 122194 584628 136614
rect 585784 132524 585836 132530
rect 585784 132466 585836 132472
rect 584588 122188 584640 122194
rect 584588 122130 584640 122136
rect 585796 112878 585824 132466
rect 585980 131170 586008 143550
rect 587164 142452 587216 142458
rect 587164 142394 587216 142400
rect 585968 131164 586020 131170
rect 585968 131106 586020 131112
rect 587176 129062 587204 142394
rect 588556 138718 588584 147591
rect 589462 146024 589518 146033
rect 589462 145959 589518 145968
rect 589476 144974 589504 145959
rect 589464 144968 589516 144974
rect 589464 144910 589516 144916
rect 589462 144392 589518 144401
rect 589462 144327 589518 144336
rect 589476 143614 589504 144327
rect 589464 143608 589516 143614
rect 589464 143550 589516 143556
rect 589830 142760 589886 142769
rect 589830 142695 589886 142704
rect 589844 142458 589872 142695
rect 589832 142452 589884 142458
rect 589832 142394 589884 142400
rect 590028 142154 590056 150855
rect 589936 142126 590056 142154
rect 589462 141128 589518 141137
rect 589462 141063 589518 141072
rect 589476 140826 589504 141063
rect 589464 140820 589516 140826
rect 589464 140762 589516 140768
rect 589462 139496 589518 139505
rect 589462 139431 589464 139440
rect 589516 139431 589518 139440
rect 589464 139402 589516 139408
rect 589936 139330 589964 142126
rect 589924 139324 589976 139330
rect 589924 139266 589976 139272
rect 588544 138712 588596 138718
rect 588544 138654 588596 138660
rect 589462 137864 589518 137873
rect 589462 137799 589518 137808
rect 589476 136678 589504 137799
rect 589464 136672 589516 136678
rect 589464 136614 589516 136620
rect 589462 136232 589518 136241
rect 589462 136167 589518 136176
rect 589476 134570 589504 136167
rect 590382 134600 590438 134609
rect 589464 134564 589516 134570
rect 590382 134535 590438 134544
rect 589464 134506 589516 134512
rect 589462 132968 589518 132977
rect 589462 132903 589518 132912
rect 589476 132530 589504 132903
rect 589464 132524 589516 132530
rect 589464 132466 589516 132472
rect 589462 131336 589518 131345
rect 589462 131271 589464 131280
rect 589516 131271 589518 131280
rect 589464 131242 589516 131248
rect 588542 129704 588598 129713
rect 588542 129639 588598 129648
rect 587164 129056 587216 129062
rect 587164 128998 587216 129004
rect 587348 118720 587400 118726
rect 587348 118662 587400 118668
rect 586152 116000 586204 116006
rect 586152 115942 586204 115948
rect 585784 112872 585836 112878
rect 585784 112814 585836 112820
rect 585968 112464 586020 112470
rect 585968 112406 586020 112412
rect 584588 109064 584640 109070
rect 584588 109006 584640 109012
rect 584404 101856 584456 101862
rect 584404 101798 584456 101804
rect 584404 100156 584456 100162
rect 584404 100098 584456 100104
rect 583208 95056 583260 95062
rect 583208 94998 583260 95004
rect 583024 82408 583076 82414
rect 583024 82350 583076 82356
rect 581642 77888 581698 77897
rect 581642 77823 581698 77832
rect 580264 75880 580316 75886
rect 580264 75822 580316 75828
rect 579066 73128 579122 73137
rect 579066 73063 579122 73072
rect 578884 72480 578936 72486
rect 578884 72422 578936 72428
rect 577504 60036 577556 60042
rect 577504 59978 577556 59984
rect 576124 58676 576176 58682
rect 576124 58618 576176 58624
rect 574928 57248 574980 57254
rect 574928 57190 574980 57196
rect 574560 56024 574612 56030
rect 574560 55966 574612 55972
rect 574572 53990 574600 55966
rect 574744 55888 574796 55894
rect 574744 55830 574796 55836
rect 574756 54126 574784 55830
rect 574744 54120 574796 54126
rect 574744 54062 574796 54068
rect 574560 53984 574612 53990
rect 574560 53926 574612 53932
rect 574940 53854 574968 57190
rect 576136 55049 576164 58618
rect 576122 55040 576178 55049
rect 576122 54975 576178 54984
rect 577516 54233 577544 59978
rect 578896 54505 578924 72422
rect 579068 71392 579120 71398
rect 579068 71334 579120 71340
rect 579080 71233 579108 71334
rect 579066 71224 579122 71233
rect 579066 71159 579122 71168
rect 580264 68332 580316 68338
rect 580264 68274 580316 68280
rect 580276 54777 580304 68274
rect 580262 54768 580318 54777
rect 580262 54703 580318 54712
rect 578882 54496 578938 54505
rect 578882 54431 578938 54440
rect 581656 54262 581684 77823
rect 584416 71398 584444 100098
rect 584600 91118 584628 109006
rect 585980 93498 586008 112406
rect 586164 99414 586192 115942
rect 587164 106344 587216 106350
rect 587164 106286 587216 106292
rect 586152 99408 586204 99414
rect 586152 99350 586204 99356
rect 585968 93492 586020 93498
rect 585968 93434 586020 93440
rect 584588 91112 584640 91118
rect 584588 91054 584640 91060
rect 585140 89004 585192 89010
rect 585140 88946 585192 88952
rect 585152 88126 585180 88946
rect 585140 88120 585192 88126
rect 585140 88062 585192 88068
rect 587176 82142 587204 106286
rect 587360 97986 587388 118662
rect 588556 103494 588584 129639
rect 590396 129198 590424 134535
rect 590384 129192 590436 129198
rect 590384 129134 590436 129140
rect 589462 128072 589518 128081
rect 589462 128007 589518 128016
rect 589476 127022 589504 128007
rect 589464 127016 589516 127022
rect 589464 126958 589516 126964
rect 589922 126440 589978 126449
rect 589922 126375 589978 126384
rect 589462 124808 589518 124817
rect 589462 124743 589518 124752
rect 589476 124234 589504 124743
rect 589464 124228 589516 124234
rect 589464 124170 589516 124176
rect 589462 123176 589518 123185
rect 589462 123111 589518 123120
rect 589476 122874 589504 123111
rect 589464 122868 589516 122874
rect 589464 122810 589516 122816
rect 589936 122058 589964 126375
rect 589924 122052 589976 122058
rect 589924 121994 589976 122000
rect 590014 121544 590070 121553
rect 590014 121479 590070 121488
rect 589646 119912 589702 119921
rect 589646 119847 589702 119856
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 589660 115258 589688 119847
rect 590028 118726 590056 121479
rect 590016 118720 590068 118726
rect 590016 118662 590068 118668
rect 590106 118280 590162 118289
rect 590106 118215 590162 118224
rect 589648 115252 589700 115258
rect 589648 115194 589700 115200
rect 589462 113384 589518 113393
rect 589462 113319 589518 113328
rect 589476 113218 589504 113319
rect 589464 113212 589516 113218
rect 589464 113154 589516 113160
rect 590120 112470 590148 118215
rect 590290 115016 590346 115025
rect 590290 114951 590346 114960
rect 590108 112464 590160 112470
rect 590108 112406 590160 112412
rect 589462 111752 589518 111761
rect 589462 111687 589518 111696
rect 589476 110498 589504 111687
rect 589464 110492 589516 110498
rect 589464 110434 589516 110440
rect 589278 110120 589334 110129
rect 589278 110055 589334 110064
rect 589292 109070 589320 110055
rect 589280 109064 589332 109070
rect 589280 109006 589332 109012
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589830 106856 589886 106865
rect 589830 106791 589886 106800
rect 589844 106350 589872 106791
rect 589832 106344 589884 106350
rect 589832 106286 589884 106292
rect 589462 105224 589518 105233
rect 589462 105159 589518 105168
rect 589476 104922 589504 105159
rect 589464 104916 589516 104922
rect 589464 104858 589516 104864
rect 588726 103592 588782 103601
rect 588726 103527 588782 103536
rect 588544 103488 588596 103494
rect 588544 103430 588596 103436
rect 587348 97980 587400 97986
rect 587348 97922 587400 97928
rect 587164 82136 587216 82142
rect 587164 82078 587216 82084
rect 588740 79354 588768 103527
rect 590304 103514 590332 114951
rect 589936 103486 590332 103514
rect 589462 101960 589518 101969
rect 589462 101895 589518 101904
rect 589476 100162 589504 101895
rect 589464 100156 589516 100162
rect 589464 100098 589516 100104
rect 589936 89010 589964 103486
rect 589924 89004 589976 89010
rect 589924 88946 589976 88952
rect 588728 79348 588780 79354
rect 588728 79290 588780 79296
rect 584404 71392 584456 71398
rect 584404 71334 584456 71340
rect 581644 54256 581696 54262
rect 577502 54224 577558 54233
rect 581644 54198 581696 54204
rect 577502 54159 577558 54168
rect 574928 53848 574980 53854
rect 574928 53790 574980 53796
rect 459834 53680 459890 53689
rect 459834 53615 459890 53624
rect 460754 53680 460810 53689
rect 460754 53615 460810 53624
rect 461674 53680 461730 53689
rect 461674 53615 461730 53624
rect 462594 53680 462650 53689
rect 463238 53680 463294 53689
rect 462594 53615 462650 53624
rect 462964 53644 463016 53650
rect 130384 53236 130436 53242
rect 130384 53178 130436 53184
rect 129004 53100 129056 53106
rect 129004 53042 129056 53048
rect 128820 51740 128872 51746
rect 128820 51682 128872 51688
rect 128832 44810 128860 51682
rect 129016 45422 129044 53042
rect 129188 51876 129240 51882
rect 129188 51818 129240 51824
rect 129556 51876 129608 51882
rect 129556 51818 129608 51824
rect 129004 45416 129056 45422
rect 129004 45358 129056 45364
rect 128820 44804 128872 44810
rect 128820 44746 128872 44752
rect 129200 44606 129228 51818
rect 129372 49156 129424 49162
rect 129372 49098 129424 49104
rect 129384 44946 129412 49098
rect 129568 45082 129596 51818
rect 130396 45966 130424 53178
rect 312360 53168 312412 53174
rect 312018 53116 312360 53122
rect 312018 53110 312412 53116
rect 313740 53168 313792 53174
rect 316316 53168 316368 53174
rect 313792 53116 314042 53122
rect 313740 53110 314042 53116
rect 312018 53094 312400 53110
rect 313752 53108 314042 53110
rect 316020 53116 316316 53122
rect 316020 53110 316368 53116
rect 317696 53168 317748 53174
rect 317748 53116 318380 53122
rect 317696 53110 318380 53116
rect 313752 53094 314056 53108
rect 316020 53094 316356 53110
rect 317708 53094 318380 53110
rect 130568 52012 130620 52018
rect 130568 51954 130620 51960
rect 130580 46102 130608 51954
rect 314028 50386 314056 53094
rect 318352 50522 318380 53094
rect 459468 53100 459520 53106
rect 459468 53042 459520 53048
rect 459480 52578 459508 53042
rect 459848 52578 459876 53615
rect 460066 52828 460118 52834
rect 460066 52770 460118 52776
rect 459172 52550 459508 52578
rect 459632 52550 459876 52578
rect 460078 52564 460106 52770
rect 460768 52578 460796 53615
rect 461308 53236 461360 53242
rect 461308 53178 461360 53184
rect 461320 52578 461348 53178
rect 461688 52578 461716 53615
rect 462228 53508 462280 53514
rect 462228 53450 462280 53456
rect 462240 52578 462268 53450
rect 462608 52578 462636 53615
rect 464250 53680 464306 53689
rect 463238 53615 463240 53624
rect 462964 53586 463016 53592
rect 463292 53615 463294 53624
rect 463516 53644 463568 53650
rect 463240 53586 463292 53592
rect 463516 53586 463568 53592
rect 463700 53644 463752 53650
rect 476026 53680 476082 53689
rect 464250 53615 464306 53624
rect 464436 53644 464488 53650
rect 463700 53586 463752 53592
rect 462976 52970 463004 53586
rect 463148 53372 463200 53378
rect 463148 53314 463200 53320
rect 462964 52964 463016 52970
rect 462964 52906 463016 52912
rect 463160 52578 463188 53314
rect 463528 52578 463556 53586
rect 463712 53106 463740 53586
rect 464066 53272 464122 53281
rect 464066 53207 464122 53216
rect 463700 53100 463752 53106
rect 463700 53042 463752 53048
rect 464080 52578 464108 53207
rect 464264 52578 464292 53615
rect 464436 53586 464488 53592
rect 464712 53644 464764 53650
rect 476578 53680 476634 53689
rect 476026 53615 476028 53624
rect 464712 53586 464764 53592
rect 476080 53615 476082 53624
rect 476212 53644 476264 53650
rect 476028 53586 476080 53592
rect 476212 53586 476264 53592
rect 476396 53644 476448 53650
rect 476578 53615 476580 53624
rect 476396 53586 476448 53592
rect 476632 53615 476634 53624
rect 477040 53644 477092 53650
rect 476580 53586 476632 53592
rect 477040 53586 477092 53592
rect 479064 53644 479116 53650
rect 479064 53586 479116 53592
rect 479432 53644 479484 53650
rect 479432 53586 479484 53592
rect 464448 53281 464476 53586
rect 464434 53272 464490 53281
rect 464434 53207 464490 53216
rect 464528 52964 464580 52970
rect 464528 52906 464580 52912
rect 460552 52550 460796 52578
rect 461012 52550 461348 52578
rect 461472 52550 461716 52578
rect 461932 52550 462268 52578
rect 462392 52550 462636 52578
rect 462852 52550 463188 52578
rect 463312 52550 463556 52578
rect 463772 52550 464108 52578
rect 464232 52550 464292 52578
rect 464540 52578 464568 52906
rect 464724 52834 464752 53586
rect 476224 53417 476252 53586
rect 476210 53408 476266 53417
rect 476210 53343 476266 53352
rect 465448 53100 465500 53106
rect 465448 53042 465500 53048
rect 464712 52828 464764 52834
rect 464712 52770 464764 52776
rect 465460 52578 465488 53042
rect 476408 52834 476436 53586
rect 477052 53417 477080 53586
rect 477038 53408 477094 53417
rect 477038 53343 477094 53352
rect 479076 53106 479104 53586
rect 479444 53514 479472 53586
rect 479616 53576 479668 53582
rect 479616 53518 479668 53524
rect 479432 53508 479484 53514
rect 479432 53450 479484 53456
rect 479628 53242 479656 53518
rect 479616 53236 479668 53242
rect 479616 53178 479668 53184
rect 479064 53100 479116 53106
rect 479064 53042 479116 53048
rect 465586 52828 465638 52834
rect 465586 52770 465638 52776
rect 476396 52828 476448 52834
rect 476396 52770 476448 52776
rect 464540 52550 464692 52578
rect 465152 52550 465488 52578
rect 465598 52564 465626 52770
rect 318340 50516 318392 50522
rect 318340 50458 318392 50464
rect 458180 50516 458232 50522
rect 458180 50458 458232 50464
rect 130844 50380 130896 50386
rect 130844 50322 130896 50328
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 130568 46096 130620 46102
rect 130568 46038 130620 46044
rect 130384 45960 130436 45966
rect 130384 45902 130436 45908
rect 129556 45076 129608 45082
rect 129556 45018 129608 45024
rect 129372 44940 129424 44946
rect 129372 44882 129424 44888
rect 129188 44600 129240 44606
rect 129188 44542 129240 44548
rect 50528 44328 50580 44334
rect 130856 44305 130884 50322
rect 131028 49020 131080 49026
rect 131028 48962 131080 48968
rect 50528 44270 50580 44276
rect 130842 44296 130898 44305
rect 130842 44231 130898 44240
rect 43444 44192 43496 44198
rect 43444 44134 43496 44140
rect 131040 44062 131068 48962
rect 458192 47025 458220 50458
rect 544028 50386 544056 53108
rect 545684 53094 546020 53122
rect 547892 53094 548044 53122
rect 458364 50380 458416 50386
rect 458364 50322 458416 50328
rect 522948 50380 523000 50386
rect 522948 50322 523000 50328
rect 544016 50380 544068 50386
rect 544016 50322 544068 50328
rect 458178 47016 458234 47025
rect 458178 46951 458234 46960
rect 458376 46753 458404 50322
rect 522960 47841 522988 50322
rect 522946 47832 523002 47841
rect 522946 47767 523002 47776
rect 459172 47654 459232 47682
rect 459632 47654 459968 47682
rect 460092 47654 460152 47682
rect 460552 47654 460888 47682
rect 461012 47654 461072 47682
rect 461472 47654 461808 47682
rect 461932 47654 461992 47682
rect 462392 47654 462728 47682
rect 462852 47654 462912 47682
rect 458362 46744 458418 46753
rect 142370 46702 142660 46730
rect 132868 46096 132920 46102
rect 132868 46038 132920 46044
rect 132592 45960 132644 45966
rect 132592 45902 132644 45908
rect 131580 44696 131632 44702
rect 131580 44638 131632 44644
rect 131592 44334 131620 44638
rect 132604 44402 132632 45902
rect 132880 44422 132908 46038
rect 132868 44416 132920 44422
rect 132592 44396 132644 44402
rect 132868 44358 132920 44364
rect 132592 44338 132644 44344
rect 131580 44328 131632 44334
rect 132776 44305 132828 44310
rect 142632 44305 142660 46702
rect 458362 46679 458418 46688
rect 131580 44270 131632 44276
rect 132774 44304 132830 44305
rect 132774 44296 132776 44304
rect 132828 44296 132830 44304
rect 132774 44231 132830 44240
rect 142618 44296 142674 44305
rect 142618 44231 142674 44240
rect 255870 44160 255926 44169
rect 255870 44095 255926 44104
rect 131028 44056 131080 44062
rect 131028 43998 131080 44004
rect 255884 42838 255912 44095
rect 361762 43888 361818 43897
rect 361762 43823 361818 43832
rect 440238 43888 440294 43897
rect 440238 43823 440240 43832
rect 187332 42832 187384 42838
rect 187332 42774 187384 42780
rect 255872 42832 255924 42838
rect 255872 42774 255924 42780
rect 187344 42092 187372 42774
rect 307300 42764 307352 42770
rect 307300 42706 307352 42712
rect 307312 42106 307340 42706
rect 310428 42628 310480 42634
rect 310428 42570 310480 42576
rect 310440 42106 310468 42570
rect 307004 42078 307340 42106
rect 310132 42078 310468 42106
rect 361776 42092 361804 43823
rect 440292 43823 440294 43832
rect 441066 43888 441122 43897
rect 441066 43823 441068 43832
rect 440240 43794 440292 43800
rect 441120 43823 441122 43832
rect 441068 43794 441120 43800
rect 431224 42764 431276 42770
rect 431224 42706 431276 42712
rect 441068 42764 441120 42770
rect 441068 42706 441120 42712
rect 449164 42764 449216 42770
rect 449164 42706 449216 42712
rect 453580 42764 453632 42770
rect 453580 42706 453632 42712
rect 427084 42628 427136 42634
rect 427084 42570 427136 42576
rect 415582 42392 415638 42401
rect 404452 42356 404504 42362
rect 404452 42298 404504 42304
rect 405188 42356 405240 42362
rect 415582 42327 415638 42336
rect 420736 42356 420788 42362
rect 405188 42298 405240 42304
rect 365074 41848 365130 41857
rect 364918 41806 365074 41834
rect 365074 41783 365130 41792
rect 404464 41478 404492 42298
rect 405200 42106 405228 42298
rect 415596 42106 415624 42327
rect 420736 42298 420788 42304
rect 426900 42356 426952 42362
rect 426900 42298 426952 42304
rect 405200 42078 405582 42106
rect 415426 42078 415624 42106
rect 416686 41848 416742 41857
rect 416622 41806 416686 41834
rect 419906 41848 419962 41857
rect 419750 41806 419906 41834
rect 416686 41783 416742 41792
rect 419906 41783 419962 41792
rect 420748 41478 420776 42298
rect 426912 41478 426940 42298
rect 427096 42022 427124 42570
rect 431236 42022 431264 42706
rect 441080 42022 441108 42706
rect 441252 42628 441304 42634
rect 441252 42570 441304 42576
rect 446404 42628 446456 42634
rect 446404 42570 446456 42576
rect 427084 42016 427136 42022
rect 427084 41958 427136 41964
rect 431224 42016 431276 42022
rect 431224 41958 431276 41964
rect 441068 42016 441120 42022
rect 441068 41958 441120 41964
rect 441264 41886 441292 42570
rect 446218 42256 446274 42265
rect 446218 42191 446274 42200
rect 441252 41880 441304 41886
rect 441252 41822 441304 41828
rect 446232 41585 446260 42191
rect 446416 42022 446444 42570
rect 446404 42016 446456 42022
rect 446404 41958 446456 41964
rect 449176 41886 449204 42706
rect 453592 41886 453620 42706
rect 454500 42492 454552 42498
rect 454500 42434 454552 42440
rect 454512 42022 454540 42434
rect 454500 42016 454552 42022
rect 454500 41958 454552 41964
rect 449164 41880 449216 41886
rect 449164 41822 449216 41828
rect 453580 41880 453632 41886
rect 453580 41822 453632 41828
rect 446218 41576 446274 41585
rect 446218 41511 446274 41520
rect 459204 41478 459232 47654
rect 459940 42106 459968 47654
rect 460124 44169 460152 47654
rect 460110 44160 460166 44169
rect 460110 44095 460166 44104
rect 460860 43489 460888 47654
rect 461044 44441 461072 47654
rect 461030 44432 461086 44441
rect 461030 44367 461086 44376
rect 460846 43480 460902 43489
rect 460846 43415 460902 43424
rect 461780 42945 461808 47654
rect 461766 42936 461822 42945
rect 461766 42871 461822 42880
rect 461964 42265 461992 47654
rect 462700 43217 462728 47654
rect 462884 44441 462912 47654
rect 463068 47654 463312 47682
rect 463772 47654 463832 47682
rect 462870 44432 462926 44441
rect 462870 44367 462926 44376
rect 462686 43208 462742 43217
rect 462686 43143 462742 43152
rect 463068 42498 463096 47654
rect 463804 44441 463832 47654
rect 464218 47410 464246 47668
rect 464172 47382 464246 47410
rect 464356 47654 464692 47682
rect 463790 44432 463846 44441
rect 463790 44367 463846 44376
rect 463974 42936 464030 42945
rect 463974 42871 464030 42880
rect 463988 42514 464016 42871
rect 464172 42770 464200 47382
rect 464356 44169 464384 47654
rect 465138 47410 465166 47668
rect 465092 47382 465166 47410
rect 465276 47654 465612 47682
rect 465092 47025 465120 47382
rect 465078 47016 465134 47025
rect 465078 46951 465134 46960
rect 465276 46753 465304 47654
rect 545684 47297 545712 53094
rect 547892 47569 547920 53094
rect 550008 48929 550036 53108
rect 549994 48920 550050 48929
rect 549994 48855 550050 48864
rect 552032 47841 552060 53108
rect 553688 53094 554024 53122
rect 553688 48113 553716 53094
rect 591316 51882 591344 212502
rect 591304 51876 591356 51882
rect 591304 51818 591356 51824
rect 592696 51746 592724 212638
rect 593984 210202 594012 222974
rect 596640 222012 596692 222018
rect 596640 221954 596692 221960
rect 596652 221610 596680 221954
rect 596836 221610 596864 245618
rect 629944 241528 629996 241534
rect 629944 241470 629996 241476
rect 629956 229094 629984 241470
rect 629956 229066 630076 229094
rect 610452 224874 611032 224890
rect 610452 224868 611044 224874
rect 610452 224862 610992 224868
rect 610452 224670 610480 224862
rect 610992 224810 611044 224816
rect 614948 224868 615000 224874
rect 614948 224810 615000 224816
rect 610808 224800 610860 224806
rect 610808 224742 610860 224748
rect 610440 224664 610492 224670
rect 610440 224606 610492 224612
rect 610624 224664 610676 224670
rect 610624 224606 610676 224612
rect 610636 224126 610664 224606
rect 610624 224120 610676 224126
rect 610624 224062 610676 224068
rect 610820 224058 610848 224742
rect 610808 224052 610860 224058
rect 610808 223994 610860 224000
rect 605012 222012 605064 222018
rect 605012 221954 605064 221960
rect 600780 221876 600832 221882
rect 600780 221818 600832 221824
rect 600964 221876 601016 221882
rect 600964 221818 601016 221824
rect 596640 221604 596692 221610
rect 596640 221546 596692 221552
rect 596824 221604 596876 221610
rect 596824 221546 596876 221552
rect 599490 221504 599546 221513
rect 599490 221439 599546 221448
rect 598572 220516 598624 220522
rect 598572 220458 598624 220464
rect 598584 220114 598612 220458
rect 598572 220108 598624 220114
rect 598572 220050 598624 220056
rect 596732 219904 596784 219910
rect 596732 219846 596784 219852
rect 594800 218340 594852 218346
rect 594800 218282 594852 218288
rect 594812 216782 594840 218282
rect 595166 217288 595222 217297
rect 595166 217223 595222 217232
rect 594800 216776 594852 216782
rect 594800 216718 594852 216724
rect 594800 213240 594852 213246
rect 594800 213182 594852 213188
rect 594812 210202 594840 213182
rect 595180 210202 595208 217223
rect 595718 217016 595774 217025
rect 595718 216951 595774 216960
rect 595732 210202 595760 216951
rect 596364 216912 596416 216918
rect 596364 216854 596416 216860
rect 596376 210202 596404 216854
rect 596744 210202 596772 219846
rect 597560 219224 597612 219230
rect 597560 219166 597612 219172
rect 597572 210202 597600 219166
rect 598848 218748 598900 218754
rect 598848 218690 598900 218696
rect 598860 217326 598888 218690
rect 598480 217320 598532 217326
rect 598480 217262 598532 217268
rect 598848 217320 598900 217326
rect 598848 217262 598900 217268
rect 597928 217184 597980 217190
rect 597928 217126 597980 217132
rect 597940 210202 597968 217126
rect 598492 210202 598520 217262
rect 599030 215656 599086 215665
rect 599030 215591 599086 215600
rect 599044 210202 599072 215591
rect 599504 210202 599532 221439
rect 600792 221354 600820 221818
rect 600976 221474 601004 221818
rect 600964 221468 601016 221474
rect 600964 221410 601016 221416
rect 600792 221338 600912 221354
rect 600792 221332 600924 221338
rect 600792 221326 600872 221332
rect 600872 221274 600924 221280
rect 604644 221332 604696 221338
rect 604644 221274 604696 221280
rect 600504 221264 600556 221270
rect 600504 221206 600556 221212
rect 600686 221232 600742 221241
rect 600320 220856 600372 220862
rect 600320 220798 600372 220804
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596376 210174 596620 210202
rect 596744 210174 597172 210202
rect 597572 210174 597724 210202
rect 597940 210174 598276 210202
rect 598492 210174 598828 210202
rect 599044 210174 599380 210202
rect 599504 210174 599932 210202
rect 600332 210118 600360 220798
rect 600516 214470 600544 221206
rect 600686 221167 600742 221176
rect 600504 214464 600556 214470
rect 600504 214406 600556 214412
rect 600700 210202 600728 221167
rect 601792 221128 601844 221134
rect 601792 221070 601844 221076
rect 600964 220516 601016 220522
rect 600964 220458 601016 220464
rect 600976 219978 601004 220458
rect 600964 219972 601016 219978
rect 600964 219914 601016 219920
rect 600872 219632 600924 219638
rect 600924 219580 601280 219586
rect 600872 219574 601280 219580
rect 600884 219558 601280 219574
rect 601252 219502 601280 219558
rect 601240 219496 601292 219502
rect 601240 219438 601292 219444
rect 601240 214464 601292 214470
rect 601240 214406 601292 214412
rect 600484 210174 600728 210202
rect 601252 210202 601280 214406
rect 601804 210202 601832 221070
rect 602252 220992 602304 220998
rect 602252 220934 602304 220940
rect 602264 210202 602292 220934
rect 603080 218884 603132 218890
rect 603080 218826 603132 218832
rect 603092 217462 603120 218826
rect 604460 218476 604512 218482
rect 604460 218418 604512 218424
rect 604000 217864 604052 217870
rect 604000 217806 604052 217812
rect 603264 217728 603316 217734
rect 603264 217670 603316 217676
rect 603080 217456 603132 217462
rect 603080 217398 603132 217404
rect 603276 210202 603304 217670
rect 603448 217184 603500 217190
rect 603448 217126 603500 217132
rect 601252 210174 601588 210202
rect 601804 210174 602140 210202
rect 602264 210174 602692 210202
rect 603244 210174 603304 210202
rect 603460 210202 603488 217126
rect 604012 210202 604040 217806
rect 604472 217734 604500 218418
rect 604460 217728 604512 217734
rect 604460 217670 604512 217676
rect 604656 210202 604684 221274
rect 605024 210202 605052 221954
rect 606668 221876 606720 221882
rect 606668 221818 606720 221824
rect 606024 219768 606076 219774
rect 606024 219710 606076 219716
rect 606036 210202 606064 219710
rect 606208 217592 606260 217598
rect 606208 217534 606260 217540
rect 603460 210174 603796 210202
rect 604012 210174 604348 210202
rect 604656 210174 604900 210202
rect 605024 210174 605452 210202
rect 606004 210174 606064 210202
rect 606220 210202 606248 217534
rect 606680 210202 606708 221818
rect 608600 221740 608652 221746
rect 608600 221682 608652 221688
rect 607312 220108 607364 220114
rect 607312 220050 607364 220056
rect 607324 210202 607352 220050
rect 607496 219496 607548 219502
rect 607496 219438 607548 219444
rect 607508 210338 607536 219438
rect 607508 210310 607812 210338
rect 607784 210202 607812 210310
rect 608612 210202 608640 221682
rect 610532 220652 610584 220658
rect 610532 220594 610584 220600
rect 609428 220380 609480 220386
rect 609428 220322 609480 220328
rect 608876 220244 608928 220250
rect 608876 220186 608928 220192
rect 608888 210202 608916 220186
rect 609440 210202 609468 220322
rect 610072 217048 610124 217054
rect 610072 216990 610124 216996
rect 610084 210202 610112 216990
rect 610544 210202 610572 220594
rect 611452 220516 611504 220522
rect 611452 220458 611504 220464
rect 610716 218612 610768 218618
rect 610716 218554 610768 218560
rect 610728 216782 610756 218554
rect 610716 216776 610768 216782
rect 610716 216718 610768 216724
rect 611464 210202 611492 220458
rect 611634 220280 611690 220289
rect 611634 220215 611690 220224
rect 611648 210202 611676 220215
rect 612922 219736 612978 219745
rect 612922 219671 612978 219680
rect 612280 218000 612332 218006
rect 612280 217942 612332 217948
rect 612292 210202 612320 217942
rect 612936 210202 612964 219671
rect 614120 219020 614172 219026
rect 614120 218962 614172 218968
rect 614132 217598 614160 218962
rect 614488 218000 614540 218006
rect 614488 217942 614540 217948
rect 614304 217728 614356 217734
rect 614304 217670 614356 217676
rect 614120 217592 614172 217598
rect 614120 217534 614172 217540
rect 613384 216912 613436 216918
rect 613384 216854 613436 216860
rect 613396 210202 613424 216854
rect 614316 210202 614344 217670
rect 606220 210174 606556 210202
rect 606680 210174 607108 210202
rect 607324 210174 607660 210202
rect 607784 210174 608212 210202
rect 608612 210174 608764 210202
rect 608888 210174 609316 210202
rect 609440 210174 609868 210202
rect 610084 210174 610420 210202
rect 610544 210174 610972 210202
rect 611464 210174 611524 210202
rect 611648 210174 612076 210202
rect 612292 210174 612628 210202
rect 612936 210174 613180 210202
rect 613396 210174 613732 210202
rect 614284 210174 614344 210202
rect 614500 210202 614528 217942
rect 614960 210202 614988 224810
rect 616052 224664 616104 224670
rect 616052 224606 616104 224612
rect 615684 216776 615736 216782
rect 615684 216718 615736 216724
rect 615696 210202 615724 216718
rect 616064 210202 616092 224606
rect 625436 224528 625488 224534
rect 625436 224470 625488 224476
rect 625252 224392 625304 224398
rect 625252 224334 625304 224340
rect 619640 224256 619692 224262
rect 619640 224198 619692 224204
rect 618258 220960 618314 220969
rect 618258 220895 618314 220904
rect 617154 220008 617210 220017
rect 617154 219943 617210 219952
rect 616880 214872 616932 214878
rect 616880 214814 616932 214820
rect 616892 210202 616920 214814
rect 617168 210202 617196 219943
rect 617798 215928 617854 215937
rect 617798 215863 617854 215872
rect 617812 210202 617840 215863
rect 618272 214606 618300 220895
rect 618442 219464 618498 219473
rect 618442 219399 618498 219408
rect 618260 214600 618312 214606
rect 618260 214542 618312 214548
rect 618456 210202 618484 219399
rect 618904 214600 618956 214606
rect 618904 214542 618956 214548
rect 618916 210202 618944 214542
rect 619652 210202 619680 224198
rect 623780 224052 623832 224058
rect 623780 223994 623832 224000
rect 622676 223916 622728 223922
rect 622676 223858 622728 223864
rect 621572 223780 621624 223786
rect 621572 223722 621624 223728
rect 620652 223168 620704 223174
rect 620652 223110 620704 223116
rect 620284 223032 620336 223038
rect 620284 222974 620336 222980
rect 620296 222766 620324 222974
rect 620284 222760 620336 222766
rect 620284 222702 620336 222708
rect 620468 222760 620520 222766
rect 620468 222702 620520 222708
rect 619916 222624 619968 222630
rect 619916 222566 619968 222572
rect 619928 214606 619956 222566
rect 620480 222222 620508 222702
rect 620664 222222 620692 223110
rect 620468 222216 620520 222222
rect 620468 222158 620520 222164
rect 620652 222216 620704 222222
rect 620652 222158 620704 222164
rect 620100 219632 620152 219638
rect 620100 219574 620152 219580
rect 619916 214600 619968 214606
rect 619916 214542 619968 214548
rect 620112 210202 620140 219574
rect 621110 215384 621166 215393
rect 621110 215319 621166 215328
rect 620560 214600 620612 214606
rect 620560 214542 620612 214548
rect 620572 210202 620600 214542
rect 621124 210202 621152 215319
rect 621584 210202 621612 223722
rect 622400 217320 622452 217326
rect 622400 217262 622452 217268
rect 622412 210202 622440 217262
rect 622688 210202 622716 223858
rect 623320 214736 623372 214742
rect 623320 214678 623372 214684
rect 623332 210202 623360 214678
rect 623792 210202 623820 223994
rect 623962 218104 624018 218113
rect 623962 218039 624018 218048
rect 623976 214606 624004 218039
rect 625264 214606 625292 224334
rect 623964 214600 624016 214606
rect 623964 214542 624016 214548
rect 625252 214600 625304 214606
rect 625252 214542 625304 214548
rect 624424 214464 624476 214470
rect 624424 214406 624476 214412
rect 624436 210202 624464 214406
rect 625448 210202 625476 224470
rect 628748 223644 628800 223650
rect 628748 223586 628800 223592
rect 625620 223032 625672 223038
rect 625620 222974 625672 222980
rect 614500 210174 614836 210202
rect 614960 210174 615388 210202
rect 615696 210174 615940 210202
rect 616064 210174 616492 210202
rect 616892 210174 617044 210202
rect 617168 210174 617596 210202
rect 617812 210174 618148 210202
rect 618456 210174 618700 210202
rect 618916 210174 619252 210202
rect 619652 210174 619804 210202
rect 620112 210174 620356 210202
rect 620572 210174 620908 210202
rect 621124 210174 621460 210202
rect 621584 210174 622012 210202
rect 622412 210174 622564 210202
rect 622688 210174 623116 210202
rect 623332 210174 623668 210202
rect 623792 210174 624220 210202
rect 624436 210174 624772 210202
rect 625324 210174 625476 210202
rect 625632 210202 625660 222974
rect 627092 222760 627144 222766
rect 627092 222702 627144 222708
rect 626632 217592 626684 217598
rect 626632 217534 626684 217540
rect 626080 214600 626132 214606
rect 626080 214542 626132 214548
rect 626092 210202 626120 214542
rect 626644 210202 626672 217534
rect 627104 210202 627132 222702
rect 627920 222488 627972 222494
rect 627920 222430 627972 222436
rect 627932 210202 627960 222430
rect 628288 217456 628340 217462
rect 628288 217398 628340 217404
rect 628300 210202 628328 217398
rect 628760 210202 628788 223586
rect 629852 222352 629904 222358
rect 629852 222294 629904 222300
rect 629392 214464 629444 214470
rect 629392 214406 629444 214412
rect 629404 210202 629432 214406
rect 629864 210202 629892 222294
rect 630048 214606 630076 229066
rect 633716 227044 633768 227050
rect 633716 226986 633768 226992
rect 630864 225004 630916 225010
rect 630864 224946 630916 224952
rect 630678 218376 630734 218385
rect 630678 218311 630734 218320
rect 630036 214600 630088 214606
rect 630036 214542 630088 214548
rect 630692 210202 630720 218311
rect 630876 210338 630904 224946
rect 632704 222896 632756 222902
rect 632704 222838 632756 222844
rect 631508 222216 631560 222222
rect 631508 222158 631560 222164
rect 630876 210310 630996 210338
rect 630968 210202 630996 210310
rect 631520 210202 631548 222158
rect 632716 213042 632744 222838
rect 633440 221604 633492 221610
rect 633440 221546 633492 221552
rect 632888 214600 632940 214606
rect 632888 214542 632940 214548
rect 632704 213036 632756 213042
rect 632704 212978 632756 212984
rect 632900 210202 632928 214542
rect 633452 210202 633480 221546
rect 633728 210202 633756 226986
rect 634360 213036 634412 213042
rect 634360 212978 634412 212984
rect 634372 210202 634400 212978
rect 635108 210202 635136 277743
rect 635568 272814 635596 278052
rect 635556 272808 635608 272814
rect 635556 272750 635608 272756
rect 636212 229094 636240 278287
rect 649264 278258 649316 278264
rect 650656 278186 650684 494702
rect 664456 491366 664484 549850
rect 664444 491360 664496 491366
rect 664444 491302 664496 491308
rect 665100 485858 665128 564538
rect 667018 562320 667074 562329
rect 667018 562255 667074 562264
rect 665824 552696 665876 552702
rect 665824 552638 665876 552644
rect 665836 491502 665864 552638
rect 665824 491496 665876 491502
rect 665824 491438 665876 491444
rect 665088 485852 665140 485858
rect 665088 485794 665140 485800
rect 667032 484430 667060 562255
rect 667216 535974 667244 596158
rect 667204 535968 667256 535974
rect 667204 535910 667256 535916
rect 667400 529990 667428 600879
rect 667570 594824 667626 594833
rect 667570 594759 667626 594768
rect 667388 529984 667440 529990
rect 667388 529926 667440 529932
rect 667584 524482 667612 594759
rect 667572 524476 667624 524482
rect 667572 524418 667624 524424
rect 667584 521626 667612 524418
rect 667572 521620 667624 521626
rect 667572 521562 667624 521568
rect 667020 484424 667072 484430
rect 667020 484366 667072 484372
rect 657544 467152 657596 467158
rect 657544 467094 657596 467100
rect 657556 460222 657584 467094
rect 653404 460216 653456 460222
rect 653404 460158 653456 460164
rect 657544 460216 657596 460222
rect 657544 460158 657596 460164
rect 652022 400888 652078 400897
rect 652022 400823 652078 400832
rect 651472 373992 651524 373998
rect 651472 373934 651524 373940
rect 651484 373289 651512 373934
rect 651470 373280 651526 373289
rect 651470 373215 651526 373224
rect 652036 372201 652064 400823
rect 652206 396672 652262 396681
rect 652206 396607 652262 396616
rect 652220 373969 652248 396607
rect 652206 373960 652262 373969
rect 652206 373895 652262 373904
rect 652022 372192 652078 372201
rect 652022 372127 652078 372136
rect 651472 371000 651524 371006
rect 651472 370942 651524 370948
rect 651484 370705 651512 370942
rect 651470 370696 651526 370705
rect 651470 370631 651526 370640
rect 652206 356688 652262 356697
rect 652206 356623 652262 356632
rect 652024 348424 652076 348430
rect 652024 348366 652076 348372
rect 651472 328296 651524 328302
rect 651472 328238 651524 328244
rect 651484 328137 651512 328238
rect 651470 328128 651526 328137
rect 651470 328063 651526 328072
rect 651746 325680 651802 325689
rect 651746 325615 651748 325624
rect 651800 325615 651802 325624
rect 651748 325586 651800 325592
rect 650828 322992 650880 322998
rect 650828 322934 650880 322940
rect 650840 278458 650868 322934
rect 651380 303408 651432 303414
rect 651378 303376 651380 303385
rect 651432 303376 651434 303385
rect 651378 303311 651434 303320
rect 651472 300824 651524 300830
rect 651472 300766 651524 300772
rect 651484 300665 651512 300766
rect 651470 300656 651526 300665
rect 651470 300591 651526 300600
rect 651470 298752 651526 298761
rect 651470 298687 651526 298696
rect 651484 298178 651512 298687
rect 651472 298172 651524 298178
rect 651472 298114 651524 298120
rect 651654 296848 651710 296857
rect 651654 296783 651656 296792
rect 651708 296783 651710 296792
rect 651656 296754 651708 296760
rect 652036 296714 652064 348366
rect 652220 326913 652248 356623
rect 652574 351112 652630 351121
rect 652574 351047 652630 351056
rect 652588 329769 652616 351047
rect 652574 329760 652630 329769
rect 652574 329695 652630 329704
rect 652206 326904 652262 326913
rect 652206 326839 652262 326848
rect 653416 322998 653444 460158
rect 667860 456618 667888 703802
rect 668398 689480 668454 689489
rect 668398 689415 668454 689424
rect 668216 661156 668268 661162
rect 668216 661098 668268 661104
rect 667848 456612 667900 456618
rect 667848 456554 667900 456560
rect 668228 455666 668256 661098
rect 668412 616894 668440 689415
rect 668596 671158 668624 733382
rect 668766 730144 668822 730153
rect 668766 730079 668822 730088
rect 668584 671152 668636 671158
rect 668584 671094 668636 671100
rect 668780 660142 668808 730079
rect 669056 709374 669084 782478
rect 669044 709368 669096 709374
rect 669044 709310 669096 709316
rect 669240 708801 669268 784110
rect 670424 777028 670476 777034
rect 670424 776970 670476 776976
rect 669964 775600 670016 775606
rect 669964 775542 670016 775548
rect 669596 738336 669648 738342
rect 669596 738278 669648 738284
rect 669410 728784 669466 728793
rect 669410 728719 669466 728728
rect 669226 708792 669282 708801
rect 669226 708727 669282 708736
rect 669228 705220 669280 705226
rect 669228 705162 669280 705168
rect 668952 693116 669004 693122
rect 668952 693058 669004 693064
rect 668768 660136 668820 660142
rect 668768 660078 668820 660084
rect 668584 640348 668636 640354
rect 668584 640290 668636 640296
rect 668400 616888 668452 616894
rect 668400 616830 668452 616836
rect 668596 580310 668624 640290
rect 668964 620294 668992 693058
rect 668952 620288 669004 620294
rect 668952 620230 669004 620236
rect 669044 608660 669096 608666
rect 669044 608602 669096 608608
rect 668858 593600 668914 593609
rect 668858 593535 668914 593544
rect 668584 580304 668636 580310
rect 668584 580246 668636 580252
rect 668872 528630 668900 593535
rect 669056 536489 669084 608602
rect 669042 536480 669098 536489
rect 669042 536415 669098 536424
rect 668860 528624 668912 528630
rect 668860 528566 668912 528572
rect 669240 456006 669268 705162
rect 669424 663950 669452 728719
rect 669608 665310 669636 738278
rect 669976 715766 670004 775542
rect 669964 715760 670016 715766
rect 669964 715702 670016 715708
rect 670436 705974 670464 776970
rect 670620 709238 670648 784246
rect 670896 728142 670924 886858
rect 670884 728136 670936 728142
rect 670884 728078 670936 728084
rect 671080 715494 671108 894270
rect 671436 773424 671488 773430
rect 671436 773366 671488 773372
rect 671448 750734 671476 773366
rect 671448 750706 671568 750734
rect 671540 736934 671568 750706
rect 671712 743912 671764 743918
rect 671712 743854 671764 743860
rect 671724 742642 671752 743854
rect 671908 743834 671936 894406
rect 672264 892900 672316 892906
rect 672264 892842 672316 892848
rect 671908 743806 672028 743834
rect 671448 736906 671568 736934
rect 671632 742614 671752 742642
rect 671250 733816 671306 733825
rect 671250 733751 671306 733760
rect 671068 715488 671120 715494
rect 671068 715430 671120 715436
rect 671068 713244 671120 713250
rect 671068 713186 671120 713192
rect 670608 709232 670660 709238
rect 670608 709174 670660 709180
rect 670424 705968 670476 705974
rect 670424 705910 670476 705916
rect 670606 687712 670662 687721
rect 670606 687647 670662 687656
rect 669964 687268 670016 687274
rect 669964 687210 670016 687216
rect 669778 685536 669834 685545
rect 669778 685471 669834 685480
rect 669596 665304 669648 665310
rect 669596 665246 669648 665252
rect 669412 663944 669464 663950
rect 669412 663886 669464 663892
rect 669594 644328 669650 644337
rect 669594 644263 669650 644272
rect 669412 623076 669464 623082
rect 669412 623018 669464 623024
rect 669424 578202 669452 623018
rect 669412 578196 669464 578202
rect 669412 578138 669464 578144
rect 669412 576972 669464 576978
rect 669412 576914 669464 576920
rect 669424 532574 669452 576914
rect 669608 572286 669636 644263
rect 669792 615670 669820 685471
rect 669976 625598 670004 687210
rect 670240 669384 670292 669390
rect 670240 669326 670292 669332
rect 669964 625592 670016 625598
rect 669964 625534 670016 625540
rect 670252 625054 670280 669326
rect 670240 625048 670292 625054
rect 670240 624990 670292 624996
rect 670424 624708 670476 624714
rect 670424 624650 670476 624656
rect 670240 623892 670292 623898
rect 670240 623834 670292 623840
rect 669780 615664 669832 615670
rect 669780 615606 669832 615612
rect 669964 597576 670016 597582
rect 669964 597518 670016 597524
rect 669596 572280 669648 572286
rect 669596 572222 669648 572228
rect 669780 568608 669832 568614
rect 669780 568550 669832 568556
rect 669412 532568 669464 532574
rect 669412 532510 669464 532516
rect 669228 456000 669280 456006
rect 669228 455942 669280 455948
rect 668216 455660 668268 455666
rect 668216 455602 668268 455608
rect 669792 455433 669820 568550
rect 669976 535702 670004 597518
rect 670252 579086 670280 623834
rect 670436 579902 670464 624650
rect 670620 617506 670648 687647
rect 670884 685976 670936 685982
rect 670884 685918 670936 685924
rect 670896 620022 670924 685918
rect 671080 668574 671108 713186
rect 671068 668568 671120 668574
rect 671068 668510 671120 668516
rect 671068 667956 671120 667962
rect 671068 667898 671120 667904
rect 671080 623558 671108 667898
rect 671264 661638 671292 733751
rect 671448 710054 671476 736906
rect 671436 710048 671488 710054
rect 671436 709990 671488 709996
rect 671436 668228 671488 668234
rect 671436 668170 671488 668176
rect 671252 661632 671304 661638
rect 671252 661574 671304 661580
rect 671448 659654 671476 668170
rect 671632 667214 671660 742614
rect 671804 742212 671856 742218
rect 671804 742154 671856 742160
rect 671816 734174 671844 742154
rect 672000 734174 672028 743806
rect 671724 734146 671844 734174
rect 671908 734146 672028 734174
rect 671724 692774 671752 734146
rect 671908 714542 671936 734146
rect 672078 732728 672134 732737
rect 672078 732663 672134 732672
rect 671896 714536 671948 714542
rect 671896 714478 671948 714484
rect 671896 712428 671948 712434
rect 671896 712370 671948 712376
rect 671724 692746 671844 692774
rect 671620 667208 671672 667214
rect 671620 667150 671672 667156
rect 671816 667026 671844 692746
rect 671724 666998 671844 667026
rect 671724 664426 671752 666998
rect 671908 666942 671936 712370
rect 671896 666936 671948 666942
rect 671896 666878 671948 666884
rect 671896 666596 671948 666602
rect 671896 666538 671948 666544
rect 671712 664420 671764 664426
rect 671712 664362 671764 664368
rect 671448 659626 671568 659654
rect 671540 640334 671568 659626
rect 671710 647864 671766 647873
rect 671710 647799 671766 647808
rect 671540 640306 671660 640334
rect 671342 638616 671398 638625
rect 671342 638551 671398 638560
rect 671356 632942 671384 638551
rect 671632 633026 671660 640306
rect 671540 633010 671660 633026
rect 671528 633004 671660 633010
rect 671580 632998 671660 633004
rect 671528 632946 671580 632952
rect 671344 632936 671396 632942
rect 671344 632878 671396 632884
rect 671344 632800 671396 632806
rect 671344 632742 671396 632748
rect 671356 627994 671384 632742
rect 671528 632664 671580 632670
rect 671528 632606 671580 632612
rect 671356 627966 671476 627994
rect 671448 624374 671476 627966
rect 671540 627914 671568 632606
rect 671540 627886 671660 627914
rect 671436 624368 671488 624374
rect 671436 624310 671488 624316
rect 671068 623552 671120 623558
rect 671068 623494 671120 623500
rect 671434 620800 671490 620809
rect 671434 620735 671490 620744
rect 670884 620016 670936 620022
rect 670884 619958 670936 619964
rect 670608 617500 670660 617506
rect 670608 617442 670660 617448
rect 670608 614168 670660 614174
rect 670608 614110 670660 614116
rect 670424 579896 670476 579902
rect 670424 579838 670476 579844
rect 670240 579080 670292 579086
rect 670240 579022 670292 579028
rect 670240 577788 670292 577794
rect 670240 577730 670292 577736
rect 669964 535696 670016 535702
rect 669964 535638 670016 535644
rect 670252 533390 670280 577730
rect 670422 549672 670478 549681
rect 670422 549607 670478 549616
rect 670240 533384 670292 533390
rect 670240 533326 670292 533332
rect 669964 500268 670016 500274
rect 669964 500210 670016 500216
rect 669976 491910 670004 500210
rect 669964 491904 670016 491910
rect 669964 491846 670016 491852
rect 670436 480758 670464 549607
rect 669964 480752 670016 480758
rect 669964 480694 670016 480700
rect 670424 480752 670476 480758
rect 670424 480694 670476 480700
rect 669976 467158 670004 480694
rect 669964 467152 670016 467158
rect 669964 467094 670016 467100
rect 669778 455424 669834 455433
rect 669778 455359 669834 455368
rect 670620 455161 670648 614110
rect 670974 607744 671030 607753
rect 670974 607679 671030 607688
rect 670792 579420 670844 579426
rect 670792 579362 670844 579368
rect 670804 534886 670832 579362
rect 670792 534880 670844 534886
rect 670792 534822 670844 534828
rect 670790 533896 670846 533905
rect 670790 533831 670846 533840
rect 670804 490958 670832 533831
rect 670988 529310 671016 607679
rect 671160 578604 671212 578610
rect 671160 578546 671212 578552
rect 671172 534614 671200 578546
rect 671448 577454 671476 620735
rect 671436 577448 671488 577454
rect 671436 577390 671488 577396
rect 671632 574598 671660 627886
rect 671724 611354 671752 647799
rect 671908 637574 671936 666538
rect 672092 663474 672120 732663
rect 672276 712910 672304 892842
rect 672736 866658 672764 895766
rect 675864 895694 675892 896679
rect 676034 896336 676090 896345
rect 676034 896271 676090 896280
rect 676048 895830 676076 896271
rect 676036 895824 676088 895830
rect 676036 895766 676088 895772
rect 675852 895688 675904 895694
rect 675852 895630 675904 895636
rect 675850 895520 675906 895529
rect 675850 895455 675906 895464
rect 675864 894334 675892 895455
rect 676034 894704 676090 894713
rect 676034 894639 676090 894648
rect 676048 894470 676076 894639
rect 676036 894464 676088 894470
rect 676036 894406 676088 894412
rect 675852 894328 675904 894334
rect 675852 894270 675904 894276
rect 675850 893888 675906 893897
rect 675850 893823 675906 893832
rect 675864 893042 675892 893823
rect 676034 893072 676090 893081
rect 673276 893036 673328 893042
rect 673276 892978 673328 892984
rect 675852 893036 675904 893042
rect 676034 893007 676090 893016
rect 675852 892978 675904 892984
rect 673090 885456 673146 885465
rect 673090 885391 673146 885400
rect 672724 866652 672776 866658
rect 672724 866594 672776 866600
rect 672906 777472 672962 777481
rect 672906 777407 672962 777416
rect 672724 775668 672776 775674
rect 672724 775610 672776 775616
rect 672448 739152 672500 739158
rect 672448 739094 672500 739100
rect 672264 712904 672316 712910
rect 672264 712846 672316 712852
rect 672262 696960 672318 696969
rect 672262 696895 672318 696904
rect 672080 663468 672132 663474
rect 672080 663410 672132 663416
rect 672078 652080 672134 652089
rect 672078 652015 672134 652024
rect 672092 647234 672120 652015
rect 672276 649994 672304 696895
rect 672460 665174 672488 739094
rect 672736 721754 672764 775610
rect 672920 760394 672948 777407
rect 672552 721726 672764 721754
rect 672828 760366 672948 760394
rect 672552 715034 672580 721726
rect 672828 717614 672856 760366
rect 673104 728346 673132 885391
rect 673288 728385 673316 892978
rect 676048 892906 676076 893007
rect 676036 892900 676088 892906
rect 676036 892842 676088 892848
rect 676034 892664 676090 892673
rect 676090 892622 676444 892650
rect 676034 892599 676090 892608
rect 676034 891440 676090 891449
rect 676034 891375 676090 891384
rect 675850 891032 675906 891041
rect 675850 890967 675906 890976
rect 674840 890384 674892 890390
rect 674840 890326 674892 890332
rect 674380 888956 674432 888962
rect 674380 888898 674432 888904
rect 674196 887324 674248 887330
rect 674196 887266 674248 887272
rect 674012 879028 674064 879034
rect 674012 878970 674064 878976
rect 674024 873730 674052 878970
rect 674012 873724 674064 873730
rect 674012 873666 674064 873672
rect 674208 872030 674236 887266
rect 674196 872024 674248 872030
rect 674196 871966 674248 871972
rect 674392 869666 674420 888898
rect 674656 888548 674708 888554
rect 674656 888490 674708 888496
rect 674668 872114 674696 888490
rect 674852 874954 674880 890326
rect 675864 888758 675892 890967
rect 676048 890390 676076 891375
rect 676036 890384 676088 890390
rect 676036 890326 676088 890332
rect 676034 890216 676090 890225
rect 676090 890186 676260 890202
rect 676090 890180 676272 890186
rect 676090 890174 676220 890180
rect 676034 890151 676090 890160
rect 676220 890122 676272 890128
rect 676034 889400 676090 889409
rect 676090 889358 676260 889386
rect 676034 889335 676090 889344
rect 676034 888992 676090 889001
rect 676034 888927 676036 888936
rect 676088 888927 676090 888936
rect 676036 888898 676088 888904
rect 676232 888758 676260 889358
rect 675024 888752 675076 888758
rect 675024 888694 675076 888700
rect 675852 888752 675904 888758
rect 675852 888694 675904 888700
rect 676220 888752 676272 888758
rect 676220 888694 676272 888700
rect 674840 874948 674892 874954
rect 674840 874890 674892 874896
rect 675036 874562 675064 888694
rect 676034 888584 676090 888593
rect 676034 888519 676036 888528
rect 676088 888519 676090 888528
rect 676036 888490 676088 888496
rect 676034 887360 676090 887369
rect 676034 887295 676036 887304
rect 676088 887295 676090 887304
rect 676036 887266 676088 887272
rect 676034 886952 676090 886961
rect 676034 886887 676036 886896
rect 676088 886887 676090 886896
rect 676036 886858 676088 886864
rect 676416 886650 676444 892622
rect 679622 891848 679678 891857
rect 679622 891783 679678 891792
rect 676864 890180 676916 890186
rect 676864 890122 676916 890128
rect 675576 886644 675628 886650
rect 675576 886586 675628 886592
rect 676404 886644 676456 886650
rect 676404 886586 676456 886592
rect 675588 881834 675616 886586
rect 675220 881806 675616 881834
rect 675220 879074 675248 881806
rect 675392 880388 675444 880394
rect 675392 880330 675444 880336
rect 675404 879322 675432 880330
rect 675576 879640 675628 879646
rect 675576 879582 675628 879588
rect 675128 879046 675248 879074
rect 675312 879294 675432 879322
rect 675128 876262 675156 879046
rect 675312 877418 675340 879294
rect 675588 879074 675616 879582
rect 676876 879374 676904 890122
rect 678242 889808 678298 889817
rect 678242 889743 678298 889752
rect 677048 888752 677100 888758
rect 677048 888694 677100 888700
rect 675760 879368 675812 879374
rect 675760 879310 675812 879316
rect 676864 879368 676916 879374
rect 676864 879310 676916 879316
rect 675404 879046 675616 879074
rect 675404 878084 675432 879046
rect 675772 878422 675800 879310
rect 675944 879232 675996 879238
rect 675944 879174 675996 879180
rect 675956 878529 675984 879174
rect 677060 879102 677088 888694
rect 678256 879238 678284 889743
rect 679636 880462 679664 891783
rect 681002 890624 681058 890633
rect 681002 890559 681058 890568
rect 681016 880705 681044 890559
rect 683118 888176 683174 888185
rect 683118 888111 683174 888120
rect 681002 880696 681058 880705
rect 681002 880631 681058 880640
rect 679624 880456 679676 880462
rect 683132 880433 683160 888111
rect 679624 880398 679676 880404
rect 683118 880424 683174 880433
rect 683118 880359 683174 880368
rect 678244 879232 678296 879238
rect 678244 879174 678296 879180
rect 677048 879096 677100 879102
rect 677048 879038 677100 879044
rect 675942 878520 675998 878529
rect 675942 878455 675998 878464
rect 675760 878416 675812 878422
rect 675760 878358 675812 878364
rect 675404 877418 675432 877540
rect 675312 877390 675432 877418
rect 675484 877260 675536 877266
rect 675484 877202 675536 877208
rect 675496 876860 675524 877202
rect 675128 876234 675418 876262
rect 675392 874948 675444 874954
rect 675392 874890 675444 874896
rect 675404 874834 675432 874890
rect 675404 874806 675524 874834
rect 675036 874534 675156 874562
rect 675128 873610 675156 874534
rect 675496 874412 675524 874806
rect 675574 874168 675630 874177
rect 675574 874103 675630 874112
rect 675588 873868 675616 874103
rect 675392 873724 675444 873730
rect 675392 873666 675444 873672
rect 675128 873582 675340 873610
rect 674930 873080 674986 873089
rect 674930 873015 674986 873024
rect 674668 872086 674880 872114
rect 674656 872024 674708 872030
rect 674708 871972 674788 871978
rect 674656 871966 674788 871972
rect 674668 871950 674788 871966
rect 674760 869802 674788 871950
rect 674852 869938 674880 872086
rect 674944 870074 674972 873015
rect 675312 870074 675340 873582
rect 675404 873188 675432 873666
rect 675758 872808 675814 872817
rect 675758 872743 675814 872752
rect 675772 872576 675800 872743
rect 674944 870046 675248 870074
rect 675312 870046 675418 870074
rect 675220 869938 675248 870046
rect 674852 869910 675156 869938
rect 675220 869910 675340 869938
rect 674760 869774 675064 869802
rect 674392 869638 674972 869666
rect 674656 869440 674708 869446
rect 674656 869382 674708 869388
rect 674668 867950 674696 869382
rect 674944 868170 674972 869638
rect 675036 868714 675064 869774
rect 675128 868889 675156 869910
rect 675312 869530 675340 869910
rect 675312 869502 675418 869530
rect 675128 868861 675418 868889
rect 675036 868686 675248 868714
rect 675220 868238 675248 868686
rect 675220 868210 675418 868238
rect 674944 868142 675064 868170
rect 674840 868080 674892 868086
rect 674840 868022 674892 868028
rect 674656 867944 674708 867950
rect 674656 867886 674708 867892
rect 674852 865858 674880 868022
rect 675036 867049 675064 868142
rect 675208 867944 675260 867950
rect 675208 867886 675260 867892
rect 675220 867694 675248 867886
rect 675220 867666 675418 867694
rect 675036 867021 675418 867049
rect 674852 865830 675418 865858
rect 675298 865736 675354 865745
rect 675298 865671 675354 865680
rect 675312 863818 675340 865671
rect 675758 865464 675814 865473
rect 675758 865399 675814 865408
rect 675772 865195 675800 865399
rect 675666 864920 675722 864929
rect 675666 864855 675722 864864
rect 675680 864552 675708 864855
rect 675312 863790 675432 863818
rect 675404 863328 675432 863790
rect 675392 790832 675444 790838
rect 675392 790774 675444 790780
rect 675404 788868 675432 790774
rect 675772 788089 675800 788324
rect 675758 788080 675814 788089
rect 675758 788015 675814 788024
rect 675128 787665 675418 787693
rect 675128 786729 675156 787665
rect 675404 786729 675432 787032
rect 675114 786720 675170 786729
rect 675114 786655 675170 786664
rect 675390 786720 675446 786729
rect 675390 786655 675446 786664
rect 674944 785182 675418 785210
rect 673920 782672 673972 782678
rect 673920 782614 673972 782620
rect 673642 780056 673698 780065
rect 673642 779991 673698 780000
rect 673656 746594 673684 779991
rect 673656 746566 673776 746594
rect 673460 738676 673512 738682
rect 673460 738618 673512 738624
rect 673472 735162 673500 738618
rect 673380 735134 673500 735162
rect 673380 734754 673408 735134
rect 673380 734726 673500 734754
rect 673274 728376 673330 728385
rect 673092 728340 673144 728346
rect 673274 728311 673330 728320
rect 673092 728282 673144 728288
rect 672998 728104 673054 728113
rect 672998 728039 673054 728048
rect 673012 723134 673040 728039
rect 673472 724418 673500 734726
rect 673748 734174 673776 746566
rect 673932 734210 673960 782614
rect 674944 779714 674972 785182
rect 675128 784638 675418 784666
rect 675128 784310 675156 784638
rect 675116 784304 675168 784310
rect 675116 784246 675168 784252
rect 675392 784168 675444 784174
rect 675392 784110 675444 784116
rect 675404 783972 675432 784110
rect 675128 783346 675418 783374
rect 675128 782678 675156 783346
rect 675116 782672 675168 782678
rect 675116 782614 675168 782620
rect 675300 782536 675352 782542
rect 675300 782478 675352 782484
rect 675312 781402 675340 782478
rect 675312 781374 675432 781402
rect 675208 781108 675260 781114
rect 675208 781050 675260 781056
rect 675220 779714 675248 781050
rect 675404 780844 675432 781374
rect 675496 780065 675524 780300
rect 675482 780056 675538 780065
rect 675482 779991 675538 780000
rect 674944 779686 675156 779714
rect 675220 779686 675340 779714
rect 674470 779240 674526 779249
rect 674470 779175 674526 779184
rect 674286 778832 674342 778841
rect 674286 778767 674342 778776
rect 674102 734496 674158 734505
rect 674102 734431 674158 734440
rect 673932 734182 674052 734210
rect 673656 734146 673776 734174
rect 673656 732794 673684 734146
rect 673564 732766 673684 732794
rect 673564 727954 673592 732766
rect 673828 730516 673880 730522
rect 673828 730458 673880 730464
rect 673564 727926 673684 727954
rect 673472 724390 673592 724418
rect 673368 724260 673420 724266
rect 673368 724202 673420 724208
rect 673380 723194 673408 724202
rect 673380 723166 673500 723194
rect 673012 723106 673316 723134
rect 673288 721754 673316 723106
rect 673104 721726 673316 721754
rect 672828 717586 672948 717614
rect 672552 715006 672856 715034
rect 672630 714912 672686 714921
rect 672630 714847 672686 714856
rect 672644 670177 672672 714847
rect 672828 711657 672856 715006
rect 672920 713538 672948 717586
rect 673104 713697 673132 721726
rect 673274 714096 673330 714105
rect 673274 714031 673330 714040
rect 673090 713688 673146 713697
rect 673090 713623 673146 713632
rect 672920 713510 673040 713538
rect 672814 711648 672870 711657
rect 672814 711583 672870 711592
rect 673012 708393 673040 713510
rect 672998 708384 673054 708393
rect 672998 708319 673054 708328
rect 673288 698294 673316 714031
rect 673196 698266 673316 698294
rect 672814 686216 672870 686225
rect 672814 686151 672870 686160
rect 672630 670168 672686 670177
rect 672630 670103 672686 670112
rect 672448 665168 672500 665174
rect 672448 665110 672500 665116
rect 672276 649966 672396 649994
rect 671816 637546 671936 637574
rect 672000 647206 672120 647234
rect 671816 630674 671844 637546
rect 672000 636206 672028 647206
rect 671988 636200 672040 636206
rect 671988 636142 672040 636148
rect 672172 636200 672224 636206
rect 672172 636142 672224 636148
rect 672184 634814 672212 636142
rect 672092 634786 672212 634814
rect 671816 630646 671936 630674
rect 671908 630086 671936 630646
rect 672092 630306 672120 634786
rect 672092 630278 672212 630306
rect 671896 630080 671948 630086
rect 671896 630022 671948 630028
rect 672184 629490 672212 630278
rect 671816 629462 672212 629490
rect 671816 615494 671844 629462
rect 672080 629400 672132 629406
rect 672080 629342 672132 629348
rect 672092 628946 672120 629342
rect 672000 628918 672120 628946
rect 672000 622849 672028 628918
rect 672172 625592 672224 625598
rect 672170 625560 672172 625569
rect 672224 625560 672226 625569
rect 672170 625495 672226 625504
rect 671986 622840 672042 622849
rect 671986 622775 672042 622784
rect 672368 621014 672396 649966
rect 672630 649224 672686 649233
rect 672630 649159 672686 649168
rect 672644 623098 672672 649159
rect 672828 626498 672856 686151
rect 673000 685976 673052 685982
rect 673000 685918 673052 685924
rect 673012 685817 673040 685918
rect 672998 685808 673054 685817
rect 672998 685743 673054 685752
rect 673196 669905 673224 698266
rect 673472 673454 673500 723166
rect 673564 692774 673592 724390
rect 673656 708914 673684 727926
rect 673840 724402 673868 730458
rect 674024 724520 674052 734182
rect 674116 724690 674144 734431
rect 674300 726510 674328 778767
rect 674484 726714 674512 779175
rect 674932 778388 674984 778394
rect 674932 778330 674984 778336
rect 674944 777073 674972 778330
rect 674930 777064 674986 777073
rect 674930 776999 674986 777008
rect 674930 775704 674986 775713
rect 674930 775639 674932 775648
rect 674984 775639 674986 775648
rect 674932 775610 674984 775616
rect 675128 746594 675156 779686
rect 675312 778478 675340 779686
rect 675496 779249 675524 779688
rect 675482 779240 675538 779249
rect 675482 779175 675538 779184
rect 675496 778841 675524 779008
rect 675482 778832 675538 778841
rect 675482 778767 675538 778776
rect 675312 778450 675418 778478
rect 675404 777481 675432 777852
rect 675390 777472 675446 777481
rect 675390 777407 675446 777416
rect 675482 777064 675538 777073
rect 675300 777028 675352 777034
rect 675482 776999 675538 777008
rect 675300 776970 675352 776976
rect 675312 776914 675340 776970
rect 675220 776886 675340 776914
rect 675220 775350 675248 776886
rect 675496 776628 675524 776999
rect 675404 775713 675432 776016
rect 675390 775704 675446 775713
rect 675390 775639 675446 775648
rect 675220 775322 675418 775350
rect 675404 773650 675432 774180
rect 675312 773622 675432 773650
rect 675312 773430 675340 773622
rect 675300 773424 675352 773430
rect 675300 773366 675352 773372
rect 674944 746566 675156 746594
rect 675392 746632 675444 746638
rect 675392 746574 675444 746580
rect 674944 739922 674972 746566
rect 675116 743912 675168 743918
rect 675116 743854 675168 743860
rect 675128 742030 675156 743854
rect 675404 743852 675432 746574
rect 675312 743294 675418 743322
rect 675312 742529 675340 743294
rect 675298 742520 675354 742529
rect 675298 742455 675354 742464
rect 675496 742218 675524 742696
rect 675484 742212 675536 742218
rect 675484 742154 675536 742160
rect 675312 742070 675432 742098
rect 675312 742030 675340 742070
rect 675128 742002 675340 742030
rect 675404 742016 675432 742070
rect 674944 739894 675064 739922
rect 674840 739832 674892 739838
rect 674840 739774 674892 739780
rect 674654 735040 674710 735049
rect 674654 734975 674710 734984
rect 674668 730522 674696 734975
rect 674852 734174 674880 739774
rect 674852 734146 674972 734174
rect 674944 733530 674972 734146
rect 674852 733502 674972 733530
rect 674656 730516 674708 730522
rect 674656 730458 674708 730464
rect 674852 730365 674880 733502
rect 674668 730337 674880 730365
rect 674668 729881 674696 730337
rect 675036 730266 675064 739894
rect 675404 739838 675432 740180
rect 675392 739832 675444 739838
rect 675392 739774 675444 739780
rect 675312 739622 675418 739650
rect 675312 739158 675340 739622
rect 675300 739152 675352 739158
rect 675300 739094 675352 739100
rect 675404 738682 675432 739024
rect 675392 738676 675444 738682
rect 675392 738618 675444 738624
rect 675312 738330 675418 738358
rect 675312 738177 675340 738330
rect 675298 738168 675354 738177
rect 675298 738103 675354 738112
rect 675300 737996 675352 738002
rect 675300 737938 675352 737944
rect 675312 735842 675340 737938
rect 675404 735842 675432 735896
rect 675312 735814 675432 735842
rect 675208 735752 675260 735758
rect 675208 735694 675260 735700
rect 675220 734346 675248 735694
rect 675404 735049 675432 735319
rect 675390 735040 675446 735049
rect 675390 734975 675446 734984
rect 675404 734505 675432 734672
rect 675390 734496 675446 734505
rect 675390 734431 675446 734440
rect 675128 734318 675248 734346
rect 675128 733493 675156 734318
rect 675300 734188 675352 734194
rect 675300 734130 675352 734136
rect 675312 733718 675340 734130
rect 675496 733825 675524 734031
rect 675482 733816 675538 733825
rect 675482 733751 675538 733760
rect 675300 733712 675352 733718
rect 675300 733654 675352 733660
rect 675128 733465 675418 733493
rect 675300 733372 675352 733378
rect 675300 733314 675352 733320
rect 675312 732034 675340 733314
rect 675496 732737 675524 732836
rect 675482 732728 675538 732737
rect 675482 732663 675538 732672
rect 675312 732006 675432 732034
rect 675404 731612 675432 732006
rect 675312 730986 675418 731014
rect 675312 730522 675340 730986
rect 675300 730516 675352 730522
rect 675300 730458 675352 730464
rect 674852 730238 675064 730266
rect 675128 730337 675418 730365
rect 674654 729872 674710 729881
rect 674654 729807 674710 729816
rect 674852 727274 674880 730238
rect 675128 730153 675156 730337
rect 675114 730144 675170 730153
rect 675114 730079 675170 730088
rect 675298 730144 675354 730153
rect 675298 730079 675354 730088
rect 675024 729904 675076 729910
rect 675024 729846 675076 729852
rect 675036 727274 675064 729846
rect 674760 727258 674880 727274
rect 674748 727252 674880 727258
rect 674800 727246 674880 727252
rect 674944 727246 675064 727274
rect 674748 727194 674800 727200
rect 674472 726708 674524 726714
rect 674472 726650 674524 726656
rect 674288 726504 674340 726510
rect 674288 726446 674340 726452
rect 674116 724662 674328 724690
rect 674024 724492 674144 724520
rect 673828 724396 673880 724402
rect 673828 724338 673880 724344
rect 673826 724160 673882 724169
rect 673826 724095 673882 724104
rect 673840 723134 673868 724095
rect 674116 723134 674144 724492
rect 674300 724169 674328 724662
rect 674286 724160 674342 724169
rect 674286 724095 674342 724104
rect 674944 723217 674972 727246
rect 674930 723208 674986 723217
rect 674930 723143 674986 723152
rect 673748 723106 673868 723134
rect 673932 723106 674144 723134
rect 673748 714854 673776 723106
rect 673932 717614 673960 723106
rect 675312 721750 675340 730079
rect 675496 728793 675524 729164
rect 675482 728784 675538 728793
rect 675482 728719 675538 728728
rect 681004 727252 681056 727258
rect 681004 727194 681056 727200
rect 675300 721744 675352 721750
rect 675300 721686 675352 721692
rect 675300 721268 675352 721274
rect 675300 721210 675352 721216
rect 675312 720866 675340 721210
rect 675300 720860 675352 720866
rect 675300 720802 675352 720808
rect 675300 720520 675352 720526
rect 675300 720462 675352 720468
rect 673932 717586 674696 717614
rect 674288 716508 674340 716514
rect 674288 716450 674340 716456
rect 674300 716394 674328 716450
rect 674024 716366 674328 716394
rect 674024 716310 674052 716366
rect 674012 716304 674064 716310
rect 674012 716246 674064 716252
rect 674012 715760 674064 715766
rect 674010 715728 674012 715737
rect 674064 715728 674066 715737
rect 674010 715663 674066 715672
rect 674012 715488 674064 715494
rect 674288 715488 674340 715494
rect 674064 715436 674288 715442
rect 674012 715430 674340 715436
rect 674024 715414 674328 715430
rect 674288 715352 674340 715358
rect 674024 715300 674288 715306
rect 674024 715294 674340 715300
rect 674024 715278 674328 715294
rect 674024 714950 674052 715278
rect 674012 714944 674064 714950
rect 674012 714886 674064 714892
rect 673748 714826 673868 714854
rect 673840 709345 673868 714826
rect 674012 714536 674064 714542
rect 674010 714504 674012 714513
rect 674064 714504 674066 714513
rect 674010 714439 674066 714448
rect 674010 713280 674066 713289
rect 674010 713215 674012 713224
rect 674064 713215 674066 713224
rect 674012 713186 674064 713192
rect 674012 712904 674064 712910
rect 674010 712872 674012 712881
rect 674064 712872 674066 712881
rect 674010 712807 674066 712816
rect 674010 712464 674066 712473
rect 674010 712399 674012 712408
rect 674064 712399 674066 712408
rect 674012 712370 674064 712376
rect 674012 710048 674064 710054
rect 674010 710016 674012 710025
rect 674064 710016 674066 710025
rect 674010 709951 674066 709960
rect 674288 709504 674340 709510
rect 674024 709452 674288 709458
rect 674024 709446 674340 709452
rect 674024 709430 674328 709446
rect 674024 709374 674052 709430
rect 674012 709368 674064 709374
rect 673826 709336 673882 709345
rect 674012 709310 674064 709316
rect 673826 709271 673882 709280
rect 674012 709232 674064 709238
rect 674010 709200 674012 709209
rect 674064 709200 674066 709209
rect 674010 709135 674066 709144
rect 673656 708886 674052 708914
rect 674024 707169 674052 708886
rect 674668 707606 674696 717586
rect 675312 712065 675340 720462
rect 676034 716544 676090 716553
rect 676034 716479 676036 716488
rect 676088 716479 676090 716488
rect 676036 716450 676088 716456
rect 676034 716136 676090 716145
rect 676034 716071 676090 716080
rect 675852 715488 675904 715494
rect 675852 715430 675904 715436
rect 675864 715329 675892 715430
rect 676048 715358 676076 716071
rect 676036 715352 676088 715358
rect 675850 715320 675906 715329
rect 676036 715294 676088 715300
rect 675850 715255 675906 715264
rect 675298 712056 675354 712065
rect 675298 711991 675354 712000
rect 681016 710841 681044 727194
rect 684132 726708 684184 726714
rect 684132 726650 684184 726656
rect 682382 726608 682438 726617
rect 682382 726543 682438 726552
rect 682396 711249 682424 726543
rect 683488 726436 683540 726442
rect 683488 726378 683540 726384
rect 683302 726336 683358 726345
rect 683302 726271 683358 726280
rect 682382 711240 682438 711249
rect 682382 711175 682438 711184
rect 681002 710832 681058 710841
rect 681002 710767 681058 710776
rect 676034 710424 676090 710433
rect 676034 710359 676090 710368
rect 676048 709510 676076 710359
rect 683316 709617 683344 726271
rect 683302 709608 683358 709617
rect 683302 709543 683358 709552
rect 676036 709504 676088 709510
rect 676036 709446 676088 709452
rect 674656 707600 674708 707606
rect 676036 707600 676088 707606
rect 674656 707542 674708 707548
rect 676034 707568 676036 707577
rect 676088 707568 676090 707577
rect 676034 707503 676090 707512
rect 674010 707160 674066 707169
rect 674010 707095 674066 707104
rect 673826 707024 673882 707033
rect 673826 706959 673882 706968
rect 673840 705194 673868 706959
rect 683500 706761 683528 726378
rect 684144 707985 684172 726650
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 684130 707976 684186 707985
rect 684130 707911 684186 707920
rect 683486 706752 683542 706761
rect 683486 706687 683542 706696
rect 676034 706344 676090 706353
rect 676034 706279 676090 706288
rect 674012 705968 674064 705974
rect 674064 705916 674512 705922
rect 674012 705910 674512 705916
rect 674024 705894 674512 705910
rect 674288 705832 674340 705838
rect 674024 705780 674288 705786
rect 674024 705774 674340 705780
rect 674024 705758 674328 705774
rect 674024 705226 674052 705758
rect 674484 705362 674512 705894
rect 676048 705838 676076 706279
rect 676036 705832 676088 705838
rect 676036 705774 676088 705780
rect 683118 705528 683174 705537
rect 683118 705463 683174 705472
rect 683132 705362 683160 705463
rect 674472 705356 674524 705362
rect 674472 705298 674524 705304
rect 683120 705356 683172 705362
rect 683120 705298 683172 705304
rect 673748 705166 673868 705194
rect 674012 705220 674064 705226
rect 673748 692774 673776 705166
rect 674012 705162 674064 705168
rect 676034 705120 676090 705129
rect 676034 705055 676090 705064
rect 676048 704070 676076 705055
rect 674288 704064 674340 704070
rect 674024 704012 674288 704018
rect 674024 704006 674340 704012
rect 676036 704064 676088 704070
rect 676036 704006 676088 704012
rect 674024 703990 674328 704006
rect 674024 703866 674052 703990
rect 674012 703860 674064 703866
rect 674012 703802 674064 703808
rect 674012 701208 674064 701214
rect 674064 701156 674328 701162
rect 674012 701150 674328 701156
rect 674024 701146 674328 701150
rect 674024 701140 674340 701146
rect 674024 701134 674288 701140
rect 674288 701082 674340 701088
rect 675392 701140 675444 701146
rect 675392 701082 675444 701088
rect 674012 701072 674064 701078
rect 674064 701020 674880 701026
rect 674012 701014 674880 701020
rect 674024 700998 674880 701014
rect 674852 698337 674880 700998
rect 675404 698875 675432 701082
rect 674852 698309 675418 698337
rect 675312 697666 675418 697694
rect 674012 696992 674064 696998
rect 674288 696992 674340 696998
rect 674064 696940 674288 696946
rect 674012 696934 674340 696940
rect 675116 696992 675168 696998
rect 675312 696969 675340 697666
rect 675116 696934 675168 696940
rect 675298 696960 675354 696969
rect 674024 696918 674328 696934
rect 675128 695209 675156 696934
rect 675298 696895 675354 696904
rect 675496 696833 675524 697035
rect 675482 696824 675538 696833
rect 675482 696759 675538 696768
rect 675128 695181 675418 695209
rect 675312 694742 675432 694770
rect 675114 694648 675170 694657
rect 675312 694634 675340 694742
rect 675170 694606 675340 694634
rect 675404 694620 675432 694742
rect 675114 694583 675170 694592
rect 674576 693994 675418 694022
rect 674288 693184 674340 693190
rect 674024 693132 674288 693138
rect 674024 693126 674340 693132
rect 674024 693122 674328 693126
rect 674012 693116 674328 693122
rect 674064 693110 674328 693116
rect 674012 693058 674064 693064
rect 674288 693048 674340 693054
rect 674288 692990 674340 692996
rect 674300 692774 674328 692990
rect 673564 692746 673684 692774
rect 673748 692746 673868 692774
rect 673656 682825 673684 692746
rect 673642 682816 673698 682825
rect 673642 682751 673698 682760
rect 673840 682666 673868 692746
rect 674208 692746 674328 692774
rect 674010 690160 674066 690169
rect 674010 690095 674012 690104
rect 674064 690095 674066 690104
rect 674012 690066 674064 690072
rect 674012 688832 674064 688838
rect 674010 688800 674012 688809
rect 674064 688800 674066 688809
rect 674010 688735 674066 688744
rect 674208 683114 674236 692746
rect 674576 690146 674604 693994
rect 675116 693184 675168 693190
rect 675496 693138 675524 693328
rect 675116 693126 675168 693132
rect 675128 690894 675156 693126
rect 675404 693110 675524 693138
rect 675404 693054 675432 693110
rect 675392 693048 675444 693054
rect 675392 692990 675444 692996
rect 675128 690866 675418 690894
rect 675128 690322 675340 690350
rect 674930 690160 674986 690169
rect 674576 690118 674696 690146
rect 674472 690056 674524 690062
rect 674472 689998 674524 690004
rect 674484 686746 674512 689998
rect 674668 689194 674696 690118
rect 674930 690095 674986 690104
rect 674944 689330 674972 690095
rect 675128 690062 675156 690322
rect 675312 690282 675340 690322
rect 675404 690282 675432 690336
rect 675312 690254 675432 690282
rect 675116 690056 675168 690062
rect 675116 689998 675168 690004
rect 675312 689710 675432 689738
rect 675312 689670 675340 689710
rect 675128 689642 675340 689670
rect 675404 689656 675432 689710
rect 675128 689489 675156 689642
rect 675114 689480 675170 689489
rect 675114 689415 675170 689424
rect 674944 689302 675064 689330
rect 673748 682638 673868 682666
rect 673932 683086 674236 683114
rect 674300 686718 674512 686746
rect 674576 689166 674696 689194
rect 673748 682009 673776 682638
rect 673734 682000 673790 682009
rect 673734 681935 673790 681944
rect 673472 673426 673592 673454
rect 673182 669896 673238 669905
rect 673182 669831 673238 669840
rect 673368 669384 673420 669390
rect 673368 669326 673420 669332
rect 673380 669225 673408 669326
rect 673366 669216 673422 669225
rect 673366 669151 673422 669160
rect 673368 665168 673420 665174
rect 673368 665110 673420 665116
rect 673380 664057 673408 665110
rect 673366 664048 673422 664057
rect 673366 663983 673422 663992
rect 673368 663468 673420 663474
rect 673368 663410 673420 663416
rect 673380 662969 673408 663410
rect 673366 662960 673422 662969
rect 673366 662895 673422 662904
rect 673564 662017 673592 673426
rect 673734 671392 673790 671401
rect 673734 671327 673736 671336
rect 673788 671327 673790 671336
rect 673736 671298 673788 671304
rect 673736 671152 673788 671158
rect 673736 671094 673788 671100
rect 673748 670993 673776 671094
rect 673734 670984 673790 670993
rect 673734 670919 673790 670928
rect 673734 670576 673790 670585
rect 673734 670511 673790 670520
rect 673748 669526 673776 670511
rect 673736 669520 673788 669526
rect 673736 669462 673788 669468
rect 673734 668944 673790 668953
rect 673734 668879 673790 668888
rect 673748 668710 673776 668879
rect 673736 668704 673788 668710
rect 673736 668646 673788 668652
rect 673736 668568 673788 668574
rect 673734 668536 673736 668545
rect 673788 668536 673790 668545
rect 673734 668471 673790 668480
rect 673734 668128 673790 668137
rect 673734 668063 673790 668072
rect 673748 667962 673776 668063
rect 673736 667956 673788 667962
rect 673736 667898 673788 667904
rect 673734 667720 673790 667729
rect 673734 667655 673790 667664
rect 673748 667350 673776 667655
rect 673736 667344 673788 667350
rect 673736 667286 673788 667292
rect 673736 667208 673788 667214
rect 673736 667150 673788 667156
rect 673748 666913 673776 667150
rect 673734 666904 673790 666913
rect 673734 666839 673790 666848
rect 673734 666632 673790 666641
rect 673734 666567 673736 666576
rect 673788 666567 673790 666576
rect 673736 666538 673788 666544
rect 673736 665304 673788 665310
rect 673734 665272 673736 665281
rect 673788 665272 673790 665281
rect 673734 665207 673790 665216
rect 673734 664456 673790 664465
rect 673734 664391 673736 664400
rect 673788 664391 673790 664400
rect 673736 664362 673788 664368
rect 673736 663944 673788 663950
rect 673736 663886 673788 663892
rect 673748 663785 673776 663886
rect 673734 663776 673790 663785
rect 673734 663711 673790 663720
rect 673550 662008 673606 662017
rect 673550 661943 673606 661952
rect 673736 661632 673788 661638
rect 673734 661600 673736 661609
rect 673788 661600 673790 661609
rect 673734 661535 673790 661544
rect 673734 661192 673790 661201
rect 673734 661127 673736 661136
rect 673788 661127 673790 661136
rect 673736 661098 673788 661104
rect 673736 660136 673788 660142
rect 673734 660104 673736 660113
rect 673788 660104 673790 660113
rect 673734 660039 673790 660048
rect 673366 659696 673422 659705
rect 673366 659631 673422 659640
rect 672998 648816 673054 648825
rect 672998 648751 673054 648760
rect 673012 630674 673040 648751
rect 673182 645280 673238 645289
rect 673182 645215 673238 645224
rect 673012 630646 673132 630674
rect 672828 626470 673040 626498
rect 672814 626376 672870 626385
rect 672814 626311 672870 626320
rect 672828 626142 672856 626311
rect 672816 626136 672868 626142
rect 672816 626078 672868 626084
rect 672814 625968 672870 625977
rect 672814 625903 672870 625912
rect 672828 625190 672856 625903
rect 672816 625184 672868 625190
rect 672816 625126 672868 625132
rect 672816 625048 672868 625054
rect 672814 625016 672816 625025
rect 672868 625016 672870 625025
rect 672814 624951 672870 624960
rect 672814 624744 672870 624753
rect 672814 624679 672816 624688
rect 672868 624679 672870 624688
rect 672816 624650 672868 624656
rect 672816 624368 672868 624374
rect 672814 624336 672816 624345
rect 672868 624336 672870 624345
rect 672814 624271 672870 624280
rect 672814 623928 672870 623937
rect 672814 623863 672816 623872
rect 672868 623863 672870 623872
rect 672816 623834 672868 623840
rect 672816 623552 672868 623558
rect 672814 623520 672816 623529
rect 672868 623520 672870 623529
rect 672814 623455 672870 623464
rect 672276 620986 672396 621014
rect 672552 623070 672672 623098
rect 672814 623112 672870 623121
rect 672552 621014 672580 623070
rect 672814 623047 672816 623056
rect 672868 623047 672870 623056
rect 672816 623018 672868 623024
rect 673012 622962 673040 626470
rect 672920 622934 673040 622962
rect 672920 621489 672948 622934
rect 672906 621480 672962 621489
rect 672906 621415 672962 621424
rect 672816 621104 672868 621110
rect 672814 621072 672816 621081
rect 672868 621072 672870 621081
rect 672552 620986 672672 621014
rect 672814 621007 672870 621016
rect 673104 621014 673132 630646
rect 672276 618497 672304 620986
rect 672262 618488 672318 618497
rect 672262 618423 672318 618432
rect 671816 615466 672028 615494
rect 671724 611326 671844 611354
rect 671620 574592 671672 574598
rect 671620 574534 671672 574540
rect 671816 571470 671844 611326
rect 672000 574190 672028 615466
rect 672446 604480 672502 604489
rect 672446 604415 672502 604424
rect 672264 584452 672316 584458
rect 672264 584394 672316 584400
rect 671988 574184 672040 574190
rect 671988 574126 672040 574132
rect 672276 574054 672304 584394
rect 672460 579614 672488 604415
rect 672644 584458 672672 620986
rect 673012 620986 673132 621014
rect 672816 620288 672868 620294
rect 672814 620256 672816 620265
rect 672868 620256 672870 620265
rect 672814 620191 672870 620200
rect 672816 620016 672868 620022
rect 672814 619984 672816 619993
rect 672868 619984 672870 619993
rect 672814 619919 672870 619928
rect 672816 619744 672868 619750
rect 672814 619712 672816 619721
rect 672868 619712 672870 619721
rect 672814 619647 672870 619656
rect 673012 611354 673040 620986
rect 673196 611354 673224 645215
rect 672920 611326 673040 611354
rect 673104 611326 673224 611354
rect 672920 606506 672948 611326
rect 672920 606478 673040 606506
rect 672814 597408 672870 597417
rect 672814 597343 672870 597352
rect 672632 584452 672684 584458
rect 672632 584394 672684 584400
rect 672828 582374 672856 597343
rect 672736 582346 672856 582374
rect 672736 581346 672764 582346
rect 672644 581318 672764 581346
rect 672460 579586 672580 579614
rect 672264 574048 672316 574054
rect 672264 573990 672316 573996
rect 672552 572714 672580 579586
rect 672644 573730 672672 581318
rect 673012 580938 673040 606478
rect 673104 601746 673132 611326
rect 673380 608594 673408 659631
rect 673734 655616 673790 655625
rect 673734 655551 673736 655560
rect 673788 655551 673790 655560
rect 673736 655522 673788 655528
rect 673734 645960 673790 645969
rect 673734 645895 673736 645904
rect 673788 645895 673790 645904
rect 673736 645866 673788 645872
rect 673550 643512 673606 643521
rect 673550 643447 673606 643456
rect 673564 642649 673592 643447
rect 673736 643136 673788 643142
rect 673734 643104 673736 643113
rect 673788 643104 673790 643113
rect 673734 643039 673790 643048
rect 673564 642621 673776 642649
rect 673550 642424 673606 642433
rect 673550 642359 673606 642368
rect 673564 615494 673592 642359
rect 673748 615494 673776 642621
rect 673932 618338 673960 683086
rect 674102 644600 674158 644609
rect 674102 644535 674158 644544
rect 674116 642433 674144 644535
rect 674102 642424 674158 642433
rect 674102 642359 674158 642368
rect 674102 641744 674158 641753
rect 674102 641679 674158 641688
rect 674116 619562 674144 641679
rect 674300 636886 674328 686718
rect 674576 683114 674604 689166
rect 674748 689036 674800 689042
rect 674748 688978 674800 688984
rect 674760 683114 674788 688978
rect 675036 688922 675064 689302
rect 675220 689042 675418 689058
rect 675208 689036 675418 689042
rect 675260 689030 675418 689036
rect 675208 688978 675260 688984
rect 675036 688894 675156 688922
rect 674930 688800 674986 688809
rect 674930 688735 674986 688744
rect 674944 686678 674972 688735
rect 675128 688514 675156 688894
rect 675128 688486 675340 688514
rect 675312 688378 675340 688486
rect 675404 688378 675432 688500
rect 675312 688350 675432 688378
rect 675128 687806 675418 687834
rect 675128 687721 675156 687806
rect 675114 687712 675170 687721
rect 675114 687647 675170 687656
rect 674944 686650 675340 686678
rect 675312 686610 675340 686650
rect 675404 686610 675432 686664
rect 675312 686582 675432 686610
rect 675114 686216 675170 686225
rect 675114 686151 675170 686160
rect 675128 685998 675156 686151
rect 675128 685970 675418 685998
rect 674930 685808 674986 685817
rect 674930 685743 674986 685752
rect 674944 684706 674972 685743
rect 675114 685536 675170 685545
rect 675114 685471 675170 685480
rect 675128 685386 675156 685471
rect 675128 685358 675340 685386
rect 675312 685250 675340 685358
rect 675404 685250 675432 685372
rect 675312 685222 675432 685250
rect 674944 684678 675432 684706
rect 675404 684148 675432 684678
rect 675114 684040 675170 684049
rect 675114 683975 675170 683984
rect 674484 683086 674604 683114
rect 674668 683086 674788 683114
rect 674484 637022 674512 683086
rect 674472 637016 674524 637022
rect 674472 636958 674524 636964
rect 674288 636880 674340 636886
rect 674288 636822 674340 636828
rect 674668 623082 674696 683086
rect 674838 682816 674894 682825
rect 674838 682751 674894 682760
rect 674852 682582 674880 682751
rect 674840 682576 674892 682582
rect 674840 682518 674892 682524
rect 674840 682440 674892 682446
rect 674840 682382 674892 682388
rect 674852 682009 674880 682382
rect 674838 682000 674894 682009
rect 674838 681935 674894 681944
rect 675128 676433 675156 683975
rect 675298 683768 675354 683777
rect 675298 683703 675354 683712
rect 675114 676424 675170 676433
rect 675114 676359 675170 676368
rect 674838 669896 674894 669905
rect 674838 669831 674840 669840
rect 674892 669831 674894 669840
rect 674840 669802 674892 669808
rect 675312 666505 675340 683703
rect 683212 682576 683264 682582
rect 683212 682518 683264 682524
rect 676496 669860 676548 669866
rect 676496 669802 676548 669808
rect 676508 669497 676536 669802
rect 676494 669488 676550 669497
rect 676494 669423 676550 669432
rect 675298 666496 675354 666505
rect 675298 666431 675354 666440
rect 676034 664864 676090 664873
rect 676034 664799 676090 664808
rect 676048 663814 676076 664799
rect 674840 663808 674892 663814
rect 674838 663776 674840 663785
rect 676036 663808 676088 663814
rect 674892 663776 674894 663785
rect 683224 663785 683252 682518
rect 683488 682440 683540 682446
rect 683488 682382 683540 682388
rect 684130 682408 684186 682417
rect 676036 663750 676088 663756
rect 683210 663776 683266 663785
rect 674838 663711 674894 663720
rect 683210 663711 683266 663720
rect 683500 662969 683528 682382
rect 684130 682343 684186 682352
rect 684144 666233 684172 682343
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 684130 666224 684186 666233
rect 684130 666159 684186 666168
rect 683486 662960 683542 662969
rect 683486 662895 683542 662904
rect 674838 660104 674894 660113
rect 674838 660039 674894 660048
rect 683118 660104 683174 660113
rect 683118 660039 683174 660048
rect 674852 659870 674880 660039
rect 683132 659870 683160 660039
rect 674840 659864 674892 659870
rect 674840 659806 674892 659812
rect 683120 659864 683172 659870
rect 683120 659806 683172 659812
rect 675114 655616 675170 655625
rect 675114 655551 675170 655560
rect 675128 653698 675156 655551
rect 675128 653670 675418 653698
rect 675404 652905 675432 653140
rect 675390 652896 675446 652905
rect 675390 652831 675446 652840
rect 675496 652089 675524 652460
rect 675482 652080 675538 652089
rect 675482 652015 675538 652024
rect 674852 651834 675418 651862
rect 674852 640422 674880 651834
rect 675404 649994 675432 650012
rect 674944 649966 675432 649994
rect 674944 643226 674972 649966
rect 675404 649233 675432 649468
rect 675390 649224 675446 649233
rect 675390 649159 675446 649168
rect 675114 648816 675170 648825
rect 675170 648774 675418 648802
rect 675114 648751 675170 648760
rect 675404 647873 675432 648176
rect 675390 647864 675446 647873
rect 675390 647799 675446 647808
rect 675114 645960 675170 645969
rect 675114 645895 675170 645904
rect 675128 643294 675156 645895
rect 675312 645646 675418 645674
rect 675312 645289 675340 645646
rect 675298 645280 675354 645289
rect 675298 645215 675354 645224
rect 675312 645102 675418 645130
rect 675312 644609 675340 645102
rect 675298 644600 675354 644609
rect 675298 644535 675354 644544
rect 675404 644337 675432 644475
rect 675390 644328 675446 644337
rect 675390 644263 675446 644272
rect 675312 643810 675418 643838
rect 675312 643521 675340 643810
rect 675298 643512 675354 643521
rect 675298 643447 675354 643456
rect 675128 643266 675418 643294
rect 674944 643198 675064 643226
rect 674840 640416 674892 640422
rect 674840 640358 674892 640364
rect 675036 640334 675064 643198
rect 675298 643104 675354 643113
rect 675128 643062 675298 643090
rect 675128 641458 675156 643062
rect 675298 643039 675354 643048
rect 675312 642621 675418 642649
rect 675312 641753 675340 642621
rect 675298 641744 675354 641753
rect 675298 641679 675354 641688
rect 675128 641430 675418 641458
rect 675312 640781 675418 640809
rect 675312 640506 675340 640781
rect 674944 640306 675064 640334
rect 675128 640478 675340 640506
rect 674944 635526 674972 640306
rect 674932 635520 674984 635526
rect 674932 635462 674984 635468
rect 674656 623076 674708 623082
rect 674656 623018 674708 623024
rect 674288 621036 674340 621042
rect 674288 620978 674340 620984
rect 674300 620809 674328 620978
rect 674286 620800 674342 620809
rect 674286 620735 674342 620744
rect 674380 619744 674432 619750
rect 674378 619712 674380 619721
rect 674432 619712 674434 619721
rect 674378 619647 674434 619656
rect 674116 619534 674512 619562
rect 674288 618520 674340 618526
rect 674286 618488 674288 618497
rect 674340 618488 674342 618497
rect 674286 618423 674342 618432
rect 673932 618310 674328 618338
rect 674300 618050 674328 618310
rect 674288 618044 674340 618050
rect 674288 617986 674340 617992
rect 674288 617908 674340 617914
rect 674288 617850 674340 617856
rect 674300 617794 674328 617850
rect 674024 617766 674328 617794
rect 674024 617506 674052 617766
rect 674012 617500 674064 617506
rect 674012 617442 674064 617448
rect 674288 617500 674340 617506
rect 674288 617442 674340 617448
rect 674300 617386 674328 617442
rect 674024 617358 674328 617386
rect 674024 616894 674052 617358
rect 674012 616888 674064 616894
rect 674012 616830 674064 616836
rect 674012 615664 674064 615670
rect 674012 615606 674064 615612
rect 674024 615516 674052 615606
rect 674288 615528 674340 615534
rect 673564 615466 673684 615494
rect 673748 615466 673868 615494
rect 674024 615488 674288 615516
rect 674288 615470 674340 615476
rect 673656 611354 673684 615466
rect 673288 608566 673408 608594
rect 673564 611326 673684 611354
rect 673288 603786 673316 608566
rect 673564 607306 673592 611326
rect 673552 607300 673604 607306
rect 673552 607242 673604 607248
rect 673552 607096 673604 607102
rect 673552 607038 673604 607044
rect 673288 603758 673500 603786
rect 673276 603560 673328 603566
rect 673276 603502 673328 603508
rect 673104 601718 673224 601746
rect 672828 580910 673040 580938
rect 672828 574818 672856 580910
rect 673196 580802 673224 601718
rect 672920 580774 673224 580802
rect 672920 579578 672948 580774
rect 673090 580680 673146 580689
rect 673090 580615 673146 580624
rect 673104 579698 673132 580615
rect 673092 579692 673144 579698
rect 673092 579634 673144 579640
rect 672920 579550 673040 579578
rect 673012 574977 673040 579550
rect 672998 574968 673054 574977
rect 672998 574903 673054 574912
rect 672828 574790 672948 574818
rect 672644 573702 672764 573730
rect 672460 572686 672580 572714
rect 672736 572714 672764 573702
rect 672920 573481 672948 574790
rect 673092 574048 673144 574054
rect 673092 573990 673144 573996
rect 673104 573753 673132 573990
rect 673090 573744 673146 573753
rect 673090 573679 673146 573688
rect 672906 573472 672962 573481
rect 672906 573407 672962 573416
rect 672736 572686 672856 572714
rect 671804 571464 671856 571470
rect 671804 571406 671856 571412
rect 671344 570444 671396 570450
rect 671344 570386 671396 570392
rect 671160 534608 671212 534614
rect 671160 534550 671212 534556
rect 671158 532128 671214 532137
rect 671158 532063 671214 532072
rect 670976 529304 671028 529310
rect 670976 529246 671028 529252
rect 670792 490952 670844 490958
rect 670792 490894 670844 490900
rect 671172 488510 671200 532063
rect 671160 488504 671212 488510
rect 671160 488446 671212 488452
rect 670606 455152 670662 455161
rect 670606 455087 670662 455096
rect 663062 403336 663118 403345
rect 663062 403271 663118 403280
rect 654782 382936 654838 382945
rect 654782 382871 654838 382880
rect 654796 371006 654824 382871
rect 663076 373998 663104 403271
rect 670514 392592 670570 392601
rect 670514 392527 670570 392536
rect 663064 373992 663116 373998
rect 663064 373934 663116 373940
rect 654784 371000 654836 371006
rect 654784 370942 654836 370948
rect 666466 365664 666522 365673
rect 666466 365599 666522 365608
rect 666480 364410 666508 365599
rect 662420 364404 662472 364410
rect 662420 364346 662472 364352
rect 666468 364404 666520 364410
rect 666468 364346 666520 364352
rect 662432 360262 662460 364346
rect 657544 360256 657596 360262
rect 657544 360198 657596 360204
rect 662420 360256 662472 360262
rect 662420 360198 662472 360204
rect 654782 358592 654838 358601
rect 654782 358527 654838 358536
rect 653586 338736 653642 338745
rect 653586 338671 653642 338680
rect 653600 325650 653628 338671
rect 654796 328302 654824 358527
rect 657556 348430 657584 360198
rect 657544 348424 657596 348430
rect 657544 348366 657596 348372
rect 669410 347304 669466 347313
rect 669410 347239 669466 347248
rect 654784 328296 654836 328302
rect 654784 328238 654836 328244
rect 653588 325644 653640 325650
rect 653588 325586 653640 325592
rect 653404 322992 653456 322998
rect 653404 322934 653456 322940
rect 653402 313304 653458 313313
rect 653402 313239 653458 313248
rect 652482 309904 652538 309913
rect 652482 309839 652538 309848
rect 652496 302161 652524 309839
rect 653416 303414 653444 313239
rect 658922 311944 658978 311953
rect 658922 311879 658978 311888
rect 653404 303408 653456 303414
rect 653404 303350 653456 303356
rect 652482 302152 652538 302161
rect 652482 302087 652538 302096
rect 658936 300830 658964 311879
rect 658924 300824 658976 300830
rect 658924 300766 658976 300772
rect 660580 298172 660632 298178
rect 660580 298114 660632 298120
rect 652298 297528 652354 297537
rect 652298 297463 652354 297472
rect 651760 296686 652064 296714
rect 651470 294264 651526 294273
rect 651470 294199 651526 294208
rect 651484 294030 651512 294199
rect 651472 294024 651524 294030
rect 651472 293966 651524 293972
rect 651470 293040 651526 293049
rect 651470 292975 651526 292984
rect 651484 292602 651512 292975
rect 651472 292596 651524 292602
rect 651472 292538 651524 292544
rect 651760 290834 651788 296686
rect 651930 295352 651986 295361
rect 651930 295287 651986 295296
rect 651944 291825 651972 295287
rect 651930 291816 651986 291825
rect 651930 291751 651986 291760
rect 652114 291544 652170 291553
rect 652114 291479 652170 291488
rect 651748 290828 651800 290834
rect 651748 290770 651800 290776
rect 651470 290456 651526 290465
rect 651470 290391 651526 290400
rect 651484 289882 651512 290391
rect 651472 289876 651524 289882
rect 651472 289818 651524 289824
rect 651654 289232 651710 289241
rect 651654 289167 651710 289176
rect 651470 288688 651526 288697
rect 651470 288623 651526 288632
rect 651484 288454 651512 288623
rect 651472 288448 651524 288454
rect 651472 288390 651524 288396
rect 651668 287745 651696 289167
rect 651654 287736 651710 287745
rect 651654 287671 651710 287680
rect 651470 287464 651526 287473
rect 651470 287399 651526 287408
rect 651484 287094 651512 287399
rect 651472 287088 651524 287094
rect 651472 287030 651524 287036
rect 652128 287054 652156 291479
rect 652312 287054 652340 297463
rect 658924 296744 658976 296750
rect 658924 296686 658976 296692
rect 652128 287026 652248 287054
rect 652312 287026 652616 287054
rect 651470 285968 651526 285977
rect 651470 285903 651526 285912
rect 651484 285734 651512 285903
rect 651472 285728 651524 285734
rect 651472 285670 651524 285676
rect 651470 284744 651526 284753
rect 651470 284679 651526 284688
rect 651484 284374 651512 284679
rect 651472 284368 651524 284374
rect 651472 284310 651524 284316
rect 651470 283384 651526 283393
rect 651470 283319 651526 283328
rect 651484 282946 651512 283319
rect 651472 282940 651524 282946
rect 651472 282882 651524 282888
rect 652022 282160 652078 282169
rect 652022 282095 652078 282104
rect 651470 280936 651526 280945
rect 651470 280871 651526 280880
rect 651484 280226 651512 280871
rect 651472 280220 651524 280226
rect 651472 280162 651524 280168
rect 650828 278452 650880 278458
rect 650828 278394 650880 278400
rect 650644 278180 650696 278186
rect 650644 278122 650696 278128
rect 636764 275466 636792 278052
rect 637684 278038 637974 278066
rect 636752 275460 636804 275466
rect 636752 275402 636804 275408
rect 637684 269822 637712 278038
rect 637856 277432 637908 277438
rect 637856 277374 637908 277380
rect 637672 269816 637724 269822
rect 637672 269758 637724 269764
rect 637868 229094 637896 277374
rect 639156 273970 639184 278052
rect 639144 273964 639196 273970
rect 639144 273906 639196 273912
rect 640352 272678 640380 278052
rect 640536 278038 641470 278066
rect 641732 278038 642666 278066
rect 640340 272672 640392 272678
rect 640340 272614 640392 272620
rect 640536 269958 640564 278038
rect 640524 269952 640576 269958
rect 640524 269894 640576 269900
rect 641732 268394 641760 278038
rect 643848 275330 643876 278052
rect 643836 275324 643888 275330
rect 643836 275266 643888 275272
rect 645044 271318 645072 278052
rect 645872 278038 646254 278066
rect 647252 278038 647450 278066
rect 645032 271312 645084 271318
rect 645032 271254 645084 271260
rect 641720 268388 641772 268394
rect 641720 268330 641772 268336
rect 645872 261526 645900 278038
rect 645860 261520 645912 261526
rect 645860 261462 645912 261468
rect 647252 246362 647280 278038
rect 647240 246356 647292 246362
rect 647240 246298 647292 246304
rect 648632 242214 648660 278052
rect 648620 242208 648672 242214
rect 648620 242150 648672 242156
rect 636212 229066 636516 229094
rect 637868 229066 638172 229094
rect 636488 210202 636516 229066
rect 638144 210202 638172 229066
rect 650642 225040 650698 225049
rect 650642 224975 650698 224984
rect 648620 220244 648672 220250
rect 648620 220186 648672 220192
rect 645858 219872 645914 219881
rect 645858 219807 645914 219816
rect 644940 215960 644992 215966
rect 644940 215902 644992 215908
rect 643836 213376 643888 213382
rect 643836 213318 643888 213324
rect 641720 212696 641772 212702
rect 641720 212638 641772 212644
rect 639880 212560 639932 212566
rect 639880 212502 639932 212508
rect 639892 210202 639920 212502
rect 641732 210202 641760 212638
rect 643848 210202 643876 213318
rect 644952 210202 644980 215902
rect 645872 213926 645900 219807
rect 648434 218648 648490 218657
rect 648434 218583 648490 218592
rect 648252 216708 648304 216714
rect 648252 216650 648304 216656
rect 646320 214600 646372 214606
rect 646320 214542 646372 214548
rect 645860 213920 645912 213926
rect 645860 213862 645912 213868
rect 645492 213172 645544 213178
rect 645492 213114 645544 213120
rect 645504 210202 645532 213114
rect 646332 210202 646360 214542
rect 646504 213920 646556 213926
rect 646504 213862 646556 213868
rect 625632 210174 625876 210202
rect 626092 210174 626428 210202
rect 626644 210174 626980 210202
rect 627104 210174 627532 210202
rect 627932 210174 628084 210202
rect 628300 210174 628636 210202
rect 628760 210174 629188 210202
rect 629404 210174 629740 210202
rect 629864 210174 630292 210202
rect 630692 210174 630844 210202
rect 630968 210174 631396 210202
rect 631520 210174 631948 210202
rect 632900 210174 633052 210202
rect 633452 210174 633604 210202
rect 633728 210174 634156 210202
rect 634372 210174 634708 210202
rect 635108 210174 635260 210202
rect 636488 210174 636916 210202
rect 638144 210174 638572 210202
rect 639892 210174 640228 210202
rect 641732 210174 641884 210202
rect 643540 210174 643876 210202
rect 644644 210174 644980 210202
rect 645196 210174 645532 210202
rect 646300 210174 646360 210202
rect 646516 210202 646544 213862
rect 648264 210202 648292 216650
rect 646516 210174 646852 210202
rect 647956 210174 648292 210202
rect 648448 210202 648476 218583
rect 648632 213450 648660 220186
rect 650656 216714 650684 224975
rect 651288 222896 651340 222902
rect 651288 222838 651340 222844
rect 651102 217832 651158 217841
rect 651102 217767 651158 217776
rect 650644 216708 650696 216714
rect 650644 216650 650696 216656
rect 648620 213444 648672 213450
rect 648620 213386 648672 213392
rect 649264 213444 649316 213450
rect 649264 213386 649316 213392
rect 649276 210202 649304 213386
rect 650460 212764 650512 212770
rect 650460 212706 650512 212712
rect 650472 210202 650500 212706
rect 648448 210174 648508 210202
rect 649276 210174 649612 210202
rect 650164 210174 650500 210202
rect 651116 210202 651144 217767
rect 651300 212770 651328 222838
rect 651470 221504 651526 221513
rect 651470 221439 651526 221448
rect 651288 212764 651340 212770
rect 651288 212706 651340 212712
rect 651484 210202 651512 221439
rect 651116 210174 651268 210202
rect 651484 210174 651820 210202
rect 600320 210112 600372 210118
rect 600320 210054 600372 210060
rect 600688 210112 600740 210118
rect 600740 210060 601036 210066
rect 600688 210054 601036 210060
rect 600700 210038 601036 210054
rect 652036 209574 652064 282095
rect 652220 233918 652248 287026
rect 652390 280392 652446 280401
rect 652390 280327 652446 280336
rect 652208 233912 652260 233918
rect 652208 233854 652260 233860
rect 652404 226953 652432 280327
rect 652588 279449 652616 287026
rect 652574 279440 652630 279449
rect 652574 279375 652630 279384
rect 658936 268161 658964 296686
rect 660592 293865 660620 298114
rect 664444 294024 664496 294030
rect 664444 293966 664496 293972
rect 660578 293856 660634 293865
rect 660578 293791 660634 293800
rect 660304 292596 660356 292602
rect 660304 292538 660356 292544
rect 658922 268152 658978 268161
rect 658922 268087 658978 268096
rect 660316 232558 660344 292538
rect 663064 289876 663116 289882
rect 663064 289818 663116 289824
rect 663076 232694 663104 289818
rect 664456 248305 664484 293966
rect 667756 287088 667808 287094
rect 667756 287030 667808 287036
rect 667572 285728 667624 285734
rect 667572 285670 667624 285676
rect 667204 282940 667256 282946
rect 667204 282882 667256 282888
rect 664442 248296 664498 248305
rect 664442 248231 664498 248240
rect 663064 232688 663116 232694
rect 663064 232630 663116 232636
rect 660304 232552 660356 232558
rect 660304 232494 660356 232500
rect 662512 231532 662564 231538
rect 662512 231474 662564 231480
rect 662328 229764 662380 229770
rect 662328 229706 662380 229712
rect 660948 229628 661000 229634
rect 660948 229570 661000 229576
rect 652390 226944 652446 226953
rect 652390 226879 652446 226888
rect 658922 226400 658978 226409
rect 658922 226335 658978 226344
rect 652758 225720 652814 225729
rect 652758 225655 652814 225664
rect 652772 220250 652800 225655
rect 656162 225312 656218 225321
rect 656162 225247 656218 225256
rect 654782 223952 654838 223961
rect 654782 223887 654838 223896
rect 653402 222864 653458 222873
rect 653402 222799 653458 222808
rect 652760 220244 652812 220250
rect 652760 220186 652812 220192
rect 653220 213784 653272 213790
rect 653220 213726 653272 213732
rect 653232 210202 653260 213726
rect 653416 213314 653444 222799
rect 654138 220416 654194 220425
rect 654138 220351 654194 220360
rect 653770 217560 653826 217569
rect 653770 217495 653826 217504
rect 653404 213308 653456 213314
rect 653404 213250 653456 213256
rect 653784 210202 653812 217495
rect 654152 213450 654180 220351
rect 654600 213920 654652 213926
rect 654600 213862 654652 213868
rect 654140 213444 654192 213450
rect 654140 213386 654192 213392
rect 654612 210202 654640 213862
rect 654796 213790 654824 223887
rect 656176 214606 656204 225247
rect 657542 223680 657598 223689
rect 657542 223615 657598 223624
rect 656806 218920 656862 218929
rect 656806 218855 656862 218864
rect 656164 214600 656216 214606
rect 656164 214542 656216 214548
rect 654784 213784 654836 213790
rect 654784 213726 654836 213732
rect 654784 213444 654836 213450
rect 654784 213386 654836 213392
rect 656532 213444 656584 213450
rect 656532 213386 656584 213392
rect 652924 210174 653260 210202
rect 653476 210174 653812 210202
rect 654580 210174 654640 210202
rect 654796 210202 654824 213386
rect 656544 210202 656572 213386
rect 656820 210202 656848 218855
rect 657556 213926 657584 223615
rect 658936 215966 658964 226335
rect 660762 221776 660818 221785
rect 660762 221711 660818 221720
rect 658924 215960 658976 215966
rect 658924 215902 658976 215908
rect 659566 215384 659622 215393
rect 659566 215319 659622 215328
rect 658188 214736 658240 214742
rect 658188 214678 658240 214684
rect 657544 213920 657596 213926
rect 657544 213862 657596 213868
rect 658200 210202 658228 214678
rect 658738 213208 658794 213217
rect 658738 213143 658794 213152
rect 658752 210202 658780 213143
rect 659580 210202 659608 215319
rect 660394 214568 660450 214577
rect 660394 214503 660450 214512
rect 660408 210202 660436 214503
rect 660776 213246 660804 221711
rect 660764 213240 660816 213246
rect 660764 213182 660816 213188
rect 660960 210202 660988 229570
rect 662142 228576 662198 228585
rect 662142 228511 662198 228520
rect 661498 213480 661554 213489
rect 661498 213415 661554 213424
rect 661512 210202 661540 213415
rect 662156 210202 662184 228511
rect 662340 210202 662368 229706
rect 662524 229634 662552 231474
rect 665088 230988 665140 230994
rect 665088 230930 665140 230936
rect 664902 230480 664958 230489
rect 664902 230415 664958 230424
rect 662512 229628 662564 229634
rect 662512 229570 662564 229576
rect 663706 229120 663762 229129
rect 663706 229055 663762 229064
rect 663432 226364 663484 226370
rect 663432 226306 663484 226312
rect 663156 213920 663208 213926
rect 663156 213862 663208 213868
rect 663168 210202 663196 213862
rect 663444 210202 663472 226306
rect 663720 213926 663748 229055
rect 664626 215656 664682 215665
rect 664626 215591 664682 215600
rect 663708 213920 663760 213926
rect 663708 213862 663760 213868
rect 664640 213450 664668 215591
rect 664628 213444 664680 213450
rect 664628 213386 664680 213392
rect 664260 212764 664312 212770
rect 664260 212706 664312 212712
rect 664272 210202 664300 212706
rect 664916 210202 664944 230415
rect 665100 212770 665128 230930
rect 665272 230648 665324 230654
rect 665272 230590 665324 230596
rect 665284 226370 665312 230590
rect 665272 226364 665324 226370
rect 665272 226306 665324 226312
rect 667018 225992 667074 226001
rect 667018 225927 667074 225936
rect 667032 225321 667060 225927
rect 667018 225312 667074 225321
rect 667018 225247 667074 225256
rect 666468 225208 666520 225214
rect 666468 225150 666520 225156
rect 666480 222902 666508 225150
rect 666468 222896 666520 222902
rect 665822 222864 665878 222873
rect 666468 222838 666520 222844
rect 665822 222799 665878 222808
rect 665836 214742 665864 222799
rect 666650 219464 666706 219473
rect 666650 219399 666706 219408
rect 665824 214736 665876 214742
rect 665824 214678 665876 214684
rect 665088 212764 665140 212770
rect 665088 212706 665140 212712
rect 654796 210174 655132 210202
rect 656236 210174 656572 210202
rect 656788 210174 656848 210202
rect 657892 210174 658228 210202
rect 658444 210174 658780 210202
rect 659548 210174 659608 210202
rect 660100 210174 660436 210202
rect 660652 210174 660988 210202
rect 661204 210174 661540 210202
rect 661756 210174 662184 210202
rect 662308 210174 662368 210202
rect 662860 210174 663196 210202
rect 663412 210174 663472 210202
rect 663964 210174 664300 210202
rect 664516 210174 664944 210202
rect 632152 209568 632204 209574
rect 652024 209568 652076 209574
rect 632204 209516 632500 209522
rect 632152 209510 632500 209516
rect 652024 209510 652076 209516
rect 632164 209494 632500 209510
rect 666664 195974 666692 219399
rect 666834 215384 666890 215393
rect 666834 215319 666890 215328
rect 666848 198529 666876 215319
rect 667020 209092 667072 209098
rect 667020 209034 667072 209040
rect 666834 198520 666890 198529
rect 666834 198455 666890 198464
rect 666664 195946 666784 195974
rect 666756 175001 666784 195946
rect 666742 174992 666798 175001
rect 666742 174927 666798 174936
rect 667032 132705 667060 209034
rect 667216 134609 667244 282882
rect 667388 280220 667440 280226
rect 667388 280162 667440 280168
rect 667202 134600 667258 134609
rect 667202 134535 667258 134544
rect 667400 133521 667428 280162
rect 667584 180305 667612 285670
rect 667768 181393 667796 287030
rect 669136 264512 669188 264518
rect 669136 264454 669188 264460
rect 668216 264376 668268 264382
rect 668216 264318 668268 264324
rect 668032 231260 668084 231266
rect 668032 231202 668084 231208
rect 668044 199209 668072 231202
rect 668030 199200 668086 199209
rect 668030 199135 668086 199144
rect 668228 184521 668256 264318
rect 668952 264240 669004 264246
rect 668952 264182 669004 264188
rect 668766 232928 668822 232937
rect 668766 232863 668822 232872
rect 668584 231532 668636 231538
rect 668584 231474 668636 231480
rect 668596 230858 668624 231474
rect 668584 230852 668636 230858
rect 668584 230794 668636 230800
rect 668400 226772 668452 226778
rect 668400 226714 668452 226720
rect 668412 219434 668440 226714
rect 668584 224664 668636 224670
rect 668584 224606 668636 224612
rect 668596 221513 668624 224606
rect 668582 221504 668638 221513
rect 668582 221439 668638 221448
rect 668412 219406 668624 219434
rect 668400 218340 668452 218346
rect 668400 218282 668452 218288
rect 668412 215665 668440 218282
rect 668398 215656 668454 215665
rect 668398 215591 668454 215600
rect 668398 198792 668454 198801
rect 668398 198727 668454 198736
rect 668214 184512 668270 184521
rect 668214 184447 668270 184456
rect 667754 181384 667810 181393
rect 667754 181319 667810 181328
rect 667570 180296 667626 180305
rect 667570 180231 667626 180240
rect 668216 178016 668268 178022
rect 668214 177984 668216 177993
rect 668268 177984 668270 177993
rect 668214 177919 668270 177928
rect 668032 175092 668084 175098
rect 668032 175034 668084 175040
rect 668044 174729 668072 175034
rect 668030 174720 668086 174729
rect 668030 174655 668086 174664
rect 667940 169720 667992 169726
rect 667938 169688 667940 169697
rect 667992 169688 667994 169697
rect 667938 169623 667994 169632
rect 667940 165096 667992 165102
rect 667940 165038 667992 165044
rect 667952 164937 667980 165038
rect 667938 164928 667994 164937
rect 667938 164863 667994 164872
rect 668216 160064 668268 160070
rect 668214 160032 668216 160041
rect 668268 160032 668270 160041
rect 668214 159967 668270 159976
rect 668216 155576 668268 155582
rect 668216 155518 668268 155524
rect 668228 155145 668256 155518
rect 668214 155136 668270 155145
rect 668214 155071 668270 155080
rect 668412 143721 668440 198727
rect 668398 143712 668454 143721
rect 668398 143647 668454 143656
rect 668596 138825 668624 219406
rect 668780 163305 668808 232863
rect 668964 189417 668992 264182
rect 669148 258074 669176 264454
rect 669056 258046 669176 258074
rect 669056 209774 669084 258046
rect 669228 227180 669280 227186
rect 669228 227122 669280 227128
rect 669240 224058 669268 227122
rect 669228 224052 669280 224058
rect 669228 223994 669280 224000
rect 669228 223780 669280 223786
rect 669228 223722 669280 223728
rect 669240 220425 669268 223722
rect 669226 220416 669282 220425
rect 669226 220351 669282 220360
rect 669424 220266 669452 347239
rect 669870 302016 669926 302025
rect 669870 301951 669926 301960
rect 669688 234864 669740 234870
rect 669688 234806 669740 234812
rect 669700 234614 669728 234806
rect 669700 234586 669820 234614
rect 669792 231854 669820 234586
rect 669700 231826 669820 231854
rect 669700 223961 669728 231826
rect 669884 227186 669912 301951
rect 670330 262168 670386 262177
rect 670330 262103 670386 262112
rect 670146 258496 670202 258505
rect 670146 258431 670202 258440
rect 670160 234614 670188 258431
rect 670344 237289 670372 262103
rect 670330 237280 670386 237289
rect 670330 237215 670386 237224
rect 669976 234586 670188 234614
rect 669976 233186 670004 234586
rect 670332 234184 670384 234190
rect 670332 234126 670384 234132
rect 669976 233158 670280 233186
rect 670056 232892 670108 232898
rect 670056 232834 670108 232840
rect 669872 227180 669924 227186
rect 669872 227122 669924 227128
rect 669872 226636 669924 226642
rect 669872 226578 669924 226584
rect 669686 223952 669742 223961
rect 669686 223887 669742 223896
rect 669884 223802 669912 226578
rect 669700 223774 669912 223802
rect 670068 223786 670096 232834
rect 670056 223780 670108 223786
rect 669700 223582 669728 223774
rect 670056 223722 670108 223728
rect 669872 223644 669924 223650
rect 669872 223586 669924 223592
rect 669688 223576 669740 223582
rect 669688 223518 669740 223524
rect 669596 223440 669648 223446
rect 669332 220238 669452 220266
rect 669516 223388 669596 223394
rect 669516 223382 669648 223388
rect 669516 223366 669636 223382
rect 669332 220153 669360 220238
rect 669318 220144 669374 220153
rect 669318 220079 669374 220088
rect 669516 218346 669544 223366
rect 669884 223174 669912 223586
rect 669872 223168 669924 223174
rect 669872 223110 669924 223116
rect 669688 223100 669740 223106
rect 669688 223042 669740 223048
rect 669700 222442 669728 223042
rect 669872 222964 669924 222970
rect 669872 222906 669924 222912
rect 669884 222714 669912 222906
rect 670056 222896 670108 222902
rect 670056 222838 670108 222844
rect 669884 222686 670004 222714
rect 669608 222414 669728 222442
rect 669608 222194 669636 222414
rect 669778 222320 669834 222329
rect 669778 222255 669834 222264
rect 669608 222166 669728 222194
rect 669504 218340 669556 218346
rect 669504 218282 669556 218288
rect 669318 218240 669374 218249
rect 669700 218226 669728 222166
rect 669374 218198 669728 218226
rect 669318 218175 669374 218184
rect 669792 217682 669820 222255
rect 669424 217654 669820 217682
rect 669226 217016 669282 217025
rect 669226 216951 669282 216960
rect 669056 209746 669176 209774
rect 669148 200002 669176 209746
rect 669240 200138 669268 216951
rect 669424 215778 669452 217654
rect 669976 217546 670004 222686
rect 670068 222442 670096 222838
rect 670068 222414 670188 222442
rect 670160 222194 670188 222414
rect 669884 217530 670004 217546
rect 669872 217524 670004 217530
rect 669924 217518 670004 217524
rect 670068 222166 670188 222194
rect 669872 217466 669924 217472
rect 669872 217116 669924 217122
rect 669872 217058 669924 217064
rect 669332 215750 669452 215778
rect 669332 215506 669360 215750
rect 669332 215478 669820 215506
rect 669594 213888 669650 213897
rect 669594 213823 669650 213832
rect 669608 202881 669636 213823
rect 669594 202872 669650 202881
rect 669594 202807 669650 202816
rect 669240 200110 669544 200138
rect 669148 199974 669360 200002
rect 669332 194313 669360 199974
rect 669318 194304 669374 194313
rect 669318 194239 669374 194248
rect 669516 191834 669544 200110
rect 669792 195974 669820 215478
rect 669148 191806 669544 191834
rect 669700 195946 669820 195974
rect 669148 191593 669176 191806
rect 669134 191584 669190 191593
rect 669134 191519 669190 191528
rect 668950 189408 669006 189417
rect 668950 189343 669006 189352
rect 669134 188456 669190 188465
rect 669134 188391 669190 188400
rect 668952 184884 669004 184890
rect 668952 184826 669004 184832
rect 668766 163296 668822 163305
rect 668766 163231 668822 163240
rect 668766 156224 668822 156233
rect 668766 156159 668822 156168
rect 668780 148617 668808 156159
rect 668766 148608 668822 148617
rect 668766 148543 668822 148552
rect 668768 145784 668820 145790
rect 668768 145726 668820 145732
rect 668780 145353 668808 145726
rect 668766 145344 668822 145353
rect 668766 145279 668822 145288
rect 668582 138816 668638 138825
rect 668582 138751 668638 138760
rect 668766 135144 668822 135153
rect 668766 135079 668822 135088
rect 667940 133816 667992 133822
rect 667938 133784 667940 133793
rect 667992 133784 667994 133793
rect 667938 133719 667994 133728
rect 667386 133512 667442 133521
rect 667386 133447 667442 133456
rect 667018 132696 667074 132705
rect 667018 132631 667074 132640
rect 668584 130824 668636 130830
rect 668584 130766 668636 130772
rect 668596 130665 668624 130766
rect 668582 130656 668638 130665
rect 668582 130591 668638 130600
rect 668032 129736 668084 129742
rect 668032 129678 668084 129684
rect 668044 129033 668072 129678
rect 668030 129024 668086 129033
rect 668030 128959 668086 128968
rect 668582 127800 668638 127809
rect 668582 127735 668638 127744
rect 667940 108860 667992 108866
rect 667940 108802 667992 108808
rect 667952 107817 667980 108802
rect 667938 107808 667994 107817
rect 667938 107743 667994 107752
rect 668400 106208 668452 106214
rect 668398 106176 668400 106185
rect 668452 106176 668454 106185
rect 668398 106111 668454 106120
rect 668596 102921 668624 127735
rect 668780 119241 668808 135079
rect 668964 125769 668992 184826
rect 669148 135561 669176 188391
rect 669502 172408 669558 172417
rect 669502 172343 669558 172352
rect 669516 166994 669544 172343
rect 669700 169726 669728 195946
rect 669688 169720 669740 169726
rect 669688 169662 669740 169668
rect 669516 166966 669636 166994
rect 669318 162888 669374 162897
rect 669318 162823 669374 162832
rect 669332 158409 669360 162823
rect 669318 158400 669374 158409
rect 669318 158335 669374 158344
rect 669608 150385 669636 166966
rect 669594 150376 669650 150385
rect 669594 150311 669650 150320
rect 669134 135552 669190 135561
rect 669134 135487 669190 135496
rect 669884 133822 669912 217058
rect 670068 165102 670096 222166
rect 670252 218770 670280 233158
rect 670344 223530 670372 234126
rect 670528 226642 670556 392527
rect 670974 295896 671030 295905
rect 670974 295831 671030 295840
rect 670988 293865 671016 295831
rect 670974 293856 671030 293865
rect 670974 293791 671030 293800
rect 671356 278730 671384 570386
rect 671988 570172 672040 570178
rect 671988 570114 672040 570120
rect 671802 559600 671858 559609
rect 671802 559535 671858 559544
rect 671618 532808 671674 532817
rect 671618 532743 671674 532752
rect 671632 489326 671660 532743
rect 671620 489320 671672 489326
rect 671620 489262 671672 489268
rect 671816 483206 671844 559535
rect 671804 483200 671856 483206
rect 671804 483142 671856 483148
rect 672000 454866 672028 570114
rect 672262 555248 672318 555257
rect 672262 555183 672318 555192
rect 672276 486062 672304 555183
rect 672460 533746 672488 572686
rect 672632 535968 672684 535974
rect 672630 535936 672632 535945
rect 672684 535936 672686 535945
rect 672630 535871 672686 535880
rect 672632 535696 672684 535702
rect 672630 535664 672632 535673
rect 672684 535664 672686 535673
rect 672630 535599 672686 535608
rect 672632 534880 672684 534886
rect 672630 534848 672632 534857
rect 672684 534848 672686 534857
rect 672630 534783 672686 534792
rect 672632 534608 672684 534614
rect 672630 534576 672632 534585
rect 672684 534576 672686 534585
rect 672630 534511 672686 534520
rect 672630 534304 672686 534313
rect 672630 534239 672632 534248
rect 672684 534239 672686 534248
rect 672632 534210 672684 534216
rect 672828 534018 672856 572686
rect 673090 560280 673146 560289
rect 673090 560215 673146 560224
rect 672828 533990 673040 534018
rect 672460 533718 672856 533746
rect 672630 533624 672686 533633
rect 672630 533559 672686 533568
rect 672448 533384 672500 533390
rect 672446 533352 672448 533361
rect 672500 533352 672502 533361
rect 672446 533287 672502 533296
rect 672448 532568 672500 532574
rect 672446 532536 672448 532545
rect 672500 532536 672502 532545
rect 672446 532471 672502 532480
rect 672448 490476 672500 490482
rect 672448 490418 672500 490424
rect 672264 486056 672316 486062
rect 672264 485998 672316 486004
rect 672000 454850 672120 454866
rect 672000 454844 672132 454850
rect 672000 454838 672080 454844
rect 672080 454786 672132 454792
rect 672264 453960 672316 453966
rect 672262 453928 672264 453937
rect 672316 453928 672318 453937
rect 672262 453863 672318 453872
rect 672460 402121 672488 490418
rect 672644 490142 672672 533559
rect 672828 533474 672856 533718
rect 672736 533446 672856 533474
rect 672736 530754 672764 533446
rect 672736 530726 672856 530754
rect 672828 528873 672856 530726
rect 672814 528864 672870 528873
rect 672814 528799 672870 528808
rect 673012 528714 673040 533990
rect 672920 528686 673040 528714
rect 672920 528057 672948 528686
rect 672906 528048 672962 528057
rect 672906 527983 672962 527992
rect 672632 490136 672684 490142
rect 672632 490078 672684 490084
rect 672632 489660 672684 489666
rect 672632 489602 672684 489608
rect 672446 402112 672502 402121
rect 672446 402047 672502 402056
rect 672644 401713 672672 489602
rect 673104 484809 673132 560215
rect 673288 530942 673316 603502
rect 673472 598934 673500 603758
rect 673380 598906 673500 598934
rect 673380 531026 673408 598906
rect 673564 596873 673592 607038
rect 673840 598934 673868 615466
rect 674288 614644 674340 614650
rect 674288 614586 674340 614592
rect 674300 614258 674328 614586
rect 674024 614230 674328 614258
rect 674024 614174 674052 614230
rect 674012 614168 674064 614174
rect 674012 614110 674064 614116
rect 674024 611386 674328 611402
rect 674012 611380 674340 611386
rect 674064 611374 674288 611380
rect 674012 611322 674064 611328
rect 674288 611322 674340 611328
rect 674484 611354 674512 619534
rect 675128 615494 675156 640478
rect 675300 640280 675352 640286
rect 675220 640228 675300 640234
rect 675220 640222 675352 640228
rect 675220 640206 675340 640222
rect 675220 630674 675248 640206
rect 675404 639826 675432 640152
rect 675312 639798 675432 639826
rect 675312 631394 675340 639798
rect 675496 638625 675524 638928
rect 675482 638616 675538 638625
rect 675482 638551 675538 638560
rect 681002 637528 681058 637537
rect 681002 637463 681058 637472
rect 675668 635520 675720 635526
rect 675668 635462 675720 635468
rect 675680 631417 675708 635462
rect 675482 631408 675538 631417
rect 675312 631366 675482 631394
rect 675482 631343 675538 631352
rect 675666 631408 675722 631417
rect 675666 631343 675722 631352
rect 675220 630646 675340 630674
rect 675312 617137 675340 630646
rect 681016 622033 681044 637463
rect 683212 637016 683264 637022
rect 683212 636958 683264 636964
rect 676218 622024 676274 622033
rect 676218 621959 676274 621968
rect 681002 622024 681058 622033
rect 681002 621959 681058 621968
rect 676232 621042 676260 621959
rect 676220 621036 676272 621042
rect 676220 620978 676272 620984
rect 676034 620664 676090 620673
rect 676034 620599 676090 620608
rect 676048 619750 676076 620599
rect 676036 619744 676088 619750
rect 676036 619686 676088 619692
rect 676218 619168 676274 619177
rect 676218 619103 676274 619112
rect 676232 618526 676260 619103
rect 683224 618769 683252 636958
rect 683396 636880 683448 636886
rect 683396 636822 683448 636828
rect 683408 634814 683436 636822
rect 683408 634786 683620 634814
rect 683396 623076 683448 623082
rect 683396 623018 683448 623024
rect 683210 618760 683266 618769
rect 683210 618695 683266 618704
rect 676220 618520 676272 618526
rect 676220 618462 676272 618468
rect 676496 618044 676548 618050
rect 676496 617986 676548 617992
rect 676218 617944 676274 617953
rect 676218 617879 676220 617888
rect 676272 617879 676274 617888
rect 676220 617850 676272 617856
rect 676508 617545 676536 617986
rect 676218 617536 676274 617545
rect 676218 617471 676220 617480
rect 676272 617471 676274 617480
rect 676494 617536 676550 617545
rect 676494 617471 676550 617480
rect 676220 617442 676272 617448
rect 675298 617128 675354 617137
rect 675298 617063 675354 617072
rect 683408 616729 683436 623018
rect 683592 617137 683620 634786
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683578 617128 683634 617137
rect 683578 617063 683634 617072
rect 683394 616720 683450 616729
rect 683394 616655 683450 616664
rect 683120 615528 683172 615534
rect 674852 615466 675156 615494
rect 683118 615496 683120 615505
rect 683172 615496 683174 615505
rect 674484 611326 674788 611354
rect 674012 608660 674064 608666
rect 674288 608660 674340 608666
rect 674064 608620 674288 608648
rect 674012 608602 674064 608608
rect 674288 608602 674340 608608
rect 674010 608016 674066 608025
rect 674010 607951 674066 607960
rect 674024 603566 674052 607951
rect 674012 603560 674064 603566
rect 674012 603502 674064 603508
rect 674288 603288 674340 603294
rect 674288 603230 674340 603236
rect 674010 600400 674066 600409
rect 674010 600335 674012 600344
rect 674064 600335 674066 600344
rect 674012 600306 674064 600312
rect 674010 599720 674066 599729
rect 674010 599655 674066 599664
rect 674024 599502 674052 599655
rect 674024 599474 674236 599502
rect 674012 599412 674064 599418
rect 674012 599354 674064 599360
rect 673748 598906 673868 598934
rect 673550 596864 673606 596873
rect 673550 596799 673606 596808
rect 673748 582374 673776 598906
rect 674024 598097 674052 599354
rect 674010 598088 674066 598097
rect 674010 598023 674066 598032
rect 673918 597136 673974 597145
rect 673918 597071 673974 597080
rect 673932 592034 673960 597071
rect 674208 592034 674236 599474
rect 673656 582346 673776 582374
rect 673840 592006 673960 592034
rect 674024 592006 674236 592034
rect 673656 581369 673684 582346
rect 673642 581360 673698 581369
rect 673642 581295 673698 581304
rect 673642 581088 673698 581097
rect 673642 581023 673644 581032
rect 673696 581023 673698 581032
rect 673644 580994 673696 581000
rect 673644 580304 673696 580310
rect 673642 580272 673644 580281
rect 673696 580272 673698 580281
rect 673642 580207 673698 580216
rect 673644 579896 673696 579902
rect 673642 579864 673644 579873
rect 673696 579864 673698 579873
rect 673642 579799 673698 579808
rect 673642 579456 673698 579465
rect 673642 579391 673644 579400
rect 673696 579391 673698 579400
rect 673644 579362 673696 579368
rect 673644 579080 673696 579086
rect 673642 579048 673644 579057
rect 673696 579048 673698 579057
rect 673642 578983 673698 578992
rect 673642 578640 673698 578649
rect 673642 578575 673644 578584
rect 673696 578575 673698 578584
rect 673644 578546 673696 578552
rect 673642 578232 673698 578241
rect 673642 578167 673644 578176
rect 673696 578167 673698 578176
rect 673644 578138 673696 578144
rect 673642 577824 673698 577833
rect 673642 577759 673644 577768
rect 673696 577759 673698 577768
rect 673644 577730 673696 577736
rect 673644 577448 673696 577454
rect 673642 577416 673644 577425
rect 673696 577416 673698 577425
rect 673642 577351 673698 577360
rect 673642 577008 673698 577017
rect 673642 576943 673644 576952
rect 673696 576943 673698 576952
rect 673644 576914 673696 576920
rect 673644 574592 673696 574598
rect 673642 574560 673644 574569
rect 673696 574560 673698 574569
rect 673642 574495 673698 574504
rect 673644 574184 673696 574190
rect 673642 574152 673644 574161
rect 673696 574152 673698 574161
rect 673642 574087 673698 574096
rect 673642 572520 673698 572529
rect 673642 572455 673698 572464
rect 673656 572286 673684 572455
rect 673644 572280 673696 572286
rect 673644 572222 673696 572228
rect 673642 572112 673698 572121
rect 673642 572047 673698 572056
rect 673656 571470 673684 572047
rect 673644 571464 673696 571470
rect 673644 571406 673696 571412
rect 673642 570888 673698 570897
rect 673642 570823 673698 570832
rect 673656 570178 673684 570823
rect 673644 570172 673696 570178
rect 673644 570114 673696 570120
rect 673644 569968 673696 569974
rect 673642 569936 673644 569945
rect 673696 569936 673698 569945
rect 673642 569871 673698 569880
rect 673642 569664 673698 569673
rect 673642 569599 673698 569608
rect 673656 568614 673684 569599
rect 673644 568608 673696 568614
rect 673644 568550 673696 568556
rect 673644 565888 673696 565894
rect 673642 565856 673644 565865
rect 673696 565856 673698 565865
rect 673642 565791 673698 565800
rect 673642 564632 673698 564641
rect 673642 564567 673644 564576
rect 673696 564567 673698 564576
rect 673644 564538 673696 564544
rect 673642 554840 673698 554849
rect 673642 554775 673644 554784
rect 673696 554775 673698 554784
rect 673644 554746 673696 554752
rect 673642 553480 673698 553489
rect 673642 553415 673644 553424
rect 673696 553415 673698 553424
rect 673644 553386 673696 553392
rect 673642 553208 673698 553217
rect 673642 553143 673698 553152
rect 673380 530998 673500 531026
rect 673276 530936 673328 530942
rect 673276 530878 673328 530884
rect 673472 530822 673500 530998
rect 673380 530794 673500 530822
rect 673090 484800 673146 484809
rect 673090 484735 673146 484744
rect 673380 455870 673408 530794
rect 673656 482361 673684 553143
rect 673840 540974 673868 592006
rect 674024 586514 674052 592006
rect 673932 586486 674052 586514
rect 673932 550634 673960 586486
rect 674102 558376 674158 558385
rect 674102 558311 674158 558320
rect 674116 553394 674144 558311
rect 674300 557534 674328 603230
rect 674564 599004 674616 599010
rect 674564 598946 674616 598952
rect 674576 598482 674604 598946
rect 674576 598454 674696 598482
rect 674472 598392 674524 598398
rect 674472 598334 674524 598340
rect 674484 597145 674512 598334
rect 674470 597136 674526 597145
rect 674470 597071 674526 597080
rect 674470 596864 674526 596873
rect 674470 596799 674526 596808
rect 674484 588606 674512 596799
rect 674668 592770 674696 598454
rect 674576 592742 674696 592770
rect 674576 592034 674604 592742
rect 674760 592618 674788 611326
rect 674852 592770 674880 615466
rect 683118 615431 683174 615440
rect 676218 614680 676274 614689
rect 676218 614615 676220 614624
rect 676272 614615 676274 614624
rect 676220 614586 676272 614592
rect 675392 611380 675444 611386
rect 675392 611322 675444 611328
rect 675404 608668 675432 611322
rect 675116 608660 675168 608666
rect 675116 608602 675168 608608
rect 675128 606846 675156 608602
rect 675404 608025 675432 608124
rect 675390 608016 675446 608025
rect 675390 607951 675446 607960
rect 675482 607744 675538 607753
rect 675482 607679 675538 607688
rect 675496 607479 675524 607679
rect 675128 606818 675418 606846
rect 674944 604982 675418 605010
rect 674944 597554 674972 604982
rect 675114 604480 675170 604489
rect 675170 604438 675418 604466
rect 675114 604415 675170 604424
rect 675312 603894 675432 603922
rect 675312 603786 675340 603894
rect 675128 603758 675340 603786
rect 675404 603772 675432 603894
rect 675128 603294 675156 603758
rect 675116 603288 675168 603294
rect 675116 603230 675168 603236
rect 675128 603146 675418 603174
rect 675128 602993 675156 603146
rect 675114 602984 675170 602993
rect 675114 602919 675170 602928
rect 675390 600944 675446 600953
rect 675390 600879 675446 600888
rect 675404 600644 675432 600879
rect 675114 600400 675170 600409
rect 675114 600335 675170 600344
rect 675128 598278 675156 600335
rect 675312 600222 675432 600250
rect 675312 599010 675340 600222
rect 675404 600100 675432 600222
rect 675482 599720 675538 599729
rect 675482 599655 675538 599664
rect 675496 599488 675524 599655
rect 675300 599004 675352 599010
rect 675300 598946 675352 598952
rect 675312 598862 675432 598890
rect 675312 598398 675340 598862
rect 675404 598808 675432 598862
rect 675300 598392 675352 598398
rect 675300 598334 675352 598340
rect 675128 598250 675418 598278
rect 675114 598088 675170 598097
rect 675114 598023 675170 598032
rect 674944 597526 675064 597554
rect 674852 592742 674972 592770
rect 674748 592612 674800 592618
rect 674748 592554 674800 592560
rect 674944 592034 674972 592742
rect 674576 592006 674696 592034
rect 674472 588600 674524 588606
rect 674472 588542 674524 588548
rect 674470 581360 674526 581369
rect 674470 581295 674526 581304
rect 674484 571606 674512 581295
rect 674472 571600 674524 571606
rect 674472 571542 674524 571548
rect 674668 560294 674696 592006
rect 674852 592006 674972 592034
rect 674852 590646 674880 592006
rect 674840 590640 674892 590646
rect 674840 590582 674892 590588
rect 675036 590322 675064 597526
rect 675128 596442 675156 598023
rect 675404 597417 675432 597652
rect 675390 597408 675446 597417
rect 675390 597343 675446 597352
rect 675128 596414 675418 596442
rect 675404 595354 675432 595816
rect 675312 595326 675432 595354
rect 675312 590442 675340 595326
rect 675496 594833 675524 595136
rect 675482 594824 675538 594833
rect 675482 594759 675538 594768
rect 675496 593609 675524 593980
rect 675482 593600 675538 593609
rect 675482 593535 675538 593544
rect 675482 593192 675538 593201
rect 675482 593127 675538 593136
rect 675300 590436 675352 590442
rect 675300 590378 675352 590384
rect 675036 590294 675340 590322
rect 675116 590232 675168 590238
rect 675116 590174 675168 590180
rect 675128 586514 675156 590174
rect 675312 587894 675340 590294
rect 675036 586486 675156 586514
rect 675220 587866 675340 587894
rect 674840 570512 674892 570518
rect 674840 570454 674892 570460
rect 674852 569945 674880 570454
rect 674838 569936 674894 569945
rect 674838 569871 674894 569880
rect 675036 567194 675064 586486
rect 675220 586265 675248 587866
rect 675206 586256 675262 586265
rect 675206 586191 675262 586200
rect 675496 570518 675524 593127
rect 683396 592680 683448 592686
rect 683396 592622 683448 592628
rect 681002 591696 681058 591705
rect 681002 591631 681058 591640
rect 681016 575657 681044 591631
rect 682384 590640 682436 590646
rect 682384 590582 682436 590588
rect 682396 576473 682424 590582
rect 682382 576464 682438 576473
rect 682382 576399 682438 576408
rect 681002 575648 681058 575657
rect 681002 575583 681058 575592
rect 683408 573209 683436 592622
rect 684222 591288 684278 591297
rect 684222 591223 684278 591232
rect 684040 588600 684092 588606
rect 684040 588542 684092 588548
rect 683394 573200 683450 573209
rect 683394 573135 683450 573144
rect 684052 571985 684080 588542
rect 684236 576065 684264 591223
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 684222 576056 684278 576065
rect 684222 575991 684278 576000
rect 684038 571976 684094 571985
rect 684038 571911 684094 571920
rect 676220 571600 676272 571606
rect 676218 571568 676220 571577
rect 676272 571568 676274 571577
rect 676218 571503 676274 571512
rect 675484 570512 675536 570518
rect 675484 570454 675536 570460
rect 683120 570512 683172 570518
rect 683120 570454 683172 570460
rect 683132 570353 683160 570454
rect 683118 570344 683174 570353
rect 683118 570279 683174 570288
rect 674944 567166 675064 567194
rect 674668 560266 674788 560294
rect 674300 557506 674420 557534
rect 674116 553366 674236 553394
rect 674208 550634 674236 553366
rect 674392 550634 674420 557506
rect 674760 552106 674788 560266
rect 674944 553330 674972 567166
rect 675390 565856 675446 565865
rect 675390 565791 675446 565800
rect 675114 564632 675170 564641
rect 675114 564567 675170 564576
rect 675128 562918 675156 564567
rect 675404 563448 675432 565791
rect 675312 562958 675432 562986
rect 675312 562918 675340 562958
rect 675128 562890 675340 562918
rect 675404 562904 675432 562958
rect 675114 562320 675170 562329
rect 675170 562278 675418 562306
rect 675114 562255 675170 562264
rect 675390 561912 675446 561921
rect 675390 561847 675446 561856
rect 675404 561612 675432 561847
rect 675312 559830 675432 559858
rect 675312 559790 675340 559830
rect 675036 559762 675340 559790
rect 675404 559776 675432 559830
rect 675036 554690 675064 559762
rect 675206 559600 675262 559609
rect 675206 559535 675262 559544
rect 675220 557954 675248 559535
rect 675574 559464 675630 559473
rect 675574 559399 675630 559408
rect 675588 559232 675616 559399
rect 675496 558385 675524 558620
rect 675482 558376 675538 558385
rect 675482 558311 675538 558320
rect 675220 557926 675418 557954
rect 675298 557560 675354 557569
rect 675298 557495 675354 557504
rect 675312 556186 675340 557495
rect 675220 556158 675340 556186
rect 675220 554933 675248 556158
rect 675404 555257 675432 555492
rect 675390 555248 675446 555257
rect 675390 555183 675446 555192
rect 675220 554905 675418 554933
rect 675298 554840 675354 554849
rect 675298 554775 675354 554784
rect 675036 554662 675248 554690
rect 674944 553302 675064 553330
rect 674760 552078 674972 552106
rect 674654 551984 674710 551993
rect 674654 551919 674710 551928
rect 674668 551562 674696 551919
rect 673932 550606 674052 550634
rect 674024 548865 674052 550606
rect 674116 550606 674236 550634
rect 674300 550606 674420 550634
rect 674484 551534 674696 551562
rect 674116 548978 674144 550606
rect 674116 548950 674236 548978
rect 674010 548856 674066 548865
rect 674010 548791 674066 548800
rect 673840 540946 674052 540974
rect 673826 536208 673882 536217
rect 673826 536143 673882 536152
rect 673840 532234 673868 536143
rect 673828 532228 673880 532234
rect 673828 532170 673880 532176
rect 674024 531978 674052 540946
rect 674208 536217 674236 548950
rect 674300 540974 674328 550606
rect 674300 540946 674420 540974
rect 674194 536208 674250 536217
rect 674194 536143 674250 536152
rect 674392 535786 674420 540946
rect 674116 535758 674420 535786
rect 674116 533746 674144 535758
rect 674288 534132 674340 534138
rect 674288 534074 674340 534080
rect 674300 533905 674328 534074
rect 674286 533896 674342 533905
rect 674286 533831 674342 533840
rect 674116 533718 674328 533746
rect 674300 533390 674328 533718
rect 674288 533384 674340 533390
rect 674288 533326 674340 533332
rect 674024 531950 674144 531978
rect 673828 531820 673880 531826
rect 673828 531762 673880 531768
rect 673840 531434 673868 531762
rect 673748 531406 673868 531434
rect 673748 518894 673776 531406
rect 674116 531314 674144 531950
rect 673840 531286 674144 531314
rect 673840 528442 673868 531286
rect 674012 530936 674064 530942
rect 674064 530884 674328 530890
rect 674012 530878 674328 530884
rect 674024 530874 674328 530878
rect 674024 530868 674340 530874
rect 674024 530862 674288 530868
rect 674288 530810 674340 530816
rect 674012 529984 674064 529990
rect 674288 529984 674340 529990
rect 674064 529932 674288 529938
rect 674012 529926 674340 529932
rect 674024 529910 674328 529926
rect 674012 529304 674064 529310
rect 674064 529252 674328 529258
rect 674012 529246 674328 529252
rect 674024 529242 674328 529246
rect 674024 529236 674340 529242
rect 674024 529230 674288 529236
rect 674288 529178 674340 529184
rect 674288 529032 674340 529038
rect 674024 528980 674288 528986
rect 674024 528974 674340 528980
rect 674024 528958 674328 528974
rect 674024 528630 674052 528958
rect 674012 528624 674064 528630
rect 674012 528566 674064 528572
rect 673840 528414 674328 528442
rect 674300 526386 674328 528414
rect 674288 526380 674340 526386
rect 674288 526322 674340 526328
rect 674024 524482 674328 524498
rect 674012 524476 674340 524482
rect 674064 524470 674288 524476
rect 674012 524418 674064 524424
rect 674288 524418 674340 524424
rect 673748 518866 674144 518894
rect 674116 499574 674144 518866
rect 674116 499546 674328 499574
rect 673826 492144 673882 492153
rect 673826 492079 673882 492088
rect 673840 491366 673868 492079
rect 674300 492046 674328 499546
rect 674288 492040 674340 492046
rect 674288 491982 674340 491988
rect 674012 491904 674064 491910
rect 674064 491852 674328 491858
rect 674012 491846 674328 491852
rect 674024 491842 674328 491846
rect 674024 491836 674340 491842
rect 674024 491830 674288 491836
rect 674288 491778 674340 491784
rect 674288 491700 674340 491706
rect 674288 491642 674340 491648
rect 674300 491586 674328 491642
rect 674024 491558 674328 491586
rect 674024 491502 674052 491558
rect 674012 491496 674064 491502
rect 674012 491438 674064 491444
rect 673828 491360 673880 491366
rect 673828 491302 673880 491308
rect 674012 490952 674064 490958
rect 674010 490920 674012 490929
rect 674064 490920 674066 490929
rect 674010 490855 674066 490864
rect 674010 490512 674066 490521
rect 674010 490447 674012 490456
rect 674064 490447 674066 490456
rect 674012 490418 674064 490424
rect 674012 490136 674064 490142
rect 674010 490104 674012 490113
rect 674064 490104 674066 490113
rect 674010 490039 674066 490048
rect 674010 489696 674066 489705
rect 674010 489631 674012 489640
rect 674064 489631 674066 489640
rect 674012 489602 674064 489608
rect 674012 489320 674064 489326
rect 674010 489288 674012 489297
rect 674064 489288 674066 489297
rect 674010 489223 674066 489232
rect 674012 488504 674064 488510
rect 674010 488472 674012 488481
rect 674064 488472 674066 488481
rect 674010 488407 674066 488416
rect 674288 486192 674340 486198
rect 674024 486140 674288 486146
rect 674024 486134 674340 486140
rect 674024 486118 674328 486134
rect 673828 486056 673880 486062
rect 673826 486024 673828 486033
rect 673880 486024 673882 486033
rect 673826 485959 673882 485968
rect 674024 485858 674052 486118
rect 674012 485852 674064 485858
rect 674012 485794 674064 485800
rect 674288 485172 674340 485178
rect 674288 485114 674340 485120
rect 674300 485058 674328 485114
rect 674024 485030 674328 485058
rect 674024 484430 674052 485030
rect 674012 484424 674064 484430
rect 674012 484366 674064 484372
rect 674484 484022 674512 551534
rect 674944 550746 674972 552078
rect 674852 550718 674972 550746
rect 674852 550662 674880 550718
rect 674656 550656 674708 550662
rect 674656 550598 674708 550604
rect 674840 550656 674892 550662
rect 674840 550598 674892 550604
rect 674668 526794 674696 550598
rect 675036 550066 675064 553302
rect 675220 552634 675248 554662
rect 675312 553466 675340 554775
rect 675772 553897 675800 554268
rect 675758 553888 675814 553897
rect 675758 553823 675814 553832
rect 675588 553489 675616 553656
rect 675574 553480 675630 553489
rect 675312 553438 675432 553466
rect 675404 553079 675432 553438
rect 675574 553415 675630 553424
rect 675208 552628 675260 552634
rect 675208 552570 675260 552576
rect 675208 552356 675260 552362
rect 675208 552298 675260 552304
rect 675220 550526 675248 552298
rect 675404 551993 675432 552432
rect 675390 551984 675446 551993
rect 675390 551919 675446 551928
rect 675390 551576 675446 551585
rect 675390 551511 675446 551520
rect 675404 551239 675432 551511
rect 675208 550520 675260 550526
rect 675208 550462 675260 550468
rect 675496 550225 675524 550596
rect 675482 550216 675538 550225
rect 675482 550151 675538 550160
rect 674852 550038 675064 550066
rect 674852 546038 674880 550038
rect 675022 549944 675078 549953
rect 675022 549879 675078 549888
rect 674840 546032 674892 546038
rect 674840 545974 674892 545980
rect 674838 545864 674894 545873
rect 674838 545799 674894 545808
rect 674656 526788 674708 526794
rect 674656 526730 674708 526736
rect 674852 500954 674880 545799
rect 675036 540974 675064 549879
rect 675300 549840 675352 549846
rect 675300 549782 675352 549788
rect 675036 540946 675156 540974
rect 675128 503674 675156 540946
rect 675116 503668 675168 503674
rect 675116 503610 675168 503616
rect 675312 503538 675340 549782
rect 675496 549681 675524 549951
rect 675482 549672 675538 549681
rect 675482 549607 675538 549616
rect 675772 548321 675800 548760
rect 675758 548312 675814 548321
rect 675758 548247 675814 548256
rect 675574 547904 675630 547913
rect 675574 547839 675630 547848
rect 675588 547194 675616 547839
rect 677414 547632 677470 547641
rect 677414 547567 677470 547576
rect 675576 547188 675628 547194
rect 675576 547130 675628 547136
rect 675482 536480 675538 536489
rect 675482 536415 675538 536424
rect 675496 532030 675524 536415
rect 676034 534508 676090 534517
rect 676034 534443 676090 534452
rect 676048 534138 676076 534443
rect 676036 534132 676088 534138
rect 676036 534074 676088 534080
rect 675484 532024 675536 532030
rect 675484 531966 675536 531972
rect 676220 532024 676272 532030
rect 676220 531966 676272 531972
rect 676232 531865 676260 531966
rect 676218 531856 676274 531865
rect 676218 531791 676274 531800
rect 676036 530868 676088 530874
rect 676034 530836 676036 530845
rect 676088 530836 676090 530845
rect 676034 530771 676090 530780
rect 676034 530020 676090 530029
rect 676034 529955 676036 529964
rect 676088 529955 676090 529964
rect 676036 529926 676088 529932
rect 676218 529408 676274 529417
rect 676218 529343 676274 529352
rect 676036 529236 676088 529242
rect 676034 529204 676036 529213
rect 676088 529204 676090 529213
rect 676034 529139 676090 529148
rect 676232 529038 676260 529343
rect 676220 529032 676272 529038
rect 676220 528974 676272 528980
rect 676036 526788 676088 526794
rect 676034 526756 676036 526765
rect 676088 526756 676090 526765
rect 676034 526691 676090 526700
rect 676036 526380 676088 526386
rect 676034 526348 676036 526357
rect 676088 526348 676090 526357
rect 676034 526283 676090 526292
rect 675484 520260 675536 520266
rect 675484 520202 675536 520208
rect 675300 503532 675352 503538
rect 675300 503474 675352 503480
rect 674840 500948 674892 500954
rect 674840 500890 674892 500896
rect 674656 492040 674708 492046
rect 674656 491982 674708 491988
rect 674668 484401 674696 491982
rect 674654 484392 674710 484401
rect 674654 484327 674710 484336
rect 674472 484016 674524 484022
rect 674472 483958 674524 483964
rect 674012 483200 674064 483206
rect 674010 483168 674012 483177
rect 674064 483168 674066 483177
rect 674010 483103 674066 483112
rect 673642 482352 673698 482361
rect 673642 482287 673698 482296
rect 674012 480752 674064 480758
rect 674012 480694 674064 480700
rect 674024 480570 674052 480694
rect 674024 480542 674328 480570
rect 674300 480418 674328 480542
rect 674288 480412 674340 480418
rect 674288 480354 674340 480360
rect 673368 455864 673420 455870
rect 673368 455806 673420 455812
rect 673274 455424 673330 455433
rect 673274 455359 673276 455368
rect 673328 455359 673330 455368
rect 673276 455330 673328 455336
rect 673386 455288 673442 455297
rect 673386 455223 673388 455232
rect 673440 455223 673442 455232
rect 673506 455252 673558 455258
rect 673388 455194 673440 455200
rect 673506 455194 673558 455200
rect 673274 455152 673330 455161
rect 673518 455138 673546 455194
rect 673330 455110 673546 455138
rect 673274 455087 673330 455096
rect 674288 454912 674340 454918
rect 672814 454880 672870 454889
rect 672814 454815 672870 454824
rect 674286 454880 674288 454889
rect 674340 454880 674342 454889
rect 674286 454815 674342 454824
rect 672828 454510 672856 454815
rect 675496 454646 675524 520202
rect 675668 518832 675720 518838
rect 675668 518774 675720 518780
rect 673046 454640 673098 454646
rect 673044 454608 673046 454617
rect 674288 454640 674340 454646
rect 673098 454608 673100 454617
rect 673044 454543 673100 454552
rect 674286 454608 674288 454617
rect 675484 454640 675536 454646
rect 674340 454608 674342 454617
rect 675484 454582 675536 454588
rect 674286 454543 674342 454552
rect 672816 454504 672868 454510
rect 672816 454446 672868 454452
rect 675680 454374 675708 518774
rect 675852 491836 675904 491842
rect 675852 491778 675904 491784
rect 675864 491337 675892 491778
rect 676034 491736 676090 491745
rect 676034 491671 676036 491680
rect 676088 491671 676090 491680
rect 676036 491642 676088 491648
rect 675850 491328 675906 491337
rect 675850 491263 675906 491272
rect 676034 486840 676090 486849
rect 676034 486775 676090 486784
rect 676048 486198 676076 486775
rect 676036 486192 676088 486198
rect 676036 486134 676088 486140
rect 676034 485208 676090 485217
rect 676034 485143 676036 485152
rect 676088 485143 676090 485152
rect 676036 485114 676088 485120
rect 676036 484016 676088 484022
rect 676034 483984 676036 483993
rect 676088 483984 676090 483993
rect 676034 483919 676090 483928
rect 677428 483002 677456 547567
rect 683212 547188 683264 547194
rect 683212 547130 683264 547136
rect 681002 546816 681058 546825
rect 681002 546751 681058 546760
rect 681016 530641 681044 546751
rect 682384 545896 682436 545902
rect 682384 545838 682436 545844
rect 682396 531457 682424 545838
rect 682382 531448 682438 531457
rect 682382 531383 682438 531392
rect 681002 530632 681058 530641
rect 681002 530567 681058 530576
rect 683224 527785 683252 547130
rect 683394 547088 683450 547097
rect 683394 547023 683450 547032
rect 683210 527776 683266 527785
rect 683210 527711 683266 527720
rect 683408 527377 683436 547023
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683580 533384 683632 533390
rect 683580 533326 683632 533332
rect 683592 528601 683620 533326
rect 683578 528592 683634 528601
rect 683578 528527 683634 528536
rect 683394 527368 683450 527377
rect 683394 527303 683450 527312
rect 677874 525736 677930 525745
rect 677874 525671 677930 525680
rect 677888 518838 677916 525671
rect 683118 524920 683174 524929
rect 683118 524855 683174 524864
rect 678978 524512 679034 524521
rect 683132 524482 683160 524855
rect 678978 524447 679034 524456
rect 683120 524476 683172 524482
rect 678992 520266 679020 524447
rect 683120 524418 683172 524424
rect 678980 520260 679032 520266
rect 678980 520202 679032 520208
rect 677876 518832 677928 518838
rect 677876 518774 677928 518780
rect 683394 503704 683450 503713
rect 679624 503668 679676 503674
rect 683394 503639 683450 503648
rect 679624 503610 679676 503616
rect 679636 487257 679664 503610
rect 681004 503532 681056 503538
rect 681004 503474 681056 503480
rect 679622 487248 679678 487257
rect 679622 487183 679678 487192
rect 681016 486441 681044 503474
rect 683210 500984 683266 500993
rect 681188 500948 681240 500954
rect 683210 500919 683266 500928
rect 681188 500890 681240 500896
rect 681200 487665 681228 500890
rect 681186 487656 681242 487665
rect 681186 487591 681242 487600
rect 681002 486432 681058 486441
rect 681002 486367 681058 486376
rect 683224 483585 683252 500919
rect 683408 485625 683436 503639
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683394 485616 683450 485625
rect 683394 485551 683450 485560
rect 683210 483576 683266 483585
rect 683210 483511 683266 483520
rect 676220 482996 676272 483002
rect 676220 482938 676272 482944
rect 677416 482996 677468 483002
rect 677416 482938 677468 482944
rect 676034 482760 676090 482769
rect 676232 482746 676260 482938
rect 676090 482718 676260 482746
rect 676034 482695 676090 482704
rect 680358 481944 680414 481953
rect 680358 481879 680414 481888
rect 675850 480720 675906 480729
rect 675850 480655 675906 480664
rect 675864 454918 675892 480655
rect 680372 476134 680400 481879
rect 683118 481128 683174 481137
rect 683118 481063 683174 481072
rect 683132 480418 683160 481063
rect 683120 480412 683172 480418
rect 683120 480354 683172 480360
rect 676036 476128 676088 476134
rect 676036 476070 676088 476076
rect 680360 476128 680412 476134
rect 680360 476070 680412 476076
rect 675852 454912 675904 454918
rect 675852 454854 675904 454860
rect 672954 454368 673006 454374
rect 672952 454336 672954 454345
rect 674288 454368 674340 454374
rect 673006 454336 673008 454345
rect 672952 454271 673008 454280
rect 674286 454336 674288 454345
rect 675668 454368 675720 454374
rect 674340 454336 674342 454345
rect 675668 454310 675720 454316
rect 674286 454271 674342 454280
rect 676048 453966 676076 476070
rect 674288 453960 674340 453966
rect 674286 453928 674288 453937
rect 676036 453960 676088 453966
rect 674340 453928 674342 453937
rect 676036 453902 676088 453908
rect 674286 453863 674342 453872
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 676218 403336 676274 403345
rect 674564 403300 674616 403306
rect 676218 403271 676220 403280
rect 674564 403242 674616 403248
rect 676272 403271 676274 403280
rect 676220 403242 676272 403248
rect 673182 402384 673238 402393
rect 673182 402319 673238 402328
rect 672630 401704 672686 401713
rect 672630 401639 672686 401648
rect 672170 399664 672226 399673
rect 672170 399599 672226 399608
rect 671894 393544 671950 393553
rect 671894 393479 671950 393488
rect 671710 348936 671766 348945
rect 671710 348871 671766 348880
rect 671724 331265 671752 348871
rect 671710 331256 671766 331265
rect 671710 331191 671766 331200
rect 671526 302288 671582 302297
rect 671526 302223 671582 302232
rect 671344 278724 671396 278730
rect 671344 278666 671396 278672
rect 671342 260536 671398 260545
rect 671342 260471 671398 260480
rect 670698 257272 670754 257281
rect 670698 257207 670754 257216
rect 670516 226636 670568 226642
rect 670516 226578 670568 226584
rect 670516 224800 670568 224806
rect 670516 224742 670568 224748
rect 670528 224505 670556 224742
rect 670514 224496 670570 224505
rect 670514 224431 670570 224440
rect 670516 224052 670568 224058
rect 670516 223994 670568 224000
rect 670528 223689 670556 223994
rect 670514 223680 670570 223689
rect 670514 223615 670570 223624
rect 670344 223502 670648 223530
rect 670620 223258 670648 223502
rect 670160 218742 670280 218770
rect 670344 223230 670648 223258
rect 670160 186314 670188 218742
rect 670344 217410 670372 223230
rect 670516 223168 670568 223174
rect 670516 223110 670568 223116
rect 670528 222873 670556 223110
rect 670514 222864 670570 222873
rect 670514 222799 670570 222808
rect 670516 222692 670568 222698
rect 670516 222634 670568 222640
rect 670528 218929 670556 222634
rect 670514 218920 670570 218929
rect 670514 218855 670570 218864
rect 670344 217382 670464 217410
rect 670436 217138 670464 217382
rect 670344 217110 670464 217138
rect 670344 186314 670372 217110
rect 670514 216744 670570 216753
rect 670514 216679 670570 216688
rect 670528 198257 670556 216679
rect 670514 198248 670570 198257
rect 670514 198183 670570 198192
rect 670160 186286 670280 186314
rect 670344 186286 670464 186314
rect 670056 165096 670108 165102
rect 670056 165038 670108 165044
rect 670252 157334 670280 186286
rect 670436 175098 670464 186286
rect 670712 184890 670740 257207
rect 671356 240281 671384 260471
rect 671342 240272 671398 240281
rect 671342 240207 671398 240216
rect 671160 236632 671212 236638
rect 671160 236574 671212 236580
rect 670976 235952 671028 235958
rect 670976 235894 671028 235900
rect 670988 234614 671016 235894
rect 670988 234586 671108 234614
rect 670884 233232 670936 233238
rect 670884 233174 670936 233180
rect 670896 186314 670924 233174
rect 670896 186286 671016 186314
rect 670700 184884 670752 184890
rect 670700 184826 670752 184832
rect 670792 178016 670844 178022
rect 670790 177984 670792 177993
rect 670844 177984 670846 177993
rect 670790 177919 670846 177928
rect 670988 176654 671016 186286
rect 670896 176626 671016 176654
rect 670424 175092 670476 175098
rect 670424 175034 670476 175040
rect 670422 171184 670478 171193
rect 670422 171119 670478 171128
rect 670160 157306 670280 157334
rect 669872 133816 669924 133822
rect 669872 133758 669924 133764
rect 669962 130928 670018 130937
rect 669962 130863 670018 130872
rect 668950 125760 669006 125769
rect 668950 125695 669006 125704
rect 668766 119232 668822 119241
rect 668766 119167 668822 119176
rect 669226 118824 669282 118833
rect 669226 118759 669282 118768
rect 668768 116748 668820 116754
rect 668768 116690 668820 116696
rect 668780 112713 668808 116690
rect 669240 114345 669268 118759
rect 669226 114336 669282 114345
rect 669226 114271 669282 114280
rect 668766 112704 668822 112713
rect 668766 112639 668822 112648
rect 669976 108866 670004 130863
rect 670160 129742 670188 157306
rect 670436 155961 670464 171119
rect 670606 170232 670662 170241
rect 670606 170167 670662 170176
rect 670422 155952 670478 155961
rect 670422 155887 670478 155896
rect 670620 147665 670648 170167
rect 670896 166994 670924 176626
rect 670804 166966 670924 166994
rect 670804 160070 670832 166966
rect 670792 160064 670844 160070
rect 670792 160006 670844 160012
rect 671080 157334 671108 234586
rect 671172 224954 671200 236574
rect 671540 234614 671568 302223
rect 671712 278520 671764 278526
rect 671710 278488 671712 278497
rect 671764 278488 671766 278497
rect 671710 278423 671766 278432
rect 671710 259720 671766 259729
rect 671710 259655 671766 259664
rect 671724 245585 671752 259655
rect 671710 245576 671766 245585
rect 671710 245511 671766 245520
rect 671908 244274 671936 393479
rect 672184 355065 672212 399599
rect 672998 394768 673054 394777
rect 672998 394703 673054 394712
rect 672814 393952 672870 393961
rect 672814 393887 672870 393896
rect 672828 376281 672856 393887
rect 673012 381041 673040 394703
rect 672998 381032 673054 381041
rect 672998 380967 673054 380976
rect 672814 376272 672870 376281
rect 672814 376207 672870 376216
rect 673196 357513 673224 402319
rect 673918 401432 673974 401441
rect 673918 401367 673974 401376
rect 673366 400480 673422 400489
rect 673366 400415 673422 400424
rect 673182 357504 673238 357513
rect 673182 357439 673238 357448
rect 672354 357096 672410 357105
rect 672354 357031 672410 357040
rect 672170 355056 672226 355065
rect 672170 354991 672226 355000
rect 672170 353424 672226 353433
rect 672170 353359 672226 353368
rect 672184 337793 672212 353359
rect 672170 337784 672226 337793
rect 672170 337719 672226 337728
rect 672368 312497 672396 357031
rect 672538 356280 672594 356289
rect 672538 356215 672594 356224
rect 672354 312488 672410 312497
rect 672354 312423 672410 312432
rect 672552 311681 672580 356215
rect 673380 355881 673408 400415
rect 673734 396128 673790 396137
rect 673734 396063 673790 396072
rect 673748 381449 673776 396063
rect 673734 381440 673790 381449
rect 673734 381375 673790 381384
rect 673932 356561 673960 401367
rect 674576 396681 674604 403242
rect 676586 402928 676642 402937
rect 676586 402863 676642 402872
rect 674838 402656 674894 402665
rect 674838 402591 674894 402600
rect 674852 402121 674880 402591
rect 674838 402112 674894 402121
rect 674838 402047 674894 402056
rect 676600 400897 676628 402863
rect 676586 400888 676642 400897
rect 676586 400823 676642 400832
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 676048 398886 676076 399327
rect 674932 398880 674984 398886
rect 674932 398822 674984 398828
rect 676036 398880 676088 398886
rect 676036 398822 676088 398828
rect 674746 397352 674802 397361
rect 674746 397287 674802 397296
rect 674562 396672 674618 396681
rect 674562 396607 674618 396616
rect 674380 395548 674432 395554
rect 674380 395490 674432 395496
rect 674392 394482 674420 395490
rect 674208 394454 674420 394482
rect 674208 378026 674236 394454
rect 674472 394324 674524 394330
rect 674472 394266 674524 394272
rect 674484 378146 674512 394266
rect 674760 393314 674788 397287
rect 674944 395842 674972 398822
rect 679622 398440 679678 398449
rect 679622 398375 679678 398384
rect 676218 398032 676274 398041
rect 676218 397967 676274 397976
rect 674668 393286 674788 393314
rect 674852 395814 674972 395842
rect 674472 378140 674524 378146
rect 674472 378082 674524 378088
rect 674208 377998 674420 378026
rect 674392 375358 674420 377998
rect 674380 375352 674432 375358
rect 674380 375294 674432 375300
rect 674668 371566 674696 393286
rect 674852 386170 674880 395814
rect 676232 395758 676260 397967
rect 678242 397624 678298 397633
rect 678242 397559 678298 397568
rect 675024 395752 675076 395758
rect 675024 395694 675076 395700
rect 676220 395752 676272 395758
rect 676220 395694 676272 395700
rect 674840 386164 674892 386170
rect 674840 386106 674892 386112
rect 675036 382582 675064 395694
rect 676218 395584 676274 395593
rect 676218 395519 676220 395528
rect 676272 395519 676274 395528
rect 676220 395490 676272 395496
rect 676218 394360 676274 394369
rect 676218 394295 676220 394304
rect 676272 394295 676274 394304
rect 676220 394266 676272 394272
rect 678256 387705 678284 397559
rect 678242 387696 678298 387705
rect 678242 387631 678298 387640
rect 679636 386782 679664 398375
rect 679624 386776 679676 386782
rect 679624 386718 679676 386724
rect 675128 386261 675418 386289
rect 675128 383654 675156 386261
rect 675300 386164 675352 386170
rect 675300 386106 675352 386112
rect 675312 384449 675340 386106
rect 675484 386028 675536 386034
rect 675484 385970 675536 385976
rect 675496 385696 675524 385970
rect 675772 384985 675800 385084
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675312 384421 675418 384449
rect 675128 383626 675248 383654
rect 675220 382945 675248 383626
rect 675206 382936 675262 382945
rect 675206 382871 675262 382880
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 675036 382554 675340 382582
rect 675404 382568 675432 382622
rect 675758 382256 675814 382265
rect 675758 382191 675814 382200
rect 675772 382024 675800 382191
rect 675114 381440 675170 381449
rect 675170 381398 675418 381426
rect 675114 381375 675170 381384
rect 675390 381032 675446 381041
rect 675390 380967 675446 380976
rect 675404 380732 675432 380967
rect 675758 378720 675814 378729
rect 675758 378655 675814 378664
rect 675772 378284 675800 378655
rect 675116 378140 675168 378146
rect 675116 378082 675168 378088
rect 675128 377754 675156 378082
rect 675128 377726 675340 377754
rect 675312 377618 675340 377726
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675758 377360 675814 377369
rect 675758 377295 675814 377304
rect 675772 377060 675800 377295
rect 675404 376281 675432 376448
rect 675390 376272 675446 376281
rect 675390 376207 675446 376216
rect 675116 375352 675168 375358
rect 675116 375294 675168 375300
rect 675128 375238 675156 375294
rect 675128 375210 675418 375238
rect 675758 373688 675814 373697
rect 675758 373623 675814 373632
rect 675772 373388 675800 373623
rect 675404 372473 675432 372776
rect 675390 372464 675446 372473
rect 675390 372399 675446 372408
rect 674668 371538 675418 371566
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 674470 358320 674526 358329
rect 674470 358255 674526 358264
rect 673918 356552 673974 356561
rect 673918 356487 673974 356496
rect 673366 355872 673422 355881
rect 673366 355807 673422 355816
rect 673182 355464 673238 355473
rect 673182 355399 673238 355408
rect 672998 349752 673054 349761
rect 672998 349687 673054 349696
rect 672722 348528 672778 348537
rect 672722 348463 672778 348472
rect 672538 311672 672594 311681
rect 672538 311607 672594 311616
rect 672538 305552 672594 305561
rect 672538 305487 672594 305496
rect 672172 288448 672224 288454
rect 672172 288390 672224 288396
rect 672184 246129 672212 288390
rect 672552 285569 672580 305487
rect 672538 285560 672594 285569
rect 672538 285495 672594 285504
rect 672356 284368 672408 284374
rect 672356 284310 672408 284316
rect 672170 246120 672226 246129
rect 672170 246055 672226 246064
rect 671816 244246 671936 244274
rect 671816 236745 671844 244246
rect 672172 237108 672224 237114
rect 672172 237050 672224 237056
rect 671802 236736 671858 236745
rect 671802 236671 671858 236680
rect 671988 236496 672040 236502
rect 671724 236456 671988 236484
rect 671540 234586 671660 234614
rect 671344 234388 671396 234394
rect 671344 234330 671396 234336
rect 671172 224926 671292 224954
rect 671264 186314 671292 224926
rect 671356 215294 671384 234330
rect 671632 224777 671660 234586
rect 671724 224954 671752 236456
rect 671988 236438 672040 236444
rect 671988 235340 672040 235346
rect 671988 235282 672040 235288
rect 672000 232898 672028 235282
rect 672184 234530 672212 237050
rect 672172 234524 672224 234530
rect 672172 234466 672224 234472
rect 671988 232892 672040 232898
rect 671988 232834 672040 232840
rect 672172 230988 672224 230994
rect 672172 230930 672224 230936
rect 672184 229770 672212 230930
rect 672172 229764 672224 229770
rect 672172 229706 672224 229712
rect 672368 227089 672396 284310
rect 672736 282914 672764 348463
rect 673012 335617 673040 349687
rect 672998 335608 673054 335617
rect 672998 335543 673054 335552
rect 672906 325000 672962 325009
rect 672906 324935 672962 324944
rect 672920 287054 672948 324935
rect 673196 310865 673224 355399
rect 673918 354648 673974 354657
rect 673918 354583 673974 354592
rect 673734 352608 673790 352617
rect 673734 352543 673790 352552
rect 673366 350160 673422 350169
rect 673366 350095 673422 350104
rect 673380 335889 673408 350095
rect 673550 349344 673606 349353
rect 673550 349279 673606 349288
rect 673366 335880 673422 335889
rect 673366 335815 673422 335824
rect 673564 332761 673592 349279
rect 673748 333985 673776 352543
rect 673734 333976 673790 333985
rect 673734 333911 673790 333920
rect 673550 332752 673606 332761
rect 673550 332687 673606 332696
rect 673182 310856 673238 310865
rect 673182 310791 673238 310800
rect 673932 310049 673960 354583
rect 674286 351384 674342 351393
rect 674286 351319 674342 351328
rect 674300 338065 674328 351319
rect 674484 351121 674512 358255
rect 675942 357912 675998 357921
rect 675942 357847 675998 357856
rect 675956 356833 675984 357847
rect 675942 356824 675998 356833
rect 675942 356759 675998 356768
rect 674654 352200 674710 352209
rect 674654 352135 674710 352144
rect 674470 351112 674526 351121
rect 674470 351047 674526 351056
rect 674470 350568 674526 350577
rect 674470 350503 674526 350512
rect 674286 338056 674342 338065
rect 674286 337991 674342 338000
rect 674484 331090 674512 350503
rect 674472 331084 674524 331090
rect 674472 331026 674524 331032
rect 674668 326913 674696 352135
rect 676034 350976 676090 350985
rect 676034 350911 676090 350920
rect 676048 346633 676076 350911
rect 676034 346624 676090 346633
rect 676034 346559 676090 346568
rect 675128 341074 675418 341102
rect 675128 338745 675156 341074
rect 675404 340082 675432 340544
rect 675758 340232 675814 340241
rect 675758 340167 675814 340176
rect 675312 340054 675432 340082
rect 675114 338736 675170 338745
rect 675114 338671 675170 338680
rect 675114 338056 675170 338065
rect 675114 337991 675170 338000
rect 675128 336857 675156 337991
rect 675312 337793 675340 340054
rect 675772 339864 675800 340167
rect 675482 339416 675538 339425
rect 675482 339351 675538 339360
rect 675496 339252 675524 339351
rect 675758 337920 675814 337929
rect 675758 337855 675814 337864
rect 675298 337784 675354 337793
rect 675298 337719 675354 337728
rect 675772 337416 675800 337855
rect 675128 336829 675418 336857
rect 675758 336560 675814 336569
rect 675758 336495 675814 336504
rect 675772 336192 675800 336495
rect 674930 335880 674986 335889
rect 674930 335815 674986 335824
rect 674944 331889 674972 335815
rect 675114 335608 675170 335617
rect 675170 335566 675340 335594
rect 675114 335543 675170 335552
rect 675312 335458 675340 335566
rect 675404 335458 675432 335580
rect 675312 335430 675432 335458
rect 675114 333976 675170 333985
rect 675114 333911 675170 333920
rect 675128 333078 675156 333911
rect 675128 333050 675418 333078
rect 675114 332752 675170 332761
rect 675114 332687 675170 332696
rect 675128 332534 675156 332687
rect 675128 332506 675418 332534
rect 674944 331861 675418 331889
rect 675114 331256 675170 331265
rect 675170 331214 675418 331242
rect 675114 331191 675170 331200
rect 675116 331084 675168 331090
rect 675116 331026 675168 331032
rect 675128 330049 675156 331026
rect 675128 330021 675418 330049
rect 675312 328222 675432 328250
rect 675312 328182 675340 328222
rect 675220 328154 675340 328182
rect 675404 328168 675432 328222
rect 675022 327992 675078 328001
rect 675022 327927 675078 327936
rect 674654 326904 674710 326913
rect 674654 326839 674710 326848
rect 675036 325009 675064 327927
rect 675220 325689 675248 328154
rect 675390 327992 675446 328001
rect 675390 327927 675446 327936
rect 675404 327556 675432 327927
rect 675390 326904 675446 326913
rect 675390 326839 675446 326848
rect 675404 326332 675432 326839
rect 675206 325680 675262 325689
rect 675206 325615 675262 325624
rect 675022 325000 675078 325009
rect 675022 324935 675078 324944
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676218 313984 676274 313993
rect 676218 313919 676274 313928
rect 674838 312896 674894 312905
rect 674838 312831 674894 312840
rect 674380 312044 674432 312050
rect 674380 311986 674432 311992
rect 674392 311894 674420 311986
rect 674852 311953 674880 312831
rect 675482 312080 675538 312089
rect 675482 312015 675484 312024
rect 675536 312015 675538 312024
rect 675484 311986 675536 311992
rect 674208 311866 674420 311894
rect 674838 311944 674894 311953
rect 674838 311879 674894 311888
rect 673918 310040 673974 310049
rect 673918 309975 673974 309984
rect 673274 309496 673330 309505
rect 673274 309431 673330 309440
rect 673090 304328 673146 304337
rect 673090 304263 673146 304272
rect 673104 287881 673132 304263
rect 673090 287872 673146 287881
rect 673090 287807 673146 287816
rect 672644 282886 672764 282914
rect 672828 287026 672948 287054
rect 672644 273254 672672 282886
rect 672828 278497 672856 287026
rect 672814 278488 672870 278497
rect 672814 278423 672870 278432
rect 672644 273226 672764 273254
rect 672538 265296 672594 265305
rect 672538 265231 672594 265240
rect 672552 228426 672580 265231
rect 672736 234614 672764 273226
rect 673090 266112 673146 266121
rect 673090 266047 673146 266056
rect 673104 263594 673132 266047
rect 673288 265033 673316 309431
rect 673826 305960 673882 305969
rect 673826 305895 673882 305904
rect 673840 291553 673868 305895
rect 674010 291816 674066 291825
rect 674010 291751 674066 291760
rect 673826 291544 673882 291553
rect 673826 291479 673882 291488
rect 673458 287600 673514 287609
rect 673458 287535 673514 287544
rect 673274 265024 673330 265033
rect 673274 264959 673330 264968
rect 673104 263566 673316 263594
rect 673090 263392 673146 263401
rect 673090 263327 673146 263336
rect 672906 259312 672962 259321
rect 672906 259247 672962 259256
rect 672920 242729 672948 259247
rect 673104 250753 673132 263327
rect 673090 250744 673146 250753
rect 673090 250679 673146 250688
rect 673090 249656 673146 249665
rect 673090 249591 673146 249600
rect 673104 245857 673132 249591
rect 673090 245848 673146 245857
rect 673090 245783 673146 245792
rect 672906 242720 672962 242729
rect 672906 242655 672962 242664
rect 673288 241777 673316 263566
rect 673472 246265 673500 287535
rect 674024 268161 674052 291751
rect 674208 282914 674236 311866
rect 674746 311264 674802 311273
rect 674746 311199 674802 311208
rect 674562 310448 674618 310457
rect 674562 310383 674618 310392
rect 674378 303920 674434 303929
rect 674378 303855 674434 303864
rect 674392 286686 674420 303855
rect 674576 292574 674604 310383
rect 674760 292574 674788 311199
rect 675942 309768 675998 309777
rect 676232 309754 676260 313919
rect 675998 309726 676260 309754
rect 675942 309703 675998 309712
rect 675114 308408 675170 308417
rect 675114 308343 675170 308352
rect 674930 306368 674986 306377
rect 674930 306303 674986 306312
rect 674944 299474 674972 306303
rect 675128 302234 675156 308343
rect 675298 308000 675354 308009
rect 675298 307935 675354 307944
rect 675312 302234 675340 307935
rect 676034 307592 676090 307601
rect 676090 307550 676444 307578
rect 676034 307527 676090 307536
rect 676034 307184 676090 307193
rect 676090 307142 676260 307170
rect 676034 307119 676090 307128
rect 676232 306406 676260 307142
rect 676220 306400 676272 306406
rect 676220 306342 676272 306348
rect 676416 304910 676444 307550
rect 678242 306776 678298 306785
rect 678242 306711 678298 306720
rect 676864 306400 676916 306406
rect 676864 306342 676916 306348
rect 675852 304904 675904 304910
rect 675852 304846 675904 304852
rect 676404 304904 676456 304910
rect 676404 304846 676456 304852
rect 675864 302234 675892 304846
rect 676586 304736 676642 304745
rect 676586 304671 676642 304680
rect 676034 303512 676090 303521
rect 676034 303447 676090 303456
rect 674852 299446 674972 299474
rect 675036 302206 675156 302234
rect 675220 302206 675340 302234
rect 675404 302206 675892 302234
rect 674852 293706 674880 299446
rect 675036 297673 675064 302206
rect 675220 299474 675248 302206
rect 675404 299474 675432 302206
rect 676048 302025 676076 303447
rect 676034 302016 676090 302025
rect 676034 301951 676090 301960
rect 676600 301617 676628 304671
rect 676586 301608 676642 301617
rect 676586 301543 676642 301552
rect 675220 299446 675340 299474
rect 675404 299446 675524 299474
rect 675022 297664 675078 297673
rect 675022 297599 675078 297608
rect 675312 296206 675340 299446
rect 675496 298217 675524 299446
rect 675482 298208 675538 298217
rect 675482 298143 675538 298152
rect 675852 298104 675904 298110
rect 675496 298052 675852 298058
rect 675496 298046 675904 298052
rect 675496 298030 675892 298046
rect 675496 296410 675524 298030
rect 676876 297401 676904 306342
rect 678256 298110 678284 306711
rect 678244 298104 678296 298110
rect 678244 298046 678296 298052
rect 676862 297392 676918 297401
rect 676862 297327 676918 297336
rect 675484 296404 675536 296410
rect 675484 296346 675536 296352
rect 675300 296200 675352 296206
rect 675300 296142 675352 296148
rect 675404 295905 675432 296072
rect 675390 295896 675446 295905
rect 675390 295831 675446 295840
rect 675574 295760 675630 295769
rect 675574 295695 675630 295704
rect 675588 295528 675616 295695
rect 675300 295452 675352 295458
rect 675300 295394 675352 295400
rect 674852 293678 675064 293706
rect 674484 292546 674604 292574
rect 674668 292546 674788 292574
rect 674484 287054 674512 292546
rect 674668 287054 674696 292546
rect 674838 292496 674894 292505
rect 674838 292431 674894 292440
rect 674852 288062 674880 292431
rect 675036 291870 675064 293678
rect 675312 292414 675340 295394
rect 675484 295248 675536 295254
rect 675484 295190 675536 295196
rect 675496 294879 675524 295190
rect 675758 294672 675814 294681
rect 675758 294607 675814 294616
rect 675772 294236 675800 294607
rect 675312 292386 675418 292414
rect 675036 291842 675418 291870
rect 675390 291544 675446 291553
rect 675390 291479 675446 291488
rect 675404 291176 675432 291479
rect 675758 291000 675814 291009
rect 675758 290935 675814 290944
rect 675772 290564 675800 290935
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 674852 288034 675340 288062
rect 675404 288048 675432 288102
rect 675114 287872 675170 287881
rect 675114 287807 675170 287816
rect 675128 287518 675156 287807
rect 675128 287490 675418 287518
rect 675758 287056 675814 287065
rect 674484 287026 674604 287054
rect 674668 287026 674788 287054
rect 674380 286680 674432 286686
rect 674380 286622 674432 286628
rect 674208 282886 674420 282914
rect 674010 268152 674066 268161
rect 674010 268087 674066 268096
rect 674392 267481 674420 282886
rect 674378 267472 674434 267481
rect 674378 267407 674434 267416
rect 673918 267064 673974 267073
rect 673918 266999 673974 267008
rect 673734 264616 673790 264625
rect 673734 264551 673790 264560
rect 673458 246256 673514 246265
rect 673458 246191 673514 246200
rect 673748 242049 673776 264551
rect 673734 242040 673790 242049
rect 673734 241975 673790 241984
rect 673274 241768 673330 241777
rect 673274 241703 673330 241712
rect 673932 239442 673960 266999
rect 674576 265849 674604 287026
rect 674760 266665 674788 287026
rect 675758 286991 675814 287000
rect 675772 286892 675800 286991
rect 675300 286680 675352 286686
rect 675300 286622 675352 286628
rect 675312 286498 675340 286622
rect 675312 286470 675432 286498
rect 675404 286212 675432 286470
rect 675114 285560 675170 285569
rect 675114 285495 675170 285504
rect 675128 285070 675156 285495
rect 675128 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675758 282704 675814 282713
rect 675758 282639 675814 282648
rect 675772 282554 675800 282639
rect 675312 282540 675800 282554
rect 675312 282526 675786 282540
rect 675312 278769 675340 282526
rect 675666 281616 675722 281625
rect 675666 281551 675722 281560
rect 675680 281355 675708 281551
rect 676862 279440 676918 279449
rect 676862 279375 676918 279384
rect 675298 278760 675354 278769
rect 675298 278695 675354 278704
rect 675482 278080 675538 278089
rect 675482 278015 675538 278024
rect 674746 266656 674802 266665
rect 674746 266591 674802 266600
rect 674562 265840 674618 265849
rect 674562 265775 674618 265784
rect 674654 262576 674710 262585
rect 674654 262511 674710 262520
rect 674102 260944 674158 260953
rect 674102 260879 674158 260888
rect 674116 246673 674144 260879
rect 674286 260128 674342 260137
rect 674286 260063 674342 260072
rect 674102 246664 674158 246673
rect 674102 246599 674158 246608
rect 674300 242321 674328 260063
rect 674470 258904 674526 258913
rect 674470 258839 674526 258848
rect 674286 242312 674342 242321
rect 674286 242247 674342 242256
rect 674484 241505 674512 258839
rect 674668 243710 674696 262511
rect 675496 258097 675524 278015
rect 676876 268569 676904 279375
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 676862 268560 676918 268569
rect 676862 268495 676918 268504
rect 676218 268152 676274 268161
rect 676218 268087 676274 268096
rect 676232 267753 676260 268087
rect 676218 267744 676274 267753
rect 676218 267679 676274 267688
rect 676402 264072 676458 264081
rect 676402 264007 676458 264016
rect 676218 262848 676274 262857
rect 676218 262783 676274 262792
rect 676232 260930 676260 262783
rect 675680 260902 676260 260930
rect 675482 258088 675538 258097
rect 675482 258023 675538 258032
rect 675680 257938 675708 260902
rect 676416 259486 676444 264007
rect 679622 263664 679678 263673
rect 679622 263599 679678 263608
rect 675852 259480 675904 259486
rect 675852 259422 675904 259428
rect 676404 259480 676456 259486
rect 676404 259422 676456 259428
rect 675128 257910 675708 257938
rect 674930 253192 674986 253201
rect 674930 253127 674986 253136
rect 674944 248962 674972 253127
rect 675128 253042 675156 257910
rect 675864 253934 675892 259422
rect 675036 253014 675156 253042
rect 675220 253906 675892 253934
rect 675036 251174 675064 253014
rect 675036 251146 675156 251174
rect 674760 248934 674972 248962
rect 674760 245834 674788 248934
rect 674930 248840 674986 248849
rect 674930 248775 674986 248784
rect 674944 246213 674972 248775
rect 675128 247398 675156 251146
rect 675220 249370 675248 253906
rect 675850 253192 675906 253201
rect 679636 253162 679664 263599
rect 675850 253127 675852 253136
rect 675904 253127 675906 253136
rect 679624 253156 679676 253162
rect 675852 253098 675904 253104
rect 679624 253098 679676 253104
rect 675312 251110 675432 251138
rect 675312 249642 675340 251110
rect 675404 251056 675432 251110
rect 675482 250744 675538 250753
rect 675482 250679 675538 250688
rect 675496 250512 675524 250679
rect 675758 250336 675814 250345
rect 675758 250271 675814 250280
rect 675772 249900 675800 250271
rect 675312 249626 675432 249642
rect 675312 249620 675444 249626
rect 675312 249614 675392 249620
rect 675392 249562 675444 249568
rect 675220 249342 675432 249370
rect 675404 249220 675432 249342
rect 675392 248532 675444 248538
rect 675392 248474 675444 248480
rect 675404 248305 675432 248474
rect 675390 248296 675446 248305
rect 675390 248231 675446 248240
rect 675128 247370 675418 247398
rect 675772 246673 675800 246840
rect 675298 246664 675354 246673
rect 675298 246599 675354 246608
rect 675758 246664 675814 246673
rect 675758 246599 675814 246608
rect 675312 246213 675340 246599
rect 674944 246185 675064 246213
rect 675312 246185 675418 246213
rect 674760 245806 674880 245834
rect 674656 243704 674708 243710
rect 674656 243646 674708 243652
rect 674852 243234 674880 245806
rect 674840 243228 674892 243234
rect 674840 243170 674892 243176
rect 674838 241768 674894 241777
rect 674838 241703 674894 241712
rect 674470 241496 674526 241505
rect 674470 241431 674526 241440
rect 673932 239414 674420 239442
rect 672952 236736 673008 236745
rect 672952 236671 672954 236680
rect 673006 236671 673008 236680
rect 674194 236736 674250 236745
rect 674194 236671 674250 236680
rect 672954 236642 673006 236648
rect 673184 236292 673236 236298
rect 673184 236234 673236 236240
rect 673196 236178 673224 236234
rect 673196 236150 673776 236178
rect 672908 235952 672960 235958
rect 672506 228410 672580 228426
rect 672494 228404 672580 228410
rect 672546 228398 672580 228404
rect 672644 234586 672764 234614
rect 672828 235900 672908 235906
rect 672828 235894 672960 235900
rect 672828 235878 672948 235894
rect 672494 228346 672546 228352
rect 672354 227080 672410 227089
rect 672644 227066 672672 234586
rect 672828 232937 672856 235878
rect 673000 235748 673052 235754
rect 673000 235690 673052 235696
rect 673012 233442 673040 235690
rect 673184 235544 673236 235550
rect 673184 235486 673236 235492
rect 673000 233436 673052 233442
rect 673000 233378 673052 233384
rect 673196 233322 673224 235486
rect 673552 234524 673604 234530
rect 673552 234466 673604 234472
rect 673104 233294 673224 233322
rect 672814 232928 672870 232937
rect 672814 232863 672870 232872
rect 673104 230330 673132 233294
rect 673564 231854 673592 234466
rect 673564 231826 673684 231854
rect 672552 227050 672672 227066
rect 672354 227015 672410 227024
rect 672540 227044 672672 227050
rect 672592 227038 672672 227044
rect 672736 230302 673132 230330
rect 672540 226986 672592 226992
rect 672736 226930 672764 230302
rect 673092 230240 673144 230246
rect 673092 230182 673144 230188
rect 672908 229628 672960 229634
rect 672908 229570 672960 229576
rect 672368 226902 672764 226930
rect 672172 225888 672224 225894
rect 672172 225830 672224 225836
rect 672184 225729 672212 225830
rect 671986 225720 672042 225729
rect 671986 225655 672042 225664
rect 672170 225720 672226 225729
rect 672368 225706 672396 226902
rect 672724 226432 672776 226438
rect 672722 226400 672724 226409
rect 672776 226400 672778 226409
rect 672722 226335 672778 226344
rect 672604 226160 672656 226166
rect 672602 226128 672604 226137
rect 672656 226128 672658 226137
rect 672602 226063 672658 226072
rect 672492 225992 672548 226001
rect 672492 225927 672494 225936
rect 672546 225927 672548 225936
rect 672494 225898 672546 225904
rect 672368 225678 672488 225706
rect 672170 225655 672226 225664
rect 672000 225298 672028 225655
rect 672264 225548 672316 225554
rect 672264 225490 672316 225496
rect 672156 225412 672208 225418
rect 672156 225354 672208 225360
rect 672000 225282 672074 225298
rect 672000 225276 672086 225282
rect 672000 225270 672034 225276
rect 672034 225218 672086 225224
rect 672168 225049 672196 225354
rect 672276 225321 672304 225490
rect 672262 225312 672318 225321
rect 672262 225247 672318 225256
rect 672168 225040 672226 225049
rect 672168 224998 672170 225040
rect 672170 224975 672226 224984
rect 672460 224954 672488 225678
rect 671724 224926 671844 224954
rect 671618 224768 671674 224777
rect 671618 224703 671674 224712
rect 671480 224496 671536 224505
rect 671480 224431 671536 224440
rect 671494 224330 671522 224431
rect 671596 224392 671648 224398
rect 671596 224334 671648 224340
rect 671482 224324 671534 224330
rect 671482 224266 671534 224272
rect 671608 224233 671636 224334
rect 671594 224224 671650 224233
rect 671594 224159 671650 224168
rect 671618 223952 671674 223961
rect 671618 223887 671674 223896
rect 671632 222194 671660 223887
rect 671632 222166 671752 222194
rect 671724 219450 671752 222166
rect 671540 219422 671752 219450
rect 671356 215266 671476 215294
rect 671448 186314 671476 215266
rect 671172 186286 671292 186314
rect 671356 186286 671476 186314
rect 671172 176654 671200 186286
rect 671356 177993 671384 186286
rect 671342 177984 671398 177993
rect 671342 177919 671398 177928
rect 671172 176626 671292 176654
rect 670988 157306 671108 157334
rect 670988 155666 671016 157306
rect 670804 155638 671016 155666
rect 670804 155582 670832 155638
rect 670792 155576 670844 155582
rect 670792 155518 670844 155524
rect 671264 151814 671292 176626
rect 670804 151786 671292 151814
rect 670606 147656 670662 147665
rect 670606 147591 670662 147600
rect 670804 145790 670832 151786
rect 670792 145784 670844 145790
rect 670792 145726 670844 145732
rect 671540 138014 671568 219422
rect 671816 215294 671844 224926
rect 672368 224926 672488 224954
rect 672078 224496 672134 224505
rect 672078 224431 672134 224440
rect 672092 217569 672120 224431
rect 672368 220130 672396 224926
rect 672538 220280 672594 220289
rect 672538 220215 672594 220224
rect 672276 220102 672396 220130
rect 672078 217560 672134 217569
rect 672078 217495 672134 217504
rect 671986 217288 672042 217297
rect 671986 217223 672042 217232
rect 672000 216753 672028 217223
rect 671986 216744 672042 216753
rect 671986 216679 672042 216688
rect 672078 216064 672134 216073
rect 672078 215999 672134 216008
rect 672092 215393 672120 215999
rect 672078 215384 672134 215393
rect 672078 215319 672134 215328
rect 671724 215266 671844 215294
rect 671724 150113 671752 215266
rect 672078 214160 672134 214169
rect 672078 214095 672134 214104
rect 672092 199753 672120 214095
rect 672078 199744 672134 199753
rect 672078 199679 672134 199688
rect 672276 176654 672304 220102
rect 672552 217818 672580 220215
rect 672368 217790 672580 217818
rect 672368 205634 672396 217790
rect 672538 216744 672594 216753
rect 672538 216679 672594 216688
rect 672552 213217 672580 216679
rect 672920 215294 672948 229570
rect 673104 228585 673132 230182
rect 673276 230036 673328 230042
rect 673276 229978 673328 229984
rect 673288 229129 673316 229978
rect 673460 229424 673512 229430
rect 673460 229366 673512 229372
rect 673274 229120 673330 229129
rect 673274 229055 673330 229064
rect 673090 228576 673146 228585
rect 673090 228511 673146 228520
rect 673092 228404 673144 228410
rect 673092 228346 673144 228352
rect 673104 220697 673132 228346
rect 673472 227089 673500 229366
rect 673458 227080 673514 227089
rect 673458 227015 673514 227024
rect 673276 226568 673328 226574
rect 673276 226510 673328 226516
rect 673288 222601 673316 226510
rect 673274 222592 673330 222601
rect 673274 222527 673330 222536
rect 673274 221096 673330 221105
rect 673274 221031 673330 221040
rect 673090 220688 673146 220697
rect 673090 220623 673146 220632
rect 673090 216200 673146 216209
rect 673090 216135 673146 216144
rect 673104 215294 673132 216135
rect 672736 215266 672948 215294
rect 673012 215266 673132 215294
rect 672736 213625 672764 215266
rect 672722 213616 672778 213625
rect 672722 213551 672778 213560
rect 672814 213344 672870 213353
rect 672814 213279 672870 213288
rect 672538 213208 672594 213217
rect 672538 213143 672594 213152
rect 672630 212120 672686 212129
rect 672630 212055 672686 212064
rect 672368 205606 672488 205634
rect 672184 176626 672304 176654
rect 671986 172000 672042 172009
rect 671986 171935 672042 171944
rect 671710 150104 671766 150113
rect 671710 150039 671766 150048
rect 672000 144945 672028 171935
rect 672184 168065 672212 176626
rect 672460 175681 672488 205606
rect 672446 175672 672502 175681
rect 672446 175607 672502 175616
rect 672354 168328 672410 168337
rect 672354 168263 672410 168272
rect 672170 168056 672226 168065
rect 672170 167991 672226 168000
rect 672368 167634 672396 168263
rect 672184 167606 672396 167634
rect 671986 144936 672042 144945
rect 671986 144871 672042 144880
rect 670804 137986 671568 138014
rect 670804 130830 670832 137986
rect 672184 135153 672212 167606
rect 672354 166968 672410 166977
rect 672354 166903 672410 166912
rect 672170 135144 672226 135153
rect 672170 135079 672226 135088
rect 671342 131744 671398 131753
rect 671342 131679 671398 131688
rect 670792 130824 670844 130830
rect 670792 130766 670844 130772
rect 670148 129736 670200 129742
rect 670148 129678 670200 129684
rect 670422 121680 670478 121689
rect 670422 121615 670478 121624
rect 670436 116754 670464 121615
rect 670424 116748 670476 116754
rect 670424 116690 670476 116696
rect 671356 109034 671384 131679
rect 671526 129296 671582 129305
rect 671526 129231 671582 129240
rect 671540 109034 671568 129231
rect 672170 124944 672226 124953
rect 672170 124879 672226 124888
rect 670804 109006 671384 109034
rect 671448 109006 671568 109034
rect 669964 108860 670016 108866
rect 669964 108802 670016 108808
rect 670804 106214 670832 109006
rect 670792 106208 670844 106214
rect 670792 106150 670844 106156
rect 671448 104802 671476 109006
rect 670804 104774 671476 104802
rect 670804 104718 670832 104774
rect 668768 104712 668820 104718
rect 668768 104654 668820 104660
rect 670792 104712 670844 104718
rect 672184 104689 672212 124879
rect 672368 115841 672396 166903
rect 672644 122834 672672 212055
rect 672828 124137 672856 213279
rect 673012 201385 673040 215266
rect 672998 201376 673054 201385
rect 672998 201311 673054 201320
rect 673090 200832 673146 200841
rect 673090 200767 673146 200776
rect 673104 181529 673132 200767
rect 673288 197985 673316 221031
rect 673458 216472 673514 216481
rect 673458 216407 673514 216416
rect 673472 213897 673500 216407
rect 673458 213888 673514 213897
rect 673458 213823 673514 213832
rect 673274 197976 673330 197985
rect 673274 197911 673330 197920
rect 673090 181520 673146 181529
rect 673090 181455 673146 181464
rect 673182 176896 673238 176905
rect 673182 176831 673238 176840
rect 673196 170626 673224 176831
rect 673458 170776 673514 170785
rect 673458 170711 673514 170720
rect 673196 170598 673316 170626
rect 672998 169144 673054 169153
rect 672998 169079 673054 169088
rect 673012 168858 673040 169079
rect 672920 168830 673040 168858
rect 672920 157334 672948 168830
rect 673090 168736 673146 168745
rect 673090 168671 673146 168680
rect 673104 166994 673132 168671
rect 673288 166994 673316 170598
rect 673472 166994 673500 170711
rect 673656 166994 673684 231826
rect 673748 171850 673776 236150
rect 673874 235136 673926 235142
rect 673874 235078 673926 235084
rect 673886 234818 673914 235078
rect 673886 234790 674052 234818
rect 673872 230208 673928 230217
rect 673872 230143 673928 230152
rect 673886 229838 673914 230143
rect 673874 229832 673926 229838
rect 673874 229774 673926 229780
rect 673874 229152 673926 229158
rect 673874 229094 673926 229100
rect 673886 228721 673914 229094
rect 673872 228712 673928 228721
rect 673872 228647 673928 228656
rect 674024 224954 674052 234790
rect 674208 234614 674236 236671
rect 674392 234614 674420 239414
rect 674852 234614 674880 241703
rect 675036 237538 675064 246185
rect 675206 245576 675262 245585
rect 675262 245534 675418 245562
rect 675206 245511 675262 245520
rect 675208 243704 675260 243710
rect 675208 243646 675260 243652
rect 675220 243085 675248 243646
rect 675220 243057 675418 243085
rect 675208 242956 675260 242962
rect 675208 242898 675260 242904
rect 675220 238218 675248 242898
rect 675390 242720 675446 242729
rect 675390 242655 675446 242664
rect 675404 242519 675432 242655
rect 675390 242312 675446 242321
rect 675390 242247 675446 242256
rect 675404 241876 675432 242247
rect 675390 241496 675446 241505
rect 675390 241431 675446 241440
rect 675404 241231 675432 241431
rect 675390 240272 675446 240281
rect 675390 240207 675446 240216
rect 675404 240040 675432 240207
rect 675220 238190 675418 238218
rect 675312 237646 675432 237674
rect 675312 237538 675340 237646
rect 675036 237510 675340 237538
rect 675404 237524 675432 237646
rect 675114 237280 675170 237289
rect 675114 237215 675170 237224
rect 675128 236382 675156 237215
rect 675128 236354 675418 236382
rect 676034 235240 676090 235249
rect 676034 235175 676090 235184
rect 674208 234586 674328 234614
rect 674392 234586 674604 234614
rect 674852 234586 675156 234614
rect 674024 224926 674144 224954
rect 673918 217696 673974 217705
rect 673918 217631 673974 217640
rect 673932 177313 673960 217631
rect 673918 177304 673974 177313
rect 673918 177239 673974 177248
rect 673918 174448 673974 174457
rect 673918 174383 673974 174392
rect 673748 171822 673868 171850
rect 673104 166966 673224 166994
rect 673288 166966 673408 166994
rect 673472 166966 673592 166994
rect 673656 166966 673776 166994
rect 673196 157334 673224 166966
rect 672920 157306 673132 157334
rect 673196 157306 673316 157334
rect 673104 152697 673132 157306
rect 673090 152688 673146 152697
rect 673090 152623 673146 152632
rect 673288 151814 673316 157306
rect 673196 151786 673316 151814
rect 673196 151337 673224 151786
rect 673182 151328 673238 151337
rect 673182 151263 673238 151272
rect 672998 133512 673054 133521
rect 672998 133447 673054 133456
rect 673012 132705 673040 133447
rect 672998 132696 673054 132705
rect 672998 132631 673054 132640
rect 673380 132161 673408 166966
rect 673564 156505 673592 166966
rect 673748 164234 673776 166966
rect 673656 164206 673776 164234
rect 673656 156618 673684 164206
rect 673840 162897 673868 171822
rect 673932 166994 673960 174383
rect 674116 172961 674144 224926
rect 674102 172952 674158 172961
rect 674102 172887 674158 172896
rect 673932 166966 674052 166994
rect 674024 164234 674052 166966
rect 674024 164206 674236 164234
rect 673826 162888 673882 162897
rect 673826 162823 673882 162832
rect 674208 162194 674236 164206
rect 673932 162166 674236 162194
rect 673656 156590 673776 156618
rect 673550 156496 673606 156505
rect 673550 156431 673606 156440
rect 673550 156224 673606 156233
rect 673748 156210 673776 156590
rect 673606 156182 673776 156210
rect 673550 156159 673606 156168
rect 673366 132152 673422 132161
rect 673366 132087 673422 132096
rect 673932 129713 673960 162166
rect 674102 162072 674158 162081
rect 674102 162007 674158 162016
rect 673918 129704 673974 129713
rect 673918 129639 673974 129648
rect 673366 126576 673422 126585
rect 673366 126511 673422 126520
rect 672814 124128 672870 124137
rect 672814 124063 672870 124072
rect 672998 123312 673054 123321
rect 672998 123247 673054 123256
rect 672552 122806 672672 122834
rect 672552 120873 672580 122806
rect 672538 120864 672594 120873
rect 673012 120850 673040 123247
rect 673182 123040 673238 123049
rect 673182 122975 673238 122984
rect 672538 120799 672594 120808
rect 672828 120822 673040 120850
rect 672828 118833 672856 120822
rect 672998 120728 673054 120737
rect 672998 120663 673054 120672
rect 672814 118824 672870 118833
rect 672814 118759 672870 118768
rect 672354 115832 672410 115841
rect 672354 115767 672410 115776
rect 673012 111081 673040 120663
rect 672998 111072 673054 111081
rect 672998 111007 673054 111016
rect 673196 106321 673224 122975
rect 673182 106312 673238 106321
rect 673182 106247 673238 106256
rect 670792 104654 670844 104660
rect 672170 104680 672226 104689
rect 668780 104553 668808 104654
rect 672170 104615 672226 104624
rect 668766 104544 668822 104553
rect 668766 104479 668822 104488
rect 668582 102912 668638 102921
rect 668582 102847 668638 102856
rect 673380 101017 673408 126511
rect 673918 124536 673974 124545
rect 673918 124471 673974 124480
rect 673932 107001 673960 124471
rect 674116 117473 674144 162007
rect 674300 153241 674328 234586
rect 674576 222329 674604 234586
rect 674840 231328 674892 231334
rect 674840 231270 674892 231276
rect 674852 230489 674880 231270
rect 674674 230480 674730 230489
rect 674674 230415 674676 230424
rect 674728 230415 674730 230424
rect 674838 230480 674894 230489
rect 674838 230415 674894 230424
rect 674676 230386 674728 230392
rect 675128 229242 675156 234586
rect 675484 233912 675536 233918
rect 675852 233912 675904 233918
rect 675536 233860 675852 233866
rect 675484 233854 675904 233860
rect 675496 233838 675892 233854
rect 675484 232688 675536 232694
rect 675852 232688 675904 232694
rect 675536 232636 675852 232642
rect 675484 232630 675904 232636
rect 675496 232614 675892 232630
rect 675484 232552 675536 232558
rect 675852 232552 675904 232558
rect 675536 232500 675852 232506
rect 675484 232494 675904 232500
rect 675496 232478 675892 232494
rect 675036 229214 675156 229242
rect 674838 226128 674894 226137
rect 674838 226063 674894 226072
rect 674562 222320 674618 222329
rect 674562 222255 674618 222264
rect 674852 221785 674880 226063
rect 674838 221776 674894 221785
rect 674838 221711 674894 221720
rect 675036 221513 675064 229214
rect 675206 225720 675262 225729
rect 675206 225655 675262 225664
rect 675022 221504 675078 221513
rect 675022 221439 675078 221448
rect 675220 219881 675248 225655
rect 675666 225040 675722 225049
rect 675666 224975 675722 224984
rect 675206 219872 675262 219881
rect 675206 219807 675262 219816
rect 674838 219056 674894 219065
rect 674838 218991 674894 219000
rect 674470 214976 674526 214985
rect 674470 214911 674526 214920
rect 674484 197169 674512 214911
rect 674654 213752 674710 213761
rect 674654 213687 674710 213696
rect 674668 205634 674696 213687
rect 674852 212534 674880 218991
rect 675482 218784 675538 218793
rect 675680 218770 675708 224975
rect 676048 224954 676076 235175
rect 678244 233912 678296 233918
rect 678244 233854 678296 233860
rect 676770 230208 676826 230217
rect 676770 230143 676826 230152
rect 676402 228576 676458 228585
rect 676402 228511 676458 228520
rect 675538 218742 675708 218770
rect 675864 224926 676076 224954
rect 675482 218719 675538 218728
rect 675864 218634 675892 224926
rect 676034 221912 676090 221921
rect 676034 221847 676090 221856
rect 675404 218606 675892 218634
rect 675404 212537 675432 218606
rect 675574 218240 675630 218249
rect 675574 218175 675630 218184
rect 674852 212506 675156 212534
rect 674576 205606 674696 205634
rect 674576 202874 674604 205606
rect 674930 204232 674986 204241
rect 674930 204167 674986 204176
rect 674944 202881 674972 204167
rect 675128 204049 675156 212506
rect 675390 212528 675446 212537
rect 675390 212463 675446 212472
rect 675588 210474 675616 218175
rect 676048 217705 676076 221847
rect 676220 220108 676272 220114
rect 676220 220050 676272 220056
rect 676034 217696 676090 217705
rect 676034 217631 676090 217640
rect 676034 216744 676090 216753
rect 676232 216730 676260 220050
rect 676090 216702 676260 216730
rect 676034 216679 676090 216688
rect 676416 215506 676444 228511
rect 675772 215478 676444 215506
rect 675772 215393 675800 215478
rect 675758 215384 675814 215393
rect 675758 215319 675814 215328
rect 676784 215218 676812 230143
rect 677322 227080 677378 227089
rect 677322 227015 677378 227024
rect 677336 220114 677364 227015
rect 678256 223825 678284 233854
rect 683120 232688 683172 232694
rect 683120 232630 683172 232636
rect 678242 223816 678298 223825
rect 678242 223751 678298 223760
rect 683132 222737 683160 232630
rect 683304 232552 683356 232558
rect 683304 232494 683356 232500
rect 683316 223145 683344 232494
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 683302 223136 683358 223145
rect 683302 223071 683358 223080
rect 683118 222728 683174 222737
rect 683118 222663 683174 222672
rect 677324 220108 677376 220114
rect 677324 220050 677376 220056
rect 675852 215212 675904 215218
rect 675852 215154 675904 215160
rect 676772 215212 676824 215218
rect 676772 215154 676824 215160
rect 675864 214713 675892 215154
rect 675850 214704 675906 214713
rect 675850 214639 675906 214648
rect 676034 214568 676090 214577
rect 676034 214503 676090 214512
rect 676048 211449 676076 214503
rect 676034 211440 676090 211449
rect 676034 211375 676090 211384
rect 675312 210446 675616 210474
rect 675312 205337 675340 210446
rect 675482 206952 675538 206961
rect 675482 206887 675538 206896
rect 675496 205875 675524 206887
rect 675312 205309 675418 205337
rect 675404 204241 675432 204680
rect 675390 204232 675446 204241
rect 675390 204167 675446 204176
rect 675128 204021 675418 204049
rect 674576 202846 674696 202874
rect 674470 197160 674526 197169
rect 674470 197095 674526 197104
rect 674668 196058 674696 202846
rect 674930 202872 674986 202881
rect 674930 202807 674986 202816
rect 675758 202736 675814 202745
rect 675758 202671 675814 202680
rect 675772 202195 675800 202671
rect 675496 201385 675524 201620
rect 675482 201376 675538 201385
rect 675482 201311 675538 201320
rect 675128 200994 675418 201022
rect 674930 199744 674986 199753
rect 674930 199679 674986 199688
rect 674944 197350 674972 199679
rect 675128 198529 675156 200994
rect 675772 200025 675800 200328
rect 675758 200016 675814 200025
rect 675758 199951 675814 199960
rect 675114 198520 675170 198529
rect 675114 198455 675170 198464
rect 675482 198248 675538 198257
rect 675482 198183 675538 198192
rect 675496 197880 675524 198183
rect 674944 197322 675248 197350
rect 675220 197282 675248 197322
rect 675404 197282 675432 197336
rect 675220 197254 675432 197282
rect 675390 197160 675446 197169
rect 675390 197095 675446 197104
rect 675404 196656 675432 197095
rect 674668 196030 675418 196058
rect 675772 194585 675800 194820
rect 675758 194576 675814 194585
rect 675758 194511 675814 194520
rect 675758 193216 675814 193225
rect 675758 193151 675814 193160
rect 675772 192984 675800 193151
rect 675666 192808 675722 192817
rect 675666 192743 675722 192752
rect 675680 192372 675708 192743
rect 675390 191584 675446 191593
rect 675390 191519 675446 191528
rect 675404 191148 675432 191519
rect 676034 190088 676090 190097
rect 676034 190023 676090 190032
rect 675850 180296 675906 180305
rect 675850 180231 675906 180240
rect 675864 177721 675892 180231
rect 675850 177712 675906 177721
rect 675850 177647 675906 177656
rect 676048 176654 676076 190023
rect 676218 181248 676274 181257
rect 676218 181183 676274 181192
rect 676232 178945 676260 181183
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 676218 178936 676274 178945
rect 676218 178871 676274 178880
rect 675680 176626 676076 176654
rect 674470 176080 674526 176089
rect 674470 176015 674526 176024
rect 674286 153232 674342 153241
rect 674286 153167 674342 153176
rect 674484 131345 674512 176015
rect 674654 175264 674710 175273
rect 674654 175199 674710 175208
rect 674470 131336 674526 131345
rect 674470 131271 674526 131280
rect 674668 130529 674696 175199
rect 674838 174040 674894 174049
rect 674838 173975 674894 173984
rect 674852 159066 674880 173975
rect 675680 167521 675708 176626
rect 681002 173632 681058 173641
rect 681002 173567 681058 173576
rect 676034 173224 676090 173233
rect 676090 173182 676260 173210
rect 676034 173159 676090 173168
rect 676232 169674 676260 173182
rect 676586 169960 676642 169969
rect 676586 169895 676642 169904
rect 675864 169646 676260 169674
rect 675666 167512 675722 167521
rect 675666 167447 675722 167456
rect 675864 166994 675892 169646
rect 675680 166966 675892 166994
rect 675206 162344 675262 162353
rect 675206 162279 675262 162288
rect 675220 159678 675248 162279
rect 675680 161786 675708 166966
rect 676600 166433 676628 169895
rect 676586 166424 676642 166433
rect 676586 166359 676642 166368
rect 675852 164212 675904 164218
rect 675852 164154 675904 164160
rect 675864 162353 675892 164154
rect 681016 162761 681044 173567
rect 682382 171592 682438 171601
rect 682382 171527 682438 171536
rect 682396 164218 682424 171527
rect 683118 167920 683174 167929
rect 683118 167855 683174 167864
rect 682384 164212 682436 164218
rect 682384 164154 682436 164160
rect 681002 162752 681058 162761
rect 681002 162687 681058 162696
rect 675850 162344 675906 162353
rect 675850 162279 675906 162288
rect 683132 162081 683160 167855
rect 683118 162072 683174 162081
rect 683118 162007 683174 162016
rect 675312 161758 675708 161786
rect 675312 160290 675340 161758
rect 675482 161528 675538 161537
rect 675482 161463 675538 161472
rect 675496 160888 675524 161463
rect 675404 160290 675432 160344
rect 675312 160262 675432 160290
rect 675220 159650 675418 159678
rect 674852 159038 675340 159066
rect 675312 158930 675340 159038
rect 675404 158930 675432 159052
rect 675312 158902 675432 158930
rect 675772 157049 675800 157216
rect 675758 157040 675814 157049
rect 675758 156975 675814 156984
rect 675128 156629 675418 156657
rect 675128 155961 675156 156629
rect 675298 156496 675354 156505
rect 675298 156431 675354 156440
rect 675312 156006 675340 156431
rect 675312 155978 675418 156006
rect 675114 155952 675170 155961
rect 675114 155887 675170 155896
rect 675758 155816 675814 155825
rect 675758 155751 675814 155760
rect 675772 155380 675800 155751
rect 674944 152850 675418 152878
rect 674944 150385 674972 152850
rect 675114 152688 675170 152697
rect 675114 152623 675170 152632
rect 675128 152334 675156 152623
rect 675128 152306 675418 152334
rect 675772 151473 675800 151675
rect 675758 151464 675814 151473
rect 675758 151399 675814 151408
rect 675114 151328 675170 151337
rect 675114 151263 675170 151272
rect 675128 151042 675156 151263
rect 675128 151014 675418 151042
rect 674930 150376 674986 150385
rect 674930 150311 674986 150320
rect 675128 149821 675418 149849
rect 675128 147665 675156 149821
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675114 147656 675170 147665
rect 675114 147591 675170 147600
rect 675390 147656 675446 147665
rect 675390 147591 675446 147600
rect 675404 147356 675432 147591
rect 675312 146254 675432 146282
rect 675312 146146 675340 146254
rect 675128 146118 675340 146146
rect 675404 146132 675432 146254
rect 675128 144945 675156 146118
rect 675114 144936 675170 144945
rect 675114 144871 675170 144880
rect 675850 134600 675906 134609
rect 675850 134535 675906 134544
rect 675864 133958 675892 134535
rect 675852 133952 675904 133958
rect 675852 133894 675904 133900
rect 676496 133952 676548 133958
rect 676496 133894 676548 133900
rect 676508 133113 676536 133894
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 676494 133104 676550 133113
rect 676494 133039 676550 133048
rect 674654 130520 674710 130529
rect 674654 130455 674710 130464
rect 676218 130248 676274 130257
rect 676218 130183 676274 130192
rect 674930 128888 674986 128897
rect 674930 128823 674986 128832
rect 674562 128480 674618 128489
rect 674562 128415 674618 128424
rect 674378 123720 674434 123729
rect 674378 123655 674434 123664
rect 674392 123049 674420 123655
rect 674378 123040 674434 123049
rect 674378 122975 674434 122984
rect 674576 122890 674604 128415
rect 674746 123040 674802 123049
rect 674746 122975 674802 122984
rect 674392 122862 674604 122890
rect 674102 117464 674158 117473
rect 674102 117399 674158 117408
rect 673918 106992 673974 107001
rect 673918 106927 673974 106936
rect 674392 102830 674420 122862
rect 674760 122834 674788 122975
rect 674944 122834 674972 128823
rect 676232 127809 676260 130183
rect 676218 127800 676274 127809
rect 676218 127735 676274 127744
rect 676402 127800 676458 127809
rect 676402 127735 676458 127744
rect 676416 125458 676444 127735
rect 679622 126168 679678 126177
rect 679622 126103 679678 126112
rect 675852 125452 675904 125458
rect 675852 125394 675904 125400
rect 676404 125452 676456 125458
rect 676404 125394 676456 125400
rect 675864 122834 675892 125394
rect 676494 123312 676550 123321
rect 676494 123247 676550 123256
rect 676508 122913 676536 123247
rect 676494 122904 676550 122913
rect 676494 122839 676550 122848
rect 674668 122806 674788 122834
rect 674852 122806 674972 122834
rect 675772 122806 675892 122834
rect 674668 105822 674696 122806
rect 674852 113846 674880 122806
rect 675022 122496 675078 122505
rect 675022 122431 675078 122440
rect 675036 121689 675064 122431
rect 675022 121680 675078 121689
rect 675022 121615 675078 121624
rect 675206 117056 675262 117065
rect 675206 116991 675262 117000
rect 675220 114493 675248 116991
rect 675772 116498 675800 122806
rect 679636 118658 679664 126103
rect 682382 125352 682438 125361
rect 682382 125287 682438 125296
rect 675944 118652 675996 118658
rect 675944 118594 675996 118600
rect 679624 118652 679676 118658
rect 679624 118594 679676 118600
rect 675956 117065 675984 118594
rect 682396 117337 682424 125287
rect 682382 117328 682438 117337
rect 682382 117263 682438 117272
rect 675942 117056 675998 117065
rect 675942 116991 675998 117000
rect 675312 116470 675800 116498
rect 675312 115138 675340 116470
rect 675482 115832 675538 115841
rect 675482 115767 675538 115776
rect 675496 115668 675524 115767
rect 675312 115110 675418 115138
rect 675220 114465 675418 114493
rect 674852 113818 675418 113846
rect 675758 112432 675814 112441
rect 675758 112367 675814 112376
rect 675772 111996 675800 112367
rect 675758 111752 675814 111761
rect 675758 111687 675814 111696
rect 675772 111452 675800 111687
rect 675758 111344 675814 111353
rect 675758 111279 675814 111288
rect 675772 110772 675800 111279
rect 675758 110392 675814 110401
rect 675758 110327 675814 110336
rect 675772 110160 675800 110327
rect 675758 108216 675814 108225
rect 675758 108151 675814 108160
rect 675772 107644 675800 108151
rect 675312 107222 675432 107250
rect 675312 107114 675340 107222
rect 675128 107086 675340 107114
rect 675404 107100 675432 107222
rect 675128 106321 675156 107086
rect 675390 106992 675446 107001
rect 675390 106927 675446 106936
rect 675404 106488 675432 106927
rect 675114 106312 675170 106321
rect 675114 106247 675170 106256
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 674668 105794 675340 105822
rect 675404 105808 675432 105862
rect 675114 104680 675170 104689
rect 675170 104638 675340 104666
rect 675114 104615 675170 104624
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 674392 102802 675340 102830
rect 675312 102762 675340 102802
rect 675404 102762 675432 102816
rect 675312 102734 675432 102762
rect 675390 102640 675446 102649
rect 675390 102575 675446 102584
rect 675404 102136 675432 102575
rect 673366 101008 673422 101017
rect 673366 100943 673422 100952
rect 675114 101008 675170 101017
rect 675170 100966 675340 100994
rect 675114 100943 675170 100952
rect 675312 100858 675340 100966
rect 675404 100858 675432 100980
rect 675312 100830 675432 100858
rect 595272 100014 595608 100042
rect 596344 100014 596496 100042
rect 595272 99142 595300 100014
rect 595260 99136 595312 99142
rect 595260 99078 595312 99084
rect 595272 93854 595300 99078
rect 596180 96960 596232 96966
rect 596180 96902 596232 96908
rect 595272 93826 595484 93854
rect 595456 80714 595484 93826
rect 595444 80708 595496 80714
rect 595444 80650 595496 80656
rect 596192 54398 596220 96902
rect 596468 55214 596496 100014
rect 596744 100014 597080 100042
rect 596744 96966 596772 100014
rect 597802 99770 597830 100028
rect 598216 100014 598552 100042
rect 598952 100014 599288 100042
rect 599504 100014 600024 100042
rect 600516 100014 600760 100042
rect 601160 100014 601496 100042
rect 601896 100014 602232 100042
rect 602632 100014 602968 100042
rect 603092 100014 603704 100042
rect 597802 99742 597876 99770
rect 596732 96960 596784 96966
rect 596732 96902 596784 96908
rect 597652 96960 597704 96966
rect 597652 96902 597704 96908
rect 596456 55208 596508 55214
rect 596456 55150 596508 55156
rect 597664 54942 597692 96902
rect 597848 55078 597876 99742
rect 598216 96966 598244 100014
rect 598204 96960 598256 96966
rect 598204 96902 598256 96908
rect 597836 55072 597888 55078
rect 597836 55014 597888 55020
rect 597652 54936 597704 54942
rect 597652 54878 597704 54884
rect 598952 54806 598980 100014
rect 599504 84194 599532 100014
rect 600320 96960 600372 96966
rect 600320 96902 600372 96908
rect 599136 84166 599532 84194
rect 599136 56030 599164 84166
rect 600332 57254 600360 96902
rect 600320 57248 600372 57254
rect 600320 57190 600372 57196
rect 599124 56024 599176 56030
rect 599124 55966 599176 55972
rect 600516 55894 600544 100014
rect 601160 96966 601188 100014
rect 601148 96960 601200 96966
rect 601148 96902 601200 96908
rect 601700 96960 601752 96966
rect 601700 96902 601752 96908
rect 601712 58682 601740 96902
rect 601896 72486 601924 100014
rect 602632 96966 602660 100014
rect 602620 96960 602672 96966
rect 602620 96902 602672 96908
rect 601884 72480 601936 72486
rect 601884 72422 601936 72428
rect 603092 60042 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 606984 100042
rect 607384 100014 607720 100042
rect 608120 100014 608548 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 604426 99742 604500 99770
rect 604472 68338 604500 99742
rect 605484 97306 605512 100014
rect 605472 97300 605524 97306
rect 605472 97242 605524 97248
rect 606220 96966 606248 100014
rect 606208 96960 606260 96966
rect 606208 96902 606260 96908
rect 606956 92886 606984 100014
rect 607128 96960 607180 96966
rect 607128 96902 607180 96908
rect 606944 92880 606996 92886
rect 606944 92822 606996 92828
rect 607140 75206 607168 96902
rect 607692 95946 607720 100014
rect 607680 95940 607732 95946
rect 607680 95882 607732 95888
rect 608520 84182 608548 100014
rect 609164 94518 609192 100014
rect 609152 94512 609204 94518
rect 609152 94454 609204 94460
rect 609900 85542 609928 100014
rect 610636 96762 610664 100014
rect 611050 99770 611078 100028
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 613272 100014 613608 100042
rect 611050 99742 611124 99770
rect 610624 96756 610676 96762
rect 610624 96698 610676 96704
rect 611096 96082 611124 99742
rect 611912 97300 611964 97306
rect 611912 97242 611964 97248
rect 611268 96756 611320 96762
rect 611268 96698 611320 96704
rect 611084 96076 611136 96082
rect 611084 96018 611136 96024
rect 611280 93158 611308 96698
rect 611924 93854 611952 97242
rect 612108 96898 612136 100014
rect 612660 97442 612688 100014
rect 612648 97436 612700 97442
rect 612648 97378 612700 97384
rect 613580 96966 613608 100014
rect 613764 100014 614008 100042
rect 614744 100014 615264 100042
rect 615480 100014 615816 100042
rect 616216 100014 616552 100042
rect 616952 100014 617288 100042
rect 617688 100014 617932 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620232 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 613568 96960 613620 96966
rect 613568 96902 613620 96908
rect 612096 96892 612148 96898
rect 612096 96834 612148 96840
rect 612648 96892 612700 96898
rect 612648 96834 612700 96840
rect 611924 93826 612044 93854
rect 611268 93152 611320 93158
rect 611268 93094 611320 93100
rect 610072 92880 610124 92886
rect 610072 92822 610124 92828
rect 610084 88330 610112 92822
rect 610072 88324 610124 88330
rect 610072 88266 610124 88272
rect 609888 85536 609940 85542
rect 609888 85478 609940 85484
rect 608508 84176 608560 84182
rect 608508 84118 608560 84124
rect 612016 76566 612044 93826
rect 612660 80850 612688 96834
rect 612648 80844 612700 80850
rect 612648 80786 612700 80792
rect 613764 79490 613792 100014
rect 613936 96960 613988 96966
rect 613936 96902 613988 96908
rect 613752 79484 613804 79490
rect 613752 79426 613804 79432
rect 613948 79354 613976 96902
rect 615236 93854 615264 100014
rect 615788 96966 615816 100014
rect 615776 96960 615828 96966
rect 615776 96902 615828 96908
rect 616524 95062 616552 100014
rect 616788 96960 616840 96966
rect 616788 96902 616840 96908
rect 616512 95056 616564 95062
rect 616512 94998 616564 95004
rect 615236 93826 615448 93854
rect 613936 79348 613988 79354
rect 613936 79290 613988 79296
rect 612004 76560 612056 76566
rect 612004 76502 612056 76508
rect 615420 75342 615448 93826
rect 616800 76702 616828 96902
rect 617260 96762 617288 100014
rect 617248 96756 617300 96762
rect 617248 96698 617300 96704
rect 617904 92478 617932 100014
rect 618732 97850 618760 100014
rect 618720 97844 618772 97850
rect 618720 97786 618772 97792
rect 618904 97436 618956 97442
rect 618904 97378 618956 97384
rect 618076 96756 618128 96762
rect 618076 96698 618128 96704
rect 617892 92472 617944 92478
rect 617892 92414 617944 92420
rect 618088 91050 618116 96698
rect 618076 91044 618128 91050
rect 618076 90986 618128 90992
rect 616788 76696 616840 76702
rect 616788 76638 616840 76644
rect 618916 75478 618944 97378
rect 619560 93838 619588 100014
rect 620204 97986 620232 100014
rect 620192 97980 620244 97986
rect 620192 97922 620244 97928
rect 620940 95198 620968 100014
rect 621676 97578 621704 100014
rect 622320 99346 622348 100014
rect 622308 99340 622360 99346
rect 622308 99282 622360 99288
rect 621664 97572 621716 97578
rect 621664 97514 621716 97520
rect 623148 97442 623176 100014
rect 623700 99210 623728 100014
rect 623688 99204 623740 99210
rect 623688 99146 623740 99152
rect 623136 97436 623188 97442
rect 623136 97378 623188 97384
rect 624620 97034 624648 100014
rect 625034 99770 625062 100028
rect 625784 100014 626120 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628328 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 632008 100042
rect 632408 100014 632744 100042
rect 633144 100014 633296 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635596 100042
rect 625034 99742 625108 99770
rect 625080 99074 625108 99742
rect 625068 99068 625120 99074
rect 625068 99010 625120 99016
rect 625804 97844 625856 97850
rect 625804 97786 625856 97792
rect 624608 97028 624660 97034
rect 624608 96970 624660 96976
rect 622308 96076 622360 96082
rect 622308 96018 622360 96024
rect 620928 95192 620980 95198
rect 620928 95134 620980 95140
rect 620284 94512 620336 94518
rect 620284 94454 620336 94460
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 619272 93152 619324 93158
rect 619272 93094 619324 93100
rect 619284 86358 619312 93094
rect 619272 86352 619324 86358
rect 619272 86294 619324 86300
rect 620296 85406 620324 94454
rect 622320 88194 622348 96018
rect 624976 95940 625028 95946
rect 624976 95882 625028 95888
rect 622952 95056 623004 95062
rect 622952 94998 623004 95004
rect 622964 89690 622992 94998
rect 622952 89684 623004 89690
rect 622952 89626 623004 89632
rect 624988 88641 625016 95882
rect 625816 92041 625844 97786
rect 626092 97170 626120 100014
rect 626264 97980 626316 97986
rect 626264 97922 626316 97928
rect 626080 97164 626132 97170
rect 626080 97106 626132 97112
rect 626276 93673 626304 97922
rect 626828 97306 626856 100014
rect 627564 97850 627592 100014
rect 628300 98938 628328 100014
rect 628288 98932 628340 98938
rect 628288 98874 628340 98880
rect 629036 98802 629064 100014
rect 629024 98796 629076 98802
rect 629024 98738 629076 98744
rect 629772 97986 629800 100014
rect 630508 98666 630536 100014
rect 630772 99340 630824 99346
rect 630772 99282 630824 99288
rect 630496 98660 630548 98666
rect 630496 98602 630548 98608
rect 629760 97980 629812 97986
rect 629760 97922 629812 97928
rect 627552 97844 627604 97850
rect 627552 97786 627604 97792
rect 629300 97572 629352 97578
rect 629300 97514 629352 97520
rect 626816 97300 626868 97306
rect 626816 97242 626868 97248
rect 629312 95826 629340 97514
rect 630784 95826 630812 99282
rect 631244 96354 631272 100014
rect 631980 97714 632008 100014
rect 632716 97850 632744 100014
rect 632704 97844 632756 97850
rect 632704 97786 632756 97792
rect 631968 97708 632020 97714
rect 631968 97650 632020 97656
rect 633268 97442 633296 100014
rect 633440 99204 633492 99210
rect 633440 99146 633492 99152
rect 632060 97436 632112 97442
rect 632060 97378 632112 97384
rect 633256 97436 633308 97442
rect 633256 97378 633308 97384
rect 631232 96348 631284 96354
rect 631232 96290 631284 96296
rect 629280 95798 629340 95826
rect 630752 95798 630812 95826
rect 632072 95826 632100 97378
rect 633452 95826 633480 99146
rect 634188 97578 634216 100014
rect 634176 97572 634228 97578
rect 634176 97514 634228 97520
rect 634740 96898 634768 100014
rect 635568 97034 635596 100014
rect 635752 100014 636088 100042
rect 636824 100014 637068 100042
rect 635004 97028 635056 97034
rect 635004 96970 635056 96976
rect 635556 97028 635608 97034
rect 635556 96970 635608 96976
rect 634728 96892 634780 96898
rect 634728 96834 634780 96840
rect 635016 95826 635044 96970
rect 632072 95798 632224 95826
rect 633452 95798 633696 95826
rect 635016 95798 635168 95826
rect 635752 95441 635780 100014
rect 636292 99068 636344 99074
rect 636292 99010 636344 99016
rect 636304 95826 636332 99010
rect 637040 96937 637068 100014
rect 637546 99770 637574 100028
rect 638296 100014 638632 100042
rect 637546 99742 637620 99770
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 96218 637620 99742
rect 637764 97164 637816 97170
rect 637764 97106 637816 97112
rect 637580 96212 637632 96218
rect 637580 96154 637632 96160
rect 637776 95826 637804 97106
rect 636304 95798 636640 95826
rect 637776 95798 638112 95826
rect 638604 95742 638632 100014
rect 639018 99770 639046 100028
rect 639768 100014 640104 100042
rect 639018 99742 639092 99770
rect 639064 96490 639092 99742
rect 639236 97300 639288 97306
rect 639236 97242 639288 97248
rect 639052 96484 639104 96490
rect 639052 96426 639104 96432
rect 639248 95826 639276 97242
rect 639248 95798 639584 95826
rect 638592 95736 638644 95742
rect 638592 95678 638644 95684
rect 640076 95606 640104 100014
rect 640490 99770 640518 100028
rect 641240 100014 641576 100042
rect 640490 99742 640564 99770
rect 640536 96626 640564 99742
rect 640708 98048 640760 98054
rect 640708 97990 640760 97996
rect 640524 96620 640576 96626
rect 640524 96562 640576 96568
rect 640720 95826 640748 97990
rect 640720 95798 641056 95826
rect 640064 95600 640116 95606
rect 640064 95542 640116 95548
rect 641548 95470 641576 100014
rect 641962 99770 641990 100028
rect 642712 100014 643048 100042
rect 641962 99742 642036 99770
rect 642008 96529 642036 99742
rect 642180 98932 642232 98938
rect 642180 98874 642232 98880
rect 641994 96520 642050 96529
rect 641994 96455 642050 96464
rect 642192 95826 642220 98874
rect 643020 97306 643048 100014
rect 643434 99770 643462 100028
rect 644184 100014 644336 100042
rect 643434 99742 643508 99770
rect 643008 97300 643060 97306
rect 643008 97242 643060 97248
rect 643480 95878 643508 99742
rect 643652 98796 643704 98802
rect 643652 98738 643704 98744
rect 643468 95872 643520 95878
rect 642192 95798 642528 95826
rect 643468 95814 643520 95820
rect 643664 95826 643692 98738
rect 644308 97170 644336 100014
rect 644906 99770 644934 100028
rect 645656 100014 645808 100042
rect 644906 99742 644980 99770
rect 644296 97164 644348 97170
rect 644296 97106 644348 97112
rect 644952 96014 644980 99742
rect 645308 98252 645360 98258
rect 645308 98194 645360 98200
rect 645124 96484 645176 96490
rect 645124 96426 645176 96432
rect 644940 96008 644992 96014
rect 644940 95950 644992 95956
rect 643664 95798 644000 95826
rect 645136 95470 645164 96426
rect 645320 95826 645348 98194
rect 645780 96626 645808 100014
rect 646378 99770 646406 100028
rect 647114 99770 647142 100028
rect 647864 100014 648476 100042
rect 648600 100014 648936 100042
rect 649336 100014 649764 100042
rect 650072 100014 650408 100042
rect 650808 100014 651328 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 655224 100014 655468 100042
rect 646378 99742 646452 99770
rect 647114 99742 647188 99770
rect 645768 96620 645820 96626
rect 645768 96562 645820 96568
rect 646424 96490 646452 99742
rect 647160 98802 647188 99742
rect 647148 98796 647200 98802
rect 647148 98738 647200 98744
rect 646596 98660 646648 98666
rect 646596 98602 646648 98608
rect 646412 96484 646464 96490
rect 646412 96426 646464 96432
rect 646608 95826 646636 98602
rect 648252 97844 648304 97850
rect 648252 97786 648304 97792
rect 647516 97708 647568 97714
rect 647516 97650 647568 97656
rect 647148 96348 647200 96354
rect 647148 96290 647200 96296
rect 645320 95798 645472 95826
rect 646608 95798 646944 95826
rect 641536 95464 641588 95470
rect 635738 95432 635794 95441
rect 641536 95406 641588 95412
rect 645124 95464 645176 95470
rect 645124 95406 645176 95412
rect 635738 95367 635794 95376
rect 626448 95192 626500 95198
rect 626448 95134 626500 95140
rect 626460 94489 626488 95134
rect 647160 95033 647188 96290
rect 647332 95736 647384 95742
rect 647332 95678 647384 95684
rect 647146 95024 647202 95033
rect 647146 94959 647202 94968
rect 626446 94480 626502 94489
rect 626446 94415 626502 94424
rect 626448 93832 626500 93838
rect 626448 93774 626500 93780
rect 626262 93664 626318 93673
rect 626262 93599 626318 93608
rect 626460 92857 626488 93774
rect 626446 92848 626502 92857
rect 626446 92783 626502 92792
rect 626448 92472 626500 92478
rect 626448 92414 626500 92420
rect 625802 92032 625858 92041
rect 625802 91967 625858 91976
rect 626460 91225 626488 92414
rect 647344 92410 647372 95678
rect 647528 92449 647556 97650
rect 647700 97028 647752 97034
rect 647700 96970 647752 96976
rect 647712 95130 647740 96970
rect 647884 96756 647936 96762
rect 647884 96698 647936 96704
rect 647896 95742 647924 96698
rect 647884 95736 647936 95742
rect 647884 95678 647936 95684
rect 647884 95600 647936 95606
rect 647884 95542 647936 95548
rect 647700 95124 647752 95130
rect 647700 95066 647752 95072
rect 647514 92440 647570 92449
rect 647332 92404 647384 92410
rect 647514 92375 647570 92384
rect 647332 92346 647384 92352
rect 626446 91216 626502 91225
rect 626446 91151 626502 91160
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90409 626488 90986
rect 626446 90400 626502 90409
rect 626446 90335 626502 90344
rect 626448 89616 626500 89622
rect 626446 89584 626448 89593
rect 626500 89584 626502 89593
rect 626446 89519 626502 89528
rect 624974 88632 625030 88641
rect 624974 88567 625030 88576
rect 626448 88324 626500 88330
rect 626448 88266 626500 88272
rect 622308 88188 622360 88194
rect 622308 88130 622360 88136
rect 626264 88188 626316 88194
rect 626264 88130 626316 88136
rect 626276 87145 626304 88130
rect 626460 87961 626488 88266
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 626262 87136 626318 87145
rect 626262 87071 626318 87080
rect 626448 86352 626500 86358
rect 626446 86320 626448 86329
rect 626500 86320 626502 86329
rect 626446 86255 626502 86264
rect 647896 86222 647924 95542
rect 648264 89593 648292 97786
rect 648250 89584 648306 89593
rect 648250 89519 648306 89528
rect 648448 87038 648476 100014
rect 648620 97436 648672 97442
rect 648620 97378 648672 97384
rect 648632 92546 648660 97378
rect 648908 96354 648936 100014
rect 648896 96348 648948 96354
rect 648896 96290 648948 96296
rect 649540 96008 649592 96014
rect 649540 95950 649592 95956
rect 649264 95872 649316 95878
rect 649264 95814 649316 95820
rect 648804 95124 648856 95130
rect 648804 95066 648856 95072
rect 648620 92540 648672 92546
rect 648620 92482 648672 92488
rect 648436 87032 648488 87038
rect 648436 86974 648488 86980
rect 647884 86216 647936 86222
rect 647884 86158 647936 86164
rect 626448 85536 626500 85542
rect 626446 85504 626448 85513
rect 626500 85504 626502 85513
rect 626446 85439 626502 85448
rect 620284 85400 620336 85406
rect 620284 85342 620336 85348
rect 625252 85400 625304 85406
rect 625252 85342 625304 85348
rect 625264 84697 625292 85342
rect 625250 84688 625306 84697
rect 625250 84623 625306 84632
rect 625804 84176 625856 84182
rect 625804 84118 625856 84124
rect 625816 83881 625844 84118
rect 625802 83872 625858 83881
rect 625802 83807 625858 83816
rect 628746 83328 628802 83337
rect 628746 83263 628802 83272
rect 628760 80986 628788 83263
rect 629206 81696 629262 81705
rect 629206 81631 629262 81640
rect 628748 80980 628800 80986
rect 628748 80922 628800 80928
rect 629220 80034 629248 81631
rect 632808 80974 633144 81002
rect 642456 80980 642508 80986
rect 629208 80028 629260 80034
rect 629208 79970 629260 79976
rect 631048 77988 631100 77994
rect 631048 77930 631100 77936
rect 628472 77784 628524 77790
rect 628472 77726 628524 77732
rect 624422 77344 624478 77353
rect 624422 77279 624478 77288
rect 625804 77308 625856 77314
rect 618904 75472 618956 75478
rect 618904 75414 618956 75420
rect 615408 75336 615460 75342
rect 615408 75278 615460 75284
rect 607128 75200 607180 75206
rect 607128 75142 607180 75148
rect 604460 68332 604512 68338
rect 604460 68274 604512 68280
rect 603080 60036 603132 60042
rect 603080 59978 603132 59984
rect 601700 58676 601752 58682
rect 601700 58618 601752 58624
rect 600504 55888 600556 55894
rect 600504 55830 600556 55836
rect 598940 54800 598992 54806
rect 598940 54742 598992 54748
rect 624436 54670 624464 77279
rect 625804 77250 625856 77256
rect 624424 54664 624476 54670
rect 624424 54606 624476 54612
rect 625816 54534 625844 77250
rect 628484 75290 628512 77726
rect 631060 77314 631088 77930
rect 632808 77790 632836 80974
rect 643080 80974 643140 81002
rect 642456 80922 642508 80928
rect 636752 80708 636804 80714
rect 636752 80650 636804 80656
rect 633440 80028 633492 80034
rect 633440 79970 633492 79976
rect 633452 78130 633480 79970
rect 633898 78568 633954 78577
rect 633898 78503 633954 78512
rect 633440 78124 633492 78130
rect 633440 78066 633492 78072
rect 632796 77784 632848 77790
rect 632796 77726 632848 77732
rect 633912 77353 633940 78503
rect 633898 77344 633954 77353
rect 631048 77308 631100 77314
rect 633898 77279 633954 77288
rect 631048 77250 631100 77256
rect 631060 75290 631088 77250
rect 633912 75290 633940 77279
rect 636764 75290 636792 80650
rect 639602 78160 639658 78169
rect 639602 78095 639658 78104
rect 639616 75290 639644 78095
rect 642468 75290 642496 80922
rect 643112 77994 643140 80974
rect 647424 80844 647476 80850
rect 647424 80786 647476 80792
rect 646044 79484 646096 79490
rect 646044 79426 646096 79432
rect 645308 78124 645360 78130
rect 645308 78066 645360 78072
rect 643100 77988 643152 77994
rect 643100 77930 643152 77936
rect 645320 75290 645348 78066
rect 628176 75262 628512 75290
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 636732 75262 636792 75290
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 646056 70530 646084 79426
rect 646504 79348 646556 79354
rect 646504 79290 646556 79296
rect 646228 75200 646280 75206
rect 646228 75142 646280 75148
rect 646240 74225 646268 75142
rect 646226 74216 646282 74225
rect 646226 74151 646282 74160
rect 646056 70502 646268 70530
rect 646240 67153 646268 70502
rect 646226 67144 646282 67153
rect 646226 67079 646282 67088
rect 646516 64433 646544 79290
rect 646688 76696 646740 76702
rect 646688 76638 646740 76644
rect 646700 71777 646728 76638
rect 646872 75336 646924 75342
rect 646872 75278 646924 75284
rect 646884 74534 646912 75278
rect 646884 74506 647280 74534
rect 646686 71768 646742 71777
rect 646686 71703 646742 71712
rect 647252 68921 647280 74506
rect 647238 68912 647294 68921
rect 647238 68847 647294 68856
rect 647436 64874 647464 80786
rect 648620 75472 648672 75478
rect 648620 75414 648672 75420
rect 647252 64846 647464 64874
rect 646502 64424 646558 64433
rect 646502 64359 646558 64368
rect 647252 59265 647280 64846
rect 648632 62121 648660 75414
rect 648618 62112 648674 62121
rect 648618 62047 648674 62056
rect 647238 59256 647294 59265
rect 647238 59191 647294 59200
rect 648816 57361 648844 95066
rect 649276 86630 649304 95814
rect 649552 93022 649580 95950
rect 649540 93016 649592 93022
rect 649540 92958 649592 92964
rect 649736 88806 649764 100014
rect 650380 97714 650408 100014
rect 650368 97708 650420 97714
rect 650368 97650 650420 97656
rect 650552 97572 650604 97578
rect 650552 97514 650604 97520
rect 650368 96892 650420 96898
rect 650368 96834 650420 96840
rect 649908 96076 649960 96082
rect 649908 96018 649960 96024
rect 649920 95334 649948 96018
rect 649908 95328 649960 95334
rect 649908 95270 649960 95276
rect 650000 92540 650052 92546
rect 650000 92482 650052 92488
rect 649724 88800 649776 88806
rect 649724 88742 649776 88748
rect 650012 87145 650040 92482
rect 649998 87136 650054 87145
rect 649998 87071 650054 87080
rect 649264 86624 649316 86630
rect 649264 86566 649316 86572
rect 650380 82249 650408 96834
rect 650564 84697 650592 97514
rect 651300 93566 651328 100014
rect 651852 97442 651880 100014
rect 651840 97436 651892 97442
rect 651840 97378 651892 97384
rect 652588 96490 652616 100014
rect 652024 96484 652076 96490
rect 652024 96426 652076 96432
rect 652576 96484 652628 96490
rect 652576 96426 652628 96432
rect 651840 95464 651892 95470
rect 651840 95406 651892 95412
rect 651288 93560 651340 93566
rect 651288 93502 651340 93508
rect 651852 90710 651880 95406
rect 651840 90704 651892 90710
rect 651840 90646 651892 90652
rect 652036 86494 652064 96426
rect 653324 95674 653352 100014
rect 653968 96898 653996 100014
rect 654796 96898 654824 100014
rect 655440 97850 655468 100014
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655428 97844 655480 97850
rect 655428 97786 655480 97792
rect 653956 96892 654008 96898
rect 653956 96834 654008 96840
rect 654600 96892 654652 96898
rect 654600 96834 654652 96840
rect 654784 96892 654836 96898
rect 654784 96834 654836 96840
rect 655428 96892 655480 96898
rect 655428 96834 655480 96840
rect 653312 95668 653364 95674
rect 653312 95610 653364 95616
rect 654612 94217 654640 96834
rect 654598 94208 654654 94217
rect 654598 94143 654654 94152
rect 655440 93854 655468 96834
rect 655256 93826 655468 93854
rect 654324 92404 654376 92410
rect 654324 92346 654376 92352
rect 654336 91497 654364 92346
rect 654322 91488 654378 91497
rect 654322 91423 654378 91432
rect 655256 88330 655284 93826
rect 655428 93560 655480 93566
rect 655428 93502 655480 93508
rect 655440 93401 655468 93502
rect 655426 93392 655482 93401
rect 655426 93327 655482 93336
rect 655428 90704 655480 90710
rect 655426 90672 655428 90681
rect 655480 90672 655482 90681
rect 655426 90607 655482 90616
rect 655808 89865 655836 100014
rect 656624 97572 656676 97578
rect 656624 97514 656676 97520
rect 656636 97306 656664 97514
rect 656820 97306 656848 100014
rect 656624 97300 656676 97306
rect 656624 97242 656676 97248
rect 656808 97300 656860 97306
rect 656808 97242 656860 97248
rect 656716 96960 656768 96966
rect 656716 96902 656768 96908
rect 656348 96620 656400 96626
rect 656348 96562 656400 96568
rect 656164 93016 656216 93022
rect 656164 92958 656216 92964
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 655244 88324 655296 88330
rect 655244 88266 655296 88272
rect 656176 86766 656204 92958
rect 656360 88670 656388 96562
rect 656348 88664 656400 88670
rect 656348 88606 656400 88612
rect 656728 86902 656756 96902
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 658108 99742 658182 99770
rect 658108 96830 658136 99742
rect 658280 97708 658332 97714
rect 658280 97650 658332 97656
rect 658096 96824 658148 96830
rect 658096 96766 658148 96772
rect 658292 95132 658320 97650
rect 659212 97578 659240 100014
rect 659948 97986 659976 100014
rect 660132 100014 660376 100042
rect 659936 97980 659988 97986
rect 659936 97922 659988 97928
rect 659844 97708 659896 97714
rect 659844 97650 659896 97656
rect 659200 97572 659252 97578
rect 659200 97514 659252 97520
rect 659568 97436 659620 97442
rect 659568 97378 659620 97384
rect 658832 97164 658884 97170
rect 658832 97106 658884 97112
rect 658844 95132 658872 97106
rect 659580 95132 659608 97378
rect 659856 95146 659884 97650
rect 660132 96966 660160 100014
rect 661960 98796 662012 98802
rect 661960 98738 662012 98744
rect 661408 97300 661460 97306
rect 661408 97242 661460 97248
rect 660120 96960 660172 96966
rect 660120 96902 660172 96908
rect 660672 96212 660724 96218
rect 660672 96154 660724 96160
rect 659856 95118 660146 95146
rect 660684 95132 660712 96154
rect 661420 95132 661448 97242
rect 661972 95132 662000 98738
rect 665548 97980 665600 97986
rect 665548 97922 665600 97928
rect 662512 97844 662564 97850
rect 662512 97786 662564 97792
rect 662524 95132 662552 97786
rect 664168 97572 664220 97578
rect 664168 97514 664220 97520
rect 663064 96824 663116 96830
rect 663064 96766 663116 96772
rect 663076 95132 663104 96766
rect 663800 96076 663852 96082
rect 663800 96018 663852 96024
rect 663812 93129 663840 96018
rect 663984 95668 664036 95674
rect 663984 95610 664036 95616
rect 663798 93120 663854 93129
rect 663798 93055 663854 93064
rect 663996 89049 664024 95610
rect 663982 89040 664038 89049
rect 663982 88975 664038 88984
rect 664180 88806 664208 97514
rect 665364 96484 665416 96490
rect 665364 96426 665416 96432
rect 664352 96348 664404 96354
rect 664352 96290 664404 96296
rect 664364 89865 664392 96290
rect 665180 95940 665232 95946
rect 665180 95882 665232 95888
rect 665192 91769 665220 95882
rect 665178 91760 665234 91769
rect 665178 91695 665234 91704
rect 665376 90681 665404 96426
rect 665560 93401 665588 97922
rect 665546 93392 665602 93401
rect 665546 93327 665602 93336
rect 665362 90672 665418 90681
rect 665362 90607 665418 90616
rect 664350 89856 664406 89865
rect 664350 89791 664406 89800
rect 658556 88800 658608 88806
rect 662328 88800 662380 88806
rect 658608 88748 658858 88754
rect 658556 88742 658858 88748
rect 658568 88726 658858 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 664168 88800 664220 88806
rect 664168 88742 664220 88748
rect 661986 88726 662368 88742
rect 657452 88664 657504 88670
rect 657504 88612 657754 88618
rect 657452 88606 657754 88612
rect 657464 88590 657754 88606
rect 658306 88330 658504 88346
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 658464 88266 658516 88272
rect 656716 86896 656768 86902
rect 656716 86838 656768 86844
rect 656164 86760 656216 86766
rect 656164 86702 656216 86708
rect 657188 86494 657216 88196
rect 659580 86902 659608 88196
rect 659568 86896 659620 86902
rect 659568 86838 659620 86844
rect 652024 86488 652076 86494
rect 652024 86430 652076 86436
rect 657176 86488 657228 86494
rect 657176 86430 657228 86436
rect 660132 86222 660160 88196
rect 660684 86766 660712 88196
rect 660672 86760 660724 86766
rect 660672 86702 660724 86708
rect 661420 86630 661448 88196
rect 662524 87038 662552 88196
rect 662512 87032 662564 87038
rect 662512 86974 662564 86980
rect 661408 86624 661460 86630
rect 661408 86566 661460 86572
rect 660120 86216 660172 86222
rect 660120 86158 660172 86164
rect 650550 84688 650606 84697
rect 650550 84623 650606 84632
rect 650366 82240 650422 82249
rect 650366 82175 650422 82184
rect 662420 76560 662472 76566
rect 662420 76502 662472 76508
rect 648802 57352 648858 57361
rect 648802 57287 648858 57296
rect 625804 54528 625856 54534
rect 625804 54470 625856 54476
rect 596180 54392 596232 54398
rect 596180 54334 596232 54340
rect 592684 51740 592736 51746
rect 592684 51682 592736 51688
rect 661590 48510 661646 48519
rect 661590 48445 661646 48454
rect 553674 48104 553730 48113
rect 553674 48039 553730 48048
rect 552018 47832 552074 47841
rect 552018 47767 552074 47776
rect 547878 47560 547934 47569
rect 547878 47495 547934 47504
rect 545670 47288 545726 47297
rect 545670 47223 545726 47232
rect 465262 46744 465318 46753
rect 465262 46679 465318 46688
rect 661604 45554 661632 48445
rect 662432 47433 662460 76502
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 661420 45526 661632 45554
rect 464342 44160 464398 44169
rect 464342 44095 464398 44104
rect 471058 43480 471114 43489
rect 471058 43415 471114 43424
rect 465814 43208 465870 43217
rect 465814 43143 465870 43152
rect 464160 42764 464212 42770
rect 464160 42706 464212 42712
rect 463056 42492 463108 42498
rect 463988 42486 464050 42514
rect 463056 42434 463108 42440
rect 461950 42256 462006 42265
rect 464022 42228 464050 42486
rect 465828 42364 465856 43143
rect 461950 42191 462006 42200
rect 471072 42106 471100 43415
rect 518806 42800 518862 42809
rect 518806 42735 518862 42744
rect 518820 42228 518848 42735
rect 661420 42187 661448 45526
rect 661408 42181 661460 42187
rect 515402 42120 515458 42129
rect 459940 42078 460368 42106
rect 471072 42078 471408 42106
rect 515154 42078 515402 42106
rect 520922 42120 520978 42129
rect 520674 42078 520922 42106
rect 515402 42055 515458 42064
rect 522026 42120 522082 42129
rect 521870 42078 522026 42106
rect 520922 42055 520978 42064
rect 526442 42120 526498 42129
rect 526194 42078 526442 42106
rect 522026 42055 522082 42064
rect 529570 42120 529626 42129
rect 661408 42123 661460 42129
rect 529322 42078 529570 42106
rect 526442 42055 526498 42064
rect 529570 42055 529626 42064
rect 404452 41472 404504 41478
rect 404452 41414 404504 41420
rect 420736 41472 420788 41478
rect 420736 41414 420788 41420
rect 426900 41472 426952 41478
rect 426900 41414 426952 41420
rect 459192 41472 459244 41478
rect 459192 41414 459244 41420
rect 141698 40352 141754 40361
rect 141698 40287 141754 40296
rect 141712 39984 141740 40287
<< via2 >>
rect 185030 1002088 185086 1002144
rect 82174 1001952 82230 1002008
rect 133694 1001972 133750 1002008
rect 133694 1001952 133696 1001972
rect 133696 1001952 133748 1001972
rect 133748 1001952 133750 1001972
rect 81346 983456 81402 983512
rect 483018 1001952 483074 1002008
rect 534998 1001952 535054 1002008
rect 232962 997328 233018 997384
rect 240138 997192 240194 997248
rect 235906 990936 235962 990992
rect 238666 984000 238722 984056
rect 285402 997328 285458 997384
rect 292578 997328 292634 997384
rect 286966 987944 287022 988000
rect 235906 983728 235962 983784
rect 240138 983728 240194 983784
rect 286966 983728 287022 983784
rect 184938 983456 184994 983512
rect 132498 982504 132554 982560
rect 387522 997328 387578 997384
rect 389178 990936 389234 990992
rect 404358 997328 404414 997384
rect 292578 983728 292634 983784
rect 391938 983456 391994 983512
rect 394422 983492 394424 983512
rect 394424 983492 394476 983512
rect 394476 983492 394478 983512
rect 394422 983456 394478 983492
rect 399758 983456 399814 983512
rect 636198 1001952 636254 1002008
rect 535458 983728 535514 983784
rect 636198 983728 636254 983784
rect 483846 982524 483902 982560
rect 483846 982504 483848 982524
rect 483848 982504 483900 982524
rect 483900 982504 483902 982524
rect 289726 980872 289782 980928
rect 30102 960200 30158 960256
rect 651378 959132 651434 959168
rect 651378 959112 651380 959132
rect 651380 959112 651432 959132
rect 651432 959112 651434 959132
rect 677414 959132 677470 959168
rect 677414 959112 677416 959132
rect 677416 959112 677468 959132
rect 677468 959112 677470 959132
rect 63406 958976 63462 959032
rect 676034 897116 676090 897152
rect 676034 897096 676036 897116
rect 676036 897096 676088 897116
rect 676088 897096 676090 897116
rect 651470 868536 651526 868592
rect 651470 867448 651526 867504
rect 651470 866224 651526 866280
rect 651378 865172 651380 865192
rect 651380 865172 651432 865192
rect 651432 865172 651434 865192
rect 651378 865136 651434 865172
rect 651470 863812 651472 863832
rect 651472 863812 651524 863832
rect 651524 863812 651526 863832
rect 651470 863776 651526 863812
rect 675850 896688 675906 896744
rect 651470 862280 651526 862336
rect 35806 817944 35862 818000
rect 35438 817264 35494 817320
rect 35622 816856 35678 816912
rect 35806 816040 35862 816096
rect 35622 815224 35678 815280
rect 35806 814408 35862 814464
rect 41326 813592 41382 813648
rect 40958 812776 41014 812832
rect 37922 811552 37978 811608
rect 34518 811144 34574 811200
rect 32586 810736 32642 810792
rect 31022 809920 31078 809976
rect 32586 802440 32642 802496
rect 36542 809512 36598 809568
rect 41326 812368 41382 812424
rect 41142 811960 41198 812016
rect 41970 810328 42026 810384
rect 41786 809920 41842 809976
rect 41326 809104 41382 809160
rect 41786 808696 41842 808752
rect 41142 808288 41198 808344
rect 41326 807492 41382 807528
rect 41326 807472 41328 807492
rect 41328 807472 41380 807492
rect 41380 807472 41382 807492
rect 41142 806656 41198 806712
rect 41326 806248 41382 806304
rect 41970 805568 42026 805624
rect 41786 805160 41842 805216
rect 42154 798088 42210 798144
rect 42062 797272 42118 797328
rect 41786 794824 41842 794880
rect 42154 794416 42210 794472
rect 42430 791968 42486 792024
rect 41786 790608 41842 790664
rect 41786 789248 41842 789304
rect 42430 788296 42486 788352
rect 42430 788024 42486 788080
rect 35806 774696 35862 774752
rect 35438 773880 35494 773936
rect 35806 773472 35862 773528
rect 39578 773472 39634 773528
rect 35806 773100 35808 773120
rect 35808 773100 35860 773120
rect 35860 773100 35862 773120
rect 35806 773064 35862 773100
rect 40314 773064 40370 773120
rect 35622 772656 35678 772712
rect 35622 772248 35678 772304
rect 40774 772248 40830 772304
rect 42890 772248 42946 772304
rect 35438 771840 35494 771896
rect 35806 771840 35862 771896
rect 35438 771024 35494 771080
rect 35622 770616 35678 770672
rect 35806 770208 35862 770264
rect 40498 770208 40554 770264
rect 43074 770208 43130 770264
rect 35622 769392 35678 769448
rect 39946 769392 40002 769448
rect 35806 768984 35862 769040
rect 35162 768168 35218 768224
rect 32402 767760 32458 767816
rect 33782 766944 33838 767000
rect 35806 767352 35862 767408
rect 35806 766128 35862 766184
rect 35806 765720 35862 765776
rect 35806 764532 35808 764552
rect 35808 764532 35860 764552
rect 35860 764532 35862 764552
rect 35806 764496 35862 764532
rect 35622 764088 35678 764144
rect 35806 763680 35862 763736
rect 35806 762864 35862 762920
rect 39762 765720 39818 765776
rect 39762 764532 39764 764552
rect 39764 764532 39816 764552
rect 39816 764532 39818 764552
rect 39762 764496 39818 764532
rect 39210 764088 39266 764144
rect 41694 763272 41750 763328
rect 41694 762864 41750 762920
rect 39302 758276 39304 758296
rect 39304 758276 39356 758296
rect 39356 758276 39358 758296
rect 39302 758240 39358 758276
rect 36542 757696 36598 757752
rect 41786 757016 41842 757072
rect 41878 756608 41934 756664
rect 42614 762864 42670 762920
rect 42338 753888 42394 753944
rect 42062 752936 42118 752992
rect 42154 751712 42210 751768
rect 42062 750896 42118 750952
rect 41786 750488 41842 750544
rect 41786 746680 41842 746736
rect 42798 758240 42854 758296
rect 42338 745592 42394 745648
rect 42890 752936 42946 752992
rect 42614 745048 42670 745104
rect 41878 743008 41934 743064
rect 42430 730496 42486 730552
rect 41326 729272 41382 729328
rect 40682 728626 40738 728682
rect 41326 728680 41382 728682
rect 41326 728628 41328 728680
rect 41328 728628 41380 728680
rect 41380 728628 41382 728680
rect 41326 728626 41382 728628
rect 40866 728048 40922 728104
rect 42982 727640 43038 727696
rect 42982 727232 43038 727288
rect 41142 726824 41198 726880
rect 40958 726416 41014 726472
rect 40958 725600 41014 725656
rect 32402 725192 32458 725248
rect 31666 723968 31722 724024
rect 35162 724784 35218 724840
rect 37278 724376 37334 724432
rect 39302 723152 39358 723208
rect 37278 716896 37334 716952
rect 41786 725600 41842 725656
rect 41786 722336 41842 722392
rect 41602 719208 41658 719264
rect 40958 718936 41014 718992
rect 42798 720296 42854 720352
rect 42246 719208 42302 719264
rect 42062 718936 42118 718992
rect 41786 718528 41842 718584
rect 40222 715808 40278 715864
rect 40590 715264 40646 715320
rect 42706 715808 42762 715864
rect 42430 715264 42486 715320
rect 41694 714448 41750 714504
rect 42062 709824 42118 709880
rect 41878 708464 41934 708520
rect 42062 708464 42118 708520
rect 42154 707648 42210 707704
rect 41786 707376 41842 707432
rect 42246 706152 42302 706208
rect 42062 703432 42118 703488
rect 42062 703024 42118 703080
rect 42706 703024 42762 703080
rect 42614 702752 42670 702808
rect 42614 702072 42670 702128
rect 42430 701800 42486 701856
rect 35438 688336 35494 688392
rect 35806 687656 35862 687712
rect 41694 687540 41750 687576
rect 41694 687520 41696 687540
rect 41696 687520 41748 687540
rect 41748 687520 41750 687540
rect 35622 687248 35678 687304
rect 35438 686840 35494 686896
rect 41694 687148 41696 687168
rect 41696 687148 41748 687168
rect 41748 687148 41750 687168
rect 41694 687112 41750 687148
rect 35806 686432 35862 686488
rect 35806 686044 35862 686080
rect 35806 686024 35808 686044
rect 35808 686024 35860 686044
rect 35860 686024 35862 686044
rect 35806 685616 35862 685672
rect 35622 685208 35678 685264
rect 35806 684800 35862 684856
rect 35622 684392 35678 684448
rect 35438 683984 35494 684040
rect 41694 685072 41750 685128
rect 41694 684256 41750 684312
rect 41694 683848 41750 683904
rect 42982 683848 43038 683904
rect 35806 683168 35862 683224
rect 35622 682760 35678 682816
rect 35162 681944 35218 682000
rect 33046 681536 33102 681592
rect 31022 680720 31078 680776
rect 33782 681128 33838 681184
rect 35806 682352 35862 682408
rect 41786 681672 41842 681728
rect 41694 680620 41696 680640
rect 41696 680620 41748 680640
rect 41748 680620 41750 680640
rect 41694 680584 41750 680620
rect 35806 680312 35862 680368
rect 35622 679904 35678 679960
rect 35438 679496 35494 679552
rect 41694 679396 41696 679416
rect 41696 679396 41748 679416
rect 41748 679396 41750 679416
rect 41694 679360 41750 679396
rect 35806 679088 35862 679144
rect 41786 678272 41842 678328
rect 40774 677748 40830 677750
rect 40774 677696 40776 677748
rect 40776 677696 40828 677748
rect 40828 677696 40830 677748
rect 40774 677694 40830 677696
rect 33782 672696 33838 672752
rect 42430 673104 42486 673160
rect 39578 670928 39634 670984
rect 42982 677864 43038 677920
rect 42798 677048 42854 677104
rect 41970 668480 42026 668536
rect 42154 667664 42210 667720
rect 42338 667392 42394 667448
rect 42062 666984 42118 667040
rect 41786 665216 41842 665272
rect 41786 664128 41842 664184
rect 41786 658280 41842 658336
rect 41786 657192 41842 657248
rect 42522 658552 42578 658608
rect 35806 644680 35862 644736
rect 38566 644272 38622 644328
rect 39578 644272 39634 644328
rect 35346 643864 35402 643920
rect 35530 643456 35586 643512
rect 35806 643492 35808 643512
rect 35808 643492 35860 643512
rect 35860 643492 35862 643512
rect 35806 643456 35862 643492
rect 35806 642640 35862 642696
rect 35622 642232 35678 642288
rect 39762 643864 39818 643920
rect 35806 641860 35808 641880
rect 35808 641860 35860 641880
rect 35860 641860 35862 641880
rect 35806 641824 35862 641860
rect 35622 641416 35678 641472
rect 35806 641008 35862 641064
rect 39302 641008 39358 641064
rect 35806 640600 35862 640656
rect 40774 642232 40830 642288
rect 40222 640192 40278 640248
rect 34426 639784 34482 639840
rect 35530 639376 35586 639432
rect 35806 639376 35862 639432
rect 40406 639376 40462 639432
rect 40866 638968 40922 639024
rect 35622 638560 35678 638616
rect 32402 637744 32458 637800
rect 35162 637336 35218 637392
rect 32402 629856 32458 629912
rect 35806 638152 35862 638208
rect 35806 636928 35862 636984
rect 35530 636520 35586 636576
rect 35806 636520 35862 636576
rect 35806 635704 35862 635760
rect 35806 634480 35862 634536
rect 35806 633664 35862 633720
rect 39946 632848 40002 632904
rect 40590 636520 40646 636576
rect 40590 634480 40646 634536
rect 40130 632440 40186 632496
rect 41510 633256 41566 633312
rect 40774 632168 40830 632224
rect 42154 633256 42210 633312
rect 40498 630536 40554 630592
rect 39302 629176 39358 629232
rect 39670 628224 39726 628280
rect 41786 627408 41842 627464
rect 41786 627136 41842 627192
rect 42522 636520 42578 636576
rect 42890 632848 42946 632904
rect 42706 628224 42762 628280
rect 42522 625912 42578 625968
rect 42154 624552 42210 624608
rect 41970 623328 42026 623384
rect 42062 622104 42118 622160
rect 41786 620880 41842 620936
rect 41970 620200 42026 620256
rect 42706 616800 42762 616856
rect 42430 616392 42486 616448
rect 42062 615848 42118 615904
rect 42614 615848 42670 615904
rect 42706 615440 42762 615496
rect 42246 612348 42248 612368
rect 42248 612348 42300 612368
rect 42300 612348 42302 612368
rect 42246 612312 42302 612348
rect 43626 797272 43682 797328
rect 43442 773472 43498 773528
rect 43442 769392 43498 769448
rect 44178 764496 44234 764552
rect 43626 764088 43682 764144
rect 43626 750896 43682 750952
rect 43626 731312 43682 731368
rect 44178 729680 44234 729736
rect 46202 773064 46258 773120
rect 44730 765720 44786 765776
rect 44914 763272 44970 763328
rect 44546 730088 44602 730144
rect 43994 723560 44050 723616
rect 43626 721112 43682 721168
rect 43442 685072 43498 685128
rect 43442 684256 43498 684312
rect 43442 644272 43498 644328
rect 43810 707648 43866 707704
rect 43994 703432 44050 703488
rect 44730 722744 44786 722800
rect 44730 708464 44786 708520
rect 43994 679360 44050 679416
rect 44362 641008 44418 641064
rect 44546 640192 44602 640248
rect 44362 634480 44418 634536
rect 43810 632440 43866 632496
rect 43534 630536 43590 630592
rect 43994 632168 44050 632224
rect 44178 624552 44234 624608
rect 44178 622104 44234 622160
rect 43534 610952 43590 611008
rect 40314 601976 40370 602032
rect 33782 601704 33838 601760
rect 33046 595176 33102 595232
rect 31022 594360 31078 594416
rect 39946 601296 40002 601352
rect 37922 595754 37978 595810
rect 35162 594768 35218 594824
rect 33782 589600 33838 589656
rect 35622 591912 35678 591968
rect 35806 591504 35862 591560
rect 35162 585928 35218 585984
rect 40130 600888 40186 600944
rect 45098 751712 45154 751768
rect 46202 730904 46258 730960
rect 45098 721520 45154 721576
rect 45098 708736 45154 708792
rect 45282 687520 45338 687576
rect 46202 687112 46258 687168
rect 45466 680584 45522 680640
rect 45834 667664 45890 667720
rect 45650 666984 45706 667040
rect 46202 643864 46258 643920
rect 45098 642232 45154 642288
rect 45098 639376 45154 639432
rect 44730 610952 44786 611008
rect 44546 600480 44602 600536
rect 44914 600072 44970 600128
rect 44638 599256 44694 599312
rect 43074 597624 43130 597680
rect 42890 596944 42946 597000
rect 42430 596808 42486 596864
rect 41326 595754 41382 595810
rect 41694 595756 41696 595776
rect 41696 595756 41748 595776
rect 41748 595756 41750 595776
rect 41694 595720 41750 595756
rect 41694 594496 41750 594552
rect 41786 593544 41842 593600
rect 41786 592320 41842 592376
rect 40774 589328 40830 589384
rect 41510 589056 41566 589112
rect 40406 585656 40462 585712
rect 39302 584568 39358 584624
rect 41786 584296 41842 584352
rect 41786 583888 41842 583944
rect 42246 582392 42302 582448
rect 42062 580624 42118 580680
rect 41878 580216 41934 580272
rect 42246 580216 42302 580272
rect 41786 579536 41842 579592
rect 42062 579264 42118 579320
rect 42154 578312 42210 578368
rect 41786 577768 41842 577824
rect 42154 575728 42210 575784
rect 41786 574640 41842 574696
rect 42614 572872 42670 572928
rect 42062 572600 42118 572656
rect 42062 571512 42118 571568
rect 42430 571376 42486 571432
rect 41786 570152 41842 570208
rect 40958 558048 41014 558104
rect 37922 553352 37978 553408
rect 29642 551928 29698 551984
rect 42798 555600 42854 555656
rect 44362 593136 44418 593192
rect 43442 589328 43498 589384
rect 43626 581168 43682 581224
rect 43626 579808 43682 579864
rect 44362 578312 44418 578368
rect 43074 554784 43130 554840
rect 41326 553352 41382 553408
rect 43074 550704 43130 550760
rect 42062 550432 42118 550488
rect 40682 549888 40738 549944
rect 39578 547440 39634 547496
rect 41326 548256 41382 548312
rect 40682 545536 40738 545592
rect 42798 549072 42854 549128
rect 39578 542544 39634 542600
rect 37922 542272 37978 542328
rect 42614 539552 42670 539608
rect 42430 538192 42486 538248
rect 42154 537920 42210 537976
rect 42430 536424 42486 536480
rect 42154 535608 42210 535664
rect 42430 533840 42486 533896
rect 42246 533296 42302 533352
rect 44362 556824 44418 556880
rect 43718 554376 43774 554432
rect 43810 552336 43866 552392
rect 43994 551112 44050 551168
rect 42614 531664 42670 531720
rect 42430 530168 42486 530224
rect 42062 529896 42118 529952
rect 42430 528944 42486 529000
rect 42614 528944 42670 529000
rect 42798 527176 42854 527232
rect 35806 430072 35862 430128
rect 35806 428440 35862 428496
rect 41786 428440 41842 428496
rect 41786 426536 41842 426592
rect 42890 426536 42946 426592
rect 41142 425992 41198 426048
rect 39302 425584 39358 425640
rect 33046 424768 33102 424824
rect 34518 424360 34574 424416
rect 33782 423952 33838 424008
rect 42706 422728 42762 422784
rect 41878 421912 41934 421968
rect 41878 418648 41934 418704
rect 39302 415248 39358 415304
rect 33782 414568 33838 414624
rect 41786 413480 41842 413536
rect 41786 413072 41842 413128
rect 42430 407904 42486 407960
rect 42062 407496 42118 407552
rect 41786 406952 41842 407008
rect 41786 406680 41842 406736
rect 42430 404912 42486 404968
rect 42246 404504 42302 404560
rect 42338 402872 42394 402928
rect 42430 402464 42486 402520
rect 42430 401920 42486 401976
rect 41786 400016 41842 400072
rect 41970 399336 42026 399392
rect 41786 398792 41842 398848
rect 42154 397432 42210 397488
rect 41326 387096 41382 387152
rect 41142 386688 41198 386744
rect 40866 385872 40922 385928
rect 41142 385872 41198 385928
rect 41050 383016 41106 383072
rect 41326 383016 41382 383072
rect 40866 382608 40922 382664
rect 40038 382200 40094 382256
rect 35530 381792 35586 381848
rect 33966 380976 34022 381032
rect 39302 381384 39358 381440
rect 35806 379344 35862 379400
rect 35806 377304 35862 377360
rect 35806 376488 35862 376544
rect 35806 376080 35862 376136
rect 35530 374584 35586 374640
rect 41050 381792 41106 381848
rect 42890 385600 42946 385656
rect 41786 381520 41842 381576
rect 42890 379888 42946 379944
rect 40038 379344 40094 379400
rect 40406 377304 40462 377360
rect 41510 376488 41566 376544
rect 41694 376488 41750 376544
rect 41510 376080 41566 376136
rect 42062 366152 42118 366208
rect 41786 364792 41842 364848
rect 41786 364112 41842 364168
rect 42062 363568 42118 363624
rect 42614 365744 42670 365800
rect 42246 362208 42302 362264
rect 41786 360032 41842 360088
rect 42430 358944 42486 359000
rect 41878 358672 41934 358728
rect 41786 356904 41842 356960
rect 42246 356088 42302 356144
rect 43074 377304 43130 377360
rect 43074 366152 43130 366208
rect 43074 364248 43130 364304
rect 42798 356632 42854 356688
rect 43258 355272 43314 355328
rect 43810 533840 43866 533896
rect 44178 550160 44234 550216
rect 44178 538192 44234 538248
rect 43994 529896 44050 529952
rect 45466 638968 45522 639024
rect 45282 599664 45338 599720
rect 45466 598848 45522 598904
rect 45098 598032 45154 598088
rect 45098 580624 45154 580680
rect 44914 558728 44970 558784
rect 44638 556416 44694 556472
rect 44546 556008 44602 556064
rect 44362 429664 44418 429720
rect 44178 429256 44234 429312
rect 43626 427216 43682 427272
rect 43994 425176 44050 425232
rect 43810 423544 43866 423600
rect 43626 420688 43682 420744
rect 43810 402464 43866 402520
rect 43994 401920 44050 401976
rect 45098 555192 45154 555248
rect 45282 551520 45338 551576
rect 45466 548664 45522 548720
rect 44730 542544 44786 542600
rect 45190 539824 45246 539880
rect 45190 537920 45246 537976
rect 45190 535608 45246 535664
rect 44822 430888 44878 430944
rect 44546 428848 44602 428904
rect 44362 427624 44418 427680
rect 44178 386416 44234 386472
rect 44638 423136 44694 423192
rect 44638 402872 44694 402928
rect 45650 536832 45706 536888
rect 45466 528944 45522 529000
rect 45282 527176 45338 527232
rect 45098 428032 45154 428088
rect 45282 426808 45338 426864
rect 45006 421096 45062 421152
rect 45006 407496 45062 407552
rect 45098 385192 45154 385248
rect 44362 384784 44418 384840
rect 44914 384376 44970 384432
rect 44546 380296 44602 380352
rect 44178 378256 44234 378312
rect 43810 376488 43866 376544
rect 44178 363568 44234 363624
rect 44730 364248 44786 364304
rect 44546 358944 44602 359000
rect 43810 355816 43866 355872
rect 43626 355544 43682 355600
rect 44638 355272 44694 355328
rect 42706 354320 42762 354376
rect 43994 354592 44050 354648
rect 43994 354320 44050 354376
rect 42706 351872 42762 351928
rect 35530 344256 35586 344312
rect 35806 344256 35862 344312
rect 45282 383968 45338 384024
rect 45282 383560 45338 383616
rect 39854 343848 39910 343904
rect 44914 343848 44970 343904
rect 33046 343440 33102 343496
rect 35806 341808 35862 341864
rect 33046 341400 33102 341456
rect 40038 343440 40094 343496
rect 45006 343440 45062 343496
rect 40222 342216 40278 342272
rect 45466 382608 45522 382664
rect 46018 355816 46074 355872
rect 45834 355544 45890 355600
rect 45650 353812 45652 353832
rect 45652 353812 45704 353832
rect 45704 353812 45706 353832
rect 45650 353776 45706 353812
rect 45650 352144 45706 352200
rect 45466 343168 45522 343224
rect 45558 342760 45614 342816
rect 45190 342488 45246 342544
rect 44822 341808 44878 341864
rect 45006 341808 45062 341864
rect 35530 341028 35532 341048
rect 35532 341028 35584 341048
rect 35584 341028 35586 341048
rect 35530 340992 35586 341028
rect 35806 340992 35862 341048
rect 40038 340584 40094 340640
rect 44822 340992 44878 341048
rect 45374 340584 45430 340640
rect 39854 340176 39910 340232
rect 40222 340176 40278 340232
rect 35530 339768 35586 339824
rect 35806 339768 35862 339824
rect 39854 339768 39910 339824
rect 35162 338544 35218 338600
rect 35806 335688 35862 335744
rect 35806 334872 35862 334928
rect 45374 338000 45430 338056
rect 38934 335688 38990 335744
rect 42062 334600 42118 334656
rect 43810 334600 43866 334656
rect 45098 334600 45154 334656
rect 37922 332832 37978 332888
rect 40222 334056 40278 334112
rect 39762 332424 39818 332480
rect 35162 331744 35218 331800
rect 42982 334056 43038 334112
rect 42798 332424 42854 332480
rect 42062 327664 42118 327720
rect 42430 326984 42486 327040
rect 41786 324808 41842 324864
rect 41786 322768 41842 322824
rect 42062 321544 42118 321600
rect 42062 321136 42118 321192
rect 42430 320728 42486 320784
rect 42982 321136 43038 321192
rect 42614 319368 42670 319424
rect 42430 318960 42486 319016
rect 42246 317464 42302 317520
rect 42062 317192 42118 317248
rect 41786 315968 41842 316024
rect 41786 315560 41842 315616
rect 42154 313656 42210 313712
rect 42430 313112 42486 313168
rect 42246 312432 42302 312488
rect 42062 311888 42118 311944
rect 41142 300872 41198 300928
rect 42798 298968 42854 299024
rect 41970 298696 42026 298752
rect 41326 296384 41382 296440
rect 39302 295976 39358 296032
rect 33046 294752 33102 294808
rect 33782 294344 33838 294400
rect 35806 291896 35862 291952
rect 35162 290264 35218 290320
rect 33782 284824 33838 284880
rect 42338 295160 42394 295216
rect 41786 293936 41842 293992
rect 40590 292544 40592 292588
rect 40592 292544 40644 292588
rect 40644 292544 40646 292588
rect 40590 292532 40646 292544
rect 41786 290400 41842 290456
rect 39302 284280 39358 284336
rect 42154 279792 42210 279848
rect 42430 279384 42486 279440
rect 41970 278432 42026 278488
rect 42062 277208 42118 277264
rect 42522 275848 42578 275904
rect 41786 274216 41842 274272
rect 41786 272992 41842 273048
rect 41786 272176 41842 272232
rect 41786 270000 41842 270056
rect 41970 269048 42026 269104
rect 42430 267688 42486 267744
rect 42154 266192 42210 266248
rect 35806 257080 35862 257136
rect 39578 257080 39634 257136
rect 35622 255856 35678 255912
rect 39946 255856 40002 255912
rect 35806 255468 35862 255504
rect 35806 255448 35808 255468
rect 35808 255448 35860 255468
rect 35860 255448 35862 255468
rect 35806 254632 35862 254688
rect 35622 254224 35678 254280
rect 43166 297200 43222 297256
rect 42982 293528 43038 293584
rect 43350 290400 43406 290456
rect 43994 334464 44050 334520
rect 44362 334328 44418 334384
rect 44178 334192 44234 334248
rect 44178 321544 44234 321600
rect 44362 317192 44418 317248
rect 44270 311208 44326 311264
rect 44270 298016 44326 298072
rect 43994 278704 44050 278760
rect 43810 278296 43866 278352
rect 43350 273808 43406 273864
rect 43258 263200 43314 263256
rect 43258 257080 43314 257136
rect 43074 255856 43130 255912
rect 40498 254632 40554 254688
rect 35806 253816 35862 253872
rect 35622 253408 35678 253464
rect 41510 253816 41566 253872
rect 35806 253000 35862 253056
rect 40682 253000 40738 253056
rect 42890 253000 42946 253056
rect 35806 252184 35862 252240
rect 35806 250552 35862 250608
rect 40314 245656 40370 245712
rect 42246 240080 42302 240136
rect 42246 238448 42302 238504
rect 41786 236544 41842 236600
rect 42338 235864 42394 235920
rect 41786 234640 41842 234696
rect 42338 231920 42394 231976
rect 42338 231240 42394 231296
rect 42154 230288 42210 230344
rect 42706 237360 42762 237416
rect 42706 232192 42762 232248
rect 41970 227296 42026 227352
rect 42154 226616 42210 226672
rect 42430 223488 42486 223544
rect 42154 223216 42210 223272
rect 35806 217912 35862 217968
rect 35806 214648 35862 214704
rect 35806 214240 35862 214296
rect 39762 214240 39818 214296
rect 39854 213016 39910 213072
rect 35806 212644 35808 212664
rect 35808 212644 35860 212664
rect 35860 212644 35862 212664
rect 35806 212608 35862 212644
rect 43074 245656 43130 245712
rect 43626 269728 43682 269784
rect 43626 263200 43682 263256
rect 44638 299648 44694 299704
rect 44454 297608 44510 297664
rect 44454 293120 44510 293176
rect 44454 279792 44510 279848
rect 44822 284280 44878 284336
rect 44730 257624 44786 257680
rect 44546 256808 44602 256864
rect 44914 256400 44970 256456
rect 44270 255176 44326 255232
rect 43810 254632 43866 254688
rect 43626 253816 43682 253872
rect 44454 251504 44510 251560
rect 44178 250280 44234 250336
rect 44638 251096 44694 251152
rect 44454 240080 44510 240136
rect 44178 230288 44234 230344
rect 44638 226616 44694 226672
rect 43442 214240 43498 214296
rect 40774 212200 40830 212256
rect 42890 212200 42946 212256
rect 35622 211792 35678 211848
rect 40130 211792 40186 211848
rect 35806 211420 35808 211440
rect 35808 211420 35860 211440
rect 35860 211420 35862 211440
rect 35806 211384 35862 211420
rect 44914 213696 44970 213752
rect 43810 213016 43866 213072
rect 43626 211792 43682 211848
rect 35806 210160 35862 210216
rect 35622 209344 35678 209400
rect 35806 208120 35862 208176
rect 35806 207304 35862 207360
rect 39210 206896 39266 206952
rect 35806 206080 35862 206136
rect 44454 208528 44510 208584
rect 44178 207984 44234 208040
rect 40958 207712 41014 207768
rect 43258 207712 43314 207768
rect 40958 207304 41014 207360
rect 43074 207304 43130 207360
rect 42890 206896 42946 206952
rect 39946 205264 40002 205320
rect 35806 204856 35862 204912
rect 41510 204856 41566 204912
rect 35806 204448 35862 204504
rect 41510 204448 41566 204504
rect 41694 204484 41696 204504
rect 41696 204484 41748 204504
rect 41748 204484 41750 204504
rect 41694 204448 41750 204484
rect 39394 204040 39450 204096
rect 42706 204040 42762 204096
rect 35806 203632 35862 203688
rect 42430 201320 42486 201376
rect 39302 197784 39358 197840
rect 41878 195744 41934 195800
rect 42338 195472 42394 195528
rect 41786 195200 41842 195256
rect 41786 193432 41842 193488
rect 42338 193160 42394 193216
rect 42246 192752 42302 192808
rect 42062 191528 42118 191584
rect 42430 190440 42486 190496
rect 42430 189896 42486 189952
rect 42430 187584 42486 187640
rect 42338 186224 42394 186280
rect 42154 185952 42210 186008
rect 43442 205264 43498 205320
rect 43810 204448 43866 204504
rect 43442 201320 43498 201376
rect 42430 183096 42486 183152
rect 42062 179288 42118 179344
rect 43810 191528 43866 191584
rect 43626 187584 43682 187640
rect 44638 205536 44694 205592
rect 44638 190440 44694 190496
rect 44454 189896 44510 189952
rect 44178 183096 44234 183152
rect 45282 326984 45338 327040
rect 45742 340992 45798 341048
rect 45558 300056 45614 300112
rect 46018 340176 46074 340232
rect 45742 299240 45798 299296
rect 46018 298424 46074 298480
rect 45282 292712 45338 292768
rect 45466 291488 45522 291544
rect 45558 284316 45560 284336
rect 45560 284316 45612 284336
rect 45612 284316 45614 284336
rect 45558 284280 45614 284316
rect 45374 278976 45430 279032
rect 45466 278704 45522 278760
rect 45374 277208 45430 277264
rect 46938 380704 46994 380760
rect 47582 376080 47638 376136
rect 46938 356088 46994 356144
rect 46570 338408 46626 338464
rect 46386 337592 46442 337648
rect 46570 318960 46626 319016
rect 46386 313112 46442 313168
rect 46938 296792 46994 296848
rect 47582 290672 47638 290728
rect 46938 267688 46994 267744
rect 46386 258032 46442 258088
rect 46938 252728 46994 252784
rect 45558 249056 45614 249112
rect 45926 248648 45982 248704
rect 45742 248240 45798 248296
rect 45742 235864 45798 235920
rect 46110 247016 46166 247072
rect 46110 238448 46166 238504
rect 45926 232192 45982 232248
rect 45558 231240 45614 231296
rect 47122 251912 47178 251968
rect 47122 231920 47178 231976
rect 46938 223488 46994 223544
rect 46202 204856 46258 204912
rect 47766 247424 47822 247480
rect 49146 291080 49202 291136
rect 62210 790472 62266 790528
rect 62118 787344 62174 787400
rect 62118 786120 62174 786176
rect 62946 789112 63002 789168
rect 62946 787072 63002 787128
rect 62762 784896 62818 784952
rect 51722 581168 51778 581224
rect 51722 539824 51778 539880
rect 50526 419872 50582 419928
rect 51078 407904 51134 407960
rect 51446 404912 51502 404968
rect 51078 397432 51134 397488
rect 51078 362208 51134 362264
rect 51722 301280 51778 301336
rect 50526 247832 50582 247888
rect 54482 558456 54538 558512
rect 54482 430480 54538 430536
rect 54482 387504 54538 387560
rect 53838 320728 53894 320784
rect 53838 312432 53894 312488
rect 54482 300464 54538 300520
rect 51722 223488 51778 223544
rect 55862 277480 55918 277536
rect 56046 266192 56102 266248
rect 62762 747632 62818 747688
rect 62118 746136 62174 746192
rect 62118 744096 62174 744152
rect 62118 743724 62120 743744
rect 62120 743724 62172 743744
rect 62172 743724 62174 743744
rect 62118 743688 62174 743724
rect 62118 742364 62120 742384
rect 62120 742364 62172 742384
rect 62172 742364 62174 742384
rect 62118 742328 62174 742364
rect 63038 741784 63094 741840
rect 57426 275848 57482 275904
rect 62118 704384 62174 704440
rect 62118 703296 62174 703352
rect 62210 701256 62266 701312
rect 62762 700848 62818 700904
rect 62302 699524 62304 699544
rect 62304 699524 62356 699544
rect 62356 699524 62358 699544
rect 62302 699488 62358 699524
rect 62118 698128 62174 698184
rect 62118 660900 62120 660920
rect 62120 660900 62172 660920
rect 62172 660900 62174 660920
rect 62118 660864 62174 660900
rect 62118 659540 62120 659560
rect 62120 659540 62172 659560
rect 62172 659540 62174 659560
rect 62118 659504 62174 659540
rect 62118 658280 62174 658336
rect 62118 656512 62174 656568
rect 63406 657600 63462 657656
rect 62302 655288 62358 655344
rect 62118 616528 62174 616584
rect 62118 614624 62174 614680
rect 62118 613808 62174 613864
rect 62118 612584 62174 612640
rect 63130 618024 63186 618080
rect 62946 612040 63002 612096
rect 62762 595720 62818 595776
rect 62578 590008 62634 590064
rect 62118 574776 62174 574832
rect 62118 573552 62174 573608
rect 63130 594088 63186 594144
rect 62946 590688 63002 590744
rect 62762 571104 62818 571160
rect 62578 569880 62634 569936
rect 62210 556688 62266 556744
rect 62762 550160 62818 550216
rect 62118 531276 62174 531312
rect 62118 531256 62120 531276
rect 62120 531256 62172 531276
rect 62172 531256 62174 531276
rect 62118 530576 62174 530632
rect 62118 528572 62120 528592
rect 62120 528572 62172 528592
rect 62172 528572 62174 528592
rect 62118 528536 62174 528572
rect 62302 527992 62358 528048
rect 62118 527076 62120 527096
rect 62120 527076 62172 527096
rect 62172 527076 62174 527096
rect 62118 527040 62174 527076
rect 62762 525680 62818 525736
rect 62394 428440 62450 428496
rect 62118 404096 62174 404152
rect 62118 402600 62174 402656
rect 62118 400560 62174 400616
rect 62394 400152 62450 400208
rect 62118 399336 62174 399392
rect 62118 398248 62174 398304
rect 62762 381520 62818 381576
rect 62118 360848 62174 360904
rect 62118 359760 62174 359816
rect 62302 357448 62358 357504
rect 62302 356632 62358 356688
rect 62118 355952 62174 356008
rect 62762 354456 62818 354512
rect 62670 341672 62726 341728
rect 62302 341400 62358 341456
rect 62486 332560 62542 332616
rect 61566 319368 61622 319424
rect 62118 317364 62120 317384
rect 62120 317364 62172 317384
rect 62172 317364 62174 317384
rect 62118 317328 62174 317364
rect 61566 315968 61622 316024
rect 62118 314764 62174 314800
rect 62118 314744 62120 314764
rect 62120 314744 62172 314764
rect 62172 314744 62174 314764
rect 62394 314064 62450 314120
rect 62302 295296 62358 295352
rect 62118 294092 62174 294128
rect 62118 294072 62120 294092
rect 62120 294072 62172 294092
rect 62172 294072 62174 294092
rect 62118 292460 62174 292496
rect 62118 292440 62120 292460
rect 62120 292440 62172 292460
rect 62172 292440 62174 292460
rect 62118 290944 62174 291000
rect 62118 288516 62174 288552
rect 62118 288496 62120 288516
rect 62120 288496 62172 288516
rect 62172 288496 62174 288516
rect 62118 285912 62174 285968
rect 62762 311752 62818 311808
rect 62762 292712 62818 292768
rect 62762 287136 62818 287192
rect 62486 282104 62542 282160
rect 62302 280880 62358 280936
rect 62118 280372 62120 280392
rect 62120 280372 62172 280392
rect 62172 280372 62174 280392
rect 62118 280336 62174 280372
rect 61934 279384 61990 279440
rect 63130 568520 63186 568576
rect 63130 385872 63186 385928
rect 63130 357176 63186 357232
rect 63222 341944 63278 342000
rect 63222 312976 63278 313032
rect 63130 298696 63186 298752
rect 63130 289720 63186 289776
rect 62946 284552 63002 284608
rect 63130 283192 63186 283248
rect 62946 280064 63002 280120
rect 62302 273808 62358 273864
rect 62486 269728 62542 269784
rect 62854 265512 62910 265568
rect 61382 264152 61438 264208
rect 54482 217912 54538 217968
rect 63406 278704 63462 278760
rect 63406 278024 63462 278080
rect 63590 278024 63646 278080
rect 63590 277480 63646 277536
rect 651470 778368 651526 778424
rect 652022 777008 652078 777064
rect 651470 776056 651526 776112
rect 651378 775276 651380 775296
rect 651380 775276 651432 775296
rect 651432 775276 651434 775296
rect 651378 775240 651434 775276
rect 651470 774172 651526 774208
rect 651470 774152 651472 774172
rect 651472 774152 651524 774172
rect 651524 774152 651526 774172
rect 651470 773336 651526 773392
rect 651470 734168 651526 734224
rect 652666 732808 652722 732864
rect 651470 731720 651526 731776
rect 651378 731076 651380 731096
rect 651380 731076 651432 731096
rect 651432 731076 651434 731096
rect 651378 731040 651434 731076
rect 651470 729816 651526 729872
rect 651470 728492 651472 728512
rect 651472 728492 651524 728512
rect 651524 728492 651526 728512
rect 651470 728456 651526 728492
rect 651470 689424 651526 689480
rect 651654 688744 651710 688800
rect 651470 687384 651526 687440
rect 651470 686704 651526 686760
rect 651470 685208 651526 685264
rect 652574 684392 652630 684448
rect 651470 643184 651526 643240
rect 651838 641824 651894 641880
rect 651470 640736 651526 640792
rect 651378 640092 651380 640112
rect 651380 640092 651432 640112
rect 651432 640092 651434 640112
rect 651378 640056 651434 640092
rect 651470 638560 651526 638616
rect 651654 638152 651710 638208
rect 651470 597896 651526 597952
rect 651470 596672 651526 596728
rect 651470 595312 651526 595368
rect 651654 595040 651710 595096
rect 651470 594088 651526 594144
rect 651470 592864 651526 592920
rect 651470 553424 651526 553480
rect 651470 552064 651526 552120
rect 652022 550976 652078 551032
rect 651654 550332 651656 550352
rect 651656 550332 651708 550352
rect 651708 550332 651710 550352
rect 651654 550296 651710 550332
rect 651470 549228 651526 549264
rect 651470 549208 651472 549228
rect 651472 549208 651524 549228
rect 651524 549208 651526 549228
rect 651470 548392 651526 548448
rect 667386 600888 667442 600944
rect 636198 278296 636254 278352
rect 460938 272312 460994 272368
rect 464802 272448 464858 272504
rect 463698 272312 463754 272368
rect 470690 272484 470692 272504
rect 470692 272484 470744 272504
rect 470744 272484 470746 272504
rect 470690 272448 470746 272484
rect 470598 271904 470654 271960
rect 478050 271904 478106 271960
rect 479522 271904 479578 271960
rect 480534 271940 480536 271960
rect 480536 271940 480588 271960
rect 480588 271940 480590 271960
rect 480534 271904 480590 271940
rect 501602 271904 501658 271960
rect 504546 271940 504548 271960
rect 504548 271940 504600 271960
rect 504600 271940 504602 271960
rect 504546 271904 504602 271940
rect 509238 269864 509294 269920
rect 509146 269456 509202 269512
rect 509882 269492 509884 269512
rect 509884 269492 509936 269512
rect 509936 269492 509938 269512
rect 509882 269456 509938 269492
rect 516414 269864 516470 269920
rect 532238 270136 532294 270192
rect 534078 270136 534134 270192
rect 536562 272448 536618 272504
rect 539322 273944 539378 274000
rect 538034 269728 538090 269784
rect 545946 273964 546002 274000
rect 545946 273944 545948 273964
rect 545948 273944 546000 273964
rect 546000 273944 546002 273964
rect 542450 269764 542452 269784
rect 542452 269764 542504 269784
rect 542504 269764 542506 269784
rect 542450 269728 542506 269764
rect 547694 272448 547750 272504
rect 547510 272076 547512 272096
rect 547512 272076 547564 272096
rect 547564 272076 547566 272096
rect 547510 272040 547566 272076
rect 547878 272040 547934 272096
rect 635094 277752 635150 277808
rect 554410 262112 554466 262168
rect 554318 259936 554374 259992
rect 553950 257760 554006 257816
rect 554502 255604 554558 255640
rect 554502 255584 554504 255604
rect 554504 255584 554556 255604
rect 554556 255584 554558 255604
rect 554410 253408 554466 253464
rect 554134 251252 554190 251288
rect 554134 251232 554136 251252
rect 554136 251232 554188 251252
rect 554188 251232 554190 251252
rect 554042 249056 554098 249112
rect 553858 246880 553914 246936
rect 553490 244704 553546 244760
rect 553674 242528 553730 242584
rect 553766 236000 553822 236056
rect 64142 231104 64198 231160
rect 63406 223488 63462 223544
rect 140042 229064 140098 229120
rect 136638 227860 136694 227896
rect 136638 227840 136640 227860
rect 136640 227840 136692 227860
rect 136692 227840 136694 227860
rect 136178 219292 136234 219328
rect 136178 219272 136180 219292
rect 136180 219272 136232 219292
rect 136232 219272 136234 219292
rect 138018 224304 138074 224360
rect 137282 224032 137338 224088
rect 138110 224068 138112 224088
rect 138112 224068 138164 224088
rect 138164 224068 138166 224088
rect 138110 224032 138166 224068
rect 138478 221584 138534 221640
rect 137282 219272 137338 219328
rect 139858 222808 139914 222864
rect 142158 230152 142214 230208
rect 141974 229880 142030 229936
rect 141514 227860 141570 227896
rect 141514 227840 141516 227860
rect 141516 227840 141568 227860
rect 141568 227840 141570 227860
rect 142618 229900 142674 229936
rect 142618 229880 142620 229900
rect 142620 229880 142672 229900
rect 142672 229880 142674 229900
rect 143538 229064 143594 229120
rect 141790 226500 141846 226536
rect 141790 226480 141792 226500
rect 141792 226480 141844 226500
rect 141844 226480 141846 226500
rect 142250 226500 142306 226536
rect 142250 226480 142252 226500
rect 142252 226480 142304 226500
rect 142304 226480 142306 226500
rect 142618 225972 142620 225992
rect 142620 225972 142672 225992
rect 142672 225972 142674 225992
rect 142618 225936 142674 225972
rect 141514 221604 141570 221640
rect 141514 221584 141516 221604
rect 141516 221584 141568 221604
rect 141568 221584 141570 221604
rect 142526 223116 142528 223136
rect 142528 223116 142580 223136
rect 142580 223116 142582 223136
rect 142526 223080 142582 223116
rect 142066 221584 142122 221640
rect 143630 223116 143632 223136
rect 143632 223116 143684 223136
rect 143684 223116 143686 223136
rect 143630 223080 143686 223116
rect 144642 229356 144698 229392
rect 144642 229336 144644 229356
rect 144644 229336 144696 229356
rect 144696 229336 144698 229356
rect 145930 227976 145986 228032
rect 143814 222808 143870 222864
rect 147126 227976 147182 228032
rect 148322 229336 148378 229392
rect 147586 221604 147642 221640
rect 147586 221584 147588 221604
rect 147588 221584 147640 221604
rect 147640 221584 147642 221604
rect 147218 220804 147220 220824
rect 147220 220804 147272 220824
rect 147272 220804 147274 220824
rect 147218 220768 147274 220804
rect 147218 220380 147274 220416
rect 147218 220360 147220 220380
rect 147220 220360 147272 220380
rect 147272 220360 147274 220380
rect 148874 225392 148930 225448
rect 148322 220360 148378 220416
rect 150530 230152 150586 230208
rect 150346 229064 150402 229120
rect 149794 225936 149850 225992
rect 151358 226208 151414 226264
rect 151174 220768 151230 220824
rect 150714 220516 150770 220552
rect 150714 220496 150716 220516
rect 150716 220496 150768 220516
rect 150768 220496 150770 220516
rect 152370 224304 152426 224360
rect 151910 220516 151966 220552
rect 151910 220496 151912 220516
rect 151912 220496 151964 220516
rect 151964 220496 151966 220516
rect 151726 220244 151782 220280
rect 151726 220224 151728 220244
rect 151728 220224 151780 220244
rect 151780 220224 151782 220244
rect 155866 227024 155922 227080
rect 154394 220244 154450 220280
rect 154394 220224 154396 220244
rect 154396 220224 154448 220244
rect 154448 220224 154450 220244
rect 154486 218612 154542 218648
rect 154486 218592 154488 218612
rect 154488 218592 154540 218612
rect 154540 218592 154542 218612
rect 157430 230172 157486 230208
rect 157430 230152 157432 230172
rect 157432 230152 157484 230172
rect 157484 230152 157486 230172
rect 157154 230036 157210 230072
rect 157154 230016 157156 230036
rect 157156 230016 157208 230036
rect 157208 230016 157210 230036
rect 157798 230152 157854 230208
rect 157614 229608 157670 229664
rect 157154 229064 157210 229120
rect 157338 227432 157394 227488
rect 157430 227180 157486 227216
rect 157430 227160 157432 227180
rect 157432 227160 157484 227180
rect 157484 227160 157486 227180
rect 157154 226208 157210 226264
rect 156602 225800 156658 225856
rect 157798 225800 157854 225856
rect 157154 225392 157210 225448
rect 158718 229628 158774 229664
rect 158718 229608 158720 229628
rect 158720 229608 158772 229628
rect 158772 229608 158774 229628
rect 158350 220904 158406 220960
rect 160006 228520 160062 228576
rect 161294 230172 161350 230208
rect 161294 230152 161296 230172
rect 161296 230152 161348 230172
rect 161348 230152 161350 230172
rect 160190 218612 160246 218648
rect 160190 218592 160192 218612
rect 160192 218592 160244 218612
rect 160244 218592 160246 218612
rect 161432 221740 161488 221776
rect 161432 221720 161434 221740
rect 161434 221720 161486 221740
rect 161486 221720 161488 221740
rect 161570 220924 161626 220960
rect 161570 220904 161572 220924
rect 161572 220904 161624 220924
rect 161624 220904 161626 220924
rect 166354 228812 166410 228848
rect 166354 228792 166356 228812
rect 166356 228792 166408 228812
rect 166408 228792 166410 228812
rect 166814 228520 166870 228576
rect 166538 227432 166594 227488
rect 167366 229200 167422 229256
rect 167550 228792 167606 228848
rect 167642 221740 167698 221776
rect 167642 221720 167644 221740
rect 167644 221720 167696 221740
rect 167696 221720 167698 221740
rect 169390 227316 169446 227352
rect 169390 227296 169392 227316
rect 169392 227296 169444 227316
rect 169444 227296 169446 227316
rect 171690 227296 171746 227352
rect 170954 219292 171010 219328
rect 170954 219272 170956 219292
rect 170956 219272 171008 219292
rect 171008 219272 171010 219292
rect 171782 219272 171838 219328
rect 173346 221876 173402 221912
rect 173346 221856 173348 221876
rect 173348 221856 173400 221876
rect 173400 221856 173402 221876
rect 174358 229200 174414 229256
rect 176290 220632 176346 220688
rect 177394 221856 177450 221912
rect 180798 220904 180854 220960
rect 180890 220652 180946 220688
rect 180890 220632 180892 220652
rect 180892 220632 180944 220652
rect 180944 220632 180946 220652
rect 185122 220904 185178 220960
rect 185950 220768 186006 220824
rect 193034 228928 193090 228984
rect 190550 220788 190606 220824
rect 190550 220768 190552 220788
rect 190552 220768 190604 220788
rect 190604 220768 190606 220788
rect 195058 229900 195114 229936
rect 195058 229880 195060 229900
rect 195060 229880 195112 229900
rect 195112 229880 195114 229900
rect 195610 228948 195666 228984
rect 195610 228928 195612 228948
rect 195612 228928 195664 228948
rect 195664 228928 195666 228948
rect 196898 229880 196954 229936
rect 204810 227568 204866 227624
rect 205638 227588 205694 227624
rect 205638 227568 205640 227588
rect 205640 227568 205692 227588
rect 205692 227568 205694 227588
rect 486974 220224 487030 220280
rect 487802 218048 487858 218104
rect 488814 217096 488870 217152
rect 492954 219680 493010 219736
rect 493690 219680 493746 219736
rect 494702 218320 494758 218376
rect 495162 217096 495218 217152
rect 502246 217232 502302 217288
rect 510986 217504 511042 217560
rect 513562 221448 513618 221504
rect 515770 221176 515826 221232
rect 515126 219952 515182 220008
rect 520186 219408 520242 219464
rect 520002 217504 520058 217560
rect 522578 220904 522634 220960
rect 531502 217504 531558 217560
rect 532514 217504 532570 217560
rect 535734 221992 535790 222048
rect 539782 222028 539784 222048
rect 539784 222028 539836 222048
rect 539836 222028 539838 222048
rect 539782 221992 539838 222028
rect 547832 221756 547834 221776
rect 547834 221756 547886 221776
rect 547886 221756 547888 221776
rect 547832 221720 547888 221756
rect 549258 224440 549314 224496
rect 549902 224440 549958 224496
rect 549258 221756 549260 221776
rect 549260 221756 549312 221776
rect 549312 221756 549314 221776
rect 549258 221720 549314 221756
rect 552846 224476 552848 224496
rect 552848 224476 552900 224496
rect 552900 224476 552902 224496
rect 552846 224440 552902 224476
rect 554502 240352 554558 240408
rect 554318 238176 554374 238232
rect 554410 233824 554466 233880
rect 554778 224868 554834 224904
rect 554778 224848 554780 224868
rect 554780 224848 554832 224868
rect 554832 224848 554834 224868
rect 553950 221856 554006 221912
rect 557998 220496 558054 220552
rect 558550 221856 558606 221912
rect 558734 220496 558790 220552
rect 559378 221892 559380 221912
rect 559380 221892 559432 221912
rect 559432 221892 559434 221912
rect 559378 221856 559434 221892
rect 561678 224848 561734 224904
rect 562138 224748 562140 224768
rect 562140 224748 562192 224768
rect 562192 224748 562194 224768
rect 562138 224712 562194 224748
rect 563794 224712 563850 224768
rect 561494 221856 561550 221912
rect 560758 217504 560814 217560
rect 563794 221720 563850 221776
rect 562874 220496 562930 220552
rect 563334 220496 563390 220552
rect 562874 219156 562930 219192
rect 562874 219136 562876 219156
rect 562876 219136 562928 219156
rect 562928 219136 562930 219156
rect 563518 219156 563574 219192
rect 563518 219136 563520 219156
rect 563520 219136 563572 219156
rect 563572 219136 563574 219156
rect 563426 218864 563482 218920
rect 563058 218592 563114 218648
rect 562874 217776 562930 217832
rect 563150 217504 563206 217560
rect 565634 220632 565690 220688
rect 564162 218864 564218 218920
rect 564806 218864 564862 218920
rect 568302 217776 568358 217832
rect 569958 220652 570014 220688
rect 569958 220632 569960 220652
rect 569960 220632 570012 220652
rect 570012 220632 570014 220652
rect 572626 221720 572682 221776
rect 572258 220496 572314 220552
rect 572074 219156 572130 219192
rect 572074 219136 572076 219156
rect 572076 219136 572128 219156
rect 572128 219136 572130 219156
rect 572074 217776 572130 217832
rect 572258 217504 572314 217560
rect 572902 217504 572958 217560
rect 574190 217504 574246 217560
rect 53286 215056 53342 215112
rect 574558 219136 574614 219192
rect 574742 218884 574798 218920
rect 574742 218864 574744 218884
rect 574744 218864 574796 218884
rect 574796 218864 574798 218884
rect 574742 218592 574798 218648
rect 574926 217776 574982 217832
rect 575478 216688 575534 216744
rect 51906 179288 51962 179344
rect 578882 213968 578938 214024
rect 578514 211656 578570 211712
rect 579526 209788 579528 209808
rect 579528 209788 579580 209808
rect 579580 209788 579582 209808
rect 579526 209752 579582 209788
rect 579526 207440 579582 207496
rect 579526 205828 579582 205864
rect 579526 205808 579528 205828
rect 579528 205808 579580 205828
rect 579580 205808 579582 205828
rect 578330 203224 578386 203280
rect 578790 200776 578846 200832
rect 579526 198872 579582 198928
rect 578514 196424 578570 196480
rect 579526 194928 579582 194984
rect 579526 192208 579582 192264
rect 579526 190712 579582 190768
rect 579526 187992 579582 188048
rect 579526 186260 579528 186280
rect 579528 186260 579580 186280
rect 579580 186260 579582 186280
rect 579526 186224 579582 186260
rect 579526 184320 579582 184376
rect 579526 181872 579582 181928
rect 578790 180104 578846 180160
rect 579526 177656 579582 177712
rect 578790 175072 578846 175128
rect 578422 173440 578478 173496
rect 578238 170992 578294 171048
rect 578698 169224 578754 169280
rect 578238 166912 578294 166968
rect 579526 164464 579582 164520
rect 579342 162696 579398 162752
rect 578238 159840 578294 159896
rect 578422 158344 578478 158400
rect 578882 155896 578938 155952
rect 578330 153992 578386 154048
rect 578238 151680 578294 151736
rect 578882 149640 578938 149696
rect 579526 147464 579582 147520
rect 578606 140528 578662 140584
rect 578606 138760 578662 138816
rect 579250 144644 579252 144664
rect 579252 144644 579304 144664
rect 579304 144644 579306 144664
rect 579250 144608 579306 144644
rect 579526 142976 579582 143032
rect 578882 136584 578938 136640
rect 579526 134408 579582 134464
rect 579066 132232 579122 132288
rect 578882 129648 578938 129704
rect 579526 127880 579582 127936
rect 578330 125296 578386 125352
rect 578422 123564 578424 123584
rect 578424 123564 578476 123584
rect 578476 123564 578478 123584
rect 578422 123528 578478 123564
rect 578882 121352 578938 121408
rect 578514 118396 578516 118416
rect 578516 118396 578568 118416
rect 578568 118396 578570 118416
rect 578514 118360 578570 118396
rect 578330 108296 578386 108352
rect 578606 99220 578608 99240
rect 578608 99220 578660 99240
rect 578660 99220 578662 99240
rect 578606 99184 578662 99220
rect 578330 97416 578386 97472
rect 578514 93064 578570 93120
rect 579526 116900 579528 116920
rect 579528 116900 579580 116920
rect 579580 116900 579582 116920
rect 579526 116864 579582 116900
rect 579250 114452 579252 114472
rect 579252 114452 579304 114472
rect 579304 114452 579306 114472
rect 579250 114416 579306 114452
rect 579526 112512 579582 112568
rect 579342 110100 579344 110120
rect 579344 110100 579396 110120
rect 579396 110100 579398 110120
rect 579342 110064 579398 110100
rect 579066 105848 579122 105904
rect 579526 103264 579582 103320
rect 579526 101632 579582 101688
rect 579526 95004 579528 95024
rect 579528 95004 579580 95024
rect 579580 95004 579582 95024
rect 579526 94968 579582 95004
rect 579066 90888 579122 90944
rect 579526 88068 579528 88088
rect 579528 88068 579580 88088
rect 579580 88068 579582 88088
rect 579526 88032 579582 88068
rect 579342 86400 579398 86456
rect 579158 83952 579214 84008
rect 579066 82184 579122 82240
rect 578882 80008 578938 80064
rect 578238 75520 578294 75576
rect 579526 77832 579582 77888
rect 589462 207984 589518 208040
rect 589462 206352 589518 206408
rect 589462 204720 589518 204776
rect 589462 203088 589518 203144
rect 589462 201456 589518 201512
rect 589462 199824 589518 199880
rect 590382 198192 590438 198248
rect 589462 196560 589518 196616
rect 589278 194928 589334 194984
rect 589462 193296 589518 193352
rect 589462 191664 589518 191720
rect 590566 190032 590622 190088
rect 589646 188400 589702 188456
rect 589462 186768 589518 186824
rect 589462 185136 589518 185192
rect 589462 183504 589518 183560
rect 590566 181872 590622 181928
rect 589646 180240 589702 180296
rect 589462 178608 589518 178664
rect 589646 176976 589702 177032
rect 589462 175364 589518 175400
rect 589462 175344 589464 175364
rect 589464 175344 589516 175364
rect 589516 175344 589518 175364
rect 589462 173712 589518 173768
rect 589462 172080 589518 172136
rect 589646 170448 589702 170504
rect 589462 168816 589518 168872
rect 589462 167184 589518 167240
rect 589462 165552 589518 165608
rect 589462 163920 589518 163976
rect 589462 162288 589518 162344
rect 589462 160656 589518 160712
rect 589462 159024 589518 159080
rect 589278 157412 589334 157448
rect 589278 157392 589280 157412
rect 589280 157392 589332 157412
rect 589332 157392 589334 157412
rect 589462 155760 589518 155816
rect 589462 154128 589518 154184
rect 589462 152496 589518 152552
rect 590014 150864 590070 150920
rect 589462 149232 589518 149288
rect 588542 147600 588598 147656
rect 589462 145968 589518 146024
rect 589462 144336 589518 144392
rect 589830 142704 589886 142760
rect 589462 141072 589518 141128
rect 589462 139460 589518 139496
rect 589462 139440 589464 139460
rect 589464 139440 589516 139460
rect 589516 139440 589518 139460
rect 589462 137808 589518 137864
rect 589462 136176 589518 136232
rect 590382 134544 590438 134600
rect 589462 132912 589518 132968
rect 589462 131300 589518 131336
rect 589462 131280 589464 131300
rect 589464 131280 589516 131300
rect 589516 131280 589518 131300
rect 588542 129648 588598 129704
rect 581642 77832 581698 77888
rect 579066 73072 579122 73128
rect 576122 54984 576178 55040
rect 579066 71168 579122 71224
rect 580262 54712 580318 54768
rect 578882 54440 578938 54496
rect 589462 128016 589518 128072
rect 589922 126384 589978 126440
rect 589462 124752 589518 124808
rect 589462 123120 589518 123176
rect 590014 121488 590070 121544
rect 589646 119856 589702 119912
rect 589462 116592 589518 116648
rect 590106 118224 590162 118280
rect 589462 113328 589518 113384
rect 590290 114960 590346 115016
rect 589462 111696 589518 111752
rect 589278 110064 589334 110120
rect 589462 108432 589518 108488
rect 589830 106800 589886 106856
rect 589462 105168 589518 105224
rect 588726 103536 588782 103592
rect 589462 101904 589518 101960
rect 577502 54168 577558 54224
rect 459834 53624 459890 53680
rect 460754 53624 460810 53680
rect 461674 53624 461730 53680
rect 462594 53624 462650 53680
rect 463238 53644 463294 53680
rect 463238 53624 463240 53644
rect 463240 53624 463292 53644
rect 463292 53624 463294 53644
rect 464250 53624 464306 53680
rect 464066 53216 464122 53272
rect 476026 53644 476082 53680
rect 476026 53624 476028 53644
rect 476028 53624 476080 53644
rect 476080 53624 476082 53644
rect 476578 53644 476634 53680
rect 476578 53624 476580 53644
rect 476580 53624 476632 53644
rect 476632 53624 476634 53644
rect 464434 53216 464490 53272
rect 476210 53352 476266 53408
rect 477038 53352 477094 53408
rect 130842 44240 130898 44296
rect 458178 46960 458234 47016
rect 522946 47776 523002 47832
rect 458362 46688 458418 46744
rect 132774 44252 132776 44296
rect 132776 44252 132828 44296
rect 132828 44252 132830 44296
rect 132774 44240 132830 44252
rect 142618 44240 142674 44296
rect 255870 44104 255926 44160
rect 361762 43832 361818 43888
rect 440238 43852 440294 43888
rect 440238 43832 440240 43852
rect 440240 43832 440292 43852
rect 440292 43832 440294 43852
rect 441066 43852 441122 43888
rect 441066 43832 441068 43852
rect 441068 43832 441120 43852
rect 441120 43832 441122 43852
rect 415582 42336 415638 42392
rect 365074 41792 365130 41848
rect 416686 41792 416742 41848
rect 419906 41792 419962 41848
rect 446218 42200 446274 42256
rect 446218 41520 446274 41576
rect 460110 44104 460166 44160
rect 461030 44376 461086 44432
rect 460846 43424 460902 43480
rect 461766 42880 461822 42936
rect 462870 44376 462926 44432
rect 462686 43152 462742 43208
rect 463790 44376 463846 44432
rect 463974 42880 464030 42936
rect 465078 46960 465134 47016
rect 549994 48864 550050 48920
rect 599490 221448 599546 221504
rect 595166 217232 595222 217288
rect 595718 216960 595774 217016
rect 599030 215600 599086 215656
rect 600686 221176 600742 221232
rect 611634 220224 611690 220280
rect 612922 219680 612978 219736
rect 618258 220904 618314 220960
rect 617154 219952 617210 220008
rect 617798 215872 617854 215928
rect 618442 219408 618498 219464
rect 621110 215328 621166 215384
rect 623962 218048 624018 218104
rect 630678 218320 630734 218376
rect 667018 562264 667074 562320
rect 667570 594768 667626 594824
rect 652022 400832 652078 400888
rect 651470 373224 651526 373280
rect 652206 396616 652262 396672
rect 652206 373904 652262 373960
rect 652022 372136 652078 372192
rect 651470 370640 651526 370696
rect 652206 356632 652262 356688
rect 651470 328072 651526 328128
rect 651746 325644 651802 325680
rect 651746 325624 651748 325644
rect 651748 325624 651800 325644
rect 651800 325624 651802 325644
rect 651378 303356 651380 303376
rect 651380 303356 651432 303376
rect 651432 303356 651434 303376
rect 651378 303320 651434 303356
rect 651470 300600 651526 300656
rect 651470 298696 651526 298752
rect 651654 296812 651710 296848
rect 651654 296792 651656 296812
rect 651656 296792 651708 296812
rect 651708 296792 651710 296812
rect 652574 351056 652630 351112
rect 652574 329704 652630 329760
rect 652206 326848 652262 326904
rect 668398 689424 668454 689480
rect 668766 730088 668822 730144
rect 669410 728728 669466 728784
rect 669226 708736 669282 708792
rect 668858 593544 668914 593600
rect 669042 536424 669098 536480
rect 671250 733760 671306 733816
rect 670606 687656 670662 687712
rect 669778 685480 669834 685536
rect 669594 644272 669650 644328
rect 672078 732672 672134 732728
rect 671710 647808 671766 647864
rect 671342 638560 671398 638616
rect 671434 620744 671490 620800
rect 670422 549616 670478 549672
rect 669778 455368 669834 455424
rect 670974 607688 671030 607744
rect 670790 533840 670846 533896
rect 676034 896280 676090 896336
rect 675850 895464 675906 895520
rect 676034 894648 676090 894704
rect 675850 893832 675906 893888
rect 676034 893016 676090 893072
rect 673090 885400 673146 885456
rect 672906 777416 672962 777472
rect 672262 696904 672318 696960
rect 672078 652024 672134 652080
rect 676034 892608 676090 892664
rect 676034 891384 676090 891440
rect 675850 890976 675906 891032
rect 676034 890160 676090 890216
rect 676034 889344 676090 889400
rect 676034 888956 676090 888992
rect 676034 888936 676036 888956
rect 676036 888936 676088 888956
rect 676088 888936 676090 888956
rect 676034 888548 676090 888584
rect 676034 888528 676036 888548
rect 676036 888528 676088 888548
rect 676088 888528 676090 888548
rect 676034 887324 676090 887360
rect 676034 887304 676036 887324
rect 676036 887304 676088 887324
rect 676088 887304 676090 887324
rect 676034 886916 676090 886952
rect 676034 886896 676036 886916
rect 676036 886896 676088 886916
rect 676088 886896 676090 886916
rect 679622 891792 679678 891848
rect 678242 889752 678298 889808
rect 681002 890568 681058 890624
rect 683118 888120 683174 888176
rect 681002 880640 681058 880696
rect 683118 880368 683174 880424
rect 675942 878464 675998 878520
rect 675574 874112 675630 874168
rect 674930 873024 674986 873080
rect 675758 872752 675814 872808
rect 675298 865680 675354 865736
rect 675758 865408 675814 865464
rect 675666 864864 675722 864920
rect 675758 788024 675814 788080
rect 675114 786664 675170 786720
rect 675390 786664 675446 786720
rect 673642 780000 673698 780056
rect 673274 728320 673330 728376
rect 672998 728048 673054 728104
rect 675482 780000 675538 780056
rect 674470 779184 674526 779240
rect 674286 778776 674342 778832
rect 674102 734440 674158 734496
rect 672630 714856 672686 714912
rect 673274 714040 673330 714096
rect 673090 713632 673146 713688
rect 672814 711592 672870 711648
rect 672998 708328 673054 708384
rect 672814 686160 672870 686216
rect 672630 670112 672686 670168
rect 672170 625540 672172 625560
rect 672172 625540 672224 625560
rect 672224 625540 672226 625560
rect 672170 625504 672226 625540
rect 671986 622784 672042 622840
rect 672630 649168 672686 649224
rect 672998 685752 673054 685808
rect 674930 777008 674986 777064
rect 674930 775668 674986 775704
rect 674930 775648 674932 775668
rect 674932 775648 674984 775668
rect 674984 775648 674986 775668
rect 675482 779184 675538 779240
rect 675482 778776 675538 778832
rect 675390 777416 675446 777472
rect 675482 777008 675538 777064
rect 675390 775648 675446 775704
rect 675298 742464 675354 742520
rect 674654 734984 674710 735040
rect 675298 738112 675354 738168
rect 675390 734984 675446 735040
rect 675390 734440 675446 734496
rect 675482 733760 675538 733816
rect 675482 732672 675538 732728
rect 674654 729816 674710 729872
rect 675114 730088 675170 730144
rect 675298 730088 675354 730144
rect 673826 724104 673882 724160
rect 674286 724104 674342 724160
rect 674930 723152 674986 723208
rect 675482 728728 675538 728784
rect 674010 715708 674012 715728
rect 674012 715708 674064 715728
rect 674064 715708 674066 715728
rect 674010 715672 674066 715708
rect 674010 714484 674012 714504
rect 674012 714484 674064 714504
rect 674064 714484 674066 714504
rect 674010 714448 674066 714484
rect 674010 713244 674066 713280
rect 674010 713224 674012 713244
rect 674012 713224 674064 713244
rect 674064 713224 674066 713244
rect 674010 712852 674012 712872
rect 674012 712852 674064 712872
rect 674064 712852 674066 712872
rect 674010 712816 674066 712852
rect 674010 712428 674066 712464
rect 674010 712408 674012 712428
rect 674012 712408 674064 712428
rect 674064 712408 674066 712428
rect 674010 709996 674012 710016
rect 674012 709996 674064 710016
rect 674064 709996 674066 710016
rect 674010 709960 674066 709996
rect 673826 709280 673882 709336
rect 674010 709180 674012 709200
rect 674012 709180 674064 709200
rect 674064 709180 674066 709200
rect 674010 709144 674066 709180
rect 676034 716508 676090 716544
rect 676034 716488 676036 716508
rect 676036 716488 676088 716508
rect 676088 716488 676090 716508
rect 676034 716080 676090 716136
rect 675850 715264 675906 715320
rect 675298 712000 675354 712056
rect 682382 726552 682438 726608
rect 683302 726280 683358 726336
rect 682382 711184 682438 711240
rect 681002 710776 681058 710832
rect 676034 710368 676090 710424
rect 683302 709552 683358 709608
rect 676034 707548 676036 707568
rect 676036 707548 676088 707568
rect 676088 707548 676090 707568
rect 676034 707512 676090 707548
rect 674010 707104 674066 707160
rect 673826 706968 673882 707024
rect 684130 707920 684186 707976
rect 683486 706696 683542 706752
rect 676034 706288 676090 706344
rect 683118 705472 683174 705528
rect 676034 705064 676090 705120
rect 675298 696904 675354 696960
rect 675482 696768 675538 696824
rect 675114 694592 675170 694648
rect 673642 682760 673698 682816
rect 674010 690124 674066 690160
rect 674010 690104 674012 690124
rect 674012 690104 674064 690124
rect 674064 690104 674066 690124
rect 674010 688780 674012 688800
rect 674012 688780 674064 688800
rect 674064 688780 674066 688800
rect 674010 688744 674066 688780
rect 674930 690104 674986 690160
rect 675114 689424 675170 689480
rect 673734 681944 673790 682000
rect 673182 669840 673238 669896
rect 673366 669160 673422 669216
rect 673366 663992 673422 664048
rect 673366 662904 673422 662960
rect 673734 671356 673790 671392
rect 673734 671336 673736 671356
rect 673736 671336 673788 671356
rect 673788 671336 673790 671356
rect 673734 670928 673790 670984
rect 673734 670520 673790 670576
rect 673734 668888 673790 668944
rect 673734 668516 673736 668536
rect 673736 668516 673788 668536
rect 673788 668516 673790 668536
rect 673734 668480 673790 668516
rect 673734 668072 673790 668128
rect 673734 667664 673790 667720
rect 673734 666848 673790 666904
rect 673734 666596 673790 666632
rect 673734 666576 673736 666596
rect 673736 666576 673788 666596
rect 673788 666576 673790 666596
rect 673734 665252 673736 665272
rect 673736 665252 673788 665272
rect 673788 665252 673790 665272
rect 673734 665216 673790 665252
rect 673734 664420 673790 664456
rect 673734 664400 673736 664420
rect 673736 664400 673788 664420
rect 673788 664400 673790 664420
rect 673734 663720 673790 663776
rect 673550 661952 673606 662008
rect 673734 661580 673736 661600
rect 673736 661580 673788 661600
rect 673788 661580 673790 661600
rect 673734 661544 673790 661580
rect 673734 661156 673790 661192
rect 673734 661136 673736 661156
rect 673736 661136 673788 661156
rect 673788 661136 673790 661156
rect 673734 660084 673736 660104
rect 673736 660084 673788 660104
rect 673788 660084 673790 660104
rect 673734 660048 673790 660084
rect 673366 659640 673422 659696
rect 672998 648760 673054 648816
rect 673182 645224 673238 645280
rect 672814 626320 672870 626376
rect 672814 625912 672870 625968
rect 672814 624996 672816 625016
rect 672816 624996 672868 625016
rect 672868 624996 672870 625016
rect 672814 624960 672870 624996
rect 672814 624708 672870 624744
rect 672814 624688 672816 624708
rect 672816 624688 672868 624708
rect 672868 624688 672870 624708
rect 672814 624316 672816 624336
rect 672816 624316 672868 624336
rect 672868 624316 672870 624336
rect 672814 624280 672870 624316
rect 672814 623892 672870 623928
rect 672814 623872 672816 623892
rect 672816 623872 672868 623892
rect 672868 623872 672870 623892
rect 672814 623500 672816 623520
rect 672816 623500 672868 623520
rect 672868 623500 672870 623520
rect 672814 623464 672870 623500
rect 672814 623076 672870 623112
rect 672814 623056 672816 623076
rect 672816 623056 672868 623076
rect 672868 623056 672870 623076
rect 672906 621424 672962 621480
rect 672814 621052 672816 621072
rect 672816 621052 672868 621072
rect 672868 621052 672870 621072
rect 672814 621016 672870 621052
rect 672262 618432 672318 618488
rect 672446 604424 672502 604480
rect 672814 620236 672816 620256
rect 672816 620236 672868 620256
rect 672868 620236 672870 620256
rect 672814 620200 672870 620236
rect 672814 619964 672816 619984
rect 672816 619964 672868 619984
rect 672868 619964 672870 619984
rect 672814 619928 672870 619964
rect 672814 619692 672816 619712
rect 672816 619692 672868 619712
rect 672868 619692 672870 619712
rect 672814 619656 672870 619692
rect 672814 597352 672870 597408
rect 673734 655580 673790 655616
rect 673734 655560 673736 655580
rect 673736 655560 673788 655580
rect 673788 655560 673790 655580
rect 673734 645924 673790 645960
rect 673734 645904 673736 645924
rect 673736 645904 673788 645924
rect 673788 645904 673790 645924
rect 673550 643456 673606 643512
rect 673734 643084 673736 643104
rect 673736 643084 673788 643104
rect 673788 643084 673790 643104
rect 673734 643048 673790 643084
rect 673550 642368 673606 642424
rect 674102 644544 674158 644600
rect 674102 642368 674158 642424
rect 674102 641688 674158 641744
rect 674930 688744 674986 688800
rect 675114 687656 675170 687712
rect 675114 686160 675170 686216
rect 674930 685752 674986 685808
rect 675114 685480 675170 685536
rect 675114 683984 675170 684040
rect 674838 682760 674894 682816
rect 674838 681944 674894 682000
rect 675298 683712 675354 683768
rect 675114 676368 675170 676424
rect 674838 669860 674894 669896
rect 674838 669840 674840 669860
rect 674840 669840 674892 669860
rect 674892 669840 674894 669860
rect 676494 669432 676550 669488
rect 675298 666440 675354 666496
rect 676034 664808 676090 664864
rect 674838 663756 674840 663776
rect 674840 663756 674892 663776
rect 674892 663756 674894 663776
rect 674838 663720 674894 663756
rect 683210 663720 683266 663776
rect 684130 682352 684186 682408
rect 684130 666168 684186 666224
rect 683486 662904 683542 662960
rect 674838 660048 674894 660104
rect 683118 660048 683174 660104
rect 675114 655560 675170 655616
rect 675390 652840 675446 652896
rect 675482 652024 675538 652080
rect 675390 649168 675446 649224
rect 675114 648760 675170 648816
rect 675390 647808 675446 647864
rect 675114 645904 675170 645960
rect 675298 645224 675354 645280
rect 675298 644544 675354 644600
rect 675390 644272 675446 644328
rect 675298 643456 675354 643512
rect 675298 643048 675354 643104
rect 675298 641688 675354 641744
rect 674286 620744 674342 620800
rect 674378 619692 674380 619712
rect 674380 619692 674432 619712
rect 674432 619692 674434 619712
rect 674378 619656 674434 619692
rect 674286 618468 674288 618488
rect 674288 618468 674340 618488
rect 674340 618468 674342 618488
rect 674286 618432 674342 618468
rect 673090 580624 673146 580680
rect 672998 574912 673054 574968
rect 673090 573688 673146 573744
rect 672906 573416 672962 573472
rect 671158 532072 671214 532128
rect 670606 455096 670662 455152
rect 663062 403280 663118 403336
rect 654782 382880 654838 382936
rect 670514 392536 670570 392592
rect 666466 365608 666522 365664
rect 654782 358536 654838 358592
rect 653586 338680 653642 338736
rect 669410 347248 669466 347304
rect 653402 313248 653458 313304
rect 652482 309848 652538 309904
rect 658922 311888 658978 311944
rect 652482 302096 652538 302152
rect 652298 297472 652354 297528
rect 651470 294208 651526 294264
rect 651470 292984 651526 293040
rect 651930 295296 651986 295352
rect 651930 291760 651986 291816
rect 652114 291488 652170 291544
rect 651470 290400 651526 290456
rect 651654 289176 651710 289232
rect 651470 288632 651526 288688
rect 651654 287680 651710 287736
rect 651470 287408 651526 287464
rect 651470 285912 651526 285968
rect 651470 284688 651526 284744
rect 651470 283328 651526 283384
rect 652022 282104 652078 282160
rect 651470 280880 651526 280936
rect 650642 224984 650698 225040
rect 645858 219816 645914 219872
rect 648434 218592 648490 218648
rect 651102 217776 651158 217832
rect 651470 221448 651526 221504
rect 652390 280336 652446 280392
rect 652574 279384 652630 279440
rect 660578 293800 660634 293856
rect 658922 268096 658978 268152
rect 664442 248240 664498 248296
rect 652390 226888 652446 226944
rect 658922 226344 658978 226400
rect 652758 225664 652814 225720
rect 656162 225256 656218 225312
rect 654782 223896 654838 223952
rect 653402 222808 653458 222864
rect 654138 220360 654194 220416
rect 653770 217504 653826 217560
rect 657542 223624 657598 223680
rect 656806 218864 656862 218920
rect 660762 221720 660818 221776
rect 659566 215328 659622 215384
rect 658738 213152 658794 213208
rect 660394 214512 660450 214568
rect 662142 228520 662198 228576
rect 661498 213424 661554 213480
rect 664902 230424 664958 230480
rect 663706 229064 663762 229120
rect 664626 215600 664682 215656
rect 667018 225936 667074 225992
rect 667018 225256 667074 225312
rect 665822 222808 665878 222864
rect 666650 219408 666706 219464
rect 666834 215328 666890 215384
rect 666834 198464 666890 198520
rect 666742 174936 666798 174992
rect 667202 134544 667258 134600
rect 668030 199144 668086 199200
rect 668766 232872 668822 232928
rect 668582 221448 668638 221504
rect 668398 215600 668454 215656
rect 668398 198736 668454 198792
rect 668214 184456 668270 184512
rect 667754 181328 667810 181384
rect 667570 180240 667626 180296
rect 668214 177964 668216 177984
rect 668216 177964 668268 177984
rect 668268 177964 668270 177984
rect 668214 177928 668270 177964
rect 668030 174664 668086 174720
rect 667938 169668 667940 169688
rect 667940 169668 667992 169688
rect 667992 169668 667994 169688
rect 667938 169632 667994 169668
rect 667938 164872 667994 164928
rect 668214 160012 668216 160032
rect 668216 160012 668268 160032
rect 668268 160012 668270 160032
rect 668214 159976 668270 160012
rect 668214 155080 668270 155136
rect 668398 143656 668454 143712
rect 669226 220360 669282 220416
rect 669870 301960 669926 302016
rect 670330 262112 670386 262168
rect 670146 258440 670202 258496
rect 670330 237224 670386 237280
rect 669686 223896 669742 223952
rect 669318 220088 669374 220144
rect 669778 222264 669834 222320
rect 669318 218184 669374 218240
rect 669226 216960 669282 217016
rect 669594 213832 669650 213888
rect 669594 202816 669650 202872
rect 669318 194248 669374 194304
rect 669134 191528 669190 191584
rect 668950 189352 669006 189408
rect 669134 188400 669190 188456
rect 668766 163240 668822 163296
rect 668766 156168 668822 156224
rect 668766 148552 668822 148608
rect 668766 145288 668822 145344
rect 668582 138760 668638 138816
rect 668766 135088 668822 135144
rect 667938 133764 667940 133784
rect 667940 133764 667992 133784
rect 667992 133764 667994 133784
rect 667938 133728 667994 133764
rect 667386 133456 667442 133512
rect 667018 132640 667074 132696
rect 668582 130600 668638 130656
rect 668030 128968 668086 129024
rect 668582 127744 668638 127800
rect 667938 107752 667994 107808
rect 668398 106156 668400 106176
rect 668400 106156 668452 106176
rect 668452 106156 668454 106176
rect 668398 106120 668454 106156
rect 669502 172352 669558 172408
rect 669318 162832 669374 162888
rect 669318 158344 669374 158400
rect 669594 150320 669650 150376
rect 669134 135496 669190 135552
rect 670974 295840 671030 295896
rect 670974 293800 671030 293856
rect 671802 559544 671858 559600
rect 671618 532752 671674 532808
rect 672262 555192 672318 555248
rect 672630 535916 672632 535936
rect 672632 535916 672684 535936
rect 672684 535916 672686 535936
rect 672630 535880 672686 535916
rect 672630 535644 672632 535664
rect 672632 535644 672684 535664
rect 672684 535644 672686 535664
rect 672630 535608 672686 535644
rect 672630 534828 672632 534848
rect 672632 534828 672684 534848
rect 672684 534828 672686 534848
rect 672630 534792 672686 534828
rect 672630 534556 672632 534576
rect 672632 534556 672684 534576
rect 672684 534556 672686 534576
rect 672630 534520 672686 534556
rect 672630 534268 672686 534304
rect 672630 534248 672632 534268
rect 672632 534248 672684 534268
rect 672684 534248 672686 534268
rect 673090 560224 673146 560280
rect 672630 533568 672686 533624
rect 672446 533332 672448 533352
rect 672448 533332 672500 533352
rect 672500 533332 672502 533352
rect 672446 533296 672502 533332
rect 672446 532516 672448 532536
rect 672448 532516 672500 532536
rect 672500 532516 672502 532536
rect 672446 532480 672502 532516
rect 672262 453908 672264 453928
rect 672264 453908 672316 453928
rect 672316 453908 672318 453928
rect 672262 453872 672318 453908
rect 672814 528808 672870 528864
rect 672906 527992 672962 528048
rect 672446 402056 672502 402112
rect 675482 638560 675538 638616
rect 681002 637472 681058 637528
rect 675482 631352 675538 631408
rect 675666 631352 675722 631408
rect 676218 621968 676274 622024
rect 681002 621968 681058 622024
rect 676034 620608 676090 620664
rect 676218 619112 676274 619168
rect 683210 618704 683266 618760
rect 676218 617908 676274 617944
rect 676218 617888 676220 617908
rect 676220 617888 676272 617908
rect 676272 617888 676274 617908
rect 676218 617500 676274 617536
rect 676218 617480 676220 617500
rect 676220 617480 676272 617500
rect 676272 617480 676274 617500
rect 676494 617480 676550 617536
rect 675298 617072 675354 617128
rect 683578 617072 683634 617128
rect 683394 616664 683450 616720
rect 683118 615476 683120 615496
rect 683120 615476 683172 615496
rect 683172 615476 683174 615496
rect 674010 607960 674066 608016
rect 674010 600364 674066 600400
rect 674010 600344 674012 600364
rect 674012 600344 674064 600364
rect 674064 600344 674066 600364
rect 674010 599664 674066 599720
rect 673550 596808 673606 596864
rect 674010 598032 674066 598088
rect 673918 597080 673974 597136
rect 673642 581304 673698 581360
rect 673642 581052 673698 581088
rect 673642 581032 673644 581052
rect 673644 581032 673696 581052
rect 673696 581032 673698 581052
rect 673642 580252 673644 580272
rect 673644 580252 673696 580272
rect 673696 580252 673698 580272
rect 673642 580216 673698 580252
rect 673642 579844 673644 579864
rect 673644 579844 673696 579864
rect 673696 579844 673698 579864
rect 673642 579808 673698 579844
rect 673642 579420 673698 579456
rect 673642 579400 673644 579420
rect 673644 579400 673696 579420
rect 673696 579400 673698 579420
rect 673642 579028 673644 579048
rect 673644 579028 673696 579048
rect 673696 579028 673698 579048
rect 673642 578992 673698 579028
rect 673642 578604 673698 578640
rect 673642 578584 673644 578604
rect 673644 578584 673696 578604
rect 673696 578584 673698 578604
rect 673642 578196 673698 578232
rect 673642 578176 673644 578196
rect 673644 578176 673696 578196
rect 673696 578176 673698 578196
rect 673642 577788 673698 577824
rect 673642 577768 673644 577788
rect 673644 577768 673696 577788
rect 673696 577768 673698 577788
rect 673642 577396 673644 577416
rect 673644 577396 673696 577416
rect 673696 577396 673698 577416
rect 673642 577360 673698 577396
rect 673642 576972 673698 577008
rect 673642 576952 673644 576972
rect 673644 576952 673696 576972
rect 673696 576952 673698 576972
rect 673642 574540 673644 574560
rect 673644 574540 673696 574560
rect 673696 574540 673698 574560
rect 673642 574504 673698 574540
rect 673642 574132 673644 574152
rect 673644 574132 673696 574152
rect 673696 574132 673698 574152
rect 673642 574096 673698 574132
rect 673642 572464 673698 572520
rect 673642 572056 673698 572112
rect 673642 570832 673698 570888
rect 673642 569916 673644 569936
rect 673644 569916 673696 569936
rect 673696 569916 673698 569936
rect 673642 569880 673698 569916
rect 673642 569608 673698 569664
rect 673642 565836 673644 565856
rect 673644 565836 673696 565856
rect 673696 565836 673698 565856
rect 673642 565800 673698 565836
rect 673642 564596 673698 564632
rect 673642 564576 673644 564596
rect 673644 564576 673696 564596
rect 673696 564576 673698 564596
rect 673642 554804 673698 554840
rect 673642 554784 673644 554804
rect 673644 554784 673696 554804
rect 673696 554784 673698 554804
rect 673642 553444 673698 553480
rect 673642 553424 673644 553444
rect 673644 553424 673696 553444
rect 673696 553424 673698 553444
rect 673642 553152 673698 553208
rect 673090 484744 673146 484800
rect 674102 558320 674158 558376
rect 674470 597080 674526 597136
rect 674470 596808 674526 596864
rect 683118 615440 683174 615476
rect 676218 614644 676274 614680
rect 676218 614624 676220 614644
rect 676220 614624 676272 614644
rect 676272 614624 676274 614644
rect 675390 607960 675446 608016
rect 675482 607688 675538 607744
rect 675114 604424 675170 604480
rect 675114 602928 675170 602984
rect 675390 600888 675446 600944
rect 675114 600344 675170 600400
rect 675482 599664 675538 599720
rect 675114 598032 675170 598088
rect 674470 581304 674526 581360
rect 675390 597352 675446 597408
rect 675482 594768 675538 594824
rect 675482 593544 675538 593600
rect 675482 593136 675538 593192
rect 674838 569880 674894 569936
rect 675206 586200 675262 586256
rect 681002 591640 681058 591696
rect 682382 576408 682438 576464
rect 681002 575592 681058 575648
rect 684222 591232 684278 591288
rect 683394 573144 683450 573200
rect 684222 576000 684278 576056
rect 684038 571920 684094 571976
rect 676218 571548 676220 571568
rect 676220 571548 676272 571568
rect 676272 571548 676274 571568
rect 676218 571512 676274 571548
rect 683118 570288 683174 570344
rect 675390 565800 675446 565856
rect 675114 564576 675170 564632
rect 675114 562264 675170 562320
rect 675390 561856 675446 561912
rect 675206 559544 675262 559600
rect 675574 559408 675630 559464
rect 675482 558320 675538 558376
rect 675298 557504 675354 557560
rect 675390 555192 675446 555248
rect 675298 554784 675354 554840
rect 674654 551928 674710 551984
rect 674010 548800 674066 548856
rect 673826 536152 673882 536208
rect 674194 536152 674250 536208
rect 674286 533840 674342 533896
rect 673826 492088 673882 492144
rect 674010 490900 674012 490920
rect 674012 490900 674064 490920
rect 674064 490900 674066 490920
rect 674010 490864 674066 490900
rect 674010 490476 674066 490512
rect 674010 490456 674012 490476
rect 674012 490456 674064 490476
rect 674064 490456 674066 490476
rect 674010 490084 674012 490104
rect 674012 490084 674064 490104
rect 674064 490084 674066 490104
rect 674010 490048 674066 490084
rect 674010 489660 674066 489696
rect 674010 489640 674012 489660
rect 674012 489640 674064 489660
rect 674064 489640 674066 489660
rect 674010 489268 674012 489288
rect 674012 489268 674064 489288
rect 674064 489268 674066 489288
rect 674010 489232 674066 489268
rect 674010 488452 674012 488472
rect 674012 488452 674064 488472
rect 674064 488452 674066 488472
rect 674010 488416 674066 488452
rect 673826 486004 673828 486024
rect 673828 486004 673880 486024
rect 673880 486004 673882 486024
rect 673826 485968 673882 486004
rect 675758 553832 675814 553888
rect 675574 553424 675630 553480
rect 675390 551928 675446 551984
rect 675390 551520 675446 551576
rect 675482 550160 675538 550216
rect 675022 549888 675078 549944
rect 674838 545808 674894 545864
rect 675482 549616 675538 549672
rect 675758 548256 675814 548312
rect 675574 547848 675630 547904
rect 677414 547576 677470 547632
rect 675482 536424 675538 536480
rect 676034 534452 676090 534508
rect 676218 531800 676274 531856
rect 676034 530816 676036 530836
rect 676036 530816 676088 530836
rect 676088 530816 676090 530836
rect 676034 530780 676090 530816
rect 676034 529984 676090 530020
rect 676034 529964 676036 529984
rect 676036 529964 676088 529984
rect 676088 529964 676090 529984
rect 676218 529352 676274 529408
rect 676034 529184 676036 529204
rect 676036 529184 676088 529204
rect 676088 529184 676090 529204
rect 676034 529148 676090 529184
rect 676034 526736 676036 526756
rect 676036 526736 676088 526756
rect 676088 526736 676090 526756
rect 676034 526700 676090 526736
rect 676034 526328 676036 526348
rect 676036 526328 676088 526348
rect 676088 526328 676090 526348
rect 676034 526292 676090 526328
rect 674654 484336 674710 484392
rect 674010 483148 674012 483168
rect 674012 483148 674064 483168
rect 674064 483148 674066 483168
rect 674010 483112 674066 483148
rect 673642 482296 673698 482352
rect 673274 455388 673330 455424
rect 673274 455368 673276 455388
rect 673276 455368 673328 455388
rect 673328 455368 673330 455388
rect 673386 455252 673442 455288
rect 673386 455232 673388 455252
rect 673388 455232 673440 455252
rect 673440 455232 673442 455252
rect 673274 455096 673330 455152
rect 672814 454824 672870 454880
rect 674286 454860 674288 454880
rect 674288 454860 674340 454880
rect 674340 454860 674342 454880
rect 674286 454824 674342 454860
rect 673044 454588 673046 454608
rect 673046 454588 673098 454608
rect 673098 454588 673100 454608
rect 673044 454552 673100 454588
rect 674286 454588 674288 454608
rect 674288 454588 674340 454608
rect 674340 454588 674342 454608
rect 674286 454552 674342 454588
rect 676034 491700 676090 491736
rect 676034 491680 676036 491700
rect 676036 491680 676088 491700
rect 676088 491680 676090 491700
rect 675850 491272 675906 491328
rect 676034 486784 676090 486840
rect 676034 485172 676090 485208
rect 676034 485152 676036 485172
rect 676036 485152 676088 485172
rect 676088 485152 676090 485172
rect 676034 483964 676036 483984
rect 676036 483964 676088 483984
rect 676088 483964 676090 483984
rect 676034 483928 676090 483964
rect 681002 546760 681058 546816
rect 682382 531392 682438 531448
rect 681002 530576 681058 530632
rect 683394 547032 683450 547088
rect 683210 527720 683266 527776
rect 683578 528536 683634 528592
rect 683394 527312 683450 527368
rect 677874 525680 677930 525736
rect 683118 524864 683174 524920
rect 678978 524456 679034 524512
rect 683394 503648 683450 503704
rect 679622 487192 679678 487248
rect 683210 500928 683266 500984
rect 681186 487600 681242 487656
rect 681002 486376 681058 486432
rect 683394 485560 683450 485616
rect 683210 483520 683266 483576
rect 676034 482704 676090 482760
rect 680358 481888 680414 481944
rect 675850 480664 675906 480720
rect 683118 481072 683174 481128
rect 672952 454316 672954 454336
rect 672954 454316 673006 454336
rect 673006 454316 673008 454336
rect 672952 454280 673008 454316
rect 674286 454316 674288 454336
rect 674288 454316 674340 454336
rect 674340 454316 674342 454336
rect 674286 454280 674342 454316
rect 674286 453908 674288 453928
rect 674288 453908 674340 453928
rect 674340 453908 674342 453928
rect 674286 453872 674342 453908
rect 676218 403300 676274 403336
rect 676218 403280 676220 403300
rect 676220 403280 676272 403300
rect 676272 403280 676274 403300
rect 673182 402328 673238 402384
rect 672630 401648 672686 401704
rect 672170 399608 672226 399664
rect 671894 393488 671950 393544
rect 671710 348880 671766 348936
rect 671710 331200 671766 331256
rect 671526 302232 671582 302288
rect 671342 260480 671398 260536
rect 670698 257216 670754 257272
rect 670514 224440 670570 224496
rect 670514 223624 670570 223680
rect 670514 222808 670570 222864
rect 670514 218864 670570 218920
rect 670514 216688 670570 216744
rect 670514 198192 670570 198248
rect 671342 240216 671398 240272
rect 670790 177964 670792 177984
rect 670792 177964 670844 177984
rect 670844 177964 670846 177984
rect 670790 177928 670846 177964
rect 670422 171128 670478 171184
rect 669962 130872 670018 130928
rect 668950 125704 669006 125760
rect 668766 119176 668822 119232
rect 669226 118768 669282 118824
rect 669226 114280 669282 114336
rect 668766 112648 668822 112704
rect 670606 170176 670662 170232
rect 670422 155896 670478 155952
rect 671710 278468 671712 278488
rect 671712 278468 671764 278488
rect 671764 278468 671766 278488
rect 671710 278432 671766 278468
rect 671710 259664 671766 259720
rect 671710 245520 671766 245576
rect 672998 394712 673054 394768
rect 672814 393896 672870 393952
rect 672998 380976 673054 381032
rect 672814 376216 672870 376272
rect 673918 401376 673974 401432
rect 673366 400424 673422 400480
rect 673182 357448 673238 357504
rect 672354 357040 672410 357096
rect 672170 355000 672226 355056
rect 672170 353368 672226 353424
rect 672170 337728 672226 337784
rect 672538 356224 672594 356280
rect 672354 312432 672410 312488
rect 673734 396072 673790 396128
rect 673734 381384 673790 381440
rect 676586 402872 676642 402928
rect 674838 402600 674894 402656
rect 674838 402056 674894 402112
rect 676586 400832 676642 400888
rect 676034 399336 676090 399392
rect 674746 397296 674802 397352
rect 674562 396616 674618 396672
rect 679622 398384 679678 398440
rect 676218 397976 676274 398032
rect 678242 397568 678298 397624
rect 676218 395548 676274 395584
rect 676218 395528 676220 395548
rect 676220 395528 676272 395548
rect 676272 395528 676274 395548
rect 676218 394324 676274 394360
rect 676218 394304 676220 394324
rect 676220 394304 676272 394324
rect 676272 394304 676274 394324
rect 678242 387640 678298 387696
rect 675758 384920 675814 384976
rect 675206 382880 675262 382936
rect 675758 382200 675814 382256
rect 675114 381384 675170 381440
rect 675390 380976 675446 381032
rect 675758 378664 675814 378720
rect 675758 377304 675814 377360
rect 675390 376216 675446 376272
rect 675758 373632 675814 373688
rect 675390 372408 675446 372464
rect 674470 358264 674526 358320
rect 673918 356496 673974 356552
rect 673366 355816 673422 355872
rect 673182 355408 673238 355464
rect 672998 349696 673054 349752
rect 672722 348472 672778 348528
rect 672538 311616 672594 311672
rect 672538 305496 672594 305552
rect 672538 285504 672594 285560
rect 672170 246064 672226 246120
rect 671802 236680 671858 236736
rect 672998 335552 673054 335608
rect 672906 324944 672962 325000
rect 673918 354592 673974 354648
rect 673734 352552 673790 352608
rect 673366 350104 673422 350160
rect 673550 349288 673606 349344
rect 673366 335824 673422 335880
rect 673734 333920 673790 333976
rect 673550 332696 673606 332752
rect 673182 310800 673238 310856
rect 674286 351328 674342 351384
rect 675942 357856 675998 357912
rect 675942 356768 675998 356824
rect 674654 352144 674710 352200
rect 674470 351056 674526 351112
rect 674470 350512 674526 350568
rect 674286 338000 674342 338056
rect 676034 350920 676090 350976
rect 676034 346568 676090 346624
rect 675758 340176 675814 340232
rect 675114 338680 675170 338736
rect 675114 338000 675170 338056
rect 675482 339360 675538 339416
rect 675758 337864 675814 337920
rect 675298 337728 675354 337784
rect 675758 336504 675814 336560
rect 674930 335824 674986 335880
rect 675114 335552 675170 335608
rect 675114 333920 675170 333976
rect 675114 332696 675170 332752
rect 675114 331200 675170 331256
rect 675022 327936 675078 327992
rect 674654 326848 674710 326904
rect 675390 327936 675446 327992
rect 675390 326848 675446 326904
rect 675206 325624 675262 325680
rect 675022 324944 675078 325000
rect 676218 313928 676274 313984
rect 674838 312840 674894 312896
rect 675482 312044 675538 312080
rect 675482 312024 675484 312044
rect 675484 312024 675536 312044
rect 675536 312024 675538 312044
rect 674838 311888 674894 311944
rect 673918 309984 673974 310040
rect 673274 309440 673330 309496
rect 673090 304272 673146 304328
rect 673090 287816 673146 287872
rect 672814 278432 672870 278488
rect 672538 265240 672594 265296
rect 673090 266056 673146 266112
rect 673826 305904 673882 305960
rect 674010 291760 674066 291816
rect 673826 291488 673882 291544
rect 673458 287544 673514 287600
rect 673274 264968 673330 265024
rect 673090 263336 673146 263392
rect 672906 259256 672962 259312
rect 673090 250688 673146 250744
rect 673090 249600 673146 249656
rect 673090 245792 673146 245848
rect 672906 242664 672962 242720
rect 674746 311208 674802 311264
rect 674562 310392 674618 310448
rect 674378 303864 674434 303920
rect 675942 309712 675998 309768
rect 675114 308352 675170 308408
rect 674930 306312 674986 306368
rect 675298 307944 675354 308000
rect 676034 307536 676090 307592
rect 676034 307128 676090 307184
rect 678242 306720 678298 306776
rect 676586 304680 676642 304736
rect 676034 303456 676090 303512
rect 676034 301960 676090 302016
rect 676586 301552 676642 301608
rect 675022 297608 675078 297664
rect 675482 298152 675538 298208
rect 676862 297336 676918 297392
rect 675390 295840 675446 295896
rect 675574 295704 675630 295760
rect 674838 292440 674894 292496
rect 675758 294616 675814 294672
rect 675390 291488 675446 291544
rect 675758 290944 675814 291000
rect 675114 287816 675170 287872
rect 674010 268096 674066 268152
rect 674378 267416 674434 267472
rect 673918 267008 673974 267064
rect 673734 264560 673790 264616
rect 673458 246200 673514 246256
rect 673734 241984 673790 242040
rect 673274 241712 673330 241768
rect 675758 287000 675814 287056
rect 675114 285504 675170 285560
rect 675758 283600 675814 283656
rect 675758 282648 675814 282704
rect 675666 281560 675722 281616
rect 676862 279384 676918 279440
rect 675298 278704 675354 278760
rect 675482 278024 675538 278080
rect 674746 266600 674802 266656
rect 674562 265784 674618 265840
rect 674654 262520 674710 262576
rect 674102 260888 674158 260944
rect 674286 260072 674342 260128
rect 674102 246608 674158 246664
rect 674470 258848 674526 258904
rect 674286 242256 674342 242312
rect 676862 268504 676918 268560
rect 676218 268096 676274 268152
rect 676218 267688 676274 267744
rect 676402 264016 676458 264072
rect 676218 262792 676274 262848
rect 675482 258032 675538 258088
rect 679622 263608 679678 263664
rect 674930 253136 674986 253192
rect 674930 248784 674986 248840
rect 675850 253156 675906 253192
rect 675850 253136 675852 253156
rect 675852 253136 675904 253156
rect 675904 253136 675906 253156
rect 675482 250688 675538 250744
rect 675758 250280 675814 250336
rect 675390 248240 675446 248296
rect 675298 246608 675354 246664
rect 675758 246608 675814 246664
rect 674838 241712 674894 241768
rect 674470 241440 674526 241496
rect 672952 236700 673008 236736
rect 672952 236680 672954 236700
rect 672954 236680 673006 236700
rect 673006 236680 673008 236700
rect 674194 236680 674250 236736
rect 672354 227024 672410 227080
rect 672814 232872 672870 232928
rect 671986 225664 672042 225720
rect 672170 225664 672226 225720
rect 672722 226380 672724 226400
rect 672724 226380 672776 226400
rect 672776 226380 672778 226400
rect 672722 226344 672778 226380
rect 672602 226108 672604 226128
rect 672604 226108 672656 226128
rect 672656 226108 672658 226128
rect 672602 226072 672658 226108
rect 672492 225956 672548 225992
rect 672492 225936 672494 225956
rect 672494 225936 672546 225956
rect 672546 225936 672548 225956
rect 672262 225256 672318 225312
rect 672170 224984 672226 225040
rect 671618 224712 671674 224768
rect 671480 224440 671536 224496
rect 671594 224168 671650 224224
rect 671618 223896 671674 223952
rect 671342 177928 671398 177984
rect 670606 147600 670662 147656
rect 672078 224440 672134 224496
rect 672538 220224 672594 220280
rect 672078 217504 672134 217560
rect 671986 217232 672042 217288
rect 671986 216688 672042 216744
rect 672078 216008 672134 216064
rect 672078 215328 672134 215384
rect 672078 214104 672134 214160
rect 672078 199688 672134 199744
rect 672538 216688 672594 216744
rect 673274 229064 673330 229120
rect 673090 228520 673146 228576
rect 673458 227024 673514 227080
rect 673274 222536 673330 222592
rect 673274 221040 673330 221096
rect 673090 220632 673146 220688
rect 673090 216144 673146 216200
rect 672722 213560 672778 213616
rect 672814 213288 672870 213344
rect 672538 213152 672594 213208
rect 672630 212064 672686 212120
rect 671986 171944 672042 172000
rect 671710 150048 671766 150104
rect 672446 175616 672502 175672
rect 672354 168272 672410 168328
rect 672170 168000 672226 168056
rect 671986 144880 672042 144936
rect 672354 166912 672410 166968
rect 672170 135088 672226 135144
rect 671342 131688 671398 131744
rect 670422 121624 670478 121680
rect 671526 129240 671582 129296
rect 672170 124888 672226 124944
rect 672998 201320 673054 201376
rect 673090 200776 673146 200832
rect 673458 216416 673514 216472
rect 673458 213832 673514 213888
rect 673274 197920 673330 197976
rect 673090 181464 673146 181520
rect 673182 176840 673238 176896
rect 673458 170720 673514 170776
rect 672998 169088 673054 169144
rect 673090 168680 673146 168736
rect 673872 230152 673928 230208
rect 673872 228656 673928 228712
rect 675206 245520 675262 245576
rect 675390 242664 675446 242720
rect 675390 242256 675446 242312
rect 675390 241440 675446 241496
rect 675390 240216 675446 240272
rect 675114 237224 675170 237280
rect 676034 235184 676090 235240
rect 673918 217640 673974 217696
rect 673918 177248 673974 177304
rect 673918 174392 673974 174448
rect 673090 152632 673146 152688
rect 673182 151272 673238 151328
rect 672998 133456 673054 133512
rect 672998 132640 673054 132696
rect 674102 172896 674158 172952
rect 673826 162832 673882 162888
rect 673550 156440 673606 156496
rect 673550 156168 673606 156224
rect 673366 132096 673422 132152
rect 674102 162016 674158 162072
rect 673918 129648 673974 129704
rect 673366 126520 673422 126576
rect 672814 124072 672870 124128
rect 672998 123256 673054 123312
rect 672538 120808 672594 120864
rect 673182 122984 673238 123040
rect 672998 120672 673054 120728
rect 672814 118768 672870 118824
rect 672354 115776 672410 115832
rect 672998 111016 673054 111072
rect 673182 106256 673238 106312
rect 672170 104624 672226 104680
rect 668766 104488 668822 104544
rect 668582 102856 668638 102912
rect 673918 124480 673974 124536
rect 674674 230444 674730 230480
rect 674674 230424 674676 230444
rect 674676 230424 674728 230444
rect 674728 230424 674730 230444
rect 674838 230424 674894 230480
rect 674838 226072 674894 226128
rect 674562 222264 674618 222320
rect 674838 221720 674894 221776
rect 675206 225664 675262 225720
rect 675022 221448 675078 221504
rect 675666 224984 675722 225040
rect 675206 219816 675262 219872
rect 674838 219000 674894 219056
rect 674470 214920 674526 214976
rect 674654 213696 674710 213752
rect 675482 218728 675538 218784
rect 676770 230152 676826 230208
rect 676402 228520 676458 228576
rect 676034 221856 676090 221912
rect 675574 218184 675630 218240
rect 674930 204176 674986 204232
rect 675390 212472 675446 212528
rect 676034 217640 676090 217696
rect 676034 216688 676090 216744
rect 675758 215328 675814 215384
rect 677322 227024 677378 227080
rect 678242 223760 678298 223816
rect 683302 223080 683358 223136
rect 683118 222672 683174 222728
rect 675850 214648 675906 214704
rect 676034 214512 676090 214568
rect 676034 211384 676090 211440
rect 675482 206896 675538 206952
rect 675390 204176 675446 204232
rect 674470 197104 674526 197160
rect 674930 202816 674986 202872
rect 675758 202680 675814 202736
rect 675482 201320 675538 201376
rect 674930 199688 674986 199744
rect 675758 199960 675814 200016
rect 675114 198464 675170 198520
rect 675482 198192 675538 198248
rect 675390 197104 675446 197160
rect 675758 194520 675814 194576
rect 675758 193160 675814 193216
rect 675666 192752 675722 192808
rect 675390 191528 675446 191584
rect 676034 190032 676090 190088
rect 675850 180240 675906 180296
rect 675850 177656 675906 177712
rect 676218 181192 676274 181248
rect 676218 178880 676274 178936
rect 674470 176024 674526 176080
rect 674286 153176 674342 153232
rect 674654 175208 674710 175264
rect 674470 131280 674526 131336
rect 674838 173984 674894 174040
rect 681002 173576 681058 173632
rect 676034 173168 676090 173224
rect 676586 169904 676642 169960
rect 675666 167456 675722 167512
rect 675206 162288 675262 162344
rect 676586 166368 676642 166424
rect 682382 171536 682438 171592
rect 683118 167864 683174 167920
rect 681002 162696 681058 162752
rect 675850 162288 675906 162344
rect 683118 162016 683174 162072
rect 675482 161472 675538 161528
rect 675758 156984 675814 157040
rect 675298 156440 675354 156496
rect 675114 155896 675170 155952
rect 675758 155760 675814 155816
rect 675114 152632 675170 152688
rect 675758 151408 675814 151464
rect 675114 151272 675170 151328
rect 674930 150320 674986 150376
rect 675758 148416 675814 148472
rect 675114 147600 675170 147656
rect 675390 147600 675446 147656
rect 675114 144880 675170 144936
rect 675850 134544 675906 134600
rect 676494 133048 676550 133104
rect 674654 130464 674710 130520
rect 676218 130192 676274 130248
rect 674930 128832 674986 128888
rect 674562 128424 674618 128480
rect 674378 123664 674434 123720
rect 674378 122984 674434 123040
rect 674746 122984 674802 123040
rect 674102 117408 674158 117464
rect 673918 106936 673974 106992
rect 676218 127744 676274 127800
rect 676402 127744 676458 127800
rect 679622 126112 679678 126168
rect 676494 123256 676550 123312
rect 676494 122848 676550 122904
rect 675022 122440 675078 122496
rect 675022 121624 675078 121680
rect 675206 117000 675262 117056
rect 682382 125296 682438 125352
rect 682382 117272 682438 117328
rect 675942 117000 675998 117056
rect 675482 115776 675538 115832
rect 675758 112376 675814 112432
rect 675758 111696 675814 111752
rect 675758 111288 675814 111344
rect 675758 110336 675814 110392
rect 675758 108160 675814 108216
rect 675390 106936 675446 106992
rect 675114 106256 675170 106312
rect 675114 104624 675170 104680
rect 675390 102584 675446 102640
rect 673366 100952 673422 101008
rect 675114 100952 675170 101008
rect 637026 96872 637082 96928
rect 641994 96464 642050 96520
rect 635738 95376 635794 95432
rect 647146 94968 647202 95024
rect 626446 94424 626502 94480
rect 626262 93608 626318 93664
rect 626446 92792 626502 92848
rect 625802 91976 625858 92032
rect 647514 92384 647570 92440
rect 626446 91160 626502 91216
rect 626446 90344 626502 90400
rect 626446 89564 626448 89584
rect 626448 89564 626500 89584
rect 626500 89564 626502 89584
rect 626446 89528 626502 89564
rect 624974 88576 625030 88632
rect 626446 87896 626502 87952
rect 626262 87080 626318 87136
rect 626446 86300 626448 86320
rect 626448 86300 626500 86320
rect 626500 86300 626502 86320
rect 626446 86264 626502 86300
rect 648250 89528 648306 89584
rect 626446 85484 626448 85504
rect 626448 85484 626500 85504
rect 626500 85484 626502 85504
rect 626446 85448 626502 85484
rect 625250 84632 625306 84688
rect 625802 83816 625858 83872
rect 628746 83272 628802 83328
rect 629206 81640 629262 81696
rect 624422 77288 624478 77344
rect 633898 78512 633954 78568
rect 633898 77288 633954 77344
rect 639602 78104 639658 78160
rect 646226 74160 646282 74216
rect 646226 67088 646282 67144
rect 646686 71712 646742 71768
rect 647238 68856 647294 68912
rect 646502 64368 646558 64424
rect 648618 62056 648674 62112
rect 647238 59200 647294 59256
rect 649998 87080 650054 87136
rect 654598 94152 654654 94208
rect 654322 91432 654378 91488
rect 655426 93336 655482 93392
rect 655426 90652 655428 90672
rect 655428 90652 655480 90672
rect 655480 90652 655482 90672
rect 655426 90616 655482 90652
rect 655794 89800 655850 89856
rect 663798 93064 663854 93120
rect 663982 88984 664038 89040
rect 665178 91704 665234 91760
rect 665546 93336 665602 93392
rect 665362 90616 665418 90672
rect 664350 89800 664406 89856
rect 650550 84632 650606 84688
rect 650366 82184 650422 82240
rect 648802 57296 648858 57352
rect 661590 48454 661646 48510
rect 553674 48048 553730 48104
rect 552018 47776 552074 47832
rect 547878 47504 547934 47560
rect 545670 47232 545726 47288
rect 465262 46688 465318 46744
rect 662418 47368 662474 47424
rect 464342 44104 464398 44160
rect 471058 43424 471114 43480
rect 465814 43152 465870 43208
rect 461950 42200 462006 42256
rect 518806 42744 518862 42800
rect 515402 42064 515458 42120
rect 520922 42064 520978 42120
rect 522026 42064 522082 42120
rect 526442 42064 526498 42120
rect 529570 42064 529626 42120
rect 141698 40296 141754 40352
<< metal3 >>
rect 185025 1002146 185091 1002149
rect 185012 1002144 185091 1002146
rect 185012 1002088 185030 1002144
rect 185086 1002088 185091 1002144
rect 185012 1002086 185091 1002088
rect 185025 1002083 185091 1002086
rect 82169 1002010 82235 1002013
rect 133689 1002010 133755 1002013
rect 82156 1002008 82235 1002010
rect 82156 1001952 82174 1002008
rect 82230 1001952 82235 1002008
rect 82156 1001950 82235 1001952
rect 133676 1002008 133755 1002010
rect 133676 1001952 133694 1002008
rect 133750 1001952 133755 1002008
rect 133676 1001950 133755 1001952
rect 82169 1001947 82235 1001950
rect 133689 1001947 133755 1001950
rect 483013 1002010 483079 1002013
rect 534993 1002010 535059 1002013
rect 636193 1002010 636259 1002013
rect 483013 1002008 483092 1002010
rect 483013 1001952 483018 1002008
rect 483074 1001952 483092 1002008
rect 483013 1001950 483092 1001952
rect 534980 1002008 535059 1002010
rect 534980 1001952 534998 1002008
rect 535054 1001952 535059 1002008
rect 534980 1001950 535059 1001952
rect 636180 1002008 636259 1002010
rect 636180 1001952 636198 1002008
rect 636254 1001952 636259 1002008
rect 636180 1001950 636259 1001952
rect 483013 1001947 483079 1001950
rect 534993 1001947 535059 1001950
rect 636193 1001947 636259 1001950
rect 232957 997388 233023 997389
rect 232957 997384 233004 997388
rect 233068 997386 233074 997388
rect 232957 997328 232962 997384
rect 232957 997324 233004 997328
rect 233068 997326 233114 997386
rect 233068 997324 233074 997326
rect 232957 997323 233023 997324
rect 240133 997250 240199 997253
rect 240550 997250 240610 997628
rect 285397 997388 285463 997389
rect 285397 997384 285444 997388
rect 285508 997386 285514 997388
rect 292573 997386 292639 997389
rect 293174 997386 293234 997628
rect 404310 997389 404370 997628
rect 285397 997328 285402 997384
rect 285397 997324 285444 997328
rect 285508 997326 285554 997386
rect 292573 997384 293234 997386
rect 292573 997328 292578 997384
rect 292634 997328 293234 997384
rect 292573 997326 293234 997328
rect 387517 997388 387583 997389
rect 387517 997384 387564 997388
rect 387628 997386 387634 997388
rect 387517 997328 387522 997384
rect 285508 997324 285514 997326
rect 285397 997323 285463 997324
rect 292573 997323 292639 997326
rect 387517 997324 387564 997328
rect 387628 997326 387674 997386
rect 404310 997384 404419 997389
rect 404310 997328 404358 997384
rect 404414 997328 404419 997384
rect 404310 997326 404419 997328
rect 387628 997324 387634 997326
rect 387517 997323 387583 997324
rect 404353 997323 404419 997326
rect 240133 997248 240610 997250
rect 240133 997192 240138 997248
rect 240194 997192 240610 997248
rect 240133 997190 240610 997192
rect 240133 997187 240199 997190
rect 232998 990932 233004 990996
rect 233068 990994 233074 990996
rect 235901 990994 235967 990997
rect 233068 990992 235967 990994
rect 233068 990936 235906 990992
rect 235962 990936 235967 990992
rect 233068 990934 235967 990936
rect 233068 990932 233074 990934
rect 235901 990931 235967 990934
rect 387558 990932 387564 990996
rect 387628 990994 387634 990996
rect 389173 990994 389239 990997
rect 387628 990992 389239 990994
rect 387628 990936 389178 990992
rect 389234 990936 389239 990992
rect 387628 990934 389239 990936
rect 387628 990932 387634 990934
rect 389173 990931 389239 990934
rect 285438 987940 285444 988004
rect 285508 988002 285514 988004
rect 286961 988002 287027 988005
rect 285508 988000 287027 988002
rect 285508 987944 286966 988000
rect 287022 987944 287027 988000
rect 285508 987942 287027 987944
rect 285508 987940 285514 987942
rect 286961 987939 287027 987942
rect 238661 984058 238727 984061
rect 238661 984056 238770 984058
rect 238661 984000 238666 984056
rect 238722 984000 238770 984056
rect 238661 983995 238770 984000
rect 235901 983786 235967 983789
rect 235901 983784 236378 983786
rect 235901 983728 235906 983784
rect 235962 983728 236378 983784
rect 235901 983726 236378 983728
rect 235901 983723 235967 983726
rect 81341 983514 81407 983517
rect 184933 983514 184999 983517
rect 81341 983512 81604 983514
rect 81341 983456 81346 983512
rect 81402 983456 81604 983512
rect 81341 983454 81604 983456
rect 184933 983512 185564 983514
rect 184933 983456 184938 983512
rect 184994 983456 185564 983512
rect 236318 983484 236378 983726
rect 238710 983484 238770 983995
rect 240133 983786 240199 983789
rect 286961 983786 287027 983789
rect 292573 983786 292639 983789
rect 535453 983786 535519 983789
rect 636193 983786 636259 983789
rect 240133 983784 241346 983786
rect 240133 983728 240138 983784
rect 240194 983728 241346 983784
rect 240133 983726 241346 983728
rect 240133 983723 240199 983726
rect 241286 983484 241346 983726
rect 286961 983784 288082 983786
rect 286961 983728 286966 983784
rect 287022 983728 288082 983784
rect 286961 983726 288082 983728
rect 286961 983723 287027 983726
rect 288022 983484 288082 983726
rect 292573 983784 293234 983786
rect 292573 983728 292578 983784
rect 292634 983728 293234 983784
rect 292573 983726 293234 983728
rect 292573 983723 292639 983726
rect 293174 983484 293234 983726
rect 535453 983784 535562 983786
rect 535453 983728 535458 983784
rect 535514 983728 535562 983784
rect 535453 983723 535562 983728
rect 391933 983514 391999 983517
rect 394417 983514 394483 983517
rect 399753 983514 399819 983517
rect 391644 983512 391999 983514
rect 184933 983454 185564 983456
rect 391644 983456 391938 983512
rect 391994 983456 391999 983512
rect 391644 983454 391999 983456
rect 394220 983512 394483 983514
rect 394220 983456 394422 983512
rect 394478 983456 394483 983512
rect 394220 983454 394483 983456
rect 399556 983512 399819 983514
rect 399556 983456 399758 983512
rect 399814 983456 399819 983512
rect 535502 983484 535562 983723
rect 636150 983784 636259 983786
rect 636150 983728 636198 983784
rect 636254 983728 636259 983784
rect 636150 983723 636259 983728
rect 636150 983484 636210 983723
rect 399556 983454 399819 983456
rect 81341 983451 81407 983454
rect 184933 983451 184999 983454
rect 391933 983451 391999 983454
rect 394417 983451 394483 983454
rect 399753 983451 399819 983454
rect 132493 982562 132559 982565
rect 483841 982562 483907 982565
rect 132493 982560 133676 982562
rect 132493 982504 132498 982560
rect 132554 982504 133676 982560
rect 132493 982502 133676 982504
rect 483644 982560 483907 982562
rect 483644 982504 483846 982560
rect 483902 982504 483907 982560
rect 483644 982502 483907 982504
rect 132493 982499 132559 982502
rect 483841 982499 483907 982502
rect 289721 980930 289787 980933
rect 290414 980930 290474 981036
rect 289721 980928 290474 980930
rect 289721 980872 289726 980928
rect 289782 980872 290474 980928
rect 289721 980870 290474 980872
rect 289721 980867 289787 980870
rect 30097 960258 30163 960261
rect 30084 960256 30163 960258
rect 30084 960200 30102 960256
rect 30158 960200 30163 960256
rect 30084 960198 30163 960200
rect 30097 960195 30163 960198
rect 651373 959170 651439 959173
rect 649980 959168 651439 959170
rect 649980 959112 651378 959168
rect 651434 959112 651439 959168
rect 649980 959110 651439 959112
rect 651373 959107 651439 959110
rect 677409 959170 677475 959173
rect 677409 959168 677764 959170
rect 677409 959112 677414 959168
rect 677470 959112 677764 959168
rect 677409 959110 677764 959112
rect 677409 959107 677475 959110
rect 63401 959034 63467 959037
rect 63401 959032 64676 959034
rect 63401 958976 63406 959032
rect 63462 958976 64676 959032
rect 63401 958974 64676 958976
rect 63401 958971 63467 958974
rect 676029 897154 676095 897157
rect 676029 897152 676292 897154
rect 676029 897096 676034 897152
rect 676090 897096 676292 897152
rect 676029 897094 676292 897096
rect 676029 897091 676095 897094
rect 675845 896746 675911 896749
rect 675845 896744 676292 896746
rect 675845 896688 675850 896744
rect 675906 896688 676292 896744
rect 675845 896686 676292 896688
rect 675845 896683 675911 896686
rect 676029 896338 676095 896341
rect 676029 896336 676292 896338
rect 676029 896280 676034 896336
rect 676090 896280 676292 896336
rect 676029 896278 676292 896280
rect 676029 896275 676095 896278
rect 675845 895522 675911 895525
rect 675845 895520 676292 895522
rect 675845 895464 675850 895520
rect 675906 895464 676292 895520
rect 675845 895462 676292 895464
rect 675845 895459 675911 895462
rect 676029 894706 676095 894709
rect 676029 894704 676292 894706
rect 676029 894648 676034 894704
rect 676090 894648 676292 894704
rect 676029 894646 676292 894648
rect 676029 894643 676095 894646
rect 675845 893890 675911 893893
rect 675845 893888 676292 893890
rect 675845 893832 675850 893888
rect 675906 893832 676292 893888
rect 675845 893830 676292 893832
rect 675845 893827 675911 893830
rect 676029 893074 676095 893077
rect 676029 893072 676292 893074
rect 676029 893016 676034 893072
rect 676090 893016 676292 893072
rect 676029 893014 676292 893016
rect 676029 893011 676095 893014
rect 676029 892666 676095 892669
rect 676029 892664 676292 892666
rect 676029 892608 676034 892664
rect 676090 892608 676292 892664
rect 676029 892606 676292 892608
rect 676029 892603 676095 892606
rect 675886 892196 675892 892260
rect 675956 892258 675962 892260
rect 675956 892198 676292 892258
rect 675956 892196 675962 892198
rect 679617 891850 679683 891853
rect 679604 891848 679683 891850
rect 679604 891792 679622 891848
rect 679678 891792 679683 891848
rect 679604 891790 679683 891792
rect 679617 891787 679683 891790
rect 676029 891442 676095 891445
rect 676029 891440 676292 891442
rect 676029 891384 676034 891440
rect 676090 891384 676292 891440
rect 676029 891382 676292 891384
rect 676029 891379 676095 891382
rect 675845 891034 675911 891037
rect 675845 891032 676292 891034
rect 675845 890976 675850 891032
rect 675906 890976 676292 891032
rect 675845 890974 676292 890976
rect 675845 890971 675911 890974
rect 680997 890626 681063 890629
rect 680997 890624 681076 890626
rect 680997 890568 681002 890624
rect 681058 890568 681076 890624
rect 680997 890566 681076 890568
rect 680997 890563 681063 890566
rect 676029 890218 676095 890221
rect 676029 890216 676292 890218
rect 676029 890160 676034 890216
rect 676090 890160 676292 890216
rect 676029 890158 676292 890160
rect 676029 890155 676095 890158
rect 678237 889810 678303 889813
rect 678237 889808 678316 889810
rect 678237 889752 678242 889808
rect 678298 889752 678316 889808
rect 678237 889750 678316 889752
rect 678237 889747 678303 889750
rect 676029 889402 676095 889405
rect 676029 889400 676292 889402
rect 676029 889344 676034 889400
rect 676090 889344 676292 889400
rect 676029 889342 676292 889344
rect 676029 889339 676095 889342
rect 676029 888994 676095 888997
rect 676029 888992 676292 888994
rect 676029 888936 676034 888992
rect 676090 888936 676292 888992
rect 676029 888934 676292 888936
rect 676029 888931 676095 888934
rect 676029 888586 676095 888589
rect 676029 888584 676292 888586
rect 676029 888528 676034 888584
rect 676090 888528 676292 888584
rect 676029 888526 676292 888528
rect 676029 888523 676095 888526
rect 683113 888178 683179 888181
rect 683100 888176 683179 888178
rect 683100 888120 683118 888176
rect 683174 888120 683179 888176
rect 683100 888118 683179 888120
rect 683113 888115 683179 888118
rect 675886 887708 675892 887772
rect 675956 887770 675962 887772
rect 675956 887710 676292 887770
rect 675956 887708 675962 887710
rect 676029 887362 676095 887365
rect 676029 887360 676292 887362
rect 676029 887304 676034 887360
rect 676090 887304 676292 887360
rect 676029 887302 676292 887304
rect 676029 887299 676095 887302
rect 676029 886954 676095 886957
rect 676029 886952 676292 886954
rect 676029 886896 676034 886952
rect 676090 886896 676292 886952
rect 676029 886894 676292 886896
rect 676029 886891 676095 886894
rect 683070 886138 683130 886516
rect 675894 886108 683130 886138
rect 675894 886078 683100 886108
rect 675702 885804 675708 885868
rect 675772 885866 675778 885868
rect 675894 885866 675954 886078
rect 675772 885806 675954 885866
rect 675772 885804 675778 885806
rect 676032 885670 676292 885730
rect 673085 885458 673151 885461
rect 676032 885458 676092 885670
rect 673085 885456 676092 885458
rect 673085 885400 673090 885456
rect 673146 885400 676092 885456
rect 673085 885398 676092 885400
rect 673085 885395 673151 885398
rect 675518 880636 675524 880700
rect 675588 880698 675594 880700
rect 680997 880698 681063 880701
rect 675588 880696 681063 880698
rect 675588 880640 681002 880696
rect 681058 880640 681063 880696
rect 675588 880638 681063 880640
rect 675588 880636 675594 880638
rect 680997 880635 681063 880638
rect 676254 880364 676260 880428
rect 676324 880426 676330 880428
rect 683113 880426 683179 880429
rect 676324 880424 683179 880426
rect 676324 880368 683118 880424
rect 683174 880368 683179 880424
rect 676324 880366 683179 880368
rect 676324 880364 676330 880366
rect 683113 880363 683179 880366
rect 675334 878460 675340 878524
rect 675404 878522 675410 878524
rect 675937 878522 676003 878525
rect 675404 878520 676003 878522
rect 675404 878464 675942 878520
rect 675998 878464 676003 878520
rect 675404 878462 676003 878464
rect 675404 878460 675410 878462
rect 675937 878459 676003 878462
rect 675334 874108 675340 874172
rect 675404 874170 675410 874172
rect 675569 874170 675635 874173
rect 675404 874168 675635 874170
rect 675404 874112 675574 874168
rect 675630 874112 675635 874168
rect 675404 874110 675635 874112
rect 675404 874108 675410 874110
rect 675569 874107 675635 874110
rect 674925 873082 674991 873085
rect 676438 873082 676444 873084
rect 674925 873080 676444 873082
rect 674925 873024 674930 873080
rect 674986 873024 676444 873080
rect 674925 873022 676444 873024
rect 674925 873019 674991 873022
rect 676438 873020 676444 873022
rect 676508 873020 676514 873084
rect 675753 872810 675819 872813
rect 676254 872810 676260 872812
rect 675753 872808 676260 872810
rect 675753 872752 675758 872808
rect 675814 872752 676260 872808
rect 675753 872750 676260 872752
rect 675753 872747 675819 872750
rect 676254 872748 676260 872750
rect 676324 872748 676330 872812
rect 651465 868594 651531 868597
rect 649950 868592 651531 868594
rect 649950 868536 651470 868592
rect 651526 868536 651531 868592
rect 649950 868534 651531 868536
rect 649950 868246 650010 868534
rect 651465 868531 651531 868534
rect 651465 867506 651531 867509
rect 649950 867504 651531 867506
rect 649950 867448 651470 867504
rect 651526 867448 651531 867504
rect 649950 867446 651531 867448
rect 649950 867064 650010 867446
rect 651465 867443 651531 867446
rect 651465 866282 651531 866285
rect 649950 866280 651531 866282
rect 649950 866224 651470 866280
rect 651526 866224 651531 866280
rect 649950 866222 651531 866224
rect 649950 865882 650010 866222
rect 651465 866219 651531 866222
rect 675293 865738 675359 865741
rect 675702 865738 675708 865740
rect 675293 865736 675708 865738
rect 675293 865680 675298 865736
rect 675354 865680 675708 865736
rect 675293 865678 675708 865680
rect 675293 865675 675359 865678
rect 675702 865676 675708 865678
rect 675772 865676 675778 865740
rect 675753 865466 675819 865469
rect 676070 865466 676076 865468
rect 675753 865464 676076 865466
rect 675753 865408 675758 865464
rect 675814 865408 676076 865464
rect 675753 865406 676076 865408
rect 675753 865403 675819 865406
rect 676070 865404 676076 865406
rect 676140 865404 676146 865468
rect 651373 865194 651439 865197
rect 649950 865192 651439 865194
rect 649950 865136 651378 865192
rect 651434 865136 651439 865192
rect 649950 865134 651439 865136
rect 649950 864700 650010 865134
rect 651373 865131 651439 865134
rect 675661 864922 675727 864925
rect 675886 864922 675892 864924
rect 675661 864920 675892 864922
rect 675661 864864 675666 864920
rect 675722 864864 675892 864920
rect 675661 864862 675892 864864
rect 675661 864859 675727 864862
rect 675886 864860 675892 864862
rect 675956 864860 675962 864924
rect 651465 863834 651531 863837
rect 649766 863832 651531 863834
rect 649766 863776 651470 863832
rect 651526 863776 651531 863832
rect 649766 863774 651531 863776
rect 649766 863518 649826 863774
rect 651465 863771 651531 863774
rect 651465 862338 651531 862341
rect 649766 862336 651531 862338
rect 649766 862280 651470 862336
rect 651526 862280 651531 862336
rect 649766 862278 651531 862280
rect 651465 862275 651531 862278
rect 35801 818002 35867 818005
rect 35758 818000 35867 818002
rect 35758 817944 35806 818000
rect 35862 817944 35867 818000
rect 35758 817939 35867 817944
rect 35758 817700 35818 817939
rect 35433 817322 35499 817325
rect 35420 817320 35499 817322
rect 35420 817264 35438 817320
rect 35494 817264 35499 817320
rect 35420 817262 35499 817264
rect 35433 817259 35499 817262
rect 35617 816914 35683 816917
rect 35604 816912 35683 816914
rect 35604 816856 35622 816912
rect 35678 816856 35683 816912
rect 35604 816854 35683 816856
rect 35617 816851 35683 816854
rect 35801 816098 35867 816101
rect 35788 816096 35867 816098
rect 35788 816040 35806 816096
rect 35862 816040 35867 816096
rect 35788 816038 35867 816040
rect 35801 816035 35867 816038
rect 35617 815282 35683 815285
rect 35604 815280 35683 815282
rect 35604 815224 35622 815280
rect 35678 815224 35683 815280
rect 35604 815222 35683 815224
rect 35617 815219 35683 815222
rect 35801 814466 35867 814469
rect 35788 814464 35867 814466
rect 35788 814408 35806 814464
rect 35862 814408 35867 814464
rect 35788 814406 35867 814408
rect 35801 814403 35867 814406
rect 41321 813650 41387 813653
rect 41308 813648 41387 813650
rect 41308 813592 41326 813648
rect 41382 813592 41387 813648
rect 41308 813590 41387 813592
rect 41321 813587 41387 813590
rect 41822 813242 41828 813244
rect 41492 813182 41828 813242
rect 41822 813180 41828 813182
rect 41892 813180 41898 813244
rect 40953 812834 41019 812837
rect 40940 812832 41019 812834
rect 40940 812776 40958 812832
rect 41014 812776 41019 812832
rect 40940 812774 41019 812776
rect 40953 812771 41019 812774
rect 41321 812426 41387 812429
rect 41308 812424 41387 812426
rect 41308 812368 41326 812424
rect 41382 812368 41387 812424
rect 41308 812366 41387 812368
rect 41321 812363 41387 812366
rect 41137 812018 41203 812021
rect 41124 812016 41203 812018
rect 41124 811960 41142 812016
rect 41198 811960 41203 812016
rect 41124 811958 41203 811960
rect 41137 811955 41203 811958
rect 37917 811610 37983 811613
rect 37917 811608 37996 811610
rect 37917 811552 37922 811608
rect 37978 811552 37996 811608
rect 37917 811550 37996 811552
rect 37917 811547 37983 811550
rect 34513 811202 34579 811205
rect 34500 811200 34579 811202
rect 34500 811144 34518 811200
rect 34574 811144 34579 811200
rect 34500 811142 34579 811144
rect 34513 811139 34579 811142
rect 32581 810794 32647 810797
rect 32581 810792 32660 810794
rect 32581 810736 32586 810792
rect 32642 810736 32660 810792
rect 32581 810734 32660 810736
rect 32581 810731 32647 810734
rect 41965 810386 42031 810389
rect 41492 810384 42031 810386
rect 41492 810328 41970 810384
rect 42026 810328 42031 810384
rect 41492 810326 42031 810328
rect 41965 810323 42031 810326
rect 31017 809978 31083 809981
rect 31004 809976 31083 809978
rect 31004 809920 31022 809976
rect 31078 809920 31083 809976
rect 31004 809918 31083 809920
rect 31017 809915 31083 809918
rect 41781 809980 41847 809981
rect 41781 809976 41828 809980
rect 41892 809978 41898 809980
rect 41781 809920 41786 809976
rect 41781 809916 41828 809920
rect 41892 809918 41938 809978
rect 41892 809916 41898 809918
rect 41781 809915 41847 809916
rect 36537 809570 36603 809573
rect 36524 809568 36603 809570
rect 36524 809512 36542 809568
rect 36598 809512 36603 809568
rect 36524 809510 36603 809512
rect 36537 809507 36603 809510
rect 41321 809162 41387 809165
rect 41308 809160 41387 809162
rect 41308 809104 41326 809160
rect 41382 809104 41387 809160
rect 41308 809102 41387 809104
rect 41321 809099 41387 809102
rect 41781 808754 41847 808757
rect 41492 808752 41847 808754
rect 41492 808696 41786 808752
rect 41842 808696 41847 808752
rect 41492 808694 41847 808696
rect 41781 808691 41847 808694
rect 41137 808346 41203 808349
rect 41124 808344 41203 808346
rect 41124 808288 41142 808344
rect 41198 808288 41203 808344
rect 41124 808286 41203 808288
rect 41137 808283 41203 808286
rect 41822 807938 41828 807940
rect 41492 807878 41828 807938
rect 41822 807876 41828 807878
rect 41892 807876 41898 807940
rect 41321 807530 41387 807533
rect 41308 807528 41387 807530
rect 41308 807472 41326 807528
rect 41382 807472 41387 807528
rect 41308 807470 41387 807472
rect 41321 807467 41387 807470
rect 41094 806717 41154 807092
rect 41094 806712 41203 806717
rect 41094 806684 41142 806712
rect 41124 806656 41142 806684
rect 41198 806656 41203 806712
rect 41124 806654 41203 806656
rect 41137 806651 41203 806654
rect 41321 806306 41387 806309
rect 41308 806304 41387 806306
rect 41308 806248 41326 806304
rect 41382 806248 41387 806304
rect 41308 806246 41387 806248
rect 41321 806243 41387 806246
rect 40534 805564 40540 805628
rect 40604 805626 40610 805628
rect 41965 805626 42031 805629
rect 40604 805624 42031 805626
rect 40604 805568 41970 805624
rect 42026 805568 42031 805624
rect 40604 805566 42031 805568
rect 40604 805564 40610 805566
rect 41965 805563 42031 805566
rect 40718 805156 40724 805220
rect 40788 805218 40794 805220
rect 41781 805218 41847 805221
rect 40788 805216 41847 805218
rect 40788 805160 41786 805216
rect 41842 805160 41847 805216
rect 40788 805158 41847 805160
rect 40788 805156 40794 805158
rect 41781 805155 41847 805158
rect 40902 804748 40908 804812
rect 40972 804810 40978 804812
rect 41822 804810 41828 804812
rect 40972 804750 41828 804810
rect 40972 804748 40978 804750
rect 41822 804748 41828 804750
rect 41892 804748 41898 804812
rect 32581 802498 32647 802501
rect 41822 802498 41828 802500
rect 32581 802496 41828 802498
rect 32581 802440 32586 802496
rect 32642 802440 41828 802496
rect 32581 802438 41828 802440
rect 32581 802435 32647 802438
rect 41822 802436 41828 802438
rect 41892 802436 41898 802500
rect 42149 798148 42215 798149
rect 42149 798144 42196 798148
rect 42260 798146 42266 798148
rect 42149 798088 42154 798144
rect 42149 798084 42196 798088
rect 42260 798086 42306 798146
rect 42260 798084 42266 798086
rect 42149 798083 42215 798084
rect 42057 797330 42123 797333
rect 43621 797330 43687 797333
rect 42057 797328 43687 797330
rect 42057 797272 42062 797328
rect 42118 797272 43626 797328
rect 43682 797272 43687 797328
rect 42057 797270 43687 797272
rect 42057 797267 42123 797270
rect 43621 797267 43687 797270
rect 40902 794820 40908 794884
rect 40972 794882 40978 794884
rect 41781 794882 41847 794885
rect 40972 794880 41847 794882
rect 40972 794824 41786 794880
rect 41842 794824 41847 794880
rect 40972 794822 41847 794824
rect 40972 794820 40978 794822
rect 41781 794819 41847 794822
rect 42149 794476 42215 794477
rect 42149 794474 42196 794476
rect 42104 794472 42196 794474
rect 42104 794416 42154 794472
rect 42104 794414 42196 794416
rect 42149 794412 42196 794414
rect 42260 794412 42266 794476
rect 42149 794411 42215 794412
rect 41638 791964 41644 792028
rect 41708 792026 41714 792028
rect 42425 792026 42491 792029
rect 41708 792024 42491 792026
rect 41708 791968 42430 792024
rect 42486 791968 42491 792024
rect 41708 791966 42491 791968
rect 41708 791964 41714 791966
rect 42425 791963 42491 791966
rect 40718 790604 40724 790668
rect 40788 790666 40794 790668
rect 41781 790666 41847 790669
rect 40788 790664 41847 790666
rect 40788 790608 41786 790664
rect 41842 790608 41847 790664
rect 40788 790606 41847 790608
rect 40788 790604 40794 790606
rect 41781 790603 41847 790606
rect 62205 790530 62271 790533
rect 62205 790528 64706 790530
rect 62205 790472 62210 790528
rect 62266 790472 64706 790528
rect 62205 790470 64706 790472
rect 62205 790467 62271 790470
rect 64646 790304 64706 790470
rect 40534 789244 40540 789308
rect 40604 789306 40610 789308
rect 41781 789306 41847 789309
rect 40604 789304 41847 789306
rect 40604 789248 41786 789304
rect 41842 789248 41847 789304
rect 40604 789246 41847 789248
rect 40604 789244 40610 789246
rect 41781 789243 41847 789246
rect 62941 789170 63007 789173
rect 62941 789168 64154 789170
rect 62941 789112 62946 789168
rect 63002 789152 64154 789168
rect 63002 789112 64676 789152
rect 62941 789110 64676 789112
rect 62941 789107 63007 789110
rect 64094 789092 64676 789110
rect 41454 788292 41460 788356
rect 41524 788354 41530 788356
rect 42425 788354 42491 788357
rect 41524 788352 42491 788354
rect 41524 788296 42430 788352
rect 42486 788296 42491 788352
rect 41524 788294 42491 788296
rect 41524 788292 41530 788294
rect 42425 788291 42491 788294
rect 41822 788020 41828 788084
rect 41892 788082 41898 788084
rect 42425 788082 42491 788085
rect 41892 788080 42491 788082
rect 41892 788024 42430 788080
rect 42486 788024 42491 788080
rect 41892 788022 42491 788024
rect 41892 788020 41898 788022
rect 42425 788019 42491 788022
rect 675753 788082 675819 788085
rect 676070 788082 676076 788084
rect 675753 788080 676076 788082
rect 675753 788024 675758 788080
rect 675814 788024 676076 788080
rect 675753 788022 676076 788024
rect 675753 788019 675819 788022
rect 676070 788020 676076 788022
rect 676140 788020 676146 788084
rect 62113 787402 62179 787405
rect 64646 787402 64706 787940
rect 62113 787400 64706 787402
rect 62113 787344 62118 787400
rect 62174 787344 64706 787400
rect 62113 787342 64706 787344
rect 62113 787339 62179 787342
rect 62941 787130 63007 787133
rect 62941 787128 64706 787130
rect 62941 787072 62946 787128
rect 63002 787072 64706 787128
rect 62941 787070 64706 787072
rect 62941 787067 63007 787070
rect 64646 786758 64706 787070
rect 674414 786660 674420 786724
rect 674484 786722 674490 786724
rect 675109 786722 675175 786725
rect 675385 786724 675451 786725
rect 675334 786722 675340 786724
rect 674484 786720 675175 786722
rect 674484 786664 675114 786720
rect 675170 786664 675175 786720
rect 674484 786662 675175 786664
rect 675294 786662 675340 786722
rect 675404 786720 675451 786724
rect 675446 786664 675451 786720
rect 674484 786660 674490 786662
rect 675109 786659 675175 786662
rect 675334 786660 675340 786662
rect 675404 786660 675451 786664
rect 675385 786659 675451 786660
rect 62113 786178 62179 786181
rect 62113 786176 64706 786178
rect 62113 786120 62118 786176
rect 62174 786120 64706 786176
rect 62113 786118 64706 786120
rect 62113 786115 62179 786118
rect 64646 785576 64706 786118
rect 62757 784954 62823 784957
rect 62757 784952 64706 784954
rect 62757 784896 62762 784952
rect 62818 784896 64706 784952
rect 62757 784894 64706 784896
rect 62757 784891 62823 784894
rect 64646 784394 64706 784894
rect 673637 780058 673703 780061
rect 675477 780058 675543 780061
rect 673637 780056 675543 780058
rect 673637 780000 673642 780056
rect 673698 780000 675482 780056
rect 675538 780000 675543 780056
rect 673637 779998 675543 780000
rect 673637 779995 673703 779998
rect 675477 779995 675543 779998
rect 674465 779242 674531 779245
rect 675477 779242 675543 779245
rect 674465 779240 675543 779242
rect 674465 779184 674470 779240
rect 674526 779184 675482 779240
rect 675538 779184 675543 779240
rect 674465 779182 675543 779184
rect 674465 779179 674531 779182
rect 675477 779179 675543 779182
rect 674281 778834 674347 778837
rect 675477 778834 675543 778837
rect 674281 778832 675543 778834
rect 649950 778426 650010 778824
rect 674281 778776 674286 778832
rect 674342 778776 675482 778832
rect 675538 778776 675543 778832
rect 674281 778774 675543 778776
rect 674281 778771 674347 778774
rect 675477 778771 675543 778774
rect 651465 778426 651531 778429
rect 649950 778424 651531 778426
rect 649950 778368 651470 778424
rect 651526 778368 651531 778424
rect 649950 778366 651531 778368
rect 651465 778363 651531 778366
rect 649950 777066 650010 777642
rect 672901 777474 672967 777477
rect 675385 777474 675451 777477
rect 672901 777472 675451 777474
rect 672901 777416 672906 777472
rect 672962 777416 675390 777472
rect 675446 777416 675451 777472
rect 672901 777414 675451 777416
rect 672901 777411 672967 777414
rect 675385 777411 675451 777414
rect 652017 777066 652083 777069
rect 649950 777064 652083 777066
rect 649950 777008 652022 777064
rect 652078 777008 652083 777064
rect 649950 777006 652083 777008
rect 652017 777003 652083 777006
rect 674925 777066 674991 777069
rect 675477 777066 675543 777069
rect 674925 777064 675543 777066
rect 674925 777008 674930 777064
rect 674986 777008 675482 777064
rect 675538 777008 675543 777064
rect 674925 777006 675543 777008
rect 674925 777003 674991 777006
rect 675477 777003 675543 777006
rect 649950 776114 650010 776460
rect 651465 776114 651531 776117
rect 649950 776112 651531 776114
rect 649950 776056 651470 776112
rect 651526 776056 651531 776112
rect 649950 776054 651531 776056
rect 651465 776051 651531 776054
rect 674925 775706 674991 775709
rect 675385 775706 675451 775709
rect 674925 775704 675451 775706
rect 674925 775648 674930 775704
rect 674986 775648 675390 775704
rect 675446 775648 675451 775704
rect 674925 775646 675451 775648
rect 674925 775643 674991 775646
rect 675385 775643 675451 775646
rect 651373 775298 651439 775301
rect 649950 775296 651439 775298
rect 649950 775240 651378 775296
rect 651434 775240 651439 775296
rect 649950 775238 651439 775240
rect 651373 775235 651439 775238
rect 35801 774754 35867 774757
rect 35758 774752 35867 774754
rect 35758 774696 35806 774752
rect 35862 774696 35867 774752
rect 35758 774691 35867 774696
rect 35758 774452 35818 774691
rect 651465 774210 651531 774213
rect 649950 774208 651531 774210
rect 649950 774152 651470 774208
rect 651526 774152 651531 774208
rect 649950 774150 651531 774152
rect 649950 774096 650010 774150
rect 651465 774147 651531 774150
rect 35390 773941 35450 774044
rect 35390 773936 35499 773941
rect 35390 773880 35438 773936
rect 35494 773880 35499 773936
rect 35390 773878 35499 773880
rect 35433 773875 35499 773878
rect 35758 773533 35818 773636
rect 35758 773528 35867 773533
rect 35758 773472 35806 773528
rect 35862 773472 35867 773528
rect 35758 773470 35867 773472
rect 35801 773467 35867 773470
rect 39573 773530 39639 773533
rect 43437 773530 43503 773533
rect 39573 773528 43503 773530
rect 39573 773472 39578 773528
rect 39634 773472 43442 773528
rect 43498 773472 43503 773528
rect 39573 773470 43503 773472
rect 39573 773467 39639 773470
rect 43437 773467 43503 773470
rect 651465 773394 651531 773397
rect 649950 773392 651531 773394
rect 649950 773336 651470 773392
rect 651526 773336 651531 773392
rect 649950 773334 651531 773336
rect 35758 773125 35818 773228
rect 35758 773120 35867 773125
rect 35758 773064 35806 773120
rect 35862 773064 35867 773120
rect 35758 773062 35867 773064
rect 35801 773059 35867 773062
rect 40309 773122 40375 773125
rect 46197 773122 46263 773125
rect 40309 773120 46263 773122
rect 40309 773064 40314 773120
rect 40370 773064 46202 773120
rect 46258 773064 46263 773120
rect 40309 773062 46263 773064
rect 40309 773059 40375 773062
rect 46197 773059 46263 773062
rect 649950 772914 650010 773334
rect 651465 773331 651531 773334
rect 35574 772717 35634 772820
rect 35574 772712 35683 772717
rect 35574 772656 35622 772712
rect 35678 772656 35683 772712
rect 35574 772654 35683 772656
rect 35617 772651 35683 772654
rect 35574 772309 35634 772412
rect 35574 772304 35683 772309
rect 35574 772248 35622 772304
rect 35678 772248 35683 772304
rect 35574 772246 35683 772248
rect 35617 772243 35683 772246
rect 40769 772306 40835 772309
rect 42885 772306 42951 772309
rect 40769 772304 42951 772306
rect 40769 772248 40774 772304
rect 40830 772248 42890 772304
rect 42946 772248 42951 772304
rect 40769 772246 42951 772248
rect 40769 772243 40835 772246
rect 42885 772243 42951 772246
rect 35390 771901 35450 772004
rect 35390 771896 35499 771901
rect 35801 771898 35867 771901
rect 35390 771840 35438 771896
rect 35494 771840 35499 771896
rect 35390 771838 35499 771840
rect 35433 771835 35499 771838
rect 35758 771896 35867 771898
rect 35758 771840 35806 771896
rect 35862 771840 35867 771896
rect 35758 771835 35867 771840
rect 35758 771596 35818 771835
rect 35390 771085 35450 771188
rect 35390 771080 35499 771085
rect 35390 771024 35438 771080
rect 35494 771024 35499 771080
rect 35390 771022 35499 771024
rect 35433 771019 35499 771022
rect 35574 770677 35634 770780
rect 35574 770672 35683 770677
rect 35574 770616 35622 770672
rect 35678 770616 35683 770672
rect 35574 770614 35683 770616
rect 35617 770611 35683 770614
rect 35758 770269 35818 770372
rect 35758 770264 35867 770269
rect 35758 770208 35806 770264
rect 35862 770208 35867 770264
rect 35758 770206 35867 770208
rect 35801 770203 35867 770206
rect 40493 770266 40559 770269
rect 43069 770266 43135 770269
rect 40493 770264 43135 770266
rect 40493 770208 40498 770264
rect 40554 770208 43074 770264
rect 43130 770208 43135 770264
rect 40493 770206 43135 770208
rect 40493 770203 40559 770206
rect 43069 770203 43135 770206
rect 41462 769858 41522 769964
rect 41638 769858 41644 769860
rect 41462 769798 41644 769858
rect 41638 769796 41644 769798
rect 41708 769796 41714 769860
rect 35574 769453 35634 769556
rect 35574 769448 35683 769453
rect 35574 769392 35622 769448
rect 35678 769392 35683 769448
rect 35574 769390 35683 769392
rect 35617 769387 35683 769390
rect 39941 769450 40007 769453
rect 43437 769450 43503 769453
rect 39941 769448 43503 769450
rect 39941 769392 39946 769448
rect 40002 769392 43442 769448
rect 43498 769392 43503 769448
rect 39941 769390 43503 769392
rect 39941 769387 40007 769390
rect 43437 769387 43503 769390
rect 35801 769042 35867 769045
rect 41462 769044 41522 769148
rect 35758 769040 35867 769042
rect 35758 768984 35806 769040
rect 35862 768984 35867 769040
rect 35758 768979 35867 768984
rect 41454 768980 41460 769044
rect 41524 768980 41530 769044
rect 35758 768740 35818 768979
rect 35206 768229 35266 768332
rect 35157 768224 35266 768229
rect 35157 768168 35162 768224
rect 35218 768168 35266 768224
rect 35157 768166 35266 768168
rect 35157 768163 35223 768166
rect 32446 767821 32506 767924
rect 32397 767816 32506 767821
rect 32397 767760 32402 767816
rect 32458 767760 32506 767816
rect 32397 767758 32506 767760
rect 32397 767755 32463 767758
rect 35758 767413 35818 767516
rect 35758 767408 35867 767413
rect 35758 767352 35806 767408
rect 35862 767352 35867 767408
rect 35758 767350 35867 767352
rect 35801 767347 35867 767350
rect 33734 767005 33794 767108
rect 33734 767000 33843 767005
rect 33734 766944 33782 767000
rect 33838 766944 33843 767000
rect 33734 766942 33843 766944
rect 33777 766939 33843 766942
rect 40542 766596 40602 766700
rect 40534 766532 40540 766596
rect 40604 766532 40610 766596
rect 35758 766189 35818 766292
rect 35758 766184 35867 766189
rect 35758 766128 35806 766184
rect 35862 766128 35867 766184
rect 35758 766126 35867 766128
rect 35801 766123 35867 766126
rect 35758 765781 35818 765884
rect 35758 765776 35867 765781
rect 35758 765720 35806 765776
rect 35862 765720 35867 765776
rect 35758 765718 35867 765720
rect 35801 765715 35867 765718
rect 39757 765778 39823 765781
rect 44725 765778 44791 765781
rect 39757 765776 44791 765778
rect 39757 765720 39762 765776
rect 39818 765720 44730 765776
rect 44786 765720 44791 765776
rect 39757 765718 44791 765720
rect 39757 765715 39823 765718
rect 44725 765715 44791 765718
rect 40726 765372 40786 765476
rect 40718 765308 40724 765372
rect 40788 765308 40794 765372
rect 40910 764964 40970 765068
rect 40902 764900 40908 764964
rect 40972 764900 40978 764964
rect 35758 764557 35818 764660
rect 35758 764552 35867 764557
rect 35758 764496 35806 764552
rect 35862 764496 35867 764552
rect 35758 764494 35867 764496
rect 35801 764491 35867 764494
rect 39757 764554 39823 764557
rect 44173 764554 44239 764557
rect 39757 764552 44239 764554
rect 39757 764496 39762 764552
rect 39818 764496 44178 764552
rect 44234 764496 44239 764552
rect 39757 764494 44239 764496
rect 39757 764491 39823 764494
rect 44173 764491 44239 764494
rect 35574 764149 35634 764252
rect 35574 764144 35683 764149
rect 35574 764088 35622 764144
rect 35678 764088 35683 764144
rect 35574 764086 35683 764088
rect 35617 764083 35683 764086
rect 39205 764146 39271 764149
rect 43621 764146 43687 764149
rect 39205 764144 43687 764146
rect 39205 764088 39210 764144
rect 39266 764088 43626 764144
rect 43682 764088 43687 764144
rect 39205 764086 43687 764088
rect 39205 764083 39271 764086
rect 43621 764083 43687 764086
rect 35801 763738 35867 763741
rect 35758 763736 35867 763738
rect 35758 763680 35806 763736
rect 35862 763680 35867 763736
rect 35758 763675 35867 763680
rect 35758 763436 35818 763675
rect 41689 763330 41755 763333
rect 44909 763330 44975 763333
rect 41689 763328 44975 763330
rect 41689 763272 41694 763328
rect 41750 763272 44914 763328
rect 44970 763272 44975 763328
rect 41689 763270 44975 763272
rect 41689 763267 41755 763270
rect 44909 763267 44975 763270
rect 35758 762925 35818 763028
rect 35758 762920 35867 762925
rect 35758 762864 35806 762920
rect 35862 762864 35867 762920
rect 35758 762862 35867 762864
rect 35801 762859 35867 762862
rect 41689 762922 41755 762925
rect 42609 762922 42675 762925
rect 41689 762920 42675 762922
rect 41689 762864 41694 762920
rect 41750 762864 42614 762920
rect 42670 762864 42675 762920
rect 41689 762862 42675 762864
rect 41689 762859 41755 762862
rect 42609 762859 42675 762862
rect 39297 758298 39363 758301
rect 42793 758298 42859 758301
rect 39297 758296 42859 758298
rect 39297 758240 39302 758296
rect 39358 758240 42798 758296
rect 42854 758240 42859 758296
rect 39297 758238 42859 758240
rect 39297 758235 39363 758238
rect 42793 758235 42859 758238
rect 36537 757754 36603 757757
rect 41822 757754 41828 757756
rect 36537 757752 41828 757754
rect 36537 757696 36542 757752
rect 36598 757696 41828 757752
rect 36537 757694 41828 757696
rect 36537 757691 36603 757694
rect 41822 757692 41828 757694
rect 41892 757692 41898 757756
rect 41781 757074 41847 757077
rect 41781 757072 41890 757074
rect 41781 757016 41786 757072
rect 41842 757016 41890 757072
rect 41781 757011 41890 757016
rect 41830 756669 41890 757011
rect 41830 756664 41939 756669
rect 41830 756608 41878 756664
rect 41934 756608 41939 756664
rect 41830 756606 41939 756608
rect 41873 756603 41939 756606
rect 40718 753884 40724 753948
rect 40788 753946 40794 753948
rect 42333 753946 42399 753949
rect 40788 753944 42399 753946
rect 40788 753888 42338 753944
rect 42394 753888 42399 753944
rect 40788 753886 42399 753888
rect 40788 753884 40794 753886
rect 42333 753883 42399 753886
rect 42057 752994 42123 752997
rect 42885 752994 42951 752997
rect 42057 752992 42951 752994
rect 42057 752936 42062 752992
rect 42118 752936 42890 752992
rect 42946 752936 42951 752992
rect 42057 752934 42951 752936
rect 42057 752931 42123 752934
rect 42885 752931 42951 752934
rect 42149 751770 42215 751773
rect 45093 751770 45159 751773
rect 42149 751768 45159 751770
rect 42149 751712 42154 751768
rect 42210 751712 45098 751768
rect 45154 751712 45159 751768
rect 42149 751710 45159 751712
rect 42149 751707 42215 751710
rect 45093 751707 45159 751710
rect 42057 750954 42123 750957
rect 43621 750954 43687 750957
rect 42057 750952 43687 750954
rect 42057 750896 42062 750952
rect 42118 750896 43626 750952
rect 43682 750896 43687 750952
rect 42057 750894 43687 750896
rect 42057 750891 42123 750894
rect 43621 750891 43687 750894
rect 40902 750484 40908 750548
rect 40972 750546 40978 750548
rect 41781 750546 41847 750549
rect 40972 750544 41847 750546
rect 40972 750488 41786 750544
rect 41842 750488 41847 750544
rect 40972 750486 41847 750488
rect 40972 750484 40978 750486
rect 41781 750483 41847 750486
rect 62757 747690 62823 747693
rect 62757 747688 64706 747690
rect 62757 747632 62762 747688
rect 62818 747632 64706 747688
rect 62757 747630 64706 747632
rect 62757 747627 62823 747630
rect 64646 747082 64706 747630
rect 40534 746676 40540 746740
rect 40604 746738 40610 746740
rect 41781 746738 41847 746741
rect 40604 746736 41847 746738
rect 40604 746680 41786 746736
rect 41842 746680 41847 746736
rect 40604 746678 41847 746680
rect 40604 746676 40610 746678
rect 41781 746675 41847 746678
rect 62113 746194 62179 746197
rect 62113 746192 64706 746194
rect 62113 746136 62118 746192
rect 62174 746136 64706 746192
rect 62113 746134 64706 746136
rect 62113 746131 62179 746134
rect 64646 745900 64706 746134
rect 41638 745588 41644 745652
rect 41708 745650 41714 745652
rect 42333 745650 42399 745653
rect 41708 745648 42399 745650
rect 41708 745592 42338 745648
rect 42394 745592 42399 745648
rect 41708 745590 42399 745592
rect 41708 745588 41714 745590
rect 42333 745587 42399 745590
rect 41454 745044 41460 745108
rect 41524 745106 41530 745108
rect 42609 745106 42675 745109
rect 41524 745104 42675 745106
rect 41524 745048 42614 745104
rect 42670 745048 42675 745104
rect 41524 745046 42675 745048
rect 41524 745044 41530 745046
rect 42609 745043 42675 745046
rect 62113 744154 62179 744157
rect 64646 744154 64706 744718
rect 62113 744152 64706 744154
rect 62113 744096 62118 744152
rect 62174 744096 64706 744152
rect 62113 744094 64706 744096
rect 62113 744091 62179 744094
rect 62113 743746 62179 743749
rect 62113 743744 64706 743746
rect 62113 743688 62118 743744
rect 62174 743688 64706 743744
rect 62113 743686 64706 743688
rect 62113 743683 62179 743686
rect 64646 743536 64706 743686
rect 41873 743068 41939 743069
rect 41822 743066 41828 743068
rect 41782 743006 41828 743066
rect 41892 743064 41939 743068
rect 41934 743008 41939 743064
rect 41822 743004 41828 743006
rect 41892 743004 41939 743008
rect 41873 743003 41939 743004
rect 674230 742460 674236 742524
rect 674300 742522 674306 742524
rect 675293 742522 675359 742525
rect 674300 742520 675359 742522
rect 674300 742464 675298 742520
rect 675354 742464 675359 742520
rect 674300 742462 675359 742464
rect 674300 742460 674306 742462
rect 675293 742459 675359 742462
rect 62113 742386 62179 742389
rect 62113 742384 64706 742386
rect 62113 742328 62118 742384
rect 62174 742328 64706 742384
rect 62113 742326 64706 742328
rect 62113 742323 62179 742326
rect 63033 741842 63099 741845
rect 63033 741840 64706 741842
rect 63033 741784 63038 741840
rect 63094 741784 64706 741840
rect 63033 741782 64706 741784
rect 63033 741779 63099 741782
rect 64646 741172 64706 741782
rect 674598 738108 674604 738172
rect 674668 738170 674674 738172
rect 675293 738170 675359 738173
rect 674668 738168 675359 738170
rect 674668 738112 675298 738168
rect 675354 738112 675359 738168
rect 674668 738110 675359 738112
rect 674668 738108 674674 738110
rect 675293 738107 675359 738110
rect 674649 735042 674715 735045
rect 675385 735042 675451 735045
rect 674649 735040 675451 735042
rect 674649 734984 674654 735040
rect 674710 734984 675390 735040
rect 675446 734984 675451 735040
rect 674649 734982 675451 734984
rect 674649 734979 674715 734982
rect 675385 734979 675451 734982
rect 674097 734498 674163 734501
rect 675385 734498 675451 734501
rect 674097 734496 675451 734498
rect 674097 734440 674102 734496
rect 674158 734440 675390 734496
rect 675446 734440 675451 734496
rect 674097 734438 675451 734440
rect 674097 734435 674163 734438
rect 675385 734435 675451 734438
rect 649950 734226 650010 734402
rect 651465 734226 651531 734229
rect 649950 734224 651531 734226
rect 649950 734168 651470 734224
rect 651526 734168 651531 734224
rect 649950 734166 651531 734168
rect 651465 734163 651531 734166
rect 671245 733818 671311 733821
rect 675477 733818 675543 733821
rect 671245 733816 675543 733818
rect 671245 733760 671250 733816
rect 671306 733760 675482 733816
rect 675538 733760 675543 733816
rect 671245 733758 675543 733760
rect 671245 733755 671311 733758
rect 675477 733755 675543 733758
rect 649950 732866 650010 733220
rect 652661 732866 652727 732869
rect 649950 732864 652727 732866
rect 649950 732808 652666 732864
rect 652722 732808 652727 732864
rect 649950 732806 652727 732808
rect 652661 732803 652727 732806
rect 672073 732730 672139 732733
rect 675477 732730 675543 732733
rect 672073 732728 675543 732730
rect 672073 732672 672078 732728
rect 672134 732672 675482 732728
rect 675538 732672 675543 732728
rect 672073 732670 675543 732672
rect 672073 732667 672139 732670
rect 675477 732667 675543 732670
rect 649950 731778 650010 732038
rect 651465 731778 651531 731781
rect 649950 731776 651531 731778
rect 649950 731720 651470 731776
rect 651526 731720 651531 731776
rect 649950 731718 651531 731720
rect 651465 731715 651531 731718
rect 43621 731370 43687 731373
rect 41492 731368 43687 731370
rect 41492 731312 43626 731368
rect 43682 731312 43687 731368
rect 41492 731310 43687 731312
rect 43621 731307 43687 731310
rect 651373 731098 651439 731101
rect 649950 731096 651439 731098
rect 649950 731040 651378 731096
rect 651434 731040 651439 731096
rect 649950 731038 651439 731040
rect 46197 730962 46263 730965
rect 41492 730960 46263 730962
rect 41492 730904 46202 730960
rect 46258 730904 46263 730960
rect 41492 730902 46263 730904
rect 46197 730899 46263 730902
rect 649950 730856 650010 731038
rect 651373 731035 651439 731038
rect 42425 730554 42491 730557
rect 41492 730552 42491 730554
rect 41492 730496 42430 730552
rect 42486 730496 42491 730552
rect 41492 730494 42491 730496
rect 42425 730491 42491 730494
rect 44541 730146 44607 730149
rect 41492 730144 44607 730146
rect 41492 730088 44546 730144
rect 44602 730088 44607 730144
rect 41492 730086 44607 730088
rect 44541 730083 44607 730086
rect 668761 730146 668827 730149
rect 675109 730146 675175 730149
rect 668761 730144 675175 730146
rect 668761 730088 668766 730144
rect 668822 730088 675114 730144
rect 675170 730088 675175 730144
rect 668761 730086 675175 730088
rect 668761 730083 668827 730086
rect 675109 730083 675175 730086
rect 675293 730148 675359 730149
rect 675293 730144 675340 730148
rect 675404 730146 675410 730148
rect 675293 730088 675298 730144
rect 675293 730084 675340 730088
rect 675404 730086 675450 730146
rect 675404 730084 675410 730086
rect 675293 730083 675359 730084
rect 651465 729874 651531 729877
rect 649950 729872 651531 729874
rect 649950 729816 651470 729872
rect 651526 729816 651531 729872
rect 649950 729814 651531 729816
rect 44173 729738 44239 729741
rect 41492 729736 44239 729738
rect 41492 729680 44178 729736
rect 44234 729680 44239 729736
rect 41492 729678 44239 729680
rect 44173 729675 44239 729678
rect 649950 729674 650010 729814
rect 651465 729811 651531 729814
rect 674649 729874 674715 729877
rect 676806 729874 676812 729876
rect 674649 729872 676812 729874
rect 674649 729816 674654 729872
rect 674710 729816 676812 729872
rect 674649 729814 676812 729816
rect 674649 729811 674715 729814
rect 676806 729812 676812 729814
rect 676876 729812 676882 729876
rect 41321 729330 41387 729333
rect 41308 729328 41387 729330
rect 41308 729272 41326 729328
rect 41382 729272 41387 729328
rect 41308 729270 41387 729272
rect 41321 729267 41387 729270
rect 41278 728687 41338 728892
rect 669405 728786 669471 728789
rect 675477 728786 675543 728789
rect 669405 728784 675543 728786
rect 669405 728728 669410 728784
rect 669466 728728 675482 728784
rect 675538 728728 675543 728784
rect 669405 728726 675543 728728
rect 669405 728723 669471 728726
rect 675477 728723 675543 728726
rect 40677 728684 40743 728687
rect 40677 728682 40786 728684
rect 40677 728626 40682 728682
rect 40738 728626 40786 728682
rect 40677 728621 40786 728626
rect 41278 728682 41387 728687
rect 41278 728626 41326 728682
rect 41382 728626 41387 728682
rect 41278 728624 41387 728626
rect 41321 728621 41387 728624
rect 40726 728484 40786 728621
rect 651465 728514 651531 728517
rect 649950 728512 651531 728514
rect 649950 728456 651470 728512
rect 651526 728456 651531 728512
rect 649950 728454 651531 728456
rect 651465 728451 651531 728454
rect 673269 728378 673335 728381
rect 673269 728376 673378 728378
rect 673269 728320 673274 728376
rect 673330 728320 673378 728376
rect 673269 728315 673378 728320
rect 40861 728106 40927 728109
rect 672993 728106 673059 728109
rect 673318 728106 673378 728315
rect 40861 728104 40940 728106
rect 40861 728048 40866 728104
rect 40922 728048 40940 728104
rect 40861 728046 40940 728048
rect 672993 728104 673378 728106
rect 672993 728048 672998 728104
rect 673054 728048 673378 728104
rect 672993 728046 673378 728048
rect 40861 728043 40927 728046
rect 672993 728043 673059 728046
rect 42977 727698 43043 727701
rect 41492 727696 43043 727698
rect 41492 727640 42982 727696
rect 43038 727640 43043 727696
rect 41492 727638 43043 727640
rect 42977 727635 43043 727638
rect 42977 727290 43043 727293
rect 41492 727288 43043 727290
rect 41492 727232 42982 727288
rect 43038 727232 43043 727288
rect 41492 727230 43043 727232
rect 42977 727227 43043 727230
rect 41137 726882 41203 726885
rect 41124 726880 41203 726882
rect 41124 726824 41142 726880
rect 41198 726824 41203 726880
rect 41124 726822 41203 726824
rect 41137 726819 41203 726822
rect 676070 726548 676076 726612
rect 676140 726610 676146 726612
rect 682377 726610 682443 726613
rect 676140 726608 682443 726610
rect 676140 726552 682382 726608
rect 682438 726552 682443 726608
rect 676140 726550 682443 726552
rect 676140 726548 676146 726550
rect 682377 726547 682443 726550
rect 40953 726474 41019 726477
rect 40940 726472 41019 726474
rect 40940 726416 40958 726472
rect 41014 726416 41019 726472
rect 40940 726414 41019 726416
rect 40953 726411 41019 726414
rect 674414 726276 674420 726340
rect 674484 726338 674490 726340
rect 683297 726338 683363 726341
rect 674484 726336 683363 726338
rect 674484 726280 683302 726336
rect 683358 726280 683363 726336
rect 674484 726278 683363 726280
rect 674484 726276 674490 726278
rect 683297 726275 683363 726278
rect 41324 726066 41844 726100
rect 41308 726040 41844 726066
rect 41308 726006 41384 726040
rect 41784 725932 41844 726040
rect 41784 725870 41828 725932
rect 41822 725868 41828 725870
rect 41892 725868 41898 725932
rect 40953 725658 41019 725661
rect 40940 725656 41019 725658
rect 40940 725600 40958 725656
rect 41014 725600 41019 725656
rect 40940 725598 41019 725600
rect 40953 725595 41019 725598
rect 41781 725660 41847 725661
rect 41781 725656 41828 725660
rect 41892 725658 41898 725660
rect 41781 725600 41786 725656
rect 41781 725596 41828 725600
rect 41892 725598 41938 725658
rect 41892 725596 41898 725598
rect 41781 725595 41847 725596
rect 32397 725250 32463 725253
rect 32397 725248 32476 725250
rect 32397 725192 32402 725248
rect 32458 725192 32476 725248
rect 32397 725190 32476 725192
rect 32397 725187 32463 725190
rect 35157 724842 35223 724845
rect 35157 724840 35236 724842
rect 35157 724784 35162 724840
rect 35218 724784 35236 724840
rect 35157 724782 35236 724784
rect 35157 724779 35223 724782
rect 37273 724434 37339 724437
rect 37260 724432 37339 724434
rect 37260 724376 37278 724432
rect 37334 724376 37339 724432
rect 37260 724374 37339 724376
rect 37273 724371 37339 724374
rect 673821 724162 673887 724165
rect 674281 724162 674347 724165
rect 673821 724160 674347 724162
rect 673821 724104 673826 724160
rect 673882 724104 674286 724160
rect 674342 724104 674347 724160
rect 673821 724102 674347 724104
rect 673821 724099 673887 724102
rect 674281 724099 674347 724102
rect 31661 724026 31727 724029
rect 31661 724024 31740 724026
rect 31661 723968 31666 724024
rect 31722 723968 31740 724024
rect 31661 723966 31740 723968
rect 31661 723963 31727 723966
rect 43989 723618 44055 723621
rect 41492 723616 44055 723618
rect 41492 723560 43994 723616
rect 44050 723560 44055 723616
rect 41492 723558 44055 723560
rect 43989 723555 44055 723558
rect 39297 723210 39363 723213
rect 39284 723208 39363 723210
rect 39284 723152 39302 723208
rect 39358 723152 39363 723208
rect 39284 723150 39363 723152
rect 39297 723147 39363 723150
rect 674925 723210 674991 723213
rect 675150 723210 675156 723212
rect 674925 723208 675156 723210
rect 674925 723152 674930 723208
rect 674986 723152 675156 723208
rect 674925 723150 675156 723152
rect 674925 723147 674991 723150
rect 675150 723148 675156 723150
rect 675220 723148 675226 723212
rect 44725 722802 44791 722805
rect 41492 722800 44791 722802
rect 41492 722744 44730 722800
rect 44786 722744 44791 722800
rect 41492 722742 44791 722744
rect 44725 722739 44791 722742
rect 41781 722394 41847 722397
rect 41492 722392 41847 722394
rect 41492 722336 41786 722392
rect 41842 722336 41847 722392
rect 41492 722334 41847 722336
rect 41781 722331 41847 722334
rect 40726 721772 40786 721956
rect 40718 721708 40724 721772
rect 40788 721708 40794 721772
rect 45093 721578 45159 721581
rect 41492 721576 45159 721578
rect 41492 721520 45098 721576
rect 45154 721520 45159 721576
rect 41492 721518 45159 721520
rect 45093 721515 45159 721518
rect 43621 721170 43687 721173
rect 41492 721168 43687 721170
rect 41492 721112 43626 721168
rect 43682 721112 43687 721168
rect 41492 721110 43687 721112
rect 43621 721107 43687 721110
rect 42793 720354 42859 720357
rect 41492 720352 42859 720354
rect 41492 720296 42798 720352
rect 42854 720296 42859 720352
rect 41492 720294 42859 720296
rect 42793 720291 42859 720294
rect 41597 719266 41663 719269
rect 42241 719266 42307 719269
rect 41597 719264 42307 719266
rect 41597 719208 41602 719264
rect 41658 719208 42246 719264
rect 42302 719208 42307 719264
rect 41597 719206 42307 719208
rect 41597 719203 41663 719206
rect 42241 719203 42307 719206
rect 40953 718994 41019 718997
rect 42057 718994 42123 718997
rect 40953 718992 42123 718994
rect 40953 718936 40958 718992
rect 41014 718936 42062 718992
rect 42118 718936 42123 718992
rect 40953 718934 42123 718936
rect 40953 718931 41019 718934
rect 42057 718931 42123 718934
rect 40534 718524 40540 718588
rect 40604 718586 40610 718588
rect 41781 718586 41847 718589
rect 40604 718584 41847 718586
rect 40604 718528 41786 718584
rect 41842 718528 41847 718584
rect 40604 718526 41847 718528
rect 40604 718524 40610 718526
rect 41781 718523 41847 718526
rect 37273 716954 37339 716957
rect 41822 716954 41828 716956
rect 37273 716952 41828 716954
rect 37273 716896 37278 716952
rect 37334 716896 41828 716952
rect 37273 716894 41828 716896
rect 37273 716891 37339 716894
rect 41822 716892 41828 716894
rect 41892 716892 41898 716956
rect 676029 716546 676095 716549
rect 676029 716544 676292 716546
rect 676029 716488 676034 716544
rect 676090 716488 676292 716544
rect 676029 716486 676292 716488
rect 676029 716483 676095 716486
rect 676029 716138 676095 716141
rect 676029 716136 676292 716138
rect 676029 716080 676034 716136
rect 676090 716080 676292 716136
rect 676029 716078 676292 716080
rect 676029 716075 676095 716078
rect 40217 715866 40283 715869
rect 42701 715866 42767 715869
rect 40217 715864 42767 715866
rect 40217 715808 40222 715864
rect 40278 715808 42706 715864
rect 42762 715808 42767 715864
rect 40217 715806 42767 715808
rect 40217 715803 40283 715806
rect 42701 715803 42767 715806
rect 674005 715730 674071 715733
rect 674005 715728 676292 715730
rect 674005 715672 674010 715728
rect 674066 715672 676292 715728
rect 674005 715670 676292 715672
rect 674005 715667 674071 715670
rect 40585 715322 40651 715325
rect 42425 715322 42491 715325
rect 40585 715320 42491 715322
rect 40585 715264 40590 715320
rect 40646 715264 42430 715320
rect 42486 715264 42491 715320
rect 40585 715262 42491 715264
rect 40585 715259 40651 715262
rect 42425 715259 42491 715262
rect 675845 715322 675911 715325
rect 675845 715320 676292 715322
rect 675845 715264 675850 715320
rect 675906 715264 676292 715320
rect 675845 715262 676292 715264
rect 675845 715259 675911 715262
rect 672625 714914 672691 714917
rect 672625 714912 676292 714914
rect 672625 714856 672630 714912
rect 672686 714856 676292 714912
rect 672625 714854 676292 714856
rect 672625 714851 672691 714854
rect 41689 714506 41755 714509
rect 42006 714506 42012 714508
rect 41689 714504 42012 714506
rect 41689 714448 41694 714504
rect 41750 714448 42012 714504
rect 41689 714446 42012 714448
rect 41689 714443 41755 714446
rect 42006 714444 42012 714446
rect 42076 714444 42082 714508
rect 674005 714506 674071 714509
rect 674005 714504 676292 714506
rect 674005 714448 674010 714504
rect 674066 714448 676292 714504
rect 674005 714446 676292 714448
rect 674005 714443 674071 714446
rect 673269 714098 673335 714101
rect 673269 714096 676292 714098
rect 673269 714040 673274 714096
rect 673330 714040 676292 714096
rect 673269 714038 676292 714040
rect 673269 714035 673335 714038
rect 673085 713690 673151 713693
rect 673085 713688 676292 713690
rect 673085 713632 673090 713688
rect 673146 713632 676292 713688
rect 673085 713630 676292 713632
rect 673085 713627 673151 713630
rect 674005 713282 674071 713285
rect 674005 713280 676292 713282
rect 674005 713224 674010 713280
rect 674066 713224 676292 713280
rect 674005 713222 676292 713224
rect 674005 713219 674071 713222
rect 674005 712874 674071 712877
rect 674005 712872 676292 712874
rect 674005 712816 674010 712872
rect 674066 712816 676292 712872
rect 674005 712814 676292 712816
rect 674005 712811 674071 712814
rect 674005 712466 674071 712469
rect 674005 712464 676292 712466
rect 674005 712408 674010 712464
rect 674066 712408 676292 712464
rect 674005 712406 676292 712408
rect 674005 712403 674071 712406
rect 675293 712058 675359 712061
rect 675293 712056 676292 712058
rect 675293 712000 675298 712056
rect 675354 712000 676292 712056
rect 675293 711998 676292 712000
rect 675293 711995 675359 711998
rect 672809 711650 672875 711653
rect 672809 711648 676292 711650
rect 672809 711592 672814 711648
rect 672870 711592 676292 711648
rect 672809 711590 676292 711592
rect 672809 711587 672875 711590
rect 682377 711242 682443 711245
rect 682364 711240 682443 711242
rect 682364 711184 682382 711240
rect 682438 711184 682443 711240
rect 682364 711182 682443 711184
rect 682377 711179 682443 711182
rect 680997 710834 681063 710837
rect 680997 710832 681076 710834
rect 680997 710776 681002 710832
rect 681058 710776 681076 710832
rect 680997 710774 681076 710776
rect 680997 710771 681063 710774
rect 676029 710426 676095 710429
rect 676029 710424 676292 710426
rect 676029 710368 676034 710424
rect 676090 710368 676292 710424
rect 676029 710366 676292 710368
rect 676029 710363 676095 710366
rect 674005 710018 674071 710021
rect 674005 710016 676292 710018
rect 674005 709960 674010 710016
rect 674066 709960 676292 710016
rect 674005 709958 676292 709960
rect 674005 709955 674071 709958
rect 42057 709884 42123 709885
rect 42006 709882 42012 709884
rect 41966 709822 42012 709882
rect 42076 709880 42123 709884
rect 42118 709824 42123 709880
rect 42006 709820 42012 709822
rect 42076 709820 42123 709824
rect 42057 709819 42123 709820
rect 683297 709610 683363 709613
rect 683284 709608 683363 709610
rect 683284 709552 683302 709608
rect 683358 709552 683363 709608
rect 683284 709550 683363 709552
rect 683297 709547 683363 709550
rect 673821 709340 673887 709341
rect 673821 709338 673868 709340
rect 673776 709336 673868 709338
rect 673776 709280 673826 709336
rect 673776 709278 673868 709280
rect 673821 709276 673868 709278
rect 673932 709276 673938 709340
rect 673821 709275 673887 709276
rect 674005 709202 674071 709205
rect 674005 709200 676292 709202
rect 674005 709144 674010 709200
rect 674066 709144 676292 709200
rect 674005 709142 676292 709144
rect 674005 709139 674071 709142
rect 45093 708794 45159 708797
rect 41830 708792 45159 708794
rect 41830 708736 45098 708792
rect 45154 708736 45159 708792
rect 41830 708734 45159 708736
rect 41830 708525 41890 708734
rect 45093 708731 45159 708734
rect 669221 708794 669287 708797
rect 669221 708792 676292 708794
rect 669221 708736 669226 708792
rect 669282 708736 676292 708792
rect 669221 708734 676292 708736
rect 669221 708731 669287 708734
rect 41830 708520 41939 708525
rect 41830 708464 41878 708520
rect 41934 708464 41939 708520
rect 41830 708462 41939 708464
rect 41873 708459 41939 708462
rect 42057 708522 42123 708525
rect 44725 708522 44791 708525
rect 42057 708520 44791 708522
rect 42057 708464 42062 708520
rect 42118 708464 44730 708520
rect 44786 708464 44791 708520
rect 42057 708462 44791 708464
rect 42057 708459 42123 708462
rect 44725 708459 44791 708462
rect 672993 708386 673059 708389
rect 672993 708384 676292 708386
rect 672993 708328 672998 708384
rect 673054 708328 676292 708384
rect 672993 708326 676292 708328
rect 672993 708323 673059 708326
rect 40534 707916 40540 707980
rect 40604 707978 40610 707980
rect 42190 707978 42196 707980
rect 40604 707918 42196 707978
rect 40604 707916 40610 707918
rect 42190 707916 42196 707918
rect 42260 707916 42266 707980
rect 684125 707978 684191 707981
rect 684125 707976 684204 707978
rect 684125 707920 684130 707976
rect 684186 707920 684204 707976
rect 684125 707918 684204 707920
rect 684125 707915 684191 707918
rect 42149 707706 42215 707709
rect 43805 707706 43871 707709
rect 42149 707704 43871 707706
rect 42149 707648 42154 707704
rect 42210 707648 43810 707704
rect 43866 707648 43871 707704
rect 42149 707646 43871 707648
rect 42149 707643 42215 707646
rect 43805 707643 43871 707646
rect 676029 707570 676095 707573
rect 676029 707568 676292 707570
rect 676029 707512 676034 707568
rect 676090 707512 676292 707568
rect 676029 707510 676292 707512
rect 676029 707507 676095 707510
rect 40718 707372 40724 707436
rect 40788 707434 40794 707436
rect 41781 707434 41847 707437
rect 40788 707432 41847 707434
rect 40788 707376 41786 707432
rect 41842 707376 41847 707432
rect 40788 707374 41847 707376
rect 40788 707372 40794 707374
rect 41781 707371 41847 707374
rect 674005 707162 674071 707165
rect 674005 707160 676292 707162
rect 674005 707104 674010 707160
rect 674066 707104 676292 707160
rect 674005 707102 676292 707104
rect 674005 707099 674071 707102
rect 673821 707028 673887 707029
rect 673821 707026 673868 707028
rect 673776 707024 673868 707026
rect 673776 706968 673826 707024
rect 673776 706966 673868 706968
rect 673821 706964 673868 706966
rect 673932 706964 673938 707028
rect 673821 706963 673887 706964
rect 683481 706754 683547 706757
rect 683468 706752 683547 706754
rect 683468 706696 683486 706752
rect 683542 706696 683547 706752
rect 683468 706694 683547 706696
rect 683481 706691 683547 706694
rect 676029 706346 676095 706349
rect 676029 706344 676292 706346
rect 676029 706288 676034 706344
rect 676090 706288 676292 706344
rect 676029 706286 676292 706288
rect 676029 706283 676095 706286
rect 42241 706212 42307 706213
rect 42190 706148 42196 706212
rect 42260 706210 42307 706212
rect 42260 706208 42352 706210
rect 42302 706152 42352 706208
rect 42260 706150 42352 706152
rect 42260 706148 42307 706150
rect 42241 706147 42307 706148
rect 677182 705530 677242 705908
rect 683113 705530 683179 705533
rect 677182 705528 683179 705530
rect 677182 705500 683118 705528
rect 677212 705472 683118 705500
rect 683174 705472 683179 705528
rect 677212 705470 683179 705472
rect 683113 705467 683179 705470
rect 676029 705122 676095 705125
rect 676029 705120 676292 705122
rect 676029 705064 676034 705120
rect 676090 705064 676292 705120
rect 676029 705062 676292 705064
rect 676029 705059 676095 705062
rect 62113 704442 62179 704445
rect 62113 704440 64706 704442
rect 62113 704384 62118 704440
rect 62174 704384 64706 704440
rect 62113 704382 64706 704384
rect 62113 704379 62179 704382
rect 64646 703860 64706 704382
rect 42057 703490 42123 703493
rect 43989 703490 44055 703493
rect 42057 703488 44055 703490
rect 42057 703432 42062 703488
rect 42118 703432 43994 703488
rect 44050 703432 44055 703488
rect 42057 703430 44055 703432
rect 42057 703427 42123 703430
rect 43989 703427 44055 703430
rect 62113 703354 62179 703357
rect 62113 703352 64706 703354
rect 62113 703296 62118 703352
rect 62174 703296 64706 703352
rect 62113 703294 64706 703296
rect 62113 703291 62179 703294
rect 42057 703082 42123 703085
rect 42701 703082 42767 703085
rect 42057 703080 42767 703082
rect 42057 703024 42062 703080
rect 42118 703024 42706 703080
rect 42762 703024 42767 703080
rect 42057 703022 42767 703024
rect 42057 703019 42123 703022
rect 42701 703019 42767 703022
rect 41638 702748 41644 702812
rect 41708 702810 41714 702812
rect 42609 702810 42675 702813
rect 41708 702808 42675 702810
rect 41708 702752 42614 702808
rect 42670 702752 42675 702808
rect 41708 702750 42675 702752
rect 41708 702748 41714 702750
rect 42609 702747 42675 702750
rect 64646 702678 64706 703294
rect 41454 702068 41460 702132
rect 41524 702130 41530 702132
rect 42609 702130 42675 702133
rect 41524 702128 42675 702130
rect 41524 702072 42614 702128
rect 42670 702072 42675 702128
rect 41524 702070 42675 702072
rect 41524 702068 41530 702070
rect 42609 702067 42675 702070
rect 41822 701796 41828 701860
rect 41892 701858 41898 701860
rect 42425 701858 42491 701861
rect 41892 701856 42491 701858
rect 41892 701800 42430 701856
rect 42486 701800 42491 701856
rect 41892 701798 42491 701800
rect 41892 701796 41898 701798
rect 42425 701795 42491 701798
rect 62205 701314 62271 701317
rect 64646 701314 64706 701496
rect 62205 701312 64706 701314
rect 62205 701256 62210 701312
rect 62266 701256 64706 701312
rect 62205 701254 64706 701256
rect 62205 701251 62271 701254
rect 62757 700906 62823 700909
rect 62757 700904 64706 700906
rect 62757 700848 62762 700904
rect 62818 700848 64706 700904
rect 62757 700846 64706 700848
rect 62757 700843 62823 700846
rect 64646 700314 64706 700846
rect 62297 699546 62363 699549
rect 62297 699544 64706 699546
rect 62297 699488 62302 699544
rect 62358 699488 64706 699544
rect 62297 699486 64706 699488
rect 62297 699483 62363 699486
rect 64646 699132 64706 699486
rect 62113 698186 62179 698189
rect 62113 698184 64706 698186
rect 62113 698128 62118 698184
rect 62174 698128 64706 698184
rect 62113 698126 64706 698128
rect 62113 698123 62179 698126
rect 64646 697950 64706 698126
rect 672257 696962 672323 696965
rect 675293 696962 675359 696965
rect 672257 696960 675359 696962
rect 672257 696904 672262 696960
rect 672318 696904 675298 696960
rect 675354 696904 675359 696960
rect 672257 696902 675359 696904
rect 672257 696899 672323 696902
rect 675293 696899 675359 696902
rect 675477 696828 675543 696829
rect 675477 696824 675524 696828
rect 675588 696826 675594 696828
rect 675477 696768 675482 696824
rect 675477 696764 675524 696768
rect 675588 696766 675634 696826
rect 675588 696764 675594 696766
rect 675477 696763 675543 696764
rect 674414 694588 674420 694652
rect 674484 694650 674490 694652
rect 675109 694650 675175 694653
rect 674484 694648 675175 694650
rect 674484 694592 675114 694648
rect 675170 694592 675175 694648
rect 674484 694590 675175 694592
rect 674484 694588 674490 694590
rect 675109 694587 675175 694590
rect 674005 690162 674071 690165
rect 674925 690162 674991 690165
rect 674005 690160 674991 690162
rect 674005 690104 674010 690160
rect 674066 690104 674930 690160
rect 674986 690104 674991 690160
rect 674005 690102 674991 690104
rect 674005 690099 674071 690102
rect 674925 690099 674991 690102
rect 649950 689482 650010 689980
rect 651465 689482 651531 689485
rect 649950 689480 651531 689482
rect 649950 689424 651470 689480
rect 651526 689424 651531 689480
rect 649950 689422 651531 689424
rect 651465 689419 651531 689422
rect 668393 689482 668459 689485
rect 675109 689482 675175 689485
rect 668393 689480 675175 689482
rect 668393 689424 668398 689480
rect 668454 689424 675114 689480
rect 675170 689424 675175 689480
rect 668393 689422 675175 689424
rect 668393 689419 668459 689422
rect 675109 689419 675175 689422
rect 649980 688802 650562 688828
rect 651649 688802 651715 688805
rect 649980 688800 651715 688802
rect 649980 688768 651654 688800
rect 650502 688744 651654 688768
rect 651710 688744 651715 688800
rect 650502 688742 651715 688744
rect 651649 688739 651715 688742
rect 674005 688802 674071 688805
rect 674925 688802 674991 688805
rect 674005 688800 674991 688802
rect 674005 688744 674010 688800
rect 674066 688744 674930 688800
rect 674986 688744 674991 688800
rect 674005 688742 674991 688744
rect 674005 688739 674071 688742
rect 674925 688739 674991 688742
rect 35433 688394 35499 688397
rect 35390 688392 35499 688394
rect 35390 688336 35438 688392
rect 35494 688336 35499 688392
rect 35390 688331 35499 688336
rect 35390 688092 35450 688331
rect 35801 687714 35867 687717
rect 35788 687712 35867 687714
rect 35788 687656 35806 687712
rect 35862 687656 35867 687712
rect 35788 687654 35867 687656
rect 35801 687651 35867 687654
rect 670601 687714 670667 687717
rect 675109 687714 675175 687717
rect 670601 687712 675175 687714
rect 670601 687656 670606 687712
rect 670662 687656 675114 687712
rect 675170 687656 675175 687712
rect 670601 687654 675175 687656
rect 670601 687651 670667 687654
rect 675109 687651 675175 687654
rect 41689 687578 41755 687581
rect 45277 687578 45343 687581
rect 41689 687576 45343 687578
rect 41689 687520 41694 687576
rect 41750 687520 45282 687576
rect 45338 687520 45343 687576
rect 41689 687518 45343 687520
rect 41689 687515 41755 687518
rect 45277 687515 45343 687518
rect 649950 687442 650010 687616
rect 651465 687442 651531 687445
rect 649950 687440 651531 687442
rect 649950 687384 651470 687440
rect 651526 687384 651531 687440
rect 649950 687382 651531 687384
rect 651465 687379 651531 687382
rect 35617 687306 35683 687309
rect 35604 687304 35683 687306
rect 35604 687248 35622 687304
rect 35678 687248 35683 687304
rect 35604 687246 35683 687248
rect 35617 687243 35683 687246
rect 41689 687170 41755 687173
rect 46197 687170 46263 687173
rect 41689 687168 46263 687170
rect 41689 687112 41694 687168
rect 41750 687112 46202 687168
rect 46258 687112 46263 687168
rect 41689 687110 46263 687112
rect 41689 687107 41755 687110
rect 46197 687107 46263 687110
rect 35433 686898 35499 686901
rect 35420 686896 35499 686898
rect 35420 686840 35438 686896
rect 35494 686840 35499 686896
rect 35420 686838 35499 686840
rect 35433 686835 35499 686838
rect 651465 686762 651531 686765
rect 649950 686760 651531 686762
rect 649950 686704 651470 686760
rect 651526 686704 651531 686760
rect 649950 686702 651531 686704
rect 35801 686490 35867 686493
rect 35788 686488 35867 686490
rect 35788 686432 35806 686488
rect 35862 686432 35867 686488
rect 649950 686434 650010 686702
rect 651465 686699 651531 686702
rect 35788 686430 35867 686432
rect 35801 686427 35867 686430
rect 672809 686218 672875 686221
rect 675109 686218 675175 686221
rect 672809 686216 675175 686218
rect 672809 686160 672814 686216
rect 672870 686160 675114 686216
rect 675170 686160 675175 686216
rect 672809 686158 675175 686160
rect 672809 686155 672875 686158
rect 675109 686155 675175 686158
rect 35801 686082 35867 686085
rect 35788 686080 35867 686082
rect 35788 686024 35806 686080
rect 35862 686024 35867 686080
rect 35788 686022 35867 686024
rect 35801 686019 35867 686022
rect 672993 685810 673059 685813
rect 674925 685810 674991 685813
rect 672993 685808 674991 685810
rect 672993 685752 672998 685808
rect 673054 685752 674930 685808
rect 674986 685752 674991 685808
rect 672993 685750 674991 685752
rect 672993 685747 673059 685750
rect 674925 685747 674991 685750
rect 35801 685674 35867 685677
rect 35788 685672 35867 685674
rect 35788 685616 35806 685672
rect 35862 685616 35867 685672
rect 35788 685614 35867 685616
rect 35801 685611 35867 685614
rect 669773 685538 669839 685541
rect 675109 685538 675175 685541
rect 669773 685536 675175 685538
rect 669773 685480 669778 685536
rect 669834 685480 675114 685536
rect 675170 685480 675175 685536
rect 669773 685478 675175 685480
rect 669773 685475 669839 685478
rect 675109 685475 675175 685478
rect 35617 685266 35683 685269
rect 651465 685266 651531 685269
rect 35604 685264 35683 685266
rect 35604 685208 35622 685264
rect 35678 685208 35683 685264
rect 35604 685206 35683 685208
rect 649950 685264 651531 685266
rect 649950 685208 651470 685264
rect 651526 685208 651531 685264
rect 649950 685206 651531 685208
rect 35617 685203 35683 685206
rect 651465 685203 651531 685206
rect 41689 685130 41755 685133
rect 43437 685130 43503 685133
rect 41689 685128 43503 685130
rect 41689 685072 41694 685128
rect 41750 685072 43442 685128
rect 43498 685072 43503 685128
rect 41689 685070 43503 685072
rect 41689 685067 41755 685070
rect 43437 685067 43503 685070
rect 35801 684858 35867 684861
rect 35788 684856 35867 684858
rect 35788 684800 35806 684856
rect 35862 684800 35867 684856
rect 35788 684798 35867 684800
rect 35801 684795 35867 684798
rect 35617 684450 35683 684453
rect 652569 684450 652635 684453
rect 35604 684448 35683 684450
rect 35604 684392 35622 684448
rect 35678 684392 35683 684448
rect 35604 684390 35683 684392
rect 35617 684387 35683 684390
rect 649950 684448 652635 684450
rect 649950 684392 652574 684448
rect 652630 684392 652635 684448
rect 649950 684390 652635 684392
rect 41689 684314 41755 684317
rect 43437 684314 43503 684317
rect 41689 684312 43503 684314
rect 41689 684256 41694 684312
rect 41750 684256 43442 684312
rect 43498 684256 43503 684312
rect 41689 684254 43503 684256
rect 41689 684251 41755 684254
rect 43437 684251 43503 684254
rect 649950 684070 650010 684390
rect 652569 684387 652635 684390
rect 35433 684042 35499 684045
rect 35420 684040 35499 684042
rect 35420 683984 35438 684040
rect 35494 683984 35499 684040
rect 35420 683982 35499 683984
rect 35433 683979 35499 683982
rect 675109 684042 675175 684045
rect 675518 684042 675524 684044
rect 675109 684040 675524 684042
rect 675109 683984 675114 684040
rect 675170 683984 675524 684040
rect 675109 683982 675524 683984
rect 675109 683979 675175 683982
rect 675518 683980 675524 683982
rect 675588 683980 675594 684044
rect 41689 683906 41755 683909
rect 42977 683906 43043 683909
rect 41689 683904 43043 683906
rect 41689 683848 41694 683904
rect 41750 683848 42982 683904
rect 43038 683848 43043 683904
rect 41689 683846 43043 683848
rect 41689 683843 41755 683846
rect 42977 683843 43043 683846
rect 675293 683772 675359 683773
rect 675293 683770 675340 683772
rect 675248 683768 675340 683770
rect 675248 683712 675298 683768
rect 675248 683710 675340 683712
rect 675293 683708 675340 683710
rect 675404 683708 675410 683772
rect 675293 683707 675359 683708
rect 41822 683634 41828 683636
rect 41492 683574 41828 683634
rect 41822 683572 41828 683574
rect 41892 683572 41898 683636
rect 35801 683226 35867 683229
rect 35788 683224 35867 683226
rect 35788 683168 35806 683224
rect 35862 683168 35867 683224
rect 35788 683166 35867 683168
rect 35801 683163 35867 683166
rect 35617 682818 35683 682821
rect 35604 682816 35683 682818
rect 35604 682760 35622 682816
rect 35678 682760 35683 682816
rect 35604 682758 35683 682760
rect 35617 682755 35683 682758
rect 673637 682818 673703 682821
rect 674833 682818 674899 682821
rect 673637 682816 674899 682818
rect 673637 682760 673642 682816
rect 673698 682760 674838 682816
rect 674894 682760 674899 682816
rect 673637 682758 674899 682760
rect 673637 682755 673703 682758
rect 674833 682755 674899 682758
rect 35801 682410 35867 682413
rect 35788 682408 35867 682410
rect 35788 682352 35806 682408
rect 35862 682352 35867 682408
rect 35788 682350 35867 682352
rect 35801 682347 35867 682350
rect 674230 682348 674236 682412
rect 674300 682410 674306 682412
rect 684125 682410 684191 682413
rect 674300 682408 684191 682410
rect 674300 682352 684130 682408
rect 684186 682352 684191 682408
rect 674300 682350 684191 682352
rect 674300 682348 674306 682350
rect 684125 682347 684191 682350
rect 35157 682002 35223 682005
rect 673729 682002 673795 682005
rect 674833 682002 674899 682005
rect 35157 682000 35236 682002
rect 35157 681944 35162 682000
rect 35218 681944 35236 682000
rect 35157 681942 35236 681944
rect 673729 682000 674899 682002
rect 673729 681944 673734 682000
rect 673790 681944 674838 682000
rect 674894 681944 674899 682000
rect 673729 681942 674899 681944
rect 35157 681939 35223 681942
rect 673729 681939 673795 681942
rect 674833 681939 674899 681942
rect 41781 681732 41847 681733
rect 41781 681728 41828 681732
rect 41892 681730 41898 681732
rect 41781 681672 41786 681728
rect 41781 681668 41828 681672
rect 41892 681670 41938 681730
rect 41892 681668 41898 681670
rect 41781 681667 41847 681668
rect 33041 681594 33107 681597
rect 33028 681592 33107 681594
rect 33028 681536 33046 681592
rect 33102 681536 33107 681592
rect 33028 681534 33107 681536
rect 33041 681531 33107 681534
rect 33777 681186 33843 681189
rect 33764 681184 33843 681186
rect 33764 681128 33782 681184
rect 33838 681128 33843 681184
rect 33764 681126 33843 681128
rect 33777 681123 33843 681126
rect 31017 680778 31083 680781
rect 31004 680776 31083 680778
rect 31004 680720 31022 680776
rect 31078 680720 31083 680776
rect 31004 680718 31083 680720
rect 31017 680715 31083 680718
rect 41689 680642 41755 680645
rect 45461 680642 45527 680645
rect 41689 680640 45527 680642
rect 41689 680584 41694 680640
rect 41750 680584 45466 680640
rect 45522 680584 45527 680640
rect 41689 680582 45527 680584
rect 41689 680579 41755 680582
rect 45461 680579 45527 680582
rect 35801 680370 35867 680373
rect 35788 680368 35867 680370
rect 35788 680312 35806 680368
rect 35862 680312 35867 680368
rect 35788 680310 35867 680312
rect 35801 680307 35867 680310
rect 35617 679962 35683 679965
rect 35604 679960 35683 679962
rect 35604 679904 35622 679960
rect 35678 679904 35683 679960
rect 35604 679902 35683 679904
rect 35617 679899 35683 679902
rect 35433 679554 35499 679557
rect 35420 679552 35499 679554
rect 35420 679496 35438 679552
rect 35494 679496 35499 679552
rect 35420 679494 35499 679496
rect 35433 679491 35499 679494
rect 41689 679418 41755 679421
rect 43989 679418 44055 679421
rect 41689 679416 44055 679418
rect 41689 679360 41694 679416
rect 41750 679360 43994 679416
rect 44050 679360 44055 679416
rect 41689 679358 44055 679360
rect 41689 679355 41755 679358
rect 43989 679355 44055 679358
rect 35801 679146 35867 679149
rect 35788 679144 35867 679146
rect 35788 679088 35806 679144
rect 35862 679088 35867 679144
rect 35788 679086 35867 679088
rect 35801 679083 35867 679086
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 40542 678708 40602 678928
rect 41781 678330 41847 678333
rect 41492 678328 41847 678330
rect 41492 678272 41786 678328
rect 41842 678272 41847 678328
rect 41492 678270 41847 678272
rect 41781 678267 41847 678270
rect 42977 677922 43043 677925
rect 41492 677920 43043 677922
rect 41492 677864 42982 677920
rect 43038 677864 43043 677920
rect 41492 677862 43043 677864
rect 42977 677859 43043 677862
rect 40769 677754 40835 677755
rect 40718 677752 40724 677754
rect 40678 677692 40724 677752
rect 40788 677750 40835 677754
rect 40830 677694 40835 677750
rect 40718 677690 40724 677692
rect 40788 677690 40835 677694
rect 40769 677689 40835 677690
rect 42793 677106 42859 677109
rect 41492 677104 42859 677106
rect 41492 677048 42798 677104
rect 42854 677048 42859 677104
rect 41492 677046 42859 677048
rect 42793 677043 42859 677046
rect 675109 676426 675175 676429
rect 676070 676426 676076 676428
rect 675109 676424 676076 676426
rect 675109 676368 675114 676424
rect 675170 676368 676076 676424
rect 675109 676366 676076 676368
rect 675109 676363 675175 676366
rect 676070 676364 676076 676366
rect 676140 676364 676146 676428
rect 42190 673100 42196 673164
rect 42260 673162 42266 673164
rect 42425 673162 42491 673165
rect 42260 673160 42491 673162
rect 42260 673104 42430 673160
rect 42486 673104 42491 673160
rect 42260 673102 42491 673104
rect 42260 673100 42266 673102
rect 42425 673099 42491 673102
rect 33777 672754 33843 672757
rect 41822 672754 41828 672756
rect 33777 672752 41828 672754
rect 33777 672696 33782 672752
rect 33838 672696 41828 672752
rect 33777 672694 41828 672696
rect 33777 672691 33843 672694
rect 41822 672692 41828 672694
rect 41892 672692 41898 672756
rect 673729 671394 673795 671397
rect 673729 671392 676292 671394
rect 673729 671336 673734 671392
rect 673790 671336 676292 671392
rect 673729 671334 676292 671336
rect 673729 671331 673795 671334
rect 39573 670986 39639 670989
rect 40350 670986 40356 670988
rect 39573 670984 40356 670986
rect 39573 670928 39578 670984
rect 39634 670928 40356 670984
rect 39573 670926 40356 670928
rect 39573 670923 39639 670926
rect 40350 670924 40356 670926
rect 40420 670924 40426 670988
rect 673729 670986 673795 670989
rect 673729 670984 676292 670986
rect 673729 670928 673734 670984
rect 673790 670928 676292 670984
rect 673729 670926 676292 670928
rect 673729 670923 673795 670926
rect 673729 670578 673795 670581
rect 673729 670576 676292 670578
rect 673729 670520 673734 670576
rect 673790 670520 676292 670576
rect 673729 670518 676292 670520
rect 673729 670515 673795 670518
rect 672625 670170 672691 670173
rect 672625 670168 676292 670170
rect 672625 670112 672630 670168
rect 672686 670112 676292 670168
rect 672625 670110 676292 670112
rect 672625 670107 672691 670110
rect 673177 669898 673243 669901
rect 674833 669898 674899 669901
rect 673177 669896 674899 669898
rect 673177 669840 673182 669896
rect 673238 669840 674838 669896
rect 674894 669840 674899 669896
rect 673177 669838 674899 669840
rect 673177 669835 673243 669838
rect 674833 669835 674899 669838
rect 676262 669490 676322 669732
rect 676489 669490 676555 669493
rect 675894 669430 676322 669490
rect 676446 669488 676555 669490
rect 676446 669432 676494 669488
rect 676550 669432 676555 669488
rect 673361 669218 673427 669221
rect 675894 669218 675954 669430
rect 676446 669427 676555 669432
rect 676446 669324 676506 669427
rect 673361 669216 675954 669218
rect 673361 669160 673366 669216
rect 673422 669160 675954 669216
rect 673361 669158 675954 669160
rect 673361 669155 673427 669158
rect 673729 668946 673795 668949
rect 673729 668944 676292 668946
rect 673729 668888 673734 668944
rect 673790 668888 676292 668944
rect 673729 668886 676292 668888
rect 673729 668883 673795 668886
rect 41965 668538 42031 668541
rect 42190 668538 42196 668540
rect 41965 668536 42196 668538
rect 41965 668480 41970 668536
rect 42026 668480 42196 668536
rect 41965 668478 42196 668480
rect 41965 668475 42031 668478
rect 42190 668476 42196 668478
rect 42260 668476 42266 668540
rect 673729 668538 673795 668541
rect 673729 668536 676292 668538
rect 673729 668480 673734 668536
rect 673790 668480 676292 668536
rect 673729 668478 676292 668480
rect 673729 668475 673795 668478
rect 673729 668130 673795 668133
rect 673729 668128 676292 668130
rect 673729 668072 673734 668128
rect 673790 668072 676292 668128
rect 673729 668070 676292 668072
rect 673729 668067 673795 668070
rect 42149 667722 42215 667725
rect 45829 667722 45895 667725
rect 42149 667720 45895 667722
rect 42149 667664 42154 667720
rect 42210 667664 45834 667720
rect 45890 667664 45895 667720
rect 42149 667662 45895 667664
rect 42149 667659 42215 667662
rect 45829 667659 45895 667662
rect 673729 667722 673795 667725
rect 673729 667720 676292 667722
rect 673729 667664 673734 667720
rect 673790 667664 676292 667720
rect 673729 667662 676292 667664
rect 673729 667659 673795 667662
rect 40350 667388 40356 667452
rect 40420 667450 40426 667452
rect 42333 667450 42399 667453
rect 40420 667448 42399 667450
rect 40420 667392 42338 667448
rect 42394 667392 42399 667448
rect 40420 667390 42399 667392
rect 40420 667388 40426 667390
rect 42333 667387 42399 667390
rect 676262 667178 676322 667284
rect 673502 667118 676322 667178
rect 42057 667042 42123 667045
rect 45645 667042 45711 667045
rect 42057 667040 45711 667042
rect 42057 666984 42062 667040
rect 42118 666984 45650 667040
rect 45706 666984 45711 667040
rect 42057 666982 45711 666984
rect 42057 666979 42123 666982
rect 45645 666979 45711 666982
rect 673502 666634 673562 667118
rect 673729 666906 673795 666909
rect 673729 666904 676292 666906
rect 673729 666848 673734 666904
rect 673790 666848 676292 666904
rect 673729 666846 676292 666848
rect 673729 666843 673795 666846
rect 673729 666634 673795 666637
rect 673502 666632 673795 666634
rect 673502 666576 673734 666632
rect 673790 666576 673795 666632
rect 673502 666574 673795 666576
rect 673729 666571 673795 666574
rect 675293 666498 675359 666501
rect 675293 666496 676292 666498
rect 675293 666440 675298 666496
rect 675354 666440 676292 666496
rect 675293 666438 676292 666440
rect 675293 666435 675359 666438
rect 684125 666226 684191 666229
rect 684125 666224 684234 666226
rect 684125 666168 684130 666224
rect 684186 666168 684234 666224
rect 684125 666163 684234 666168
rect 684174 666060 684234 666163
rect 676806 665756 676812 665820
rect 676876 665756 676882 665820
rect 676814 665652 676874 665756
rect 40718 665212 40724 665276
rect 40788 665274 40794 665276
rect 41781 665274 41847 665277
rect 40788 665272 41847 665274
rect 40788 665216 41786 665272
rect 41842 665216 41847 665272
rect 40788 665214 41847 665216
rect 40788 665212 40794 665214
rect 41781 665211 41847 665214
rect 673729 665274 673795 665277
rect 673729 665272 676292 665274
rect 673729 665216 673734 665272
rect 673790 665216 676292 665272
rect 673729 665214 676292 665216
rect 673729 665211 673795 665214
rect 676029 664866 676095 664869
rect 676029 664864 676292 664866
rect 676029 664808 676034 664864
rect 676090 664808 676292 664864
rect 676029 664806 676292 664808
rect 676029 664803 676095 664806
rect 673729 664458 673795 664461
rect 673729 664456 676292 664458
rect 673729 664400 673734 664456
rect 673790 664400 676292 664456
rect 673729 664398 676292 664400
rect 673729 664395 673795 664398
rect 40534 664124 40540 664188
rect 40604 664186 40610 664188
rect 41781 664186 41847 664189
rect 40604 664184 41847 664186
rect 40604 664128 41786 664184
rect 41842 664128 41847 664184
rect 40604 664126 41847 664128
rect 40604 664124 40610 664126
rect 41781 664123 41847 664126
rect 673361 664050 673427 664053
rect 673361 664048 676292 664050
rect 673361 663992 673366 664048
rect 673422 663992 676292 664048
rect 673361 663990 676292 663992
rect 673361 663987 673427 663990
rect 673729 663778 673795 663781
rect 674833 663778 674899 663781
rect 673729 663776 674899 663778
rect 673729 663720 673734 663776
rect 673790 663720 674838 663776
rect 674894 663720 674899 663776
rect 673729 663718 674899 663720
rect 673729 663715 673795 663718
rect 674833 663715 674899 663718
rect 683205 663778 683271 663781
rect 683205 663776 683314 663778
rect 683205 663720 683210 663776
rect 683266 663720 683314 663776
rect 683205 663715 683314 663720
rect 683254 663612 683314 663715
rect 673361 662962 673427 662965
rect 676262 662962 676322 663204
rect 683481 662962 683547 662965
rect 673361 662960 676322 662962
rect 673361 662904 673366 662960
rect 673422 662904 676322 662960
rect 673361 662902 676322 662904
rect 683438 662960 683547 662962
rect 683438 662904 683486 662960
rect 683542 662904 683547 662960
rect 673361 662899 673427 662902
rect 683438 662899 683547 662904
rect 683438 662796 683498 662899
rect 674598 662356 674604 662420
rect 674668 662418 674674 662420
rect 674668 662358 676292 662418
rect 674668 662356 674674 662358
rect 673545 662010 673611 662013
rect 673545 662008 676292 662010
rect 673545 661952 673550 662008
rect 673606 661952 676292 662008
rect 673545 661950 676292 661952
rect 673545 661947 673611 661950
rect 673729 661602 673795 661605
rect 673729 661600 676292 661602
rect 673729 661544 673734 661600
rect 673790 661544 676292 661600
rect 673729 661542 676292 661544
rect 673729 661539 673795 661542
rect 673729 661194 673795 661197
rect 673729 661192 676292 661194
rect 673729 661136 673734 661192
rect 673790 661136 676292 661192
rect 673729 661134 676292 661136
rect 673729 661131 673795 661134
rect 62113 660922 62179 660925
rect 62113 660920 64706 660922
rect 62113 660864 62118 660920
rect 62174 660864 64706 660920
rect 62113 660862 64706 660864
rect 62113 660859 62179 660862
rect 64646 660638 64706 660862
rect 683070 660109 683130 660756
rect 673729 660106 673795 660109
rect 674833 660106 674899 660109
rect 673729 660104 674899 660106
rect 673729 660048 673734 660104
rect 673790 660048 674838 660104
rect 674894 660048 674899 660104
rect 673729 660046 674899 660048
rect 683070 660104 683179 660109
rect 683070 660048 683118 660104
rect 683174 660048 683179 660104
rect 683070 660046 683179 660048
rect 673729 660043 673795 660046
rect 674833 660043 674899 660046
rect 683113 660043 683179 660046
rect 673361 659698 673427 659701
rect 676262 659698 676322 659940
rect 673361 659696 676322 659698
rect 673361 659640 673366 659696
rect 673422 659640 676322 659696
rect 673361 659638 676322 659640
rect 673361 659635 673427 659638
rect 62113 659562 62179 659565
rect 62113 659560 64706 659562
rect 62113 659504 62118 659560
rect 62174 659504 64706 659560
rect 62113 659502 64706 659504
rect 62113 659499 62179 659502
rect 64646 659456 64706 659502
rect 41638 658548 41644 658612
rect 41708 658610 41714 658612
rect 42517 658610 42583 658613
rect 41708 658608 42583 658610
rect 41708 658552 42522 658608
rect 42578 658552 42583 658608
rect 41708 658550 42583 658552
rect 41708 658548 41714 658550
rect 42517 658547 42583 658550
rect 41781 658340 41847 658341
rect 41781 658336 41828 658340
rect 41892 658338 41898 658340
rect 62113 658338 62179 658341
rect 41781 658280 41786 658336
rect 41781 658276 41828 658280
rect 41892 658278 41938 658338
rect 62113 658336 64706 658338
rect 62113 658280 62118 658336
rect 62174 658280 64706 658336
rect 62113 658278 64706 658280
rect 41892 658276 41898 658278
rect 41781 658275 41847 658276
rect 62113 658275 62179 658278
rect 64646 658274 64706 658278
rect 63401 657658 63467 657661
rect 63401 657656 64706 657658
rect 63401 657600 63406 657656
rect 63462 657600 64706 657656
rect 63401 657598 64706 657600
rect 63401 657595 63467 657598
rect 41454 657188 41460 657252
rect 41524 657250 41530 657252
rect 41781 657250 41847 657253
rect 41524 657248 41847 657250
rect 41524 657192 41786 657248
rect 41842 657192 41847 657248
rect 41524 657190 41847 657192
rect 41524 657188 41530 657190
rect 41781 657187 41847 657190
rect 64646 657092 64706 657598
rect 62113 656570 62179 656573
rect 62113 656568 64706 656570
rect 62113 656512 62118 656568
rect 62174 656512 64706 656568
rect 62113 656510 64706 656512
rect 62113 656507 62179 656510
rect 64646 655910 64706 656510
rect 673729 655618 673795 655621
rect 675109 655618 675175 655621
rect 673729 655616 675175 655618
rect 673729 655560 673734 655616
rect 673790 655560 675114 655616
rect 675170 655560 675175 655616
rect 673729 655558 675175 655560
rect 673729 655555 673795 655558
rect 675109 655555 675175 655558
rect 62297 655346 62363 655349
rect 62297 655344 64706 655346
rect 62297 655288 62302 655344
rect 62358 655288 64706 655344
rect 62297 655286 64706 655288
rect 62297 655283 62363 655286
rect 64646 654728 64706 655286
rect 674230 652836 674236 652900
rect 674300 652898 674306 652900
rect 675385 652898 675451 652901
rect 674300 652896 675451 652898
rect 674300 652840 675390 652896
rect 675446 652840 675451 652896
rect 674300 652838 675451 652840
rect 674300 652836 674306 652838
rect 675385 652835 675451 652838
rect 672073 652082 672139 652085
rect 675477 652082 675543 652085
rect 672073 652080 675543 652082
rect 672073 652024 672078 652080
rect 672134 652024 675482 652080
rect 675538 652024 675543 652080
rect 672073 652022 675543 652024
rect 672073 652019 672139 652022
rect 675477 652019 675543 652022
rect 672625 649226 672691 649229
rect 675385 649226 675451 649229
rect 672625 649224 675451 649226
rect 672625 649168 672630 649224
rect 672686 649168 675390 649224
rect 675446 649168 675451 649224
rect 672625 649166 675451 649168
rect 672625 649163 672691 649166
rect 675385 649163 675451 649166
rect 672993 648818 673059 648821
rect 675109 648818 675175 648821
rect 672993 648816 675175 648818
rect 672993 648760 672998 648816
rect 673054 648760 675114 648816
rect 675170 648760 675175 648816
rect 672993 648758 675175 648760
rect 672993 648755 673059 648758
rect 675109 648755 675175 648758
rect 671705 647866 671771 647869
rect 675385 647866 675451 647869
rect 671705 647864 675451 647866
rect 671705 647808 671710 647864
rect 671766 647808 675390 647864
rect 675446 647808 675451 647864
rect 671705 647806 675451 647808
rect 671705 647803 671771 647806
rect 675385 647803 675451 647806
rect 673729 645962 673795 645965
rect 675109 645962 675175 645965
rect 673729 645960 675175 645962
rect 673729 645904 673734 645960
rect 673790 645904 675114 645960
rect 675170 645904 675175 645960
rect 673729 645902 675175 645904
rect 673729 645899 673795 645902
rect 675109 645899 675175 645902
rect 673177 645282 673243 645285
rect 675293 645282 675359 645285
rect 673177 645280 675359 645282
rect 673177 645224 673182 645280
rect 673238 645224 675298 645280
rect 675354 645224 675359 645280
rect 673177 645222 675359 645224
rect 673177 645219 673243 645222
rect 675293 645219 675359 645222
rect 35758 644741 35818 644912
rect 35758 644736 35867 644741
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644678 35867 644680
rect 35801 644675 35867 644678
rect 674097 644602 674163 644605
rect 675293 644602 675359 644605
rect 674097 644600 675359 644602
rect 674097 644544 674102 644600
rect 674158 644544 675298 644600
rect 675354 644544 675359 644600
rect 674097 644542 675359 644544
rect 674097 644539 674163 644542
rect 675293 644539 675359 644542
rect 38518 644333 38578 644504
rect 38518 644328 38627 644333
rect 38518 644272 38566 644328
rect 38622 644272 38627 644328
rect 38518 644270 38627 644272
rect 38561 644267 38627 644270
rect 39573 644330 39639 644333
rect 43437 644330 43503 644333
rect 39573 644328 43503 644330
rect 39573 644272 39578 644328
rect 39634 644272 43442 644328
rect 43498 644272 43503 644328
rect 39573 644270 43503 644272
rect 39573 644267 39639 644270
rect 43437 644267 43503 644270
rect 669589 644330 669655 644333
rect 675385 644330 675451 644333
rect 669589 644328 675451 644330
rect 669589 644272 669594 644328
rect 669650 644272 675390 644328
rect 675446 644272 675451 644328
rect 669589 644270 675451 644272
rect 669589 644267 669655 644270
rect 675385 644267 675451 644270
rect 35390 643925 35450 644096
rect 35341 643920 35450 643925
rect 35341 643864 35346 643920
rect 35402 643864 35450 643920
rect 35341 643862 35450 643864
rect 39757 643922 39823 643925
rect 46197 643922 46263 643925
rect 39757 643920 46263 643922
rect 39757 643864 39762 643920
rect 39818 643864 46202 643920
rect 46258 643864 46263 643920
rect 39757 643862 46263 643864
rect 35341 643859 35407 643862
rect 39757 643859 39823 643862
rect 46197 643859 46263 643862
rect 35574 643517 35634 643688
rect 35525 643512 35634 643517
rect 35801 643514 35867 643517
rect 35525 643456 35530 643512
rect 35586 643456 35634 643512
rect 35525 643454 35634 643456
rect 35758 643512 35867 643514
rect 35758 643456 35806 643512
rect 35862 643456 35867 643512
rect 35525 643451 35591 643454
rect 35758 643451 35867 643456
rect 35758 643280 35818 643451
rect 649950 643242 650010 643558
rect 673545 643514 673611 643517
rect 675293 643514 675359 643517
rect 673545 643512 675359 643514
rect 673545 643456 673550 643512
rect 673606 643456 675298 643512
rect 675354 643456 675359 643512
rect 673545 643454 675359 643456
rect 673545 643451 673611 643454
rect 675293 643451 675359 643454
rect 651465 643242 651531 643245
rect 649950 643240 651531 643242
rect 649950 643184 651470 643240
rect 651526 643184 651531 643240
rect 649950 643182 651531 643184
rect 651465 643179 651531 643182
rect 673729 643106 673795 643109
rect 675293 643106 675359 643109
rect 673729 643104 675359 643106
rect 673729 643048 673734 643104
rect 673790 643048 675298 643104
rect 675354 643048 675359 643104
rect 673729 643046 675359 643048
rect 673729 643043 673795 643046
rect 675293 643043 675359 643046
rect 35758 642701 35818 642872
rect 35758 642696 35867 642701
rect 35758 642640 35806 642696
rect 35862 642640 35867 642696
rect 35758 642638 35867 642640
rect 35801 642635 35867 642638
rect 35574 642293 35634 642464
rect 673545 642426 673611 642429
rect 674097 642426 674163 642429
rect 673545 642424 674163 642426
rect 35574 642288 35683 642293
rect 35574 642232 35622 642288
rect 35678 642232 35683 642288
rect 35574 642230 35683 642232
rect 35617 642227 35683 642230
rect 40769 642290 40835 642293
rect 45093 642290 45159 642293
rect 40769 642288 45159 642290
rect 40769 642232 40774 642288
rect 40830 642232 45098 642288
rect 45154 642232 45159 642288
rect 40769 642230 45159 642232
rect 40769 642227 40835 642230
rect 45093 642227 45159 642230
rect 35758 641885 35818 642056
rect 35758 641880 35867 641885
rect 35758 641824 35806 641880
rect 35862 641824 35867 641880
rect 35758 641822 35867 641824
rect 649950 641882 650010 642376
rect 673545 642368 673550 642424
rect 673606 642368 674102 642424
rect 674158 642368 674163 642424
rect 673545 642366 674163 642368
rect 673545 642363 673611 642366
rect 674097 642363 674163 642366
rect 651833 641882 651899 641885
rect 649950 641880 651899 641882
rect 649950 641824 651838 641880
rect 651894 641824 651899 641880
rect 649950 641822 651899 641824
rect 35801 641819 35867 641822
rect 651833 641819 651899 641822
rect 674097 641746 674163 641749
rect 675293 641746 675359 641749
rect 674097 641744 675359 641746
rect 674097 641688 674102 641744
rect 674158 641688 675298 641744
rect 675354 641688 675359 641744
rect 674097 641686 675359 641688
rect 674097 641683 674163 641686
rect 675293 641683 675359 641686
rect 35574 641477 35634 641648
rect 35574 641472 35683 641477
rect 35574 641416 35622 641472
rect 35678 641416 35683 641472
rect 35574 641414 35683 641416
rect 35617 641411 35683 641414
rect 35758 641069 35818 641240
rect 35758 641064 35867 641069
rect 35758 641008 35806 641064
rect 35862 641008 35867 641064
rect 35758 641006 35867 641008
rect 35801 641003 35867 641006
rect 39297 641066 39363 641069
rect 44357 641066 44423 641069
rect 39297 641064 44423 641066
rect 39297 641008 39302 641064
rect 39358 641008 44362 641064
rect 44418 641008 44423 641064
rect 39297 641006 44423 641008
rect 39297 641003 39363 641006
rect 44357 641003 44423 641006
rect 35758 640661 35818 640832
rect 649950 640794 650010 641194
rect 651465 640794 651531 640797
rect 649950 640792 651531 640794
rect 649950 640736 651470 640792
rect 651526 640736 651531 640792
rect 649950 640734 651531 640736
rect 651465 640731 651531 640734
rect 35758 640656 35867 640661
rect 35758 640600 35806 640656
rect 35862 640600 35867 640656
rect 35758 640598 35867 640600
rect 35801 640595 35867 640598
rect 41454 640596 41460 640660
rect 41524 640596 41530 640660
rect 41462 640424 41522 640596
rect 40217 640250 40283 640253
rect 44541 640250 44607 640253
rect 40217 640248 44607 640250
rect 40217 640192 40222 640248
rect 40278 640192 44546 640248
rect 44602 640192 44607 640248
rect 40217 640190 44607 640192
rect 40217 640187 40283 640190
rect 44541 640187 44607 640190
rect 651373 640114 651439 640117
rect 649950 640112 651439 640114
rect 649950 640056 651378 640112
rect 651434 640056 651439 640112
rect 649950 640054 651439 640056
rect 34470 639845 34530 640016
rect 649950 640012 650010 640054
rect 651373 640051 651439 640054
rect 34421 639840 34530 639845
rect 34421 639784 34426 639840
rect 34482 639784 34530 639840
rect 34421 639782 34530 639784
rect 34421 639779 34487 639782
rect 35574 639437 35634 639608
rect 35525 639432 35634 639437
rect 35801 639434 35867 639437
rect 35525 639376 35530 639432
rect 35586 639376 35634 639432
rect 35525 639374 35634 639376
rect 35758 639432 35867 639434
rect 35758 639376 35806 639432
rect 35862 639376 35867 639432
rect 35525 639371 35591 639374
rect 35758 639371 35867 639376
rect 40401 639434 40467 639437
rect 45093 639434 45159 639437
rect 40401 639432 45159 639434
rect 40401 639376 40406 639432
rect 40462 639376 45098 639432
rect 45154 639376 45159 639432
rect 40401 639374 45159 639376
rect 40401 639371 40467 639374
rect 45093 639371 45159 639374
rect 35758 639200 35818 639371
rect 40861 639026 40927 639029
rect 45461 639026 45527 639029
rect 40861 639024 45527 639026
rect 40861 638968 40866 639024
rect 40922 638968 45466 639024
rect 45522 638968 45527 639024
rect 40861 638966 45527 638968
rect 40861 638963 40927 638966
rect 45461 638963 45527 638966
rect 35574 638621 35634 638792
rect 35574 638616 35683 638621
rect 35574 638560 35622 638616
rect 35678 638560 35683 638616
rect 35574 638558 35683 638560
rect 649766 638618 649826 638830
rect 651465 638618 651531 638621
rect 649766 638616 651531 638618
rect 649766 638560 651470 638616
rect 651526 638560 651531 638616
rect 649766 638558 651531 638560
rect 35617 638555 35683 638558
rect 651465 638555 651531 638558
rect 671337 638618 671403 638621
rect 675477 638618 675543 638621
rect 671337 638616 675543 638618
rect 671337 638560 671342 638616
rect 671398 638560 675482 638616
rect 675538 638560 675543 638616
rect 671337 638558 675543 638560
rect 671337 638555 671403 638558
rect 675477 638555 675543 638558
rect 35758 638213 35818 638384
rect 35758 638208 35867 638213
rect 651649 638210 651715 638213
rect 35758 638152 35806 638208
rect 35862 638152 35867 638208
rect 35758 638150 35867 638152
rect 35801 638147 35867 638150
rect 649950 638208 651715 638210
rect 649950 638152 651654 638208
rect 651710 638152 651715 638208
rect 649950 638150 651715 638152
rect 32446 637805 32506 637976
rect 32397 637800 32506 637805
rect 32397 637744 32402 637800
rect 32458 637744 32506 637800
rect 32397 637742 32506 637744
rect 32397 637739 32463 637742
rect 649950 637648 650010 638150
rect 651649 638147 651715 638150
rect 35206 637397 35266 637568
rect 676070 637468 676076 637532
rect 676140 637530 676146 637532
rect 680997 637530 681063 637533
rect 676140 637528 681063 637530
rect 676140 637472 681002 637528
rect 681058 637472 681063 637528
rect 676140 637470 681063 637472
rect 676140 637468 676146 637470
rect 680997 637467 681063 637470
rect 35157 637392 35266 637397
rect 35157 637336 35162 637392
rect 35218 637336 35266 637392
rect 35157 637334 35266 637336
rect 35157 637331 35223 637334
rect 35758 636989 35818 637160
rect 35758 636984 35867 636989
rect 35758 636928 35806 636984
rect 35862 636928 35867 636984
rect 35758 636926 35867 636928
rect 35801 636923 35867 636926
rect 35574 636581 35634 636752
rect 35525 636576 35634 636581
rect 35801 636578 35867 636581
rect 35525 636520 35530 636576
rect 35586 636520 35634 636576
rect 35525 636518 35634 636520
rect 35758 636576 35867 636578
rect 35758 636520 35806 636576
rect 35862 636520 35867 636576
rect 35525 636515 35591 636518
rect 35758 636515 35867 636520
rect 40585 636578 40651 636581
rect 42517 636578 42583 636581
rect 40585 636576 42583 636578
rect 40585 636520 40590 636576
rect 40646 636520 42522 636576
rect 42578 636520 42583 636576
rect 40585 636518 42583 636520
rect 40585 636515 40651 636518
rect 42517 636515 42583 636518
rect 35758 636344 35818 636515
rect 35758 635765 35818 635936
rect 35758 635760 35867 635765
rect 35758 635704 35806 635760
rect 35862 635704 35867 635760
rect 35758 635702 35867 635704
rect 35801 635699 35867 635702
rect 40542 635356 40602 635528
rect 40534 635292 40540 635356
rect 40604 635292 40610 635356
rect 40726 634948 40786 635120
rect 40718 634884 40724 634948
rect 40788 634884 40794 634948
rect 35758 634541 35818 634712
rect 35758 634536 35867 634541
rect 35758 634480 35806 634536
rect 35862 634480 35867 634536
rect 35758 634478 35867 634480
rect 35801 634475 35867 634478
rect 40585 634538 40651 634541
rect 44357 634538 44423 634541
rect 40585 634536 44423 634538
rect 40585 634480 40590 634536
rect 40646 634480 44362 634536
rect 44418 634480 44423 634536
rect 40585 634478 44423 634480
rect 40585 634475 40651 634478
rect 44357 634475 44423 634478
rect 35758 633725 35818 633896
rect 35758 633720 35867 633725
rect 35758 633664 35806 633720
rect 35862 633664 35867 633720
rect 35758 633662 35867 633664
rect 35801 633659 35867 633662
rect 41505 633314 41571 633317
rect 42149 633314 42215 633317
rect 41505 633312 42215 633314
rect 41505 633256 41510 633312
rect 41566 633256 42154 633312
rect 42210 633256 42215 633312
rect 41505 633254 42215 633256
rect 41505 633251 41571 633254
rect 42149 633251 42215 633254
rect 39941 632906 40007 632909
rect 42885 632906 42951 632909
rect 39941 632904 42951 632906
rect 39941 632848 39946 632904
rect 40002 632848 42890 632904
rect 42946 632848 42951 632904
rect 39941 632846 42951 632848
rect 39941 632843 40007 632846
rect 42885 632843 42951 632846
rect 40125 632498 40191 632501
rect 43805 632498 43871 632501
rect 40125 632496 43871 632498
rect 40125 632440 40130 632496
rect 40186 632440 43810 632496
rect 43866 632440 43871 632496
rect 40125 632438 43871 632440
rect 40125 632435 40191 632438
rect 43805 632435 43871 632438
rect 40769 632226 40835 632229
rect 43989 632226 44055 632229
rect 40769 632224 44055 632226
rect 40769 632168 40774 632224
rect 40830 632168 43994 632224
rect 44050 632168 44055 632224
rect 40769 632166 44055 632168
rect 40769 632163 40835 632166
rect 43989 632163 44055 632166
rect 675150 631348 675156 631412
rect 675220 631410 675226 631412
rect 675477 631410 675543 631413
rect 675220 631408 675543 631410
rect 675220 631352 675482 631408
rect 675538 631352 675543 631408
rect 675220 631350 675543 631352
rect 675220 631348 675226 631350
rect 675477 631347 675543 631350
rect 675661 631410 675727 631413
rect 676070 631410 676076 631412
rect 675661 631408 676076 631410
rect 675661 631352 675666 631408
rect 675722 631352 676076 631408
rect 675661 631350 676076 631352
rect 675661 631347 675727 631350
rect 676070 631348 676076 631350
rect 676140 631348 676146 631412
rect 40493 630594 40559 630597
rect 43529 630594 43595 630597
rect 40493 630592 43595 630594
rect 40493 630536 40498 630592
rect 40554 630536 43534 630592
rect 43590 630536 43595 630592
rect 40493 630534 43595 630536
rect 40493 630531 40559 630534
rect 43529 630531 43595 630534
rect 32397 629914 32463 629917
rect 41638 629914 41644 629916
rect 32397 629912 41644 629914
rect 32397 629856 32402 629912
rect 32458 629856 41644 629912
rect 32397 629854 41644 629856
rect 32397 629851 32463 629854
rect 41638 629852 41644 629854
rect 41708 629852 41714 629916
rect 39297 629234 39363 629237
rect 41822 629234 41828 629236
rect 39297 629232 41828 629234
rect 39297 629176 39302 629232
rect 39358 629176 41828 629232
rect 39297 629174 41828 629176
rect 39297 629171 39363 629174
rect 41822 629172 41828 629174
rect 41892 629172 41898 629236
rect 39665 628282 39731 628285
rect 42701 628282 42767 628285
rect 39665 628280 42767 628282
rect 39665 628224 39670 628280
rect 39726 628224 42706 628280
rect 42762 628224 42767 628280
rect 39665 628222 42767 628224
rect 39665 628219 39731 628222
rect 42701 628219 42767 628222
rect 41781 627464 41847 627469
rect 41781 627408 41786 627464
rect 41842 627408 41847 627464
rect 41781 627403 41847 627408
rect 41784 627197 41844 627403
rect 41781 627192 41847 627197
rect 41781 627136 41786 627192
rect 41842 627136 41847 627192
rect 41781 627131 41847 627136
rect 672809 626378 672875 626381
rect 672809 626376 676292 626378
rect 672809 626320 672814 626376
rect 672870 626320 676292 626376
rect 672809 626318 676292 626320
rect 672809 626315 672875 626318
rect 42190 625908 42196 625972
rect 42260 625970 42266 625972
rect 42517 625970 42583 625973
rect 42260 625968 42583 625970
rect 42260 625912 42522 625968
rect 42578 625912 42583 625968
rect 42260 625910 42583 625912
rect 42260 625908 42266 625910
rect 42517 625907 42583 625910
rect 672809 625970 672875 625973
rect 672809 625968 676292 625970
rect 672809 625912 672814 625968
rect 672870 625912 676292 625968
rect 672809 625910 676292 625912
rect 672809 625907 672875 625910
rect 672165 625562 672231 625565
rect 672165 625560 676292 625562
rect 672165 625504 672170 625560
rect 672226 625504 676292 625560
rect 672165 625502 676292 625504
rect 672165 625499 672231 625502
rect 674054 625094 676292 625154
rect 672809 625018 672875 625021
rect 674054 625018 674114 625094
rect 672809 625016 674114 625018
rect 672809 624960 672814 625016
rect 672870 624960 674114 625016
rect 672809 624958 674114 624960
rect 672809 624955 672875 624958
rect 672809 624746 672875 624749
rect 672809 624744 676292 624746
rect 672809 624688 672814 624744
rect 672870 624688 676292 624744
rect 672809 624686 676292 624688
rect 672809 624683 672875 624686
rect 42149 624610 42215 624613
rect 44173 624610 44239 624613
rect 42149 624608 44239 624610
rect 42149 624552 42154 624608
rect 42210 624552 44178 624608
rect 44234 624552 44239 624608
rect 42149 624550 44239 624552
rect 42149 624547 42215 624550
rect 44173 624547 44239 624550
rect 672809 624338 672875 624341
rect 672809 624336 676292 624338
rect 672809 624280 672814 624336
rect 672870 624280 676292 624336
rect 672809 624278 676292 624280
rect 672809 624275 672875 624278
rect 672809 623930 672875 623933
rect 672809 623928 676292 623930
rect 672809 623872 672814 623928
rect 672870 623872 676292 623928
rect 672809 623870 676292 623872
rect 672809 623867 672875 623870
rect 40718 623732 40724 623796
rect 40788 623794 40794 623796
rect 40788 623734 42074 623794
rect 40788 623732 40794 623734
rect 42014 623389 42074 623734
rect 672809 623522 672875 623525
rect 672809 623520 676292 623522
rect 672809 623464 672814 623520
rect 672870 623464 676292 623520
rect 672809 623462 676292 623464
rect 672809 623459 672875 623462
rect 41965 623384 42074 623389
rect 41965 623328 41970 623384
rect 42026 623328 42074 623384
rect 41965 623326 42074 623328
rect 41965 623323 42031 623326
rect 672809 623114 672875 623117
rect 672809 623112 676292 623114
rect 672809 623056 672814 623112
rect 672870 623056 676292 623112
rect 672809 623054 676292 623056
rect 672809 623051 672875 623054
rect 671981 622842 672047 622845
rect 671981 622840 676230 622842
rect 671981 622784 671986 622840
rect 672042 622784 676230 622840
rect 671981 622782 676230 622784
rect 671981 622779 672047 622782
rect 676170 622706 676230 622782
rect 676170 622646 676292 622706
rect 42057 622162 42123 622165
rect 44173 622162 44239 622165
rect 42057 622160 44239 622162
rect 42057 622104 42062 622160
rect 42118 622104 44178 622160
rect 44234 622104 44239 622160
rect 42057 622102 44239 622104
rect 42057 622099 42123 622102
rect 44173 622099 44239 622102
rect 676262 622029 676322 622268
rect 676213 622024 676322 622029
rect 676213 621968 676218 622024
rect 676274 621968 676322 622024
rect 676213 621966 676322 621968
rect 680997 622026 681063 622029
rect 680997 622024 681106 622026
rect 680997 621968 681002 622024
rect 681058 621968 681106 622024
rect 676213 621963 676279 621966
rect 680997 621963 681106 621968
rect 681046 621860 681106 621963
rect 672901 621482 672967 621485
rect 672901 621480 676292 621482
rect 672901 621424 672906 621480
rect 672962 621424 676292 621480
rect 672901 621422 676292 621424
rect 672901 621419 672967 621422
rect 672809 621074 672875 621077
rect 672809 621072 676292 621074
rect 672809 621016 672814 621072
rect 672870 621016 676292 621072
rect 672809 621014 676292 621016
rect 672809 621011 672875 621014
rect 40534 620876 40540 620940
rect 40604 620938 40610 620940
rect 41781 620938 41847 620941
rect 40604 620936 41847 620938
rect 40604 620880 41786 620936
rect 41842 620880 41847 620936
rect 40604 620878 41847 620880
rect 40604 620876 40610 620878
rect 41781 620875 41847 620878
rect 671429 620802 671495 620805
rect 674281 620802 674347 620805
rect 671429 620800 674347 620802
rect 671429 620744 671434 620800
rect 671490 620744 674286 620800
rect 674342 620744 674347 620800
rect 671429 620742 674347 620744
rect 671429 620739 671495 620742
rect 674281 620739 674347 620742
rect 676029 620666 676095 620669
rect 676029 620664 676292 620666
rect 676029 620608 676034 620664
rect 676090 620608 676292 620664
rect 676029 620606 676292 620608
rect 676029 620603 676095 620606
rect 41965 620258 42031 620261
rect 42190 620258 42196 620260
rect 41965 620256 42196 620258
rect 41965 620200 41970 620256
rect 42026 620200 42196 620256
rect 41965 620198 42196 620200
rect 41965 620195 42031 620198
rect 42190 620196 42196 620198
rect 42260 620196 42266 620260
rect 672809 620258 672875 620261
rect 672809 620256 676292 620258
rect 672809 620200 672814 620256
rect 672870 620200 676292 620256
rect 672809 620198 676292 620200
rect 672809 620195 672875 620198
rect 672809 619986 672875 619989
rect 672809 619984 676322 619986
rect 672809 619928 672814 619984
rect 672870 619928 676322 619984
rect 672809 619926 676322 619928
rect 672809 619923 672875 619926
rect 676262 619820 676322 619926
rect 672809 619714 672875 619717
rect 674373 619714 674439 619717
rect 672809 619712 674439 619714
rect 672809 619656 672814 619712
rect 672870 619656 674378 619712
rect 674434 619656 674439 619712
rect 672809 619654 674439 619656
rect 672809 619651 672875 619654
rect 674373 619651 674439 619654
rect 676262 619173 676322 619412
rect 676213 619168 676322 619173
rect 676213 619112 676218 619168
rect 676274 619112 676322 619168
rect 676213 619110 676322 619112
rect 676213 619107 676279 619110
rect 674414 618700 674420 618764
rect 674484 618762 674490 618764
rect 676446 618762 676506 619004
rect 674484 618702 676506 618762
rect 683205 618762 683271 618765
rect 683205 618760 683314 618762
rect 683205 618704 683210 618760
rect 683266 618704 683314 618760
rect 674484 618700 674490 618702
rect 683205 618699 683314 618704
rect 683254 618596 683314 618699
rect 672257 618490 672323 618493
rect 674281 618490 674347 618493
rect 672257 618488 674347 618490
rect 672257 618432 672262 618488
rect 672318 618432 674286 618488
rect 674342 618432 674347 618488
rect 672257 618430 674347 618432
rect 672257 618427 672323 618430
rect 674281 618427 674347 618430
rect 63125 618082 63191 618085
rect 63125 618080 64706 618082
rect 63125 618024 63130 618080
rect 63186 618024 64706 618080
rect 63125 618022 64706 618024
rect 63125 618019 63191 618022
rect 64646 617416 64706 618022
rect 676262 617949 676322 618188
rect 676213 617944 676322 617949
rect 676213 617888 676218 617944
rect 676274 617888 676322 617944
rect 676213 617886 676322 617888
rect 676213 617883 676279 617886
rect 676262 617541 676322 617780
rect 676213 617536 676322 617541
rect 676489 617538 676555 617541
rect 676213 617480 676218 617536
rect 676274 617480 676322 617536
rect 676213 617478 676322 617480
rect 676446 617536 676555 617538
rect 676446 617480 676494 617536
rect 676550 617480 676555 617536
rect 676213 617475 676279 617478
rect 676446 617475 676555 617480
rect 676446 617372 676506 617475
rect 675293 617130 675359 617133
rect 676254 617130 676260 617132
rect 675293 617128 676260 617130
rect 675293 617072 675298 617128
rect 675354 617072 676260 617128
rect 675293 617070 676260 617072
rect 675293 617067 675359 617070
rect 676254 617068 676260 617070
rect 676324 617068 676330 617132
rect 683573 617130 683639 617133
rect 683573 617128 683682 617130
rect 683573 617072 683578 617128
rect 683634 617072 683682 617128
rect 683573 617067 683682 617072
rect 683622 616964 683682 617067
rect 41638 616796 41644 616860
rect 41708 616858 41714 616860
rect 42701 616858 42767 616861
rect 41708 616856 42767 616858
rect 41708 616800 42706 616856
rect 42762 616800 42767 616856
rect 41708 616798 42767 616800
rect 41708 616796 41714 616798
rect 42701 616795 42767 616798
rect 683389 616722 683455 616725
rect 683389 616720 683498 616722
rect 683389 616664 683394 616720
rect 683450 616664 683498 616720
rect 683389 616659 683498 616664
rect 62113 616586 62179 616589
rect 62113 616584 64706 616586
rect 62113 616528 62118 616584
rect 62174 616528 64706 616584
rect 683438 616556 683498 616659
rect 62113 616526 64706 616528
rect 62113 616523 62179 616526
rect 41454 616388 41460 616452
rect 41524 616450 41530 616452
rect 42425 616450 42491 616453
rect 41524 616448 42491 616450
rect 41524 616392 42430 616448
rect 42486 616392 42491 616448
rect 41524 616390 42491 616392
rect 41524 616388 41530 616390
rect 42425 616387 42491 616390
rect 64646 616234 64706 616526
rect 673862 616116 673868 616180
rect 673932 616178 673938 616180
rect 673932 616118 676292 616178
rect 673932 616116 673938 616118
rect 42057 615906 42123 615909
rect 42609 615906 42675 615909
rect 42057 615904 42675 615906
rect 42057 615848 42062 615904
rect 42118 615848 42614 615904
rect 42670 615848 42675 615904
rect 42057 615846 42675 615848
rect 42057 615843 42123 615846
rect 42609 615843 42675 615846
rect 683070 615501 683130 615740
rect 41822 615436 41828 615500
rect 41892 615498 41898 615500
rect 42701 615498 42767 615501
rect 41892 615496 42767 615498
rect 41892 615440 42706 615496
rect 42762 615440 42767 615496
rect 41892 615438 42767 615440
rect 41892 615436 41898 615438
rect 42701 615435 42767 615438
rect 683070 615498 683179 615501
rect 683070 615496 683260 615498
rect 683070 615440 683118 615496
rect 683174 615440 683260 615496
rect 683070 615438 683260 615440
rect 683070 615435 683179 615438
rect 683070 615332 683130 615435
rect 62113 614682 62179 614685
rect 64646 614682 64706 615052
rect 676262 614685 676322 614924
rect 62113 614680 64706 614682
rect 62113 614624 62118 614680
rect 62174 614624 64706 614680
rect 62113 614622 64706 614624
rect 676213 614680 676322 614685
rect 676213 614624 676218 614680
rect 676274 614624 676322 614680
rect 676213 614622 676322 614624
rect 62113 614619 62179 614622
rect 676213 614619 676279 614622
rect 62113 613866 62179 613869
rect 64646 613866 64706 613870
rect 62113 613864 64706 613866
rect 62113 613808 62118 613864
rect 62174 613808 64706 613864
rect 62113 613806 64706 613808
rect 62113 613803 62179 613806
rect 62113 612642 62179 612645
rect 64646 612642 64706 612688
rect 62113 612640 64706 612642
rect 62113 612584 62118 612640
rect 62174 612584 64706 612640
rect 62113 612582 64706 612584
rect 62113 612579 62179 612582
rect 40534 612308 40540 612372
rect 40604 612370 40610 612372
rect 42241 612370 42307 612373
rect 40604 612368 42307 612370
rect 40604 612312 42246 612368
rect 42302 612312 42307 612368
rect 40604 612310 42307 612312
rect 40604 612308 40610 612310
rect 42241 612307 42307 612310
rect 62941 612098 63007 612101
rect 62941 612096 64706 612098
rect 62941 612040 62946 612096
rect 63002 612040 64706 612096
rect 62941 612038 64706 612040
rect 62941 612035 63007 612038
rect 64646 611506 64706 612038
rect 43529 611010 43595 611013
rect 44725 611010 44791 611013
rect 43529 611008 44791 611010
rect 43529 610952 43534 611008
rect 43590 610952 44730 611008
rect 44786 610952 44791 611008
rect 43529 610950 44791 610952
rect 43529 610947 43595 610950
rect 44725 610947 44791 610950
rect 674005 608018 674071 608021
rect 675385 608018 675451 608021
rect 674005 608016 675451 608018
rect 674005 607960 674010 608016
rect 674066 607960 675390 608016
rect 675446 607960 675451 608016
rect 674005 607958 675451 607960
rect 674005 607955 674071 607958
rect 675385 607955 675451 607958
rect 670969 607746 671035 607749
rect 675477 607746 675543 607749
rect 670969 607744 675543 607746
rect 670969 607688 670974 607744
rect 671030 607688 675482 607744
rect 675538 607688 675543 607744
rect 670969 607686 675543 607688
rect 670969 607683 671035 607686
rect 675477 607683 675543 607686
rect 672441 604482 672507 604485
rect 675109 604482 675175 604485
rect 672441 604480 675175 604482
rect 672441 604424 672446 604480
rect 672502 604424 675114 604480
rect 675170 604424 675175 604480
rect 672441 604422 675175 604424
rect 672441 604419 672507 604422
rect 675109 604419 675175 604422
rect 674414 602924 674420 602988
rect 674484 602986 674490 602988
rect 675109 602986 675175 602989
rect 674484 602984 675175 602986
rect 674484 602928 675114 602984
rect 675170 602928 675175 602984
rect 674484 602926 675175 602928
rect 674484 602924 674490 602926
rect 675109 602923 675175 602926
rect 40309 602034 40375 602037
rect 40534 602034 40540 602036
rect 40309 602032 40540 602034
rect 40309 601976 40314 602032
rect 40370 601976 40540 602032
rect 40309 601974 40540 601976
rect 40309 601971 40375 601974
rect 40534 601972 40540 601974
rect 40604 601972 40610 602036
rect 33777 601762 33843 601765
rect 33764 601760 33843 601762
rect 33764 601704 33782 601760
rect 33838 601704 33843 601760
rect 33764 601702 33843 601704
rect 33777 601699 33843 601702
rect 39941 601354 40007 601357
rect 39941 601352 40020 601354
rect 39941 601296 39946 601352
rect 40002 601296 40020 601352
rect 39941 601294 40020 601296
rect 39941 601291 40007 601294
rect 40125 600946 40191 600949
rect 667381 600946 667447 600949
rect 675385 600946 675451 600949
rect 40125 600944 40204 600946
rect 40125 600888 40130 600944
rect 40186 600888 40204 600944
rect 40125 600886 40204 600888
rect 667381 600944 675451 600946
rect 667381 600888 667386 600944
rect 667442 600888 675390 600944
rect 675446 600888 675451 600944
rect 667381 600886 675451 600888
rect 40125 600883 40191 600886
rect 667381 600883 667447 600886
rect 675385 600883 675451 600886
rect 44541 600538 44607 600541
rect 41492 600536 44607 600538
rect 41492 600480 44546 600536
rect 44602 600480 44607 600536
rect 41492 600478 44607 600480
rect 44541 600475 44607 600478
rect 674005 600402 674071 600405
rect 675109 600402 675175 600405
rect 674005 600400 675175 600402
rect 674005 600344 674010 600400
rect 674066 600344 675114 600400
rect 675170 600344 675175 600400
rect 674005 600342 675175 600344
rect 674005 600339 674071 600342
rect 675109 600339 675175 600342
rect 44909 600130 44975 600133
rect 41492 600128 44975 600130
rect 41492 600072 44914 600128
rect 44970 600072 44975 600128
rect 41492 600070 44975 600072
rect 44909 600067 44975 600070
rect 45277 599722 45343 599725
rect 41492 599720 45343 599722
rect 41492 599664 45282 599720
rect 45338 599664 45343 599720
rect 41492 599662 45343 599664
rect 45277 599659 45343 599662
rect 674005 599722 674071 599725
rect 675477 599722 675543 599725
rect 674005 599720 675543 599722
rect 674005 599664 674010 599720
rect 674066 599664 675482 599720
rect 675538 599664 675543 599720
rect 674005 599662 675543 599664
rect 674005 599659 674071 599662
rect 675477 599659 675543 599662
rect 44633 599314 44699 599317
rect 41492 599312 44699 599314
rect 41492 599256 44638 599312
rect 44694 599256 44699 599312
rect 41492 599254 44699 599256
rect 44633 599251 44699 599254
rect 45461 598906 45527 598909
rect 41492 598904 45527 598906
rect 41492 598848 45466 598904
rect 45522 598848 45527 598904
rect 41492 598846 45527 598848
rect 45461 598843 45527 598846
rect 42926 598498 42932 598500
rect 41492 598438 42932 598498
rect 42926 598436 42932 598438
rect 42996 598436 43002 598500
rect 45093 598090 45159 598093
rect 41492 598088 45159 598090
rect 41492 598032 45098 598088
rect 45154 598032 45159 598088
rect 41492 598030 45159 598032
rect 45093 598027 45159 598030
rect 649950 597954 650010 598336
rect 674005 598090 674071 598093
rect 675109 598090 675175 598093
rect 674005 598088 675175 598090
rect 674005 598032 674010 598088
rect 674066 598032 675114 598088
rect 675170 598032 675175 598088
rect 674005 598030 675175 598032
rect 674005 598027 674071 598030
rect 675109 598027 675175 598030
rect 651465 597954 651531 597957
rect 649950 597952 651531 597954
rect 649950 597896 651470 597952
rect 651526 597896 651531 597952
rect 649950 597894 651531 597896
rect 651465 597891 651531 597894
rect 43069 597682 43135 597685
rect 41492 597680 43135 597682
rect 41492 597624 43074 597680
rect 43130 597624 43135 597680
rect 41492 597622 43135 597624
rect 43069 597619 43135 597622
rect 672809 597410 672875 597413
rect 675385 597410 675451 597413
rect 672809 597408 675451 597410
rect 672809 597352 672814 597408
rect 672870 597352 675390 597408
rect 675446 597352 675451 597408
rect 672809 597350 675451 597352
rect 672809 597347 672875 597350
rect 675385 597347 675451 597350
rect 40358 597038 40418 597244
rect 40350 596974 40356 597038
rect 40420 596974 40426 597038
rect 42885 597004 42951 597005
rect 42885 597000 42932 597004
rect 42996 597002 43002 597004
rect 42885 596944 42890 597000
rect 42885 596940 42932 596944
rect 42996 596942 43042 597002
rect 42996 596940 43002 596942
rect 42885 596939 42951 596940
rect 42425 596866 42491 596869
rect 41492 596864 42491 596866
rect 41492 596808 42430 596864
rect 42486 596808 42491 596864
rect 41492 596806 42491 596808
rect 42425 596803 42491 596806
rect 649950 596730 650010 597154
rect 673913 597138 673979 597141
rect 674465 597138 674531 597141
rect 673913 597136 674531 597138
rect 673913 597080 673918 597136
rect 673974 597080 674470 597136
rect 674526 597080 674531 597136
rect 673913 597078 674531 597080
rect 673913 597075 673979 597078
rect 674465 597075 674531 597078
rect 673545 596866 673611 596869
rect 674465 596866 674531 596869
rect 673545 596864 674531 596866
rect 673545 596808 673550 596864
rect 673606 596808 674470 596864
rect 674526 596808 674531 596864
rect 673545 596806 674531 596808
rect 673545 596803 673611 596806
rect 674465 596803 674531 596806
rect 651465 596730 651531 596733
rect 649950 596728 651531 596730
rect 649950 596672 651470 596728
rect 651526 596672 651531 596728
rect 649950 596670 651531 596672
rect 651465 596667 651531 596670
rect 42006 596458 42012 596460
rect 41492 596398 42012 596458
rect 42006 596396 42012 596398
rect 42076 596396 42082 596460
rect 41278 595815 41338 596020
rect 37917 595812 37983 595815
rect 37917 595810 38026 595812
rect 37917 595754 37922 595810
rect 37978 595754 38026 595810
rect 37917 595749 38026 595754
rect 41278 595810 41387 595815
rect 41278 595754 41326 595810
rect 41382 595754 41387 595810
rect 41278 595752 41387 595754
rect 41321 595749 41387 595752
rect 41689 595778 41755 595781
rect 62757 595778 62823 595781
rect 41689 595776 62823 595778
rect 37966 595612 38026 595749
rect 41689 595720 41694 595776
rect 41750 595720 62762 595776
rect 62818 595720 62823 595776
rect 41689 595718 62823 595720
rect 41689 595715 41755 595718
rect 62757 595715 62823 595718
rect 649950 595370 650010 595972
rect 651465 595370 651531 595373
rect 649950 595368 651531 595370
rect 649950 595312 651470 595368
rect 651526 595312 651531 595368
rect 649950 595310 651531 595312
rect 651465 595307 651531 595310
rect 33041 595234 33107 595237
rect 33028 595232 33107 595234
rect 33028 595176 33046 595232
rect 33102 595176 33107 595232
rect 33028 595174 33107 595176
rect 33041 595171 33107 595174
rect 651649 595098 651715 595101
rect 649950 595096 651715 595098
rect 649950 595040 651654 595096
rect 651710 595040 651715 595096
rect 649950 595038 651715 595040
rect 35157 594826 35223 594829
rect 35157 594824 35236 594826
rect 35157 594768 35162 594824
rect 35218 594768 35236 594824
rect 649950 594790 650010 595038
rect 651649 595035 651715 595038
rect 667565 594826 667631 594829
rect 675477 594826 675543 594829
rect 667565 594824 675543 594826
rect 35157 594766 35236 594768
rect 667565 594768 667570 594824
rect 667626 594768 675482 594824
rect 675538 594768 675543 594824
rect 667565 594766 675543 594768
rect 35157 594763 35223 594766
rect 667565 594763 667631 594766
rect 675477 594763 675543 594766
rect 41689 594554 41755 594557
rect 41689 594552 48330 594554
rect 41689 594496 41694 594552
rect 41750 594496 48330 594552
rect 41689 594494 48330 594496
rect 41689 594491 41755 594494
rect 31017 594418 31083 594421
rect 31004 594416 31083 594418
rect 31004 594360 31022 594416
rect 31078 594360 31083 594416
rect 31004 594358 31083 594360
rect 31017 594355 31083 594358
rect 48270 594146 48330 594494
rect 63125 594146 63191 594149
rect 651465 594146 651531 594149
rect 48270 594144 63191 594146
rect 48270 594088 63130 594144
rect 63186 594088 63191 594144
rect 48270 594086 63191 594088
rect 63125 594083 63191 594086
rect 649950 594144 651531 594146
rect 649950 594088 651470 594144
rect 651526 594088 651531 594144
rect 649950 594086 651531 594088
rect 41776 594010 41782 594012
rect 41492 593950 41782 594010
rect 41776 593948 41782 593950
rect 41846 593948 41852 594012
rect 649950 593608 650010 594086
rect 651465 594083 651531 594086
rect 41781 593602 41847 593605
rect 41492 593600 41847 593602
rect 41492 593544 41786 593600
rect 41842 593544 41847 593600
rect 41492 593542 41847 593544
rect 41781 593539 41847 593542
rect 668853 593602 668919 593605
rect 675477 593602 675543 593605
rect 668853 593600 675543 593602
rect 668853 593544 668858 593600
rect 668914 593544 675482 593600
rect 675538 593544 675543 593600
rect 668853 593542 675543 593544
rect 668853 593539 668919 593542
rect 675477 593539 675543 593542
rect 44357 593194 44423 593197
rect 41492 593192 44423 593194
rect 41492 593136 44362 593192
rect 44418 593136 44423 593192
rect 41492 593134 44423 593136
rect 44357 593131 44423 593134
rect 675150 593132 675156 593196
rect 675220 593194 675226 593196
rect 675477 593194 675543 593197
rect 675220 593192 675543 593194
rect 675220 593136 675482 593192
rect 675538 593136 675543 593192
rect 675220 593134 675543 593136
rect 675220 593132 675226 593134
rect 675477 593131 675543 593134
rect 651465 592922 651531 592925
rect 649950 592920 651531 592922
rect 649950 592864 651470 592920
rect 651526 592864 651531 592920
rect 649950 592862 651531 592864
rect 41776 592786 41782 592788
rect 41492 592726 41782 592786
rect 41776 592724 41782 592726
rect 41846 592724 41852 592788
rect 649950 592426 650010 592862
rect 651465 592859 651531 592862
rect 41781 592378 41847 592381
rect 41492 592376 41847 592378
rect 41492 592320 41786 592376
rect 41842 592320 41847 592376
rect 41492 592318 41847 592320
rect 41781 592315 41847 592318
rect 35617 591970 35683 591973
rect 35604 591968 35683 591970
rect 35604 591912 35622 591968
rect 35678 591912 35683 591968
rect 35604 591910 35683 591912
rect 35617 591907 35683 591910
rect 676070 591636 676076 591700
rect 676140 591698 676146 591700
rect 680997 591698 681063 591701
rect 676140 591696 681063 591698
rect 676140 591640 681002 591696
rect 681058 591640 681063 591696
rect 676140 591638 681063 591640
rect 676140 591636 676146 591638
rect 680997 591635 681063 591638
rect 35801 591562 35867 591565
rect 35788 591560 35867 591562
rect 35788 591504 35806 591560
rect 35862 591504 35867 591560
rect 35788 591502 35867 591504
rect 35801 591499 35867 591502
rect 674230 591228 674236 591292
rect 674300 591290 674306 591292
rect 684217 591290 684283 591293
rect 674300 591288 684283 591290
rect 674300 591232 684222 591288
rect 684278 591232 684283 591288
rect 674300 591230 684283 591232
rect 674300 591228 674306 591230
rect 684217 591227 684283 591230
rect 41462 590746 41522 591124
rect 62941 590746 63007 590749
rect 41462 590744 63007 590746
rect 41462 590716 62946 590744
rect 41492 590688 62946 590716
rect 63002 590688 63007 590744
rect 41492 590686 63007 590688
rect 62941 590683 63007 590686
rect 62573 590066 62639 590069
rect 51030 590064 62639 590066
rect 51030 590008 62578 590064
rect 62634 590008 62639 590064
rect 51030 590006 62639 590008
rect 33777 589658 33843 589661
rect 51030 589658 51090 590006
rect 62573 590003 62639 590006
rect 33777 589656 51090 589658
rect 33777 589600 33782 589656
rect 33838 589600 51090 589656
rect 33777 589598 51090 589600
rect 33777 589595 33843 589598
rect 40769 589386 40835 589389
rect 43437 589386 43503 589389
rect 40769 589384 43503 589386
rect 40769 589328 40774 589384
rect 40830 589328 43442 589384
rect 43498 589328 43503 589384
rect 40769 589326 43503 589328
rect 40769 589323 40835 589326
rect 43437 589323 43503 589326
rect 40902 589052 40908 589116
rect 40972 589114 40978 589116
rect 41505 589114 41571 589117
rect 40972 589112 41571 589114
rect 40972 589056 41510 589112
rect 41566 589056 41571 589112
rect 40972 589054 41571 589056
rect 40972 589052 40978 589054
rect 41505 589051 41571 589054
rect 40350 588780 40356 588844
rect 40420 588842 40426 588844
rect 41454 588842 41460 588844
rect 40420 588782 41460 588842
rect 40420 588780 40426 588782
rect 41454 588780 41460 588782
rect 41524 588780 41530 588844
rect 675201 586258 675267 586261
rect 676070 586258 676076 586260
rect 675201 586256 676076 586258
rect 675201 586200 675206 586256
rect 675262 586200 676076 586256
rect 675201 586198 676076 586200
rect 675201 586195 675267 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 35157 585986 35223 585989
rect 41822 585986 41828 585988
rect 35157 585984 41828 585986
rect 35157 585928 35162 585984
rect 35218 585928 41828 585984
rect 35157 585926 41828 585928
rect 35157 585923 35223 585926
rect 41822 585924 41828 585926
rect 41892 585924 41898 585988
rect 40401 585714 40467 585717
rect 62062 585714 62068 585716
rect 40401 585712 62068 585714
rect 40401 585656 40406 585712
rect 40462 585656 62068 585712
rect 40401 585654 62068 585656
rect 40401 585651 40467 585654
rect 62062 585652 62068 585654
rect 62132 585652 62138 585716
rect 39297 584626 39363 584629
rect 40350 584626 40356 584628
rect 39297 584624 40356 584626
rect 39297 584568 39302 584624
rect 39358 584568 40356 584624
rect 39297 584566 40356 584568
rect 39297 584563 39363 584566
rect 40350 584564 40356 584566
rect 40420 584564 40426 584628
rect 41781 584352 41847 584357
rect 41781 584296 41786 584352
rect 41842 584296 41847 584352
rect 41781 584291 41847 584296
rect 41784 583949 41844 584291
rect 41781 583944 41847 583949
rect 41781 583888 41786 583944
rect 41842 583888 41847 583944
rect 41781 583883 41847 583888
rect 42241 582452 42307 582453
rect 42190 582450 42196 582452
rect 42150 582390 42196 582450
rect 42260 582448 42307 582452
rect 42302 582392 42307 582448
rect 42190 582388 42196 582390
rect 42260 582388 42307 582392
rect 42241 582387 42307 582388
rect 673637 581362 673703 581365
rect 674465 581362 674531 581365
rect 673637 581360 674531 581362
rect 673637 581304 673642 581360
rect 673698 581304 674470 581360
rect 674526 581304 674531 581360
rect 673637 581302 674531 581304
rect 673637 581299 673703 581302
rect 674465 581299 674531 581302
rect 43621 581226 43687 581229
rect 51717 581226 51783 581229
rect 43621 581224 51783 581226
rect 43621 581168 43626 581224
rect 43682 581168 51722 581224
rect 51778 581168 51783 581224
rect 43621 581166 51783 581168
rect 43621 581163 43687 581166
rect 51717 581163 51783 581166
rect 673637 581090 673703 581093
rect 673637 581088 676292 581090
rect 673637 581032 673642 581088
rect 673698 581032 676292 581088
rect 673637 581030 676292 581032
rect 673637 581027 673703 581030
rect 42057 580682 42123 580685
rect 45093 580682 45159 580685
rect 42057 580680 45159 580682
rect 42057 580624 42062 580680
rect 42118 580624 45098 580680
rect 45154 580624 45159 580680
rect 42057 580622 45159 580624
rect 42057 580619 42123 580622
rect 45093 580619 45159 580622
rect 673085 580682 673151 580685
rect 673085 580680 676292 580682
rect 673085 580624 673090 580680
rect 673146 580624 676292 580680
rect 673085 580622 676292 580624
rect 673085 580619 673151 580622
rect 40350 580212 40356 580276
rect 40420 580274 40426 580276
rect 41873 580274 41939 580277
rect 42241 580276 42307 580277
rect 40420 580272 41939 580274
rect 40420 580216 41878 580272
rect 41934 580216 41939 580272
rect 40420 580214 41939 580216
rect 40420 580212 40426 580214
rect 41873 580211 41939 580214
rect 42190 580212 42196 580276
rect 42260 580274 42307 580276
rect 673637 580274 673703 580277
rect 42260 580272 42352 580274
rect 42302 580216 42352 580272
rect 42260 580214 42352 580216
rect 673637 580272 676292 580274
rect 673637 580216 673642 580272
rect 673698 580216 676292 580272
rect 673637 580214 676292 580216
rect 42260 580212 42307 580214
rect 42241 580211 42307 580212
rect 673637 580211 673703 580214
rect 43621 579866 43687 579869
rect 41830 579864 43687 579866
rect 41830 579808 43626 579864
rect 43682 579808 43687 579864
rect 41830 579806 43687 579808
rect 41830 579597 41890 579806
rect 43621 579803 43687 579806
rect 673637 579866 673703 579869
rect 673637 579864 676292 579866
rect 673637 579808 673642 579864
rect 673698 579808 676292 579864
rect 673637 579806 676292 579808
rect 673637 579803 673703 579806
rect 41781 579592 41890 579597
rect 41781 579536 41786 579592
rect 41842 579536 41890 579592
rect 41781 579534 41890 579536
rect 41781 579531 41847 579534
rect 673637 579458 673703 579461
rect 673637 579456 676292 579458
rect 673637 579400 673642 579456
rect 673698 579400 676292 579456
rect 673637 579398 676292 579400
rect 673637 579395 673703 579398
rect 42057 579324 42123 579325
rect 42006 579322 42012 579324
rect 41966 579262 42012 579322
rect 42076 579320 42123 579324
rect 42118 579264 42123 579320
rect 42006 579260 42012 579262
rect 42076 579260 42123 579264
rect 42057 579259 42123 579260
rect 673637 579050 673703 579053
rect 673637 579048 676292 579050
rect 673637 578992 673642 579048
rect 673698 578992 676292 579048
rect 673637 578990 676292 578992
rect 673637 578987 673703 578990
rect 673637 578642 673703 578645
rect 673637 578640 676292 578642
rect 673637 578584 673642 578640
rect 673698 578584 676292 578640
rect 673637 578582 676292 578584
rect 673637 578579 673703 578582
rect 42149 578370 42215 578373
rect 44357 578370 44423 578373
rect 42149 578368 44423 578370
rect 42149 578312 42154 578368
rect 42210 578312 44362 578368
rect 44418 578312 44423 578368
rect 42149 578310 44423 578312
rect 42149 578307 42215 578310
rect 44357 578307 44423 578310
rect 673637 578234 673703 578237
rect 673637 578232 676292 578234
rect 673637 578176 673642 578232
rect 673698 578176 676292 578232
rect 673637 578174 676292 578176
rect 673637 578171 673703 578174
rect 40902 577764 40908 577828
rect 40972 577826 40978 577828
rect 41781 577826 41847 577829
rect 40972 577824 41847 577826
rect 40972 577768 41786 577824
rect 41842 577768 41847 577824
rect 40972 577766 41847 577768
rect 40972 577764 40978 577766
rect 41781 577763 41847 577766
rect 673637 577826 673703 577829
rect 673637 577824 676292 577826
rect 673637 577768 673642 577824
rect 673698 577768 676292 577824
rect 673637 577766 676292 577768
rect 673637 577763 673703 577766
rect 673637 577418 673703 577421
rect 673637 577416 676292 577418
rect 673637 577360 673642 577416
rect 673698 577360 676292 577416
rect 673637 577358 676292 577360
rect 673637 577355 673703 577358
rect 673637 577010 673703 577013
rect 673637 577008 676292 577010
rect 673637 576952 673642 577008
rect 673698 576952 676292 577008
rect 673637 576950 676292 576952
rect 673637 576947 673703 576950
rect 676806 576812 676812 576876
rect 676876 576812 676882 576876
rect 676814 576572 676874 576812
rect 682377 576466 682443 576469
rect 682334 576464 682443 576466
rect 682334 576408 682382 576464
rect 682438 576408 682443 576464
rect 682334 576403 682443 576408
rect 682334 576164 682394 576403
rect 684217 576058 684283 576061
rect 684174 576056 684283 576058
rect 684174 576000 684222 576056
rect 684278 576000 684283 576056
rect 684174 575995 684283 576000
rect 40534 575724 40540 575788
rect 40604 575786 40610 575788
rect 42149 575786 42215 575789
rect 40604 575784 42215 575786
rect 40604 575728 42154 575784
rect 42210 575728 42215 575784
rect 684174 575756 684234 575995
rect 40604 575726 42215 575728
rect 40604 575724 40610 575726
rect 42149 575723 42215 575726
rect 680997 575650 681063 575653
rect 680997 575648 681106 575650
rect 680997 575592 681002 575648
rect 681058 575592 681106 575648
rect 680997 575587 681106 575592
rect 681046 575348 681106 575587
rect 672993 574970 673059 574973
rect 672993 574968 676292 574970
rect 672993 574912 672998 574968
rect 673054 574912 676292 574968
rect 672993 574910 676292 574912
rect 672993 574907 673059 574910
rect 62113 574834 62179 574837
rect 62113 574832 64706 574834
rect 62113 574776 62118 574832
rect 62174 574776 64706 574832
rect 62113 574774 64706 574776
rect 62113 574771 62179 574774
rect 40718 574636 40724 574700
rect 40788 574698 40794 574700
rect 41781 574698 41847 574701
rect 40788 574696 41847 574698
rect 40788 574640 41786 574696
rect 41842 574640 41847 574696
rect 40788 574638 41847 574640
rect 40788 574636 40794 574638
rect 41781 574635 41847 574638
rect 64646 574194 64706 574774
rect 673637 574562 673703 574565
rect 673637 574560 676292 574562
rect 673637 574504 673642 574560
rect 673698 574504 676292 574560
rect 673637 574502 676292 574504
rect 673637 574499 673703 574502
rect 673637 574154 673703 574157
rect 673637 574152 676292 574154
rect 673637 574096 673642 574152
rect 673698 574096 676292 574152
rect 673637 574094 676292 574096
rect 673637 574091 673703 574094
rect 673085 573746 673151 573749
rect 673085 573744 676292 573746
rect 673085 573688 673090 573744
rect 673146 573688 676292 573744
rect 673085 573686 676292 573688
rect 673085 573683 673151 573686
rect 62113 573610 62179 573613
rect 62113 573608 64706 573610
rect 62113 573552 62118 573608
rect 62174 573552 64706 573608
rect 62113 573550 64706 573552
rect 62113 573547 62179 573550
rect 64646 573012 64706 573550
rect 672901 573474 672967 573477
rect 672901 573472 676230 573474
rect 672901 573416 672906 573472
rect 672962 573416 676230 573472
rect 672901 573414 676230 573416
rect 672901 573411 672967 573414
rect 676170 573338 676230 573414
rect 676170 573278 676292 573338
rect 683389 573202 683455 573205
rect 683389 573200 683498 573202
rect 683389 573144 683394 573200
rect 683450 573144 683498 573200
rect 683389 573139 683498 573144
rect 41454 572868 41460 572932
rect 41524 572930 41530 572932
rect 42609 572930 42675 572933
rect 41524 572928 42675 572930
rect 41524 572872 42614 572928
rect 42670 572872 42675 572928
rect 683438 572900 683498 573139
rect 41524 572870 42675 572872
rect 41524 572868 41530 572870
rect 42609 572867 42675 572870
rect 42057 572660 42123 572661
rect 42006 572596 42012 572660
rect 42076 572658 42123 572660
rect 42076 572656 42168 572658
rect 42118 572600 42168 572656
rect 42076 572598 42168 572600
rect 42076 572596 42123 572598
rect 42057 572595 42123 572596
rect 673637 572522 673703 572525
rect 673637 572520 676292 572522
rect 673637 572464 673642 572520
rect 673698 572464 676292 572520
rect 673637 572462 676292 572464
rect 673637 572459 673703 572462
rect 673637 572114 673703 572117
rect 673637 572112 676292 572114
rect 673637 572056 673642 572112
rect 673698 572056 676292 572112
rect 673637 572054 676292 572056
rect 673637 572051 673703 572054
rect 684033 571978 684099 571981
rect 683990 571976 684099 571978
rect 683990 571920 684038 571976
rect 684094 571920 684099 571976
rect 683990 571915 684099 571920
rect 41638 571508 41644 571572
rect 41708 571570 41714 571572
rect 42057 571570 42123 571573
rect 41708 571568 42123 571570
rect 41708 571512 42062 571568
rect 42118 571512 42123 571568
rect 41708 571510 42123 571512
rect 41708 571508 41714 571510
rect 42057 571507 42123 571510
rect 42425 571434 42491 571437
rect 64646 571434 64706 571830
rect 683990 571676 684050 571915
rect 676213 571570 676279 571573
rect 676213 571568 676322 571570
rect 676213 571512 676218 571568
rect 676274 571512 676322 571568
rect 676213 571507 676322 571512
rect 42425 571432 64706 571434
rect 42425 571376 42430 571432
rect 42486 571376 64706 571432
rect 42425 571374 64706 571376
rect 42425 571371 42491 571374
rect 676262 571268 676322 571507
rect 62757 571162 62823 571165
rect 62757 571160 64706 571162
rect 62757 571104 62762 571160
rect 62818 571104 64706 571160
rect 62757 571102 64706 571104
rect 62757 571099 62823 571102
rect 64646 570648 64706 571102
rect 673637 570890 673703 570893
rect 673637 570888 676292 570890
rect 673637 570832 673642 570888
rect 673698 570832 676292 570888
rect 673637 570830 676292 570832
rect 673637 570827 673703 570830
rect 682886 570346 682946 570452
rect 683113 570346 683179 570349
rect 682886 570344 683179 570346
rect 682886 570288 683118 570344
rect 683174 570288 683179 570344
rect 682886 570286 683179 570288
rect 41781 570212 41847 570213
rect 41781 570208 41828 570212
rect 41892 570210 41898 570212
rect 41781 570152 41786 570208
rect 41781 570148 41828 570152
rect 41892 570150 41938 570210
rect 41892 570148 41898 570150
rect 41781 570147 41847 570148
rect 682886 570044 682946 570286
rect 683113 570283 683179 570286
rect 62573 569938 62639 569941
rect 673637 569938 673703 569941
rect 674833 569938 674899 569941
rect 62573 569936 64706 569938
rect 62573 569880 62578 569936
rect 62634 569880 64706 569936
rect 62573 569878 64706 569880
rect 62573 569875 62639 569878
rect 64646 569466 64706 569878
rect 673637 569936 674899 569938
rect 673637 569880 673642 569936
rect 673698 569880 674838 569936
rect 674894 569880 674899 569936
rect 673637 569878 674899 569880
rect 673637 569875 673703 569878
rect 674833 569875 674899 569878
rect 673637 569666 673703 569669
rect 673637 569664 676292 569666
rect 673637 569608 673642 569664
rect 673698 569608 676292 569664
rect 673637 569606 676292 569608
rect 673637 569603 673703 569606
rect 63125 568578 63191 568581
rect 63125 568576 64706 568578
rect 63125 568520 63130 568576
rect 63186 568520 64706 568576
rect 63125 568518 64706 568520
rect 63125 568515 63191 568518
rect 64646 568284 64706 568518
rect 673637 565858 673703 565861
rect 675385 565858 675451 565861
rect 673637 565856 675451 565858
rect 673637 565800 673642 565856
rect 673698 565800 675390 565856
rect 675446 565800 675451 565856
rect 673637 565798 675451 565800
rect 673637 565795 673703 565798
rect 675385 565795 675451 565798
rect 673637 564634 673703 564637
rect 675109 564634 675175 564637
rect 673637 564632 675175 564634
rect 673637 564576 673642 564632
rect 673698 564576 675114 564632
rect 675170 564576 675175 564632
rect 673637 564574 675175 564576
rect 673637 564571 673703 564574
rect 675109 564571 675175 564574
rect 667013 562322 667079 562325
rect 675109 562322 675175 562325
rect 667013 562320 675175 562322
rect 667013 562264 667018 562320
rect 667074 562264 675114 562320
rect 675170 562264 675175 562320
rect 667013 562262 675175 562264
rect 667013 562259 667079 562262
rect 675109 562259 675175 562262
rect 675385 561916 675451 561917
rect 675334 561914 675340 561916
rect 675294 561854 675340 561914
rect 675404 561912 675451 561916
rect 675446 561856 675451 561912
rect 675334 561852 675340 561854
rect 675404 561852 675451 561856
rect 675385 561851 675451 561852
rect 673085 560282 673151 560285
rect 673085 560280 675586 560282
rect 673085 560224 673090 560280
rect 673146 560224 675586 560280
rect 673085 560222 675586 560224
rect 673085 560219 673151 560222
rect 671797 559602 671863 559605
rect 675201 559602 675267 559605
rect 671797 559600 675267 559602
rect 671797 559544 671802 559600
rect 671858 559544 675206 559600
rect 675262 559544 675267 559600
rect 671797 559542 675267 559544
rect 671797 559539 671863 559542
rect 675201 559539 675267 559542
rect 675526 559469 675586 560222
rect 675526 559464 675635 559469
rect 675526 559408 675574 559464
rect 675630 559408 675635 559464
rect 675526 559406 675635 559408
rect 675569 559403 675635 559406
rect 41086 558724 41092 558788
rect 41156 558786 41162 558788
rect 44909 558786 44975 558789
rect 41156 558784 44975 558786
rect 41156 558728 44914 558784
rect 44970 558728 44975 558784
rect 41156 558726 44975 558728
rect 41156 558724 41162 558726
rect 44909 558723 44975 558726
rect 54477 558514 54543 558517
rect 41492 558512 54543 558514
rect 41492 558456 54482 558512
rect 54538 558456 54543 558512
rect 41492 558454 54543 558456
rect 54477 558451 54543 558454
rect 674097 558378 674163 558381
rect 675477 558378 675543 558381
rect 674097 558376 675543 558378
rect 674097 558320 674102 558376
rect 674158 558320 675482 558376
rect 675538 558320 675543 558376
rect 674097 558318 675543 558320
rect 674097 558315 674163 558318
rect 675477 558315 675543 558318
rect 40953 558106 41019 558109
rect 40940 558104 41019 558106
rect 40940 558048 40958 558104
rect 41014 558048 41019 558104
rect 40940 558046 41019 558048
rect 40953 558043 41019 558046
rect 41086 557488 41092 557552
rect 41156 557488 41162 557552
rect 41278 557550 41338 557668
rect 675293 557562 675359 557565
rect 676254 557562 676260 557564
rect 675293 557560 676260 557562
rect 41278 557490 41890 557550
rect 675293 557504 675298 557560
rect 675354 557504 676260 557560
rect 675293 557502 676260 557504
rect 675293 557499 675359 557502
rect 676254 557500 676260 557502
rect 676324 557500 676330 557564
rect 41094 557260 41154 557488
rect 41830 557426 41890 557490
rect 41830 557366 51090 557426
rect 44357 556882 44423 556885
rect 41492 556880 44423 556882
rect 41492 556824 44362 556880
rect 44418 556824 44423 556880
rect 41492 556822 44423 556824
rect 44357 556819 44423 556822
rect 51030 556746 51090 557366
rect 62205 556746 62271 556749
rect 51030 556744 62271 556746
rect 51030 556688 62210 556744
rect 62266 556688 62271 556744
rect 51030 556686 62271 556688
rect 62205 556683 62271 556686
rect 44633 556474 44699 556477
rect 41492 556472 44699 556474
rect 41492 556416 44638 556472
rect 44694 556416 44699 556472
rect 41492 556414 44699 556416
rect 44633 556411 44699 556414
rect 44541 556066 44607 556069
rect 41492 556064 44607 556066
rect 41492 556008 44546 556064
rect 44602 556008 44607 556064
rect 41492 556006 44607 556008
rect 44541 556003 44607 556006
rect 42793 555658 42859 555661
rect 41492 555656 42859 555658
rect 41492 555600 42798 555656
rect 42854 555600 42859 555656
rect 41492 555598 42859 555600
rect 42793 555595 42859 555598
rect 45093 555250 45159 555253
rect 41492 555248 45159 555250
rect 41492 555192 45098 555248
rect 45154 555192 45159 555248
rect 41492 555190 45159 555192
rect 45093 555187 45159 555190
rect 672257 555250 672323 555253
rect 675385 555250 675451 555253
rect 672257 555248 675451 555250
rect 672257 555192 672262 555248
rect 672318 555192 675390 555248
rect 675446 555192 675451 555248
rect 672257 555190 675451 555192
rect 672257 555187 672323 555190
rect 675385 555187 675451 555190
rect 43069 554842 43135 554845
rect 41492 554840 43135 554842
rect 41492 554784 43074 554840
rect 43130 554784 43135 554840
rect 41492 554782 43135 554784
rect 43069 554779 43135 554782
rect 673637 554842 673703 554845
rect 675293 554842 675359 554845
rect 673637 554840 675359 554842
rect 673637 554784 673642 554840
rect 673698 554784 675298 554840
rect 675354 554784 675359 554840
rect 673637 554782 675359 554784
rect 673637 554779 673703 554782
rect 675293 554779 675359 554782
rect 43713 554434 43779 554437
rect 41492 554432 43779 554434
rect 41492 554376 43718 554432
rect 43774 554376 43779 554432
rect 41492 554374 43779 554376
rect 43713 554371 43779 554374
rect 41822 554026 41828 554028
rect 41492 553966 41828 554026
rect 41822 553964 41828 553966
rect 41892 553964 41898 554028
rect 41278 553413 41338 553588
rect 649950 553482 650010 553914
rect 675753 553890 675819 553893
rect 676806 553890 676812 553892
rect 675753 553888 676812 553890
rect 675753 553832 675758 553888
rect 675814 553832 676812 553888
rect 675753 553830 676812 553832
rect 675753 553827 675819 553830
rect 676806 553828 676812 553830
rect 676876 553828 676882 553892
rect 651465 553482 651531 553485
rect 673637 553484 673703 553485
rect 673637 553482 673684 553484
rect 649950 553480 651531 553482
rect 649950 553424 651470 553480
rect 651526 553424 651531 553480
rect 649950 553422 651531 553424
rect 673592 553480 673684 553482
rect 673592 553424 673642 553480
rect 673592 553422 673684 553424
rect 651465 553419 651531 553422
rect 673637 553420 673684 553422
rect 673748 553420 673754 553484
rect 675569 553482 675635 553485
rect 675526 553480 675635 553482
rect 675526 553424 675574 553480
rect 675630 553424 675635 553480
rect 673637 553419 673703 553420
rect 675526 553419 675635 553424
rect 37917 553410 37983 553413
rect 37917 553408 38026 553410
rect 37917 553352 37922 553408
rect 37978 553352 38026 553408
rect 37917 553347 38026 553352
rect 41278 553408 41387 553413
rect 41278 553352 41326 553408
rect 41382 553352 41387 553408
rect 41278 553350 41387 553352
rect 41321 553347 41387 553350
rect 37966 553180 38026 553347
rect 673637 553210 673703 553213
rect 675526 553210 675586 553419
rect 673637 553208 675586 553210
rect 673637 553152 673642 553208
rect 673698 553152 675586 553208
rect 673637 553150 675586 553152
rect 673637 553147 673703 553150
rect 41822 552802 41828 552804
rect 41492 552742 41828 552802
rect 41822 552740 41828 552742
rect 41892 552740 41898 552804
rect 43805 552394 43871 552397
rect 41492 552392 43871 552394
rect 41492 552336 43810 552392
rect 43866 552336 43871 552392
rect 41492 552334 43871 552336
rect 43805 552331 43871 552334
rect 649950 552122 650010 552732
rect 651465 552122 651531 552125
rect 649950 552120 651531 552122
rect 649950 552064 651470 552120
rect 651526 552064 651531 552120
rect 649950 552062 651531 552064
rect 651465 552059 651531 552062
rect 29637 551986 29703 551989
rect 674649 551986 674715 551989
rect 675385 551986 675451 551989
rect 29637 551984 29716 551986
rect 29637 551928 29642 551984
rect 29698 551928 29716 551984
rect 29637 551926 29716 551928
rect 674649 551984 675451 551986
rect 674649 551928 674654 551984
rect 674710 551928 675390 551984
rect 675446 551928 675451 551984
rect 674649 551926 675451 551928
rect 29637 551923 29703 551926
rect 674649 551923 674715 551926
rect 675385 551923 675451 551926
rect 45277 551578 45343 551581
rect 41492 551576 45343 551578
rect 41492 551520 45282 551576
rect 45338 551520 45343 551576
rect 41492 551518 45343 551520
rect 45277 551515 45343 551518
rect 43989 551170 44055 551173
rect 41492 551168 44055 551170
rect 41492 551112 43994 551168
rect 44050 551112 44055 551168
rect 41492 551110 44055 551112
rect 43989 551107 44055 551110
rect 649950 551034 650010 551550
rect 673678 551516 673684 551580
rect 673748 551578 673754 551580
rect 675385 551578 675451 551581
rect 673748 551576 675451 551578
rect 673748 551520 675390 551576
rect 675446 551520 675451 551576
rect 673748 551518 675451 551520
rect 673748 551516 673754 551518
rect 675385 551515 675451 551518
rect 652017 551034 652083 551037
rect 649950 551032 652083 551034
rect 649950 550976 652022 551032
rect 652078 550976 652083 551032
rect 649950 550974 652083 550976
rect 652017 550971 652083 550974
rect 43069 550762 43135 550765
rect 41492 550760 43135 550762
rect 41492 550704 43074 550760
rect 43130 550704 43135 550760
rect 41492 550702 43135 550704
rect 43069 550699 43135 550702
rect 42057 550490 42123 550493
rect 42057 550488 48330 550490
rect 42057 550432 42062 550488
rect 42118 550432 48330 550488
rect 42057 550430 48330 550432
rect 42057 550427 42123 550430
rect 41492 550294 41890 550354
rect 41830 550218 41890 550294
rect 44173 550218 44239 550221
rect 41830 550216 44239 550218
rect 41830 550160 44178 550216
rect 44234 550160 44239 550216
rect 41830 550158 44239 550160
rect 48270 550218 48330 550430
rect 649950 550354 650010 550368
rect 651649 550354 651715 550357
rect 649950 550352 651715 550354
rect 649950 550296 651654 550352
rect 651710 550296 651715 550352
rect 649950 550294 651715 550296
rect 651649 550291 651715 550294
rect 62757 550218 62823 550221
rect 48270 550216 62823 550218
rect 48270 550160 62762 550216
rect 62818 550160 62823 550216
rect 48270 550158 62823 550160
rect 44173 550155 44239 550158
rect 62757 550155 62823 550158
rect 675477 550216 675543 550221
rect 675477 550160 675482 550216
rect 675538 550160 675543 550216
rect 675477 550155 675543 550160
rect 40677 549946 40743 549949
rect 675017 549946 675083 549949
rect 675480 549946 675540 550155
rect 40677 549944 40756 549946
rect 40677 549888 40682 549944
rect 40738 549888 40756 549944
rect 40677 549886 40756 549888
rect 675017 549944 675540 549946
rect 675017 549888 675022 549944
rect 675078 549888 675540 549944
rect 675017 549886 675540 549888
rect 40677 549883 40743 549886
rect 675017 549883 675083 549886
rect 670417 549674 670483 549677
rect 675477 549674 675543 549677
rect 670417 549672 675543 549674
rect 670417 549616 670422 549672
rect 670478 549616 675482 549672
rect 675538 549616 675543 549672
rect 670417 549614 675543 549616
rect 670417 549611 670483 549614
rect 675477 549611 675543 549614
rect 42006 549538 42012 549540
rect 41492 549478 42012 549538
rect 42006 549476 42012 549478
rect 42076 549476 42082 549540
rect 651465 549266 651531 549269
rect 649950 549264 651531 549266
rect 649950 549208 651470 549264
rect 651526 549208 651531 549264
rect 649950 549206 651531 549208
rect 649950 549186 650010 549206
rect 651465 549203 651531 549206
rect 42793 549130 42859 549133
rect 41492 549128 42859 549130
rect 41492 549072 42798 549128
rect 42854 549072 42859 549128
rect 41492 549070 42859 549072
rect 42793 549067 42859 549070
rect 674005 548858 674071 548861
rect 674966 548858 674972 548860
rect 674005 548856 674972 548858
rect 674005 548800 674010 548856
rect 674066 548800 674972 548856
rect 674005 548798 674972 548800
rect 674005 548795 674071 548798
rect 674966 548796 674972 548798
rect 675036 548796 675042 548860
rect 45461 548722 45527 548725
rect 41492 548720 45527 548722
rect 41492 548664 45466 548720
rect 45522 548664 45527 548720
rect 41492 548662 45527 548664
rect 45461 548659 45527 548662
rect 651465 548450 651531 548453
rect 649950 548448 651531 548450
rect 649950 548392 651470 548448
rect 651526 548392 651531 548448
rect 649950 548390 651531 548392
rect 41321 548314 41387 548317
rect 41308 548312 41387 548314
rect 41308 548256 41326 548312
rect 41382 548256 41387 548312
rect 41308 548254 41387 548256
rect 41321 548251 41387 548254
rect 649950 548004 650010 548390
rect 651465 548387 651531 548390
rect 675753 548314 675819 548317
rect 676990 548314 676996 548316
rect 675753 548312 676996 548314
rect 675753 548256 675758 548312
rect 675814 548256 676996 548312
rect 675753 548254 676996 548256
rect 675753 548251 675819 548254
rect 676990 548252 676996 548254
rect 677060 548252 677066 548316
rect 674966 547844 674972 547908
rect 675036 547906 675042 547908
rect 675569 547906 675635 547909
rect 675036 547904 675635 547906
rect 675036 547848 675574 547904
rect 675630 547848 675635 547904
rect 675036 547846 675635 547848
rect 675036 547844 675042 547846
rect 675569 547843 675635 547846
rect 676254 547572 676260 547636
rect 676324 547634 676330 547636
rect 677409 547634 677475 547637
rect 676324 547632 677475 547634
rect 676324 547576 677414 547632
rect 677470 547576 677475 547632
rect 676324 547574 677475 547576
rect 676324 547572 676330 547574
rect 677409 547571 677475 547574
rect 39573 547498 39639 547501
rect 39573 547496 39652 547498
rect 39573 547440 39578 547496
rect 39634 547440 39652 547496
rect 39573 547438 39652 547440
rect 39573 547435 39639 547438
rect 674414 547028 674420 547092
rect 674484 547090 674490 547092
rect 683389 547090 683455 547093
rect 674484 547088 683455 547090
rect 674484 547032 683394 547088
rect 683450 547032 683455 547088
rect 674484 547030 683455 547032
rect 674484 547028 674490 547030
rect 683389 547027 683455 547030
rect 676070 546756 676076 546820
rect 676140 546818 676146 546820
rect 680997 546818 681063 546821
rect 676140 546816 681063 546818
rect 676140 546760 681002 546816
rect 681058 546760 681063 546816
rect 676140 546758 681063 546760
rect 676140 546756 676146 546758
rect 680997 546755 681063 546758
rect 674833 545866 674899 545869
rect 675334 545866 675340 545868
rect 674833 545864 675340 545866
rect 674833 545808 674838 545864
rect 674894 545808 675340 545864
rect 674833 545806 675340 545808
rect 674833 545803 674899 545806
rect 675334 545804 675340 545806
rect 675404 545804 675410 545868
rect 40677 545596 40743 545597
rect 40677 545592 40724 545596
rect 40788 545594 40794 545596
rect 40677 545536 40682 545592
rect 40677 545532 40724 545536
rect 40788 545534 40834 545594
rect 40788 545532 40794 545534
rect 40677 545531 40743 545532
rect 40534 545260 40540 545324
rect 40604 545322 40610 545324
rect 42006 545322 42012 545324
rect 40604 545262 42012 545322
rect 40604 545260 40610 545262
rect 42006 545260 42012 545262
rect 42076 545260 42082 545324
rect 39573 542602 39639 542605
rect 44725 542602 44791 542605
rect 39573 542600 44791 542602
rect 39573 542544 39578 542600
rect 39634 542544 44730 542600
rect 44786 542544 44791 542600
rect 39573 542542 44791 542544
rect 39573 542539 39639 542542
rect 44725 542539 44791 542542
rect 37917 542330 37983 542333
rect 41822 542330 41828 542332
rect 37917 542328 41828 542330
rect 37917 542272 37922 542328
rect 37978 542272 41828 542328
rect 37917 542270 41828 542272
rect 37917 542267 37983 542270
rect 41822 542268 41828 542270
rect 41892 542268 41898 542332
rect 45185 539882 45251 539885
rect 51717 539882 51783 539885
rect 45185 539880 51783 539882
rect 45185 539824 45190 539880
rect 45246 539824 51722 539880
rect 51778 539824 51783 539880
rect 45185 539822 51783 539824
rect 45185 539819 45251 539822
rect 51717 539819 51783 539822
rect 40718 539548 40724 539612
rect 40788 539610 40794 539612
rect 42609 539610 42675 539613
rect 40788 539608 42675 539610
rect 40788 539552 42614 539608
rect 42670 539552 42675 539608
rect 40788 539550 42675 539552
rect 40788 539548 40794 539550
rect 42609 539547 42675 539550
rect 42425 538250 42491 538253
rect 44173 538250 44239 538253
rect 42425 538248 44239 538250
rect 42425 538192 42430 538248
rect 42486 538192 44178 538248
rect 44234 538192 44239 538248
rect 42425 538190 44239 538192
rect 42425 538187 42491 538190
rect 44173 538187 44239 538190
rect 42149 537978 42215 537981
rect 45185 537978 45251 537981
rect 42149 537976 45251 537978
rect 42149 537920 42154 537976
rect 42210 537920 45190 537976
rect 45246 537920 45251 537976
rect 42149 537918 45251 537920
rect 42149 537915 42215 537918
rect 45185 537915 45251 537918
rect 45645 536890 45711 536893
rect 42428 536888 45711 536890
rect 42428 536832 45650 536888
rect 45706 536832 45711 536888
rect 42428 536830 45711 536832
rect 42428 536485 42488 536830
rect 45645 536827 45711 536830
rect 42425 536480 42491 536485
rect 42425 536424 42430 536480
rect 42486 536424 42491 536480
rect 42425 536419 42491 536424
rect 669037 536482 669103 536485
rect 675477 536482 675543 536485
rect 669037 536480 675543 536482
rect 669037 536424 669042 536480
rect 669098 536424 675482 536480
rect 675538 536424 675543 536480
rect 669037 536422 675543 536424
rect 669037 536419 669103 536422
rect 675477 536419 675543 536422
rect 673821 536210 673887 536213
rect 674189 536210 674255 536213
rect 673821 536208 674255 536210
rect 673821 536152 673826 536208
rect 673882 536152 674194 536208
rect 674250 536152 674255 536208
rect 673821 536150 674255 536152
rect 673821 536147 673887 536150
rect 674189 536147 674255 536150
rect 672625 535938 672691 535941
rect 676262 535938 676322 536112
rect 672625 535936 676322 535938
rect 672625 535880 672630 535936
rect 672686 535880 676322 535936
rect 672625 535878 676322 535880
rect 672625 535875 672691 535878
rect 42149 535666 42215 535669
rect 45185 535666 45251 535669
rect 42149 535664 45251 535666
rect 42149 535608 42154 535664
rect 42210 535608 45190 535664
rect 45246 535608 45251 535664
rect 42149 535606 45251 535608
rect 42149 535603 42215 535606
rect 45185 535603 45251 535606
rect 672625 535666 672691 535669
rect 676262 535666 676322 535704
rect 672625 535664 676322 535666
rect 672625 535608 672630 535664
rect 672686 535608 676322 535664
rect 672625 535606 676322 535608
rect 672625 535603 672691 535606
rect 673494 535060 673500 535124
rect 673564 535122 673570 535124
rect 676262 535122 676322 535296
rect 673564 535062 676322 535122
rect 673564 535060 673570 535062
rect 672625 534850 672691 534853
rect 676262 534850 676322 534888
rect 672625 534848 676322 534850
rect 672625 534792 672630 534848
rect 672686 534792 676322 534848
rect 672625 534790 676322 534792
rect 672625 534787 672691 534790
rect 672625 534578 672691 534581
rect 672625 534576 673930 534578
rect 672625 534520 672630 534576
rect 672686 534520 673930 534576
rect 672625 534518 673930 534520
rect 672625 534515 672691 534518
rect 672625 534306 672691 534309
rect 673494 534306 673500 534308
rect 672625 534304 673500 534306
rect 672625 534248 672630 534304
rect 672686 534248 673500 534304
rect 672625 534246 673500 534248
rect 672625 534243 672691 534246
rect 673494 534244 673500 534246
rect 673564 534244 673570 534308
rect 673870 534306 673930 534518
rect 676029 534510 676095 534513
rect 676029 534508 676292 534510
rect 676029 534452 676034 534508
rect 676090 534452 676292 534508
rect 676029 534450 676292 534452
rect 676029 534447 676095 534450
rect 673870 534246 676322 534306
rect 676262 534072 676322 534246
rect 42425 533898 42491 533901
rect 43805 533898 43871 533901
rect 42425 533896 43871 533898
rect 42425 533840 42430 533896
rect 42486 533840 43810 533896
rect 43866 533840 43871 533896
rect 42425 533838 43871 533840
rect 42425 533835 42491 533838
rect 43805 533835 43871 533838
rect 670785 533898 670851 533901
rect 674281 533898 674347 533901
rect 670785 533896 674347 533898
rect 670785 533840 670790 533896
rect 670846 533840 674286 533896
rect 674342 533840 674347 533896
rect 670785 533838 674347 533840
rect 670785 533835 670851 533838
rect 674281 533835 674347 533838
rect 672625 533626 672691 533629
rect 676262 533626 676322 533664
rect 672625 533624 676322 533626
rect 672625 533568 672630 533624
rect 672686 533568 676322 533624
rect 672625 533566 676322 533568
rect 672625 533563 672691 533566
rect 40534 533292 40540 533356
rect 40604 533354 40610 533356
rect 42241 533354 42307 533357
rect 40604 533352 42307 533354
rect 40604 533296 42246 533352
rect 42302 533296 42307 533352
rect 40604 533294 42307 533296
rect 40604 533292 40610 533294
rect 42241 533291 42307 533294
rect 672441 533354 672507 533357
rect 672441 533352 676322 533354
rect 672441 533296 672446 533352
rect 672502 533296 676322 533352
rect 672441 533294 676322 533296
rect 672441 533291 672507 533294
rect 676262 533256 676322 533294
rect 671613 532810 671679 532813
rect 676262 532810 676322 532848
rect 671613 532808 676322 532810
rect 671613 532752 671618 532808
rect 671674 532752 676322 532808
rect 671613 532750 676322 532752
rect 671613 532747 671679 532750
rect 672441 532538 672507 532541
rect 672441 532536 676322 532538
rect 672441 532480 672446 532536
rect 672502 532480 676322 532536
rect 672441 532478 676322 532480
rect 672441 532475 672507 532478
rect 676262 532440 676322 532478
rect 671153 532130 671219 532133
rect 671153 532128 676230 532130
rect 671153 532072 671158 532128
rect 671214 532072 676230 532128
rect 671153 532070 676230 532072
rect 671153 532067 671219 532070
rect 676170 532062 676230 532070
rect 676170 532002 676292 532062
rect 676213 531858 676279 531861
rect 676213 531856 676322 531858
rect 676213 531800 676218 531856
rect 676274 531800 676322 531856
rect 676213 531795 676322 531800
rect 41638 531660 41644 531724
rect 41708 531722 41714 531724
rect 42609 531722 42675 531725
rect 41708 531720 42675 531722
rect 41708 531664 42614 531720
rect 42670 531664 42675 531720
rect 41708 531662 42675 531664
rect 41708 531660 41714 531662
rect 42609 531659 42675 531662
rect 676262 531624 676322 531795
rect 682377 531450 682443 531453
rect 682334 531448 682443 531450
rect 682334 531392 682382 531448
rect 682438 531392 682443 531448
rect 682334 531387 682443 531392
rect 62113 531314 62179 531317
rect 62113 531312 64154 531314
rect 62113 531256 62118 531312
rect 62174 531256 64154 531312
rect 62113 531254 64154 531256
rect 62113 531251 62179 531254
rect 64094 531202 64154 531254
rect 682334 531216 682394 531387
rect 64094 531142 64676 531202
rect 676029 530838 676095 530841
rect 676029 530836 676292 530838
rect 676029 530780 676034 530836
rect 676090 530780 676292 530836
rect 676029 530778 676292 530780
rect 676029 530775 676095 530778
rect 62113 530634 62179 530637
rect 680997 530634 681063 530637
rect 62113 530632 64706 530634
rect 62113 530576 62118 530632
rect 62174 530576 64706 530632
rect 62113 530574 64706 530576
rect 62113 530571 62179 530574
rect 41454 530164 41460 530228
rect 41524 530226 41530 530228
rect 42425 530226 42491 530229
rect 41524 530224 42491 530226
rect 41524 530168 42430 530224
rect 42486 530168 42491 530224
rect 41524 530166 42491 530168
rect 41524 530164 41530 530166
rect 42425 530163 42491 530166
rect 64646 529990 64706 530574
rect 680997 530632 681106 530634
rect 680997 530576 681002 530632
rect 681058 530576 681106 530632
rect 680997 530571 681106 530576
rect 681046 530400 681106 530571
rect 676029 530022 676095 530025
rect 676029 530020 676292 530022
rect 676029 529964 676034 530020
rect 676090 529964 676292 530020
rect 676029 529962 676292 529964
rect 676029 529959 676095 529962
rect 42057 529954 42123 529957
rect 43989 529954 44055 529957
rect 42057 529952 44055 529954
rect 42057 529896 42062 529952
rect 42118 529896 43994 529952
rect 44050 529896 44055 529952
rect 42057 529894 44055 529896
rect 42057 529891 42123 529894
rect 43989 529891 44055 529894
rect 676262 529413 676322 529584
rect 676213 529408 676322 529413
rect 676213 529352 676218 529408
rect 676274 529352 676322 529408
rect 676213 529350 676322 529352
rect 676213 529347 676279 529350
rect 676029 529206 676095 529209
rect 676029 529204 676292 529206
rect 676029 529148 676034 529204
rect 676090 529148 676292 529204
rect 676029 529146 676292 529148
rect 676029 529143 676095 529146
rect 41822 528940 41828 529004
rect 41892 529002 41898 529004
rect 42425 529002 42491 529005
rect 41892 529000 42491 529002
rect 41892 528944 42430 529000
rect 42486 528944 42491 529000
rect 41892 528942 42491 528944
rect 41892 528940 41898 528942
rect 42425 528939 42491 528942
rect 42609 529002 42675 529005
rect 45461 529002 45527 529005
rect 42609 529000 45527 529002
rect 42609 528944 42614 529000
rect 42670 528944 45466 529000
rect 45522 528944 45527 529000
rect 42609 528942 45527 528944
rect 42609 528939 42675 528942
rect 45461 528939 45527 528942
rect 672809 528866 672875 528869
rect 672809 528864 676322 528866
rect 672809 528808 672814 528864
rect 672870 528808 676322 528864
rect 62113 528594 62179 528597
rect 64646 528594 64706 528808
rect 672809 528806 676322 528808
rect 672809 528803 672875 528806
rect 676262 528768 676322 528806
rect 62113 528592 64706 528594
rect 62113 528536 62118 528592
rect 62174 528536 64706 528592
rect 62113 528534 64706 528536
rect 683573 528594 683639 528597
rect 683573 528592 683682 528594
rect 683573 528536 683578 528592
rect 683634 528536 683682 528592
rect 62113 528531 62179 528534
rect 683573 528531 683682 528536
rect 683622 528360 683682 528531
rect 62297 528050 62363 528053
rect 672901 528050 672967 528053
rect 62297 528048 64706 528050
rect 62297 527992 62302 528048
rect 62358 527992 64706 528048
rect 62297 527990 64706 527992
rect 62297 527987 62363 527990
rect 64646 527626 64706 527990
rect 672901 528048 676322 528050
rect 672901 527992 672906 528048
rect 672962 527992 676322 528048
rect 672901 527990 676322 527992
rect 672901 527987 672967 527990
rect 676262 527952 676322 527990
rect 683205 527778 683271 527781
rect 683205 527776 683314 527778
rect 683205 527720 683210 527776
rect 683266 527720 683314 527776
rect 683205 527715 683314 527720
rect 683254 527544 683314 527715
rect 683389 527370 683455 527373
rect 683389 527368 683498 527370
rect 683389 527312 683394 527368
rect 683450 527312 683498 527368
rect 683389 527307 683498 527312
rect 42793 527234 42859 527237
rect 45277 527234 45343 527237
rect 42793 527232 45343 527234
rect 42793 527176 42798 527232
rect 42854 527176 45282 527232
rect 45338 527176 45343 527232
rect 42793 527174 45343 527176
rect 42793 527171 42859 527174
rect 45277 527171 45343 527174
rect 683438 527136 683498 527307
rect 62113 527098 62179 527101
rect 62113 527096 64706 527098
rect 62113 527040 62118 527096
rect 62174 527040 64706 527096
rect 62113 527038 64706 527040
rect 62113 527035 62179 527038
rect 64646 526444 64706 527038
rect 676029 526758 676095 526761
rect 676029 526756 676292 526758
rect 676029 526700 676034 526756
rect 676090 526700 676292 526756
rect 676029 526698 676292 526700
rect 676029 526695 676095 526698
rect 676029 526350 676095 526353
rect 676029 526348 676292 526350
rect 676029 526292 676034 526348
rect 676090 526292 676292 526348
rect 676029 526290 676292 526292
rect 676029 526287 676095 526290
rect 677918 525741 677978 525912
rect 62757 525738 62823 525741
rect 62757 525736 64706 525738
rect 62757 525680 62762 525736
rect 62818 525680 64706 525736
rect 62757 525678 64706 525680
rect 62757 525675 62823 525678
rect 64646 525262 64706 525678
rect 677869 525736 677978 525741
rect 677869 525680 677874 525736
rect 677930 525680 677978 525736
rect 677869 525678 677978 525680
rect 677869 525675 677935 525678
rect 683070 524925 683130 525504
rect 683070 524920 683179 524925
rect 683070 524864 683118 524920
rect 683174 524864 683179 524920
rect 683070 524862 683179 524864
rect 683113 524859 683179 524862
rect 679022 524517 679082 524688
rect 678973 524512 679082 524517
rect 678973 524456 678978 524512
rect 679034 524456 679082 524512
rect 678973 524454 679082 524456
rect 678973 524451 679039 524454
rect 676990 503644 676996 503708
rect 677060 503706 677066 503708
rect 683389 503706 683455 503709
rect 677060 503704 683455 503706
rect 677060 503648 683394 503704
rect 683450 503648 683455 503704
rect 677060 503646 683455 503648
rect 677060 503644 677066 503646
rect 683389 503643 683455 503646
rect 676806 500924 676812 500988
rect 676876 500986 676882 500988
rect 683205 500986 683271 500989
rect 676876 500984 683271 500986
rect 676876 500928 683210 500984
rect 683266 500928 683271 500984
rect 676876 500926 683271 500928
rect 676876 500924 676882 500926
rect 683205 500923 683271 500926
rect 673821 492146 673887 492149
rect 673821 492144 676292 492146
rect 673821 492088 673826 492144
rect 673882 492088 676292 492144
rect 673821 492086 676292 492088
rect 673821 492083 673887 492086
rect 676029 491738 676095 491741
rect 676029 491736 676292 491738
rect 676029 491680 676034 491736
rect 676090 491680 676292 491736
rect 676029 491678 676292 491680
rect 676029 491675 676095 491678
rect 675845 491330 675911 491333
rect 675845 491328 676292 491330
rect 675845 491272 675850 491328
rect 675906 491272 676292 491328
rect 675845 491270 676292 491272
rect 675845 491267 675911 491270
rect 674005 490922 674071 490925
rect 674005 490920 676292 490922
rect 674005 490864 674010 490920
rect 674066 490864 676292 490920
rect 674005 490862 676292 490864
rect 674005 490859 674071 490862
rect 674005 490514 674071 490517
rect 674005 490512 676292 490514
rect 674005 490456 674010 490512
rect 674066 490456 676292 490512
rect 674005 490454 676292 490456
rect 674005 490451 674071 490454
rect 674005 490106 674071 490109
rect 674005 490104 676292 490106
rect 674005 490048 674010 490104
rect 674066 490048 676292 490104
rect 674005 490046 676292 490048
rect 674005 490043 674071 490046
rect 674005 489698 674071 489701
rect 674005 489696 676292 489698
rect 674005 489640 674010 489696
rect 674066 489640 676292 489696
rect 674005 489638 676292 489640
rect 674005 489635 674071 489638
rect 674005 489290 674071 489293
rect 674005 489288 676292 489290
rect 674005 489232 674010 489288
rect 674066 489232 676292 489288
rect 674005 489230 676292 489232
rect 674005 489227 674071 489230
rect 675886 488820 675892 488884
rect 675956 488882 675962 488884
rect 675956 488822 676292 488882
rect 675956 488820 675962 488822
rect 674005 488474 674071 488477
rect 674005 488472 676292 488474
rect 674005 488416 674010 488472
rect 674066 488416 676292 488472
rect 674005 488414 676292 488416
rect 674005 488411 674071 488414
rect 676170 488006 676292 488066
rect 675886 487868 675892 487932
rect 675956 487930 675962 487932
rect 676170 487930 676230 488006
rect 675956 487870 676230 487930
rect 675956 487868 675962 487870
rect 681181 487658 681247 487661
rect 681181 487656 681260 487658
rect 681181 487600 681186 487656
rect 681242 487600 681260 487656
rect 681181 487598 681260 487600
rect 681181 487595 681247 487598
rect 679617 487250 679683 487253
rect 679604 487248 679683 487250
rect 679604 487192 679622 487248
rect 679678 487192 679683 487248
rect 679604 487190 679683 487192
rect 679617 487187 679683 487190
rect 676029 486842 676095 486845
rect 676029 486840 676292 486842
rect 676029 486784 676034 486840
rect 676090 486784 676292 486840
rect 676029 486782 676292 486784
rect 676029 486779 676095 486782
rect 680997 486434 681063 486437
rect 680997 486432 681076 486434
rect 680997 486376 681002 486432
rect 681058 486376 681076 486432
rect 680997 486374 681076 486376
rect 680997 486371 681063 486374
rect 673821 486026 673887 486029
rect 673821 486024 676292 486026
rect 673821 485968 673826 486024
rect 673882 485968 676292 486024
rect 673821 485966 676292 485968
rect 673821 485963 673887 485966
rect 683389 485618 683455 485621
rect 683389 485616 683468 485618
rect 683389 485560 683394 485616
rect 683450 485560 683468 485616
rect 683389 485558 683468 485560
rect 683389 485555 683455 485558
rect 676029 485210 676095 485213
rect 676029 485208 676292 485210
rect 676029 485152 676034 485208
rect 676090 485152 676292 485208
rect 676029 485150 676292 485152
rect 676029 485147 676095 485150
rect 673085 484802 673151 484805
rect 673085 484800 676292 484802
rect 673085 484744 673090 484800
rect 673146 484744 676292 484800
rect 673085 484742 676292 484744
rect 673085 484739 673151 484742
rect 674649 484394 674715 484397
rect 674649 484392 676292 484394
rect 674649 484336 674654 484392
rect 674710 484336 676292 484392
rect 674649 484334 676292 484336
rect 674649 484331 674715 484334
rect 676029 483986 676095 483989
rect 676029 483984 676292 483986
rect 676029 483928 676034 483984
rect 676090 483928 676292 483984
rect 676029 483926 676292 483928
rect 676029 483923 676095 483926
rect 683205 483578 683271 483581
rect 683205 483576 683284 483578
rect 683205 483520 683210 483576
rect 683266 483520 683284 483576
rect 683205 483518 683284 483520
rect 683205 483515 683271 483518
rect 674005 483170 674071 483173
rect 674005 483168 676292 483170
rect 674005 483112 674010 483168
rect 674066 483112 676292 483168
rect 674005 483110 676292 483112
rect 674005 483107 674071 483110
rect 676029 482762 676095 482765
rect 676029 482760 676292 482762
rect 676029 482704 676034 482760
rect 676090 482704 676292 482760
rect 676029 482702 676292 482704
rect 676029 482699 676095 482702
rect 673637 482354 673703 482357
rect 673637 482352 676292 482354
rect 673637 482296 673642 482352
rect 673698 482296 676292 482352
rect 673637 482294 676292 482296
rect 673637 482291 673703 482294
rect 680353 481946 680419 481949
rect 680340 481944 680419 481946
rect 680340 481888 680358 481944
rect 680414 481888 680419 481944
rect 680340 481886 680419 481888
rect 680353 481883 680419 481886
rect 677182 481130 677242 481508
rect 683113 481130 683179 481133
rect 677182 481128 683179 481130
rect 677182 481100 683118 481128
rect 677212 481072 683118 481100
rect 683174 481072 683179 481128
rect 677212 481070 683179 481072
rect 683113 481067 683179 481070
rect 675845 480722 675911 480725
rect 675845 480720 676292 480722
rect 675845 480664 675850 480720
rect 675906 480664 676292 480720
rect 675845 480662 676292 480664
rect 675845 480659 675911 480662
rect 669773 455426 669839 455429
rect 673269 455426 673335 455429
rect 669773 455424 673335 455426
rect 669773 455368 669778 455424
rect 669834 455368 673274 455424
rect 673330 455368 673335 455424
rect 669773 455366 673335 455368
rect 669773 455363 669839 455366
rect 673269 455363 673335 455366
rect 673381 455290 673447 455293
rect 673862 455290 673868 455292
rect 673381 455288 673868 455290
rect 673381 455232 673386 455288
rect 673442 455232 673868 455288
rect 673381 455230 673868 455232
rect 673381 455227 673447 455230
rect 673862 455228 673868 455230
rect 673932 455228 673938 455292
rect 670601 455154 670667 455157
rect 673269 455154 673335 455157
rect 670601 455152 673335 455154
rect 670601 455096 670606 455152
rect 670662 455096 673274 455152
rect 673330 455096 673335 455152
rect 670601 455094 673335 455096
rect 670601 455091 670667 455094
rect 673269 455091 673335 455094
rect 672809 454882 672875 454885
rect 674281 454882 674347 454885
rect 672809 454880 674347 454882
rect 672809 454824 672814 454880
rect 672870 454824 674286 454880
rect 674342 454824 674347 454880
rect 672809 454822 674347 454824
rect 672809 454819 672875 454822
rect 674281 454819 674347 454822
rect 673039 454610 673105 454613
rect 674281 454610 674347 454613
rect 673039 454608 674347 454610
rect 673039 454552 673044 454608
rect 673100 454552 674286 454608
rect 674342 454552 674347 454608
rect 673039 454550 674347 454552
rect 673039 454547 673105 454550
rect 674281 454547 674347 454550
rect 672947 454338 673013 454341
rect 674281 454338 674347 454341
rect 672947 454336 674347 454338
rect 672947 454280 672952 454336
rect 673008 454280 674286 454336
rect 674342 454280 674347 454336
rect 672947 454278 674347 454280
rect 672947 454275 673013 454278
rect 674281 454275 674347 454278
rect 672257 453930 672323 453933
rect 674281 453930 674347 453933
rect 672257 453928 674347 453930
rect 672257 453872 672262 453928
rect 672318 453872 674286 453928
rect 674342 453872 674347 453928
rect 672257 453870 674347 453872
rect 672257 453867 672323 453870
rect 674281 453867 674347 453870
rect 44817 430946 44883 430949
rect 41492 430944 44883 430946
rect 41492 430888 44822 430944
rect 44878 430888 44883 430944
rect 41492 430886 44883 430888
rect 44817 430883 44883 430886
rect 54477 430538 54543 430541
rect 41492 430536 54543 430538
rect 41492 430480 54482 430536
rect 54538 430480 54543 430536
rect 41492 430478 54543 430480
rect 54477 430475 54543 430478
rect 35801 430130 35867 430133
rect 35788 430128 35867 430130
rect 35788 430072 35806 430128
rect 35862 430072 35867 430128
rect 35788 430070 35867 430072
rect 35801 430067 35867 430070
rect 44357 429722 44423 429725
rect 41492 429720 44423 429722
rect 41492 429664 44362 429720
rect 44418 429664 44423 429720
rect 41492 429662 44423 429664
rect 44357 429659 44423 429662
rect 44173 429314 44239 429317
rect 41492 429312 44239 429314
rect 41492 429256 44178 429312
rect 44234 429256 44239 429312
rect 41492 429254 44239 429256
rect 44173 429251 44239 429254
rect 44541 428906 44607 428909
rect 41492 428904 44607 428906
rect 41492 428848 44546 428904
rect 44602 428848 44607 428904
rect 41492 428846 44607 428848
rect 44541 428843 44607 428846
rect 35801 428498 35867 428501
rect 35788 428496 35867 428498
rect 35788 428440 35806 428496
rect 35862 428440 35867 428496
rect 35788 428438 35867 428440
rect 35801 428435 35867 428438
rect 41781 428498 41847 428501
rect 62389 428498 62455 428501
rect 41781 428496 62455 428498
rect 41781 428440 41786 428496
rect 41842 428440 62394 428496
rect 62450 428440 62455 428496
rect 41781 428438 62455 428440
rect 41781 428435 41847 428438
rect 62389 428435 62455 428438
rect 45093 428090 45159 428093
rect 41492 428088 45159 428090
rect 41492 428032 45098 428088
rect 45154 428032 45159 428088
rect 41492 428030 45159 428032
rect 45093 428027 45159 428030
rect 44357 427682 44423 427685
rect 41492 427680 44423 427682
rect 41492 427624 44362 427680
rect 44418 427624 44423 427680
rect 41492 427622 44423 427624
rect 44357 427619 44423 427622
rect 43621 427274 43687 427277
rect 41492 427272 43687 427274
rect 41492 427216 43626 427272
rect 43682 427216 43687 427272
rect 41492 427214 43687 427216
rect 43621 427211 43687 427214
rect 45277 426866 45343 426869
rect 41492 426864 45343 426866
rect 41492 426808 45282 426864
rect 45338 426808 45343 426864
rect 41492 426806 45343 426808
rect 45277 426803 45343 426806
rect 41454 426566 41460 426630
rect 41524 426566 41530 426630
rect 41781 426594 41847 426597
rect 42885 426594 42951 426597
rect 41781 426592 42951 426594
rect 41462 426428 41522 426566
rect 41781 426536 41786 426592
rect 41842 426536 42890 426592
rect 42946 426536 42951 426592
rect 41781 426534 42951 426536
rect 41781 426531 41847 426534
rect 42885 426531 42951 426534
rect 41137 426050 41203 426053
rect 41124 426048 41203 426050
rect 41124 425992 41142 426048
rect 41198 425992 41203 426048
rect 41124 425990 41203 425992
rect 41137 425987 41203 425990
rect 39297 425642 39363 425645
rect 39284 425640 39363 425642
rect 39284 425584 39302 425640
rect 39358 425584 39363 425640
rect 39284 425582 39363 425584
rect 39297 425579 39363 425582
rect 43989 425234 44055 425237
rect 41492 425232 44055 425234
rect 41492 425176 43994 425232
rect 44050 425176 44055 425232
rect 41492 425174 44055 425176
rect 43989 425171 44055 425174
rect 33041 424826 33107 424829
rect 33028 424824 33107 424826
rect 33028 424768 33046 424824
rect 33102 424768 33107 424824
rect 33028 424766 33107 424768
rect 33041 424763 33107 424766
rect 34513 424418 34579 424421
rect 34500 424416 34579 424418
rect 34500 424360 34518 424416
rect 34574 424360 34579 424416
rect 34500 424358 34579 424360
rect 34513 424355 34579 424358
rect 33777 424010 33843 424013
rect 33764 424008 33843 424010
rect 33764 423952 33782 424008
rect 33838 423952 33843 424008
rect 33764 423950 33843 423952
rect 33777 423947 33843 423950
rect 43805 423602 43871 423605
rect 41492 423600 43871 423602
rect 41492 423544 43810 423600
rect 43866 423544 43871 423600
rect 41492 423542 43871 423544
rect 43805 423539 43871 423542
rect 44633 423194 44699 423197
rect 41492 423192 44699 423194
rect 41492 423136 44638 423192
rect 44694 423136 44699 423192
rect 41492 423134 44699 423136
rect 44633 423131 44699 423134
rect 42701 422786 42767 422789
rect 41492 422784 42767 422786
rect 41492 422728 42706 422784
rect 42762 422728 42767 422784
rect 41492 422726 42767 422728
rect 42701 422723 42767 422726
rect 40910 422312 40970 422348
rect 40902 422248 40908 422312
rect 40972 422248 40978 422312
rect 41873 421970 41939 421973
rect 41492 421968 41939 421970
rect 41492 421912 41878 421968
rect 41934 421912 41939 421968
rect 41492 421910 41939 421912
rect 41873 421907 41939 421910
rect 41822 421562 41828 421564
rect 41492 421502 41828 421562
rect 41822 421500 41828 421502
rect 41892 421500 41898 421564
rect 45001 421154 45067 421157
rect 41492 421152 45067 421154
rect 41492 421096 45006 421152
rect 45062 421096 45067 421152
rect 41492 421094 45067 421096
rect 45001 421091 45067 421094
rect 43621 420746 43687 420749
rect 41492 420744 43687 420746
rect 41492 420688 43626 420744
rect 43682 420688 43687 420744
rect 41492 420686 43687 420688
rect 43621 420683 43687 420686
rect 41462 419930 41522 420308
rect 50521 419930 50587 419933
rect 41462 419928 50587 419930
rect 41462 419900 50526 419928
rect 41492 419872 50526 419900
rect 50582 419872 50587 419928
rect 41492 419870 50587 419872
rect 50521 419867 50587 419870
rect 40718 418644 40724 418708
rect 40788 418706 40794 418708
rect 41873 418706 41939 418709
rect 40788 418704 41939 418706
rect 40788 418648 41878 418704
rect 41934 418648 41939 418704
rect 40788 418646 41939 418648
rect 40788 418644 40794 418646
rect 41873 418643 41939 418646
rect 40534 418372 40540 418436
rect 40604 418434 40610 418436
rect 41822 418434 41828 418436
rect 40604 418374 41828 418434
rect 40604 418372 40610 418374
rect 41822 418372 41828 418374
rect 41892 418372 41898 418436
rect 39297 415306 39363 415309
rect 41638 415306 41644 415308
rect 39297 415304 41644 415306
rect 39297 415248 39302 415304
rect 39358 415248 41644 415304
rect 39297 415246 41644 415248
rect 39297 415243 39363 415246
rect 41638 415244 41644 415246
rect 41708 415244 41714 415308
rect 33777 414626 33843 414629
rect 42006 414626 42012 414628
rect 33777 414624 42012 414626
rect 33777 414568 33782 414624
rect 33838 414568 42012 414624
rect 33777 414566 42012 414568
rect 33777 414563 33843 414566
rect 42006 414564 42012 414566
rect 42076 414564 42082 414628
rect 41781 413538 41847 413541
rect 41781 413536 41890 413538
rect 41781 413480 41786 413536
rect 41842 413480 41890 413536
rect 41781 413475 41890 413480
rect 41830 413133 41890 413475
rect 41781 413128 41890 413133
rect 41781 413072 41786 413128
rect 41842 413072 41890 413128
rect 41781 413070 41890 413072
rect 41781 413067 41847 413070
rect 42425 407962 42491 407965
rect 51073 407962 51139 407965
rect 42425 407960 51139 407962
rect 42425 407904 42430 407960
rect 42486 407904 51078 407960
rect 51134 407904 51139 407960
rect 42425 407902 51139 407904
rect 42425 407899 42491 407902
rect 51073 407899 51139 407902
rect 42057 407554 42123 407557
rect 45001 407554 45067 407557
rect 42057 407552 45067 407554
rect 42057 407496 42062 407552
rect 42118 407496 45006 407552
rect 45062 407496 45067 407552
rect 42057 407494 45067 407496
rect 42057 407491 42123 407494
rect 45001 407491 45067 407494
rect 40902 406948 40908 407012
rect 40972 407010 40978 407012
rect 41781 407010 41847 407013
rect 40972 407008 41847 407010
rect 40972 406952 41786 407008
rect 41842 406952 41847 407008
rect 40972 406950 41847 406952
rect 40972 406948 40978 406950
rect 41781 406947 41847 406950
rect 40534 406676 40540 406740
rect 40604 406738 40610 406740
rect 41781 406738 41847 406741
rect 40604 406736 41847 406738
rect 40604 406680 41786 406736
rect 41842 406680 41847 406736
rect 40604 406678 41847 406680
rect 40604 406676 40610 406678
rect 41781 406675 41847 406678
rect 42425 404970 42491 404973
rect 51441 404970 51507 404973
rect 42425 404968 51507 404970
rect 42425 404912 42430 404968
rect 42486 404912 51446 404968
rect 51502 404912 51507 404968
rect 42425 404910 51507 404912
rect 42425 404907 42491 404910
rect 51441 404907 51507 404910
rect 40718 404500 40724 404564
rect 40788 404562 40794 404564
rect 42241 404562 42307 404565
rect 40788 404560 42307 404562
rect 40788 404504 42246 404560
rect 42302 404504 42307 404560
rect 40788 404502 42307 404504
rect 40788 404500 40794 404502
rect 42241 404499 42307 404502
rect 62113 404154 62179 404157
rect 62113 404152 64706 404154
rect 62113 404096 62118 404152
rect 62174 404096 64706 404152
rect 62113 404094 64706 404096
rect 62113 404091 62179 404094
rect 64646 403550 64706 404094
rect 676262 403746 676322 403852
rect 663750 403686 676322 403746
rect 663057 403338 663123 403341
rect 663750 403338 663810 403686
rect 676262 403341 676322 403444
rect 663057 403336 663810 403338
rect 663057 403280 663062 403336
rect 663118 403280 663810 403336
rect 663057 403278 663810 403280
rect 676213 403336 676322 403341
rect 676213 403280 676218 403336
rect 676274 403280 676322 403336
rect 676213 403278 676322 403280
rect 663057 403275 663123 403278
rect 676213 403275 676279 403278
rect 676630 402933 676690 403036
rect 42333 402930 42399 402933
rect 44633 402930 44699 402933
rect 42333 402928 44699 402930
rect 42333 402872 42338 402928
rect 42394 402872 44638 402928
rect 44694 402872 44699 402928
rect 42333 402870 44699 402872
rect 42333 402867 42399 402870
rect 44633 402867 44699 402870
rect 676581 402928 676690 402933
rect 676581 402872 676586 402928
rect 676642 402872 676690 402928
rect 676581 402870 676690 402872
rect 676581 402867 676647 402870
rect 62113 402658 62179 402661
rect 674833 402658 674899 402661
rect 62113 402656 64706 402658
rect 62113 402600 62118 402656
rect 62174 402600 64706 402656
rect 62113 402598 64706 402600
rect 62113 402595 62179 402598
rect 42425 402522 42491 402525
rect 43805 402522 43871 402525
rect 42425 402520 43871 402522
rect 42425 402464 42430 402520
rect 42486 402464 43810 402520
rect 43866 402464 43871 402520
rect 42425 402462 43871 402464
rect 42425 402459 42491 402462
rect 43805 402459 43871 402462
rect 64646 402368 64706 402598
rect 674833 402656 676292 402658
rect 674833 402600 674838 402656
rect 674894 402600 676292 402656
rect 674833 402598 676292 402600
rect 674833 402595 674899 402598
rect 673177 402386 673243 402389
rect 673177 402384 676322 402386
rect 673177 402328 673182 402384
rect 673238 402328 676322 402384
rect 673177 402326 676322 402328
rect 673177 402323 673243 402326
rect 676262 402220 676322 402326
rect 672441 402114 672507 402117
rect 674833 402114 674899 402117
rect 672441 402112 674899 402114
rect 672441 402056 672446 402112
rect 672502 402056 674838 402112
rect 674894 402056 674899 402112
rect 672441 402054 674899 402056
rect 672441 402051 672507 402054
rect 674833 402051 674899 402054
rect 42425 401978 42491 401981
rect 43989 401978 44055 401981
rect 42425 401976 44055 401978
rect 42425 401920 42430 401976
rect 42486 401920 43994 401976
rect 44050 401920 44055 401976
rect 42425 401918 44055 401920
rect 42425 401915 42491 401918
rect 43989 401915 44055 401918
rect 672625 401706 672691 401709
rect 676262 401706 676322 401812
rect 672625 401704 676322 401706
rect 672625 401648 672630 401704
rect 672686 401648 676322 401704
rect 672625 401646 676322 401648
rect 672625 401643 672691 401646
rect 673913 401434 673979 401437
rect 673913 401432 676292 401434
rect 673913 401376 673918 401432
rect 673974 401376 676292 401432
rect 673913 401374 676292 401376
rect 673913 401371 673979 401374
rect 677174 401236 677180 401300
rect 677244 401236 677250 401300
rect 62113 400618 62179 400621
rect 64646 400618 64706 401186
rect 677182 400996 677242 401236
rect 652017 400890 652083 400893
rect 676581 400890 676647 400893
rect 652017 400888 676647 400890
rect 652017 400832 652022 400888
rect 652078 400832 676586 400888
rect 676642 400832 676647 400888
rect 652017 400830 676647 400832
rect 652017 400827 652083 400830
rect 676581 400827 676647 400830
rect 62113 400616 64706 400618
rect 62113 400560 62118 400616
rect 62174 400560 64706 400616
rect 62113 400558 64706 400560
rect 62113 400555 62179 400558
rect 673361 400482 673427 400485
rect 676262 400482 676322 400588
rect 673361 400480 676322 400482
rect 673361 400424 673366 400480
rect 673422 400424 676322 400480
rect 673361 400422 676322 400424
rect 673361 400419 673427 400422
rect 676806 400420 676812 400484
rect 676876 400420 676882 400484
rect 62389 400210 62455 400213
rect 62389 400208 64706 400210
rect 62389 400152 62394 400208
rect 62450 400152 64706 400208
rect 676814 400180 676874 400420
rect 62389 400150 64706 400152
rect 62389 400147 62455 400150
rect 41454 400012 41460 400076
rect 41524 400074 41530 400076
rect 41781 400074 41847 400077
rect 41524 400072 41847 400074
rect 41524 400016 41786 400072
rect 41842 400016 41847 400072
rect 41524 400014 41847 400016
rect 41524 400012 41530 400014
rect 41781 400011 41847 400014
rect 64646 400004 64706 400150
rect 672165 399666 672231 399669
rect 676262 399666 676322 399772
rect 672165 399664 676322 399666
rect 672165 399608 672170 399664
rect 672226 399608 676322 399664
rect 672165 399606 676322 399608
rect 672165 399603 672231 399606
rect 41965 399396 42031 399397
rect 41965 399392 42012 399396
rect 42076 399394 42082 399396
rect 62113 399394 62179 399397
rect 676029 399394 676095 399397
rect 41965 399336 41970 399392
rect 41965 399332 42012 399336
rect 42076 399334 42122 399394
rect 62113 399392 64706 399394
rect 62113 399336 62118 399392
rect 62174 399336 64706 399392
rect 62113 399334 64706 399336
rect 42076 399332 42082 399334
rect 41965 399331 42031 399332
rect 62113 399331 62179 399334
rect 41781 398852 41847 398853
rect 41781 398848 41828 398852
rect 41892 398850 41898 398852
rect 41781 398792 41786 398848
rect 41781 398788 41828 398792
rect 41892 398790 41938 398850
rect 64646 398822 64706 399334
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 41892 398788 41898 398790
rect 676070 398788 676076 398852
rect 676140 398850 676146 398852
rect 676262 398850 676322 398956
rect 676140 398790 676322 398850
rect 676140 398788 676146 398790
rect 41781 398787 41847 398788
rect 679574 398445 679634 398548
rect 679574 398440 679683 398445
rect 679574 398384 679622 398440
rect 679678 398384 679683 398440
rect 679574 398382 679683 398384
rect 679617 398379 679683 398382
rect 62113 398306 62179 398309
rect 62113 398304 64706 398306
rect 62113 398248 62118 398304
rect 62174 398248 64706 398304
rect 62113 398246 64706 398248
rect 62113 398243 62179 398246
rect 64646 397640 64706 398246
rect 676262 398037 676322 398140
rect 676213 398032 676322 398037
rect 676213 397976 676218 398032
rect 676274 397976 676322 398032
rect 676213 397974 676322 397976
rect 676213 397971 676279 397974
rect 678286 397629 678346 397732
rect 678237 397624 678346 397629
rect 678237 397568 678242 397624
rect 678298 397568 678346 397624
rect 678237 397566 678346 397568
rect 678237 397563 678303 397566
rect 42149 397490 42215 397493
rect 51073 397490 51139 397493
rect 42149 397488 51139 397490
rect 42149 397432 42154 397488
rect 42210 397432 51078 397488
rect 51134 397432 51139 397488
rect 42149 397430 51139 397432
rect 42149 397427 42215 397430
rect 51073 397427 51139 397430
rect 674741 397354 674807 397357
rect 674741 397352 676292 397354
rect 674741 397296 674746 397352
rect 674802 397296 676292 397352
rect 674741 397294 676292 397296
rect 674741 397291 674807 397294
rect 676262 396812 676322 396916
rect 676254 396748 676260 396812
rect 676324 396748 676330 396812
rect 652201 396674 652267 396677
rect 674557 396674 674623 396677
rect 652201 396672 674623 396674
rect 652201 396616 652206 396672
rect 652262 396616 674562 396672
rect 674618 396616 674623 396672
rect 652201 396614 674623 396616
rect 652201 396611 652267 396614
rect 674557 396611 674623 396614
rect 676446 396404 676506 396508
rect 676438 396340 676444 396404
rect 676508 396340 676514 396404
rect 673729 396130 673795 396133
rect 673729 396128 676292 396130
rect 673729 396072 673734 396128
rect 673790 396072 676292 396128
rect 673729 396070 676292 396072
rect 673729 396067 673795 396070
rect 676262 395589 676322 395692
rect 676213 395584 676322 395589
rect 676213 395528 676218 395584
rect 676274 395528 676322 395584
rect 676213 395526 676322 395528
rect 676213 395523 676279 395526
rect 676630 395180 676690 395284
rect 676622 395116 676628 395180
rect 676692 395116 676698 395180
rect 672993 394770 673059 394773
rect 676262 394770 676322 394876
rect 672993 394768 676322 394770
rect 672993 394712 672998 394768
rect 673054 394712 676322 394768
rect 672993 394710 676322 394712
rect 672993 394707 673059 394710
rect 676262 394365 676322 394468
rect 676213 394360 676322 394365
rect 676213 394304 676218 394360
rect 676274 394304 676322 394360
rect 676213 394302 676322 394304
rect 676213 394299 676279 394302
rect 672809 393954 672875 393957
rect 676262 393954 676322 394060
rect 672809 393952 676322 393954
rect 672809 393896 672814 393952
rect 672870 393896 676322 393952
rect 672809 393894 676322 393896
rect 672809 393891 672875 393894
rect 671889 393546 671955 393549
rect 676262 393546 676322 393652
rect 671889 393544 676322 393546
rect 671889 393488 671894 393544
rect 671950 393488 676322 393544
rect 671889 393486 676322 393488
rect 671889 393483 671955 393486
rect 675886 392804 675892 392868
rect 675956 392866 675962 392868
rect 676262 392866 676322 393244
rect 675956 392836 676322 392866
rect 675956 392806 676292 392836
rect 675956 392804 675962 392806
rect 670509 392594 670575 392597
rect 670509 392592 676322 392594
rect 670509 392536 670514 392592
rect 670570 392536 676322 392592
rect 670509 392534 676322 392536
rect 670509 392531 670575 392534
rect 676262 392428 676322 392534
rect 41462 387562 41522 387668
rect 675702 387636 675708 387700
rect 675772 387698 675778 387700
rect 678237 387698 678303 387701
rect 675772 387696 678303 387698
rect 675772 387640 678242 387696
rect 678298 387640 678303 387696
rect 675772 387638 678303 387640
rect 675772 387636 675778 387638
rect 678237 387635 678303 387638
rect 54477 387562 54543 387565
rect 41462 387560 54543 387562
rect 41462 387504 54482 387560
rect 54538 387504 54543 387560
rect 41462 387502 54543 387504
rect 54477 387499 54543 387502
rect 41278 387157 41338 387260
rect 41278 387152 41387 387157
rect 41278 387096 41326 387152
rect 41382 387096 41387 387152
rect 41278 387094 41387 387096
rect 41321 387091 41387 387094
rect 41094 386749 41154 386852
rect 41094 386744 41203 386749
rect 41094 386688 41142 386744
rect 41198 386688 41203 386744
rect 41094 386686 41203 386688
rect 41137 386683 41203 386686
rect 44173 386474 44239 386477
rect 41492 386472 44239 386474
rect 41492 386416 44178 386472
rect 44234 386416 44239 386472
rect 41492 386414 44239 386416
rect 44173 386411 44239 386414
rect 40910 385933 40970 386036
rect 40861 385928 40970 385933
rect 40861 385872 40866 385928
rect 40922 385872 40970 385928
rect 40861 385870 40970 385872
rect 41137 385930 41203 385933
rect 63125 385930 63191 385933
rect 41137 385928 63191 385930
rect 41137 385872 41142 385928
rect 41198 385872 63130 385928
rect 63186 385872 63191 385928
rect 41137 385870 63191 385872
rect 40861 385867 40927 385870
rect 41137 385867 41203 385870
rect 63125 385867 63191 385870
rect 42885 385658 42951 385661
rect 41492 385656 42951 385658
rect 41492 385600 42890 385656
rect 42946 385600 42951 385656
rect 41492 385598 42951 385600
rect 42885 385595 42951 385598
rect 45093 385250 45159 385253
rect 41492 385248 45159 385250
rect 41492 385192 45098 385248
rect 45154 385192 45159 385248
rect 41492 385190 45159 385192
rect 45093 385187 45159 385190
rect 675753 384978 675819 384981
rect 676254 384978 676260 384980
rect 675753 384976 676260 384978
rect 675753 384920 675758 384976
rect 675814 384920 676260 384976
rect 675753 384918 676260 384920
rect 675753 384915 675819 384918
rect 676254 384916 676260 384918
rect 676324 384916 676330 384980
rect 44357 384842 44423 384845
rect 41492 384840 44423 384842
rect 41492 384784 44362 384840
rect 44418 384784 44423 384840
rect 41492 384782 44423 384784
rect 44357 384779 44423 384782
rect 44909 384434 44975 384437
rect 41492 384432 44975 384434
rect 41492 384376 44914 384432
rect 44970 384376 44975 384432
rect 41492 384374 44975 384376
rect 44909 384371 44975 384374
rect 45277 384026 45343 384029
rect 41492 384024 45343 384026
rect 41492 383968 45282 384024
rect 45338 383968 45343 384024
rect 41492 383966 45343 383968
rect 45277 383963 45343 383966
rect 45277 383618 45343 383621
rect 41492 383616 45343 383618
rect 41492 383560 45282 383616
rect 45338 383560 45343 383616
rect 41492 383558 45343 383560
rect 45277 383555 45343 383558
rect 41094 383077 41154 383180
rect 41045 383072 41154 383077
rect 41321 383074 41387 383077
rect 41045 383016 41050 383072
rect 41106 383016 41154 383072
rect 41045 383014 41154 383016
rect 41278 383072 41387 383074
rect 41278 383016 41326 383072
rect 41382 383016 41387 383072
rect 41045 383011 41111 383014
rect 41278 383011 41387 383016
rect 41278 382772 41338 383011
rect 654777 382938 654843 382941
rect 675201 382938 675267 382941
rect 654777 382936 675267 382938
rect 654777 382880 654782 382936
rect 654838 382880 675206 382936
rect 675262 382880 675267 382936
rect 654777 382878 675267 382880
rect 654777 382875 654843 382878
rect 675201 382875 675267 382878
rect 40861 382666 40927 382669
rect 45461 382666 45527 382669
rect 40861 382664 45527 382666
rect 40861 382608 40866 382664
rect 40922 382608 45466 382664
rect 45522 382608 45527 382664
rect 40861 382606 45527 382608
rect 40861 382603 40927 382606
rect 45461 382603 45527 382606
rect 39990 382261 40050 382364
rect 39990 382256 40099 382261
rect 39990 382200 40038 382256
rect 40094 382200 40099 382256
rect 39990 382198 40099 382200
rect 40033 382195 40099 382198
rect 675753 382258 675819 382261
rect 676438 382258 676444 382260
rect 675753 382256 676444 382258
rect 675753 382200 675758 382256
rect 675814 382200 676444 382256
rect 675753 382198 676444 382200
rect 675753 382195 675819 382198
rect 676438 382196 676444 382198
rect 676508 382196 676514 382260
rect 35574 381853 35634 381956
rect 35525 381848 35634 381853
rect 35525 381792 35530 381848
rect 35586 381792 35634 381848
rect 35525 381790 35634 381792
rect 41045 381850 41111 381853
rect 41454 381850 41460 381852
rect 41045 381848 41460 381850
rect 41045 381792 41050 381848
rect 41106 381792 41460 381848
rect 41045 381790 41460 381792
rect 35525 381787 35591 381790
rect 41045 381787 41111 381790
rect 41454 381788 41460 381790
rect 41524 381788 41530 381852
rect 41781 381578 41847 381581
rect 62757 381578 62823 381581
rect 41781 381576 62823 381578
rect 39254 381445 39314 381548
rect 41781 381520 41786 381576
rect 41842 381520 62762 381576
rect 62818 381520 62823 381576
rect 41781 381518 62823 381520
rect 41781 381515 41847 381518
rect 62757 381515 62823 381518
rect 39254 381440 39363 381445
rect 39254 381384 39302 381440
rect 39358 381384 39363 381440
rect 39254 381382 39363 381384
rect 39297 381379 39363 381382
rect 673729 381442 673795 381445
rect 675109 381442 675175 381445
rect 673729 381440 675175 381442
rect 673729 381384 673734 381440
rect 673790 381384 675114 381440
rect 675170 381384 675175 381440
rect 673729 381382 675175 381384
rect 673729 381379 673795 381382
rect 675109 381379 675175 381382
rect 33918 381037 33978 381140
rect 33918 381032 34027 381037
rect 33918 380976 33966 381032
rect 34022 380976 34027 381032
rect 33918 380974 34027 380976
rect 33961 380971 34027 380974
rect 672993 381034 673059 381037
rect 675385 381034 675451 381037
rect 672993 381032 675451 381034
rect 672993 380976 672998 381032
rect 673054 380976 675390 381032
rect 675446 380976 675451 381032
rect 672993 380974 675451 380976
rect 672993 380971 673059 380974
rect 675385 380971 675451 380974
rect 46933 380762 46999 380765
rect 41492 380760 46999 380762
rect 41492 380704 46938 380760
rect 46994 380704 46999 380760
rect 41492 380702 46999 380704
rect 46933 380699 46999 380702
rect 44541 380354 44607 380357
rect 41492 380352 44607 380354
rect 41492 380296 44546 380352
rect 44602 380296 44607 380352
rect 41492 380294 44607 380296
rect 44541 380291 44607 380294
rect 42885 379946 42951 379949
rect 41492 379944 42951 379946
rect 41492 379888 42890 379944
rect 42946 379888 42951 379944
rect 41492 379886 42951 379888
rect 42885 379883 42951 379886
rect 35758 379405 35818 379530
rect 35758 379400 35867 379405
rect 35758 379344 35806 379400
rect 35862 379344 35867 379400
rect 35758 379342 35867 379344
rect 35801 379339 35867 379342
rect 40033 379402 40099 379405
rect 41822 379402 41828 379404
rect 40033 379400 41828 379402
rect 40033 379344 40038 379400
rect 40094 379344 41828 379400
rect 40033 379342 41828 379344
rect 40033 379339 40099 379342
rect 41822 379340 41828 379342
rect 41892 379340 41898 379404
rect 40726 378996 40786 379100
rect 40718 378932 40724 378996
rect 40788 378932 40794 378996
rect 675753 378724 675819 378725
rect 675702 378722 675708 378724
rect 40542 378588 40602 378692
rect 675662 378662 675708 378722
rect 675772 378720 675819 378724
rect 675814 378664 675819 378720
rect 675702 378660 675708 378662
rect 675772 378660 675819 378664
rect 675753 378659 675819 378660
rect 40534 378524 40540 378588
rect 40604 378524 40610 378588
rect 44173 378314 44239 378317
rect 41492 378312 44239 378314
rect 41492 378256 44178 378312
rect 44234 378256 44239 378312
rect 41492 378254 44239 378256
rect 44173 378251 44239 378254
rect 40910 377772 40970 377876
rect 40902 377708 40908 377772
rect 40972 377708 40978 377772
rect 35758 377365 35818 377468
rect 35758 377360 35867 377365
rect 35758 377304 35806 377360
rect 35862 377304 35867 377360
rect 35758 377302 35867 377304
rect 35801 377299 35867 377302
rect 40401 377362 40467 377365
rect 43069 377362 43135 377365
rect 40401 377360 43135 377362
rect 40401 377304 40406 377360
rect 40462 377304 43074 377360
rect 43130 377304 43135 377360
rect 40401 377302 43135 377304
rect 40401 377299 40467 377302
rect 43069 377299 43135 377302
rect 675753 377362 675819 377365
rect 676622 377362 676628 377364
rect 675753 377360 676628 377362
rect 675753 377304 675758 377360
rect 675814 377304 676628 377360
rect 675753 377302 676628 377304
rect 675753 377299 675819 377302
rect 676622 377300 676628 377302
rect 676692 377300 676698 377364
rect 35758 376549 35818 377060
rect 41462 376549 41522 376652
rect 35758 376544 35867 376549
rect 35758 376488 35806 376544
rect 35862 376488 35867 376544
rect 35758 376486 35867 376488
rect 41462 376544 41571 376549
rect 41462 376488 41510 376544
rect 41566 376488 41571 376544
rect 41462 376486 41571 376488
rect 35801 376483 35867 376486
rect 41505 376483 41571 376486
rect 41689 376546 41755 376549
rect 43805 376546 43871 376549
rect 41689 376544 43871 376546
rect 41689 376488 41694 376544
rect 41750 376488 43810 376544
rect 43866 376488 43871 376544
rect 41689 376486 43871 376488
rect 41689 376483 41755 376486
rect 43805 376483 43871 376486
rect 672809 376274 672875 376277
rect 675385 376274 675451 376277
rect 672809 376272 675451 376274
rect 672809 376216 672814 376272
rect 672870 376216 675390 376272
rect 675446 376216 675451 376272
rect 672809 376214 675451 376216
rect 672809 376211 672875 376214
rect 675385 376211 675451 376214
rect 35801 376138 35867 376141
rect 41505 376138 41571 376141
rect 47577 376138 47643 376141
rect 35801 376136 47643 376138
rect 35801 376080 35806 376136
rect 35862 376080 41510 376136
rect 41566 376080 47582 376136
rect 47638 376080 47643 376136
rect 35801 376078 47643 376080
rect 35801 376075 35867 376078
rect 41505 376075 41571 376078
rect 47577 376075 47643 376078
rect 35525 374642 35591 374645
rect 41638 374642 41644 374644
rect 35525 374640 41644 374642
rect 35525 374584 35530 374640
rect 35586 374584 41644 374640
rect 35525 374582 41644 374584
rect 35525 374579 35591 374582
rect 41638 374580 41644 374582
rect 41708 374580 41714 374644
rect 652201 373962 652267 373965
rect 649950 373960 652267 373962
rect 649950 373904 652206 373960
rect 652262 373904 652267 373960
rect 649950 373902 652267 373904
rect 649950 373892 650010 373902
rect 652201 373899 652267 373902
rect 675753 373690 675819 373693
rect 676070 373690 676076 373692
rect 675753 373688 676076 373690
rect 675753 373632 675758 373688
rect 675814 373632 676076 373688
rect 675753 373630 676076 373632
rect 675753 373627 675819 373630
rect 676070 373628 676076 373630
rect 676140 373628 676146 373692
rect 651465 373282 651531 373285
rect 649950 373280 651531 373282
rect 649950 373224 651470 373280
rect 651526 373224 651531 373280
rect 649950 373222 651531 373224
rect 649950 372710 650010 373222
rect 651465 373219 651531 373222
rect 675385 372468 675451 372469
rect 675334 372404 675340 372468
rect 675404 372466 675451 372468
rect 675404 372464 675496 372466
rect 675446 372408 675496 372464
rect 675404 372406 675496 372408
rect 675404 372404 675451 372406
rect 675385 372403 675451 372404
rect 652017 372194 652083 372197
rect 649950 372192 652083 372194
rect 649950 372136 652022 372192
rect 652078 372136 652083 372192
rect 649950 372134 652083 372136
rect 649950 371528 650010 372134
rect 652017 372131 652083 372134
rect 651465 370698 651531 370701
rect 649950 370696 651531 370698
rect 649950 370640 651470 370696
rect 651526 370640 651531 370696
rect 649950 370638 651531 370640
rect 649950 370346 650010 370638
rect 651465 370635 651531 370638
rect 42057 366210 42123 366213
rect 43069 366210 43135 366213
rect 42057 366208 43135 366210
rect 42057 366152 42062 366208
rect 42118 366152 43074 366208
rect 43130 366152 43135 366208
rect 42057 366150 43135 366152
rect 42057 366147 42123 366150
rect 43069 366147 43135 366150
rect 41822 365740 41828 365804
rect 41892 365802 41898 365804
rect 42609 365802 42675 365805
rect 41892 365800 42675 365802
rect 41892 365744 42614 365800
rect 42670 365744 42675 365800
rect 41892 365742 42675 365744
rect 41892 365740 41898 365742
rect 42609 365739 42675 365742
rect 666461 365666 666527 365669
rect 675334 365666 675340 365668
rect 666461 365664 675340 365666
rect 666461 365608 666466 365664
rect 666522 365608 675340 365664
rect 666461 365606 675340 365608
rect 666461 365603 666527 365606
rect 675334 365604 675340 365606
rect 675404 365604 675410 365668
rect 40902 364788 40908 364852
rect 40972 364850 40978 364852
rect 41781 364850 41847 364853
rect 40972 364848 41847 364850
rect 40972 364792 41786 364848
rect 41842 364792 41847 364848
rect 40972 364790 41847 364792
rect 40972 364788 40978 364790
rect 41781 364787 41847 364790
rect 43069 364306 43135 364309
rect 44725 364306 44791 364309
rect 43069 364304 44791 364306
rect 43069 364248 43074 364304
rect 43130 364248 44730 364304
rect 44786 364248 44791 364304
rect 43069 364246 44791 364248
rect 43069 364243 43135 364246
rect 44725 364243 44791 364246
rect 40718 364108 40724 364172
rect 40788 364170 40794 364172
rect 41781 364170 41847 364173
rect 40788 364168 41847 364170
rect 40788 364112 41786 364168
rect 41842 364112 41847 364168
rect 40788 364110 41847 364112
rect 40788 364108 40794 364110
rect 41781 364107 41847 364110
rect 42057 363626 42123 363629
rect 44173 363626 44239 363629
rect 42057 363624 44239 363626
rect 42057 363568 42062 363624
rect 42118 363568 44178 363624
rect 44234 363568 44239 363624
rect 42057 363566 44239 363568
rect 42057 363563 42123 363566
rect 44173 363563 44239 363566
rect 42241 362266 42307 362269
rect 51073 362266 51139 362269
rect 42241 362264 51139 362266
rect 42241 362208 42246 362264
rect 42302 362208 51078 362264
rect 51134 362208 51139 362264
rect 42241 362206 51139 362208
rect 42241 362203 42307 362206
rect 51073 362203 51139 362206
rect 62113 360906 62179 360909
rect 62113 360904 64706 360906
rect 62113 360848 62118 360904
rect 62174 360848 64706 360904
rect 62113 360846 64706 360848
rect 62113 360843 62179 360846
rect 64646 360328 64706 360846
rect 40534 360028 40540 360092
rect 40604 360090 40610 360092
rect 41781 360090 41847 360093
rect 40604 360088 41847 360090
rect 40604 360032 41786 360088
rect 41842 360032 41847 360088
rect 40604 360030 41847 360032
rect 40604 360028 40610 360030
rect 41781 360027 41847 360030
rect 62113 359818 62179 359821
rect 62113 359816 64706 359818
rect 62113 359760 62118 359816
rect 62174 359760 64706 359816
rect 62113 359758 64706 359760
rect 62113 359755 62179 359758
rect 64646 359146 64706 359758
rect 42425 359002 42491 359005
rect 44541 359002 44607 359005
rect 42425 359000 44607 359002
rect 42425 358944 42430 359000
rect 42486 358944 44546 359000
rect 44602 358944 44607 359000
rect 42425 358942 44607 358944
rect 42425 358939 42491 358942
rect 44541 358939 44607 358942
rect 41873 358732 41939 358733
rect 41822 358730 41828 358732
rect 41782 358670 41828 358730
rect 41892 358728 41939 358732
rect 41934 358672 41939 358728
rect 41822 358668 41828 358670
rect 41892 358668 41939 358672
rect 41873 358667 41939 358668
rect 663750 358670 676292 358730
rect 654777 358594 654843 358597
rect 663750 358594 663810 358670
rect 654777 358592 663810 358594
rect 654777 358536 654782 358592
rect 654838 358536 663810 358592
rect 654777 358534 663810 358536
rect 654777 358531 654843 358534
rect 674465 358322 674531 358325
rect 674465 358320 676292 358322
rect 674465 358264 674470 358320
rect 674526 358264 676292 358320
rect 674465 358262 676292 358264
rect 674465 358259 674531 358262
rect 62297 357506 62363 357509
rect 64646 357506 64706 357964
rect 675937 357914 676003 357917
rect 675937 357912 676292 357914
rect 675937 357856 675942 357912
rect 675998 357856 676292 357912
rect 675937 357854 676292 357856
rect 675937 357851 676003 357854
rect 62297 357504 64706 357506
rect 62297 357448 62302 357504
rect 62358 357448 64706 357504
rect 62297 357446 64706 357448
rect 673177 357506 673243 357509
rect 673177 357504 676292 357506
rect 673177 357448 673182 357504
rect 673238 357448 676292 357504
rect 673177 357446 676292 357448
rect 62297 357443 62363 357446
rect 673177 357443 673243 357446
rect 63125 357234 63191 357237
rect 63125 357232 64706 357234
rect 63125 357176 63130 357232
rect 63186 357176 64706 357232
rect 63125 357174 64706 357176
rect 63125 357171 63191 357174
rect 41454 356900 41460 356964
rect 41524 356962 41530 356964
rect 41781 356962 41847 356965
rect 41524 356960 41847 356962
rect 41524 356904 41786 356960
rect 41842 356904 41847 356960
rect 41524 356902 41847 356904
rect 41524 356900 41530 356902
rect 41781 356899 41847 356902
rect 64646 356782 64706 357174
rect 672349 357098 672415 357101
rect 672349 357096 676292 357098
rect 672349 357040 672354 357096
rect 672410 357040 676292 357096
rect 672349 357038 676292 357040
rect 672349 357035 672415 357038
rect 675937 356826 676003 356829
rect 669270 356824 676003 356826
rect 669270 356768 675942 356824
rect 675998 356768 676003 356824
rect 669270 356766 676003 356768
rect 42793 356690 42859 356693
rect 62297 356690 62363 356693
rect 42793 356688 62363 356690
rect 42793 356632 42798 356688
rect 42854 356632 62302 356688
rect 62358 356632 62363 356688
rect 42793 356630 62363 356632
rect 42793 356627 42859 356630
rect 62297 356627 62363 356630
rect 652201 356690 652267 356693
rect 669270 356690 669330 356766
rect 675937 356763 676003 356766
rect 652201 356688 669330 356690
rect 652201 356632 652206 356688
rect 652262 356632 669330 356688
rect 652201 356630 669330 356632
rect 676170 356630 676292 356690
rect 652201 356627 652267 356630
rect 673913 356554 673979 356557
rect 676170 356554 676230 356630
rect 673913 356552 676230 356554
rect 673913 356496 673918 356552
rect 673974 356496 676230 356552
rect 673913 356494 676230 356496
rect 673913 356491 673979 356494
rect 672533 356282 672599 356285
rect 672533 356280 676292 356282
rect 672533 356224 672538 356280
rect 672594 356224 676292 356280
rect 672533 356222 676292 356224
rect 672533 356219 672599 356222
rect 42241 356146 42307 356149
rect 46933 356146 46999 356149
rect 42241 356144 46999 356146
rect 42241 356088 42246 356144
rect 42302 356088 46938 356144
rect 46994 356088 46999 356144
rect 42241 356086 46999 356088
rect 42241 356083 42307 356086
rect 46933 356083 46999 356086
rect 62113 356010 62179 356013
rect 62113 356008 64706 356010
rect 62113 355952 62118 356008
rect 62174 355952 64706 356008
rect 62113 355950 64706 355952
rect 62113 355947 62179 355950
rect 43805 355874 43871 355877
rect 46013 355874 46079 355877
rect 43805 355872 46079 355874
rect 43805 355816 43810 355872
rect 43866 355816 46018 355872
rect 46074 355816 46079 355872
rect 43805 355814 46079 355816
rect 43805 355811 43871 355814
rect 46013 355811 46079 355814
rect 43621 355602 43687 355605
rect 45829 355602 45895 355605
rect 43621 355600 45895 355602
rect 64646 355600 64706 355950
rect 673361 355874 673427 355877
rect 673361 355872 676292 355874
rect 673361 355816 673366 355872
rect 673422 355816 676292 355872
rect 673361 355814 676292 355816
rect 673361 355811 673427 355814
rect 43621 355544 43626 355600
rect 43682 355544 45834 355600
rect 45890 355544 45895 355600
rect 43621 355542 45895 355544
rect 43621 355539 43687 355542
rect 45829 355539 45895 355542
rect 673177 355466 673243 355469
rect 673177 355464 676292 355466
rect 673177 355408 673182 355464
rect 673238 355408 676292 355464
rect 673177 355406 676292 355408
rect 673177 355403 673243 355406
rect 43253 355330 43319 355333
rect 44633 355330 44699 355333
rect 43253 355328 44699 355330
rect 43253 355272 43258 355328
rect 43314 355272 44638 355328
rect 44694 355272 44699 355328
rect 43253 355270 44699 355272
rect 43253 355267 43319 355270
rect 44633 355267 44699 355270
rect 672165 355058 672231 355061
rect 672165 355056 676292 355058
rect 672165 355000 672170 355056
rect 672226 355000 676292 355056
rect 672165 354998 676292 355000
rect 672165 354995 672231 354998
rect 43662 354588 43668 354652
rect 43732 354650 43738 354652
rect 43989 354650 44055 354653
rect 43732 354648 44055 354650
rect 43732 354592 43994 354648
rect 44050 354592 44055 354648
rect 43732 354590 44055 354592
rect 43732 354588 43738 354590
rect 43989 354587 44055 354590
rect 673913 354650 673979 354653
rect 673913 354648 676292 354650
rect 673913 354592 673918 354648
rect 673974 354592 676292 354648
rect 673913 354590 676292 354592
rect 673913 354587 673979 354590
rect 62757 354514 62823 354517
rect 62757 354512 64706 354514
rect 62757 354456 62762 354512
rect 62818 354456 64706 354512
rect 62757 354454 64706 354456
rect 62757 354451 62823 354454
rect 64646 354418 64706 354454
rect 42701 354378 42767 354381
rect 43989 354378 44055 354381
rect 42701 354376 44055 354378
rect 42701 354320 42706 354376
rect 42762 354320 43994 354376
rect 44050 354320 44055 354376
rect 42701 354318 44055 354320
rect 42701 354315 42767 354318
rect 43989 354315 44055 354318
rect 675518 354180 675524 354244
rect 675588 354242 675594 354244
rect 675588 354182 676292 354242
rect 675588 354180 675594 354182
rect 45645 353834 45711 353837
rect 45142 353832 45711 353834
rect 45142 353776 45650 353832
rect 45706 353776 45711 353832
rect 45142 353774 45711 353776
rect 44766 353636 44772 353700
rect 44836 353698 44842 353700
rect 45142 353698 45202 353774
rect 45645 353771 45711 353774
rect 675886 353772 675892 353836
rect 675956 353834 675962 353836
rect 675956 353774 676292 353834
rect 675956 353772 675962 353774
rect 44836 353638 45202 353698
rect 44836 353636 44842 353638
rect 672165 353426 672231 353429
rect 672165 353424 676292 353426
rect 672165 353368 672170 353424
rect 672226 353368 676292 353424
rect 672165 353366 676292 353368
rect 672165 353363 672231 353366
rect 675702 352956 675708 353020
rect 675772 353018 675778 353020
rect 675772 352958 676292 353018
rect 675772 352956 675778 352958
rect 673729 352610 673795 352613
rect 673729 352608 676292 352610
rect 673729 352552 673734 352608
rect 673790 352552 676292 352608
rect 673729 352550 676292 352552
rect 673729 352547 673795 352550
rect 44030 352140 44036 352204
rect 44100 352202 44106 352204
rect 45645 352202 45711 352205
rect 44100 352200 45711 352202
rect 44100 352144 45650 352200
rect 45706 352144 45711 352200
rect 44100 352142 45711 352144
rect 44100 352140 44106 352142
rect 45645 352139 45711 352142
rect 674649 352202 674715 352205
rect 674649 352200 676292 352202
rect 674649 352144 674654 352200
rect 674710 352144 676292 352200
rect 674649 352142 676292 352144
rect 674649 352139 674715 352142
rect 42006 351868 42012 351932
rect 42076 351930 42082 351932
rect 42701 351930 42767 351933
rect 42076 351928 42767 351930
rect 42076 351872 42706 351928
rect 42762 351872 42767 351928
rect 42076 351870 42767 351872
rect 42076 351868 42082 351870
rect 42701 351867 42767 351870
rect 675886 351732 675892 351796
rect 675956 351794 675962 351796
rect 675956 351734 676292 351794
rect 675956 351732 675962 351734
rect 674281 351386 674347 351389
rect 674281 351384 676292 351386
rect 674281 351328 674286 351384
rect 674342 351328 676292 351384
rect 674281 351326 676292 351328
rect 674281 351323 674347 351326
rect 652569 351114 652635 351117
rect 674465 351114 674531 351117
rect 652569 351112 674531 351114
rect 652569 351056 652574 351112
rect 652630 351056 674470 351112
rect 674526 351056 674531 351112
rect 652569 351054 674531 351056
rect 652569 351051 652635 351054
rect 674465 351051 674531 351054
rect 676029 350978 676095 350981
rect 676029 350976 676292 350978
rect 676029 350920 676034 350976
rect 676090 350920 676292 350976
rect 676029 350918 676292 350920
rect 676029 350915 676095 350918
rect 674465 350570 674531 350573
rect 674465 350568 676292 350570
rect 674465 350512 674470 350568
rect 674526 350512 676292 350568
rect 674465 350510 676292 350512
rect 674465 350507 674531 350510
rect 673361 350162 673427 350165
rect 673361 350160 676292 350162
rect 673361 350104 673366 350160
rect 673422 350104 676292 350160
rect 673361 350102 676292 350104
rect 673361 350099 673427 350102
rect 672993 349754 673059 349757
rect 672993 349752 676292 349754
rect 672993 349696 672998 349752
rect 673054 349696 676292 349752
rect 672993 349694 676292 349696
rect 672993 349691 673059 349694
rect 673545 349346 673611 349349
rect 673545 349344 676292 349346
rect 673545 349288 673550 349344
rect 673606 349288 676292 349344
rect 673545 349286 676292 349288
rect 673545 349283 673611 349286
rect 671705 348938 671771 348941
rect 671705 348936 676292 348938
rect 671705 348880 671710 348936
rect 671766 348880 676292 348936
rect 671705 348878 676292 348880
rect 671705 348875 671771 348878
rect 672717 348530 672783 348533
rect 672717 348528 676292 348530
rect 672717 348472 672722 348528
rect 672778 348472 676292 348528
rect 672717 348470 676292 348472
rect 672717 348467 672783 348470
rect 675334 347652 675340 347716
rect 675404 347714 675410 347716
rect 683070 347714 683130 348092
rect 675404 347684 683130 347714
rect 675404 347654 683100 347684
rect 675404 347652 675410 347654
rect 669405 347306 669471 347309
rect 669405 347304 676292 347306
rect 669405 347248 669410 347304
rect 669466 347248 676292 347304
rect 669405 347246 676292 347248
rect 669405 347243 669471 347246
rect 676029 346626 676095 346629
rect 676438 346626 676444 346628
rect 676029 346624 676444 346626
rect 676029 346568 676034 346624
rect 676090 346568 676444 346624
rect 676029 346566 676444 346568
rect 676029 346563 676095 346566
rect 676438 346564 676444 346566
rect 676508 346564 676514 346628
rect 35574 344317 35634 344556
rect 35525 344312 35634 344317
rect 35801 344314 35867 344317
rect 35525 344256 35530 344312
rect 35586 344256 35634 344312
rect 35525 344254 35634 344256
rect 35758 344312 35867 344314
rect 35758 344256 35806 344312
rect 35862 344256 35867 344312
rect 35525 344251 35591 344254
rect 35758 344251 35867 344256
rect 35758 344148 35818 344251
rect 39849 343906 39915 343909
rect 44909 343906 44975 343909
rect 39849 343904 44975 343906
rect 39849 343848 39854 343904
rect 39910 343848 44914 343904
rect 44970 343848 44975 343904
rect 39849 343846 44975 343848
rect 39849 343843 39915 343846
rect 44909 343843 44975 343846
rect 32998 343501 33058 343740
rect 32998 343496 33107 343501
rect 32998 343440 33046 343496
rect 33102 343440 33107 343496
rect 32998 343438 33107 343440
rect 33041 343435 33107 343438
rect 40033 343498 40099 343501
rect 45001 343498 45067 343501
rect 40033 343496 45067 343498
rect 40033 343440 40038 343496
rect 40094 343440 45006 343496
rect 45062 343440 45067 343496
rect 40033 343438 45067 343440
rect 40033 343435 40099 343438
rect 45001 343435 45067 343438
rect 41462 343226 41522 343332
rect 45461 343226 45527 343229
rect 41462 343224 45527 343226
rect 41462 343168 45466 343224
rect 45522 343168 45527 343224
rect 41462 343166 45527 343168
rect 45461 343163 45527 343166
rect 41462 342818 41522 342924
rect 45553 342818 45619 342821
rect 41462 342816 45619 342818
rect 41462 342760 45558 342816
rect 45614 342760 45619 342816
rect 41462 342758 45619 342760
rect 45553 342755 45619 342758
rect 45185 342546 45251 342549
rect 41492 342544 45251 342546
rect 41492 342488 45190 342544
rect 45246 342488 45251 342544
rect 41492 342486 45251 342488
rect 45185 342483 45251 342486
rect 40217 342274 40283 342277
rect 40217 342272 42074 342274
rect 40217 342216 40222 342272
rect 40278 342216 42074 342272
rect 40217 342214 42074 342216
rect 40217 342211 40283 342214
rect 42014 342138 42074 342214
rect 50102 342138 50108 342140
rect 35801 341866 35867 341869
rect 35758 341864 35867 341866
rect 35758 341808 35806 341864
rect 35862 341808 35867 341864
rect 35758 341803 35867 341808
rect 41462 341866 41522 342108
rect 42014 342078 50108 342138
rect 50102 342076 50108 342078
rect 50172 342076 50178 342140
rect 63217 342002 63283 342005
rect 50294 342000 63283 342002
rect 50294 341944 63222 342000
rect 63278 341944 63283 342000
rect 50294 341942 63283 341944
rect 44817 341866 44883 341869
rect 41462 341864 44883 341866
rect 41462 341808 44822 341864
rect 44878 341808 44883 341864
rect 41462 341806 44883 341808
rect 44817 341803 44883 341806
rect 45001 341866 45067 341869
rect 50294 341866 50354 341942
rect 63217 341939 63283 341942
rect 45001 341864 50354 341866
rect 45001 341808 45006 341864
rect 45062 341808 50354 341864
rect 45001 341806 50354 341808
rect 45001 341803 45067 341806
rect 35758 341700 35818 341803
rect 50470 341668 50476 341732
rect 50540 341730 50546 341732
rect 62665 341730 62731 341733
rect 50540 341728 62731 341730
rect 50540 341672 62670 341728
rect 62726 341672 62731 341728
rect 50540 341670 62731 341672
rect 50540 341668 50546 341670
rect 62665 341667 62731 341670
rect 33041 341458 33107 341461
rect 62297 341458 62363 341461
rect 33041 341456 62363 341458
rect 33041 341400 33046 341456
rect 33102 341400 62302 341456
rect 62358 341400 62363 341456
rect 33041 341398 62363 341400
rect 33041 341395 33107 341398
rect 62297 341395 62363 341398
rect 35758 341053 35818 341292
rect 35525 341050 35591 341053
rect 35525 341048 35634 341050
rect 35525 340992 35530 341048
rect 35586 340992 35634 341048
rect 35525 340987 35634 340992
rect 35758 341048 35867 341053
rect 35758 340992 35806 341048
rect 35862 340992 35867 341048
rect 35758 340990 35867 340992
rect 35801 340987 35867 340990
rect 44817 341050 44883 341053
rect 45737 341050 45803 341053
rect 44817 341048 45803 341050
rect 44817 340992 44822 341048
rect 44878 340992 45742 341048
rect 45798 340992 45803 341048
rect 44817 340990 45803 340992
rect 44817 340987 44883 340990
rect 45737 340987 45803 340990
rect 35574 340884 35634 340987
rect 40033 340642 40099 340645
rect 45369 340642 45435 340645
rect 40033 340640 45435 340642
rect 40033 340584 40038 340640
rect 40094 340584 45374 340640
rect 45430 340584 45435 340640
rect 40033 340582 45435 340584
rect 40033 340579 40099 340582
rect 45369 340579 45435 340582
rect 39806 340237 39866 340476
rect 39806 340232 39915 340237
rect 39806 340176 39854 340232
rect 39910 340176 39915 340232
rect 39806 340174 39915 340176
rect 39849 340171 39915 340174
rect 40217 340234 40283 340237
rect 46013 340234 46079 340237
rect 40217 340232 46079 340234
rect 40217 340176 40222 340232
rect 40278 340176 46018 340232
rect 46074 340176 46079 340232
rect 40217 340174 46079 340176
rect 40217 340171 40283 340174
rect 46013 340171 46079 340174
rect 675753 340234 675819 340237
rect 676254 340234 676260 340236
rect 675753 340232 676260 340234
rect 675753 340176 675758 340232
rect 675814 340176 676260 340232
rect 675753 340174 676260 340176
rect 675753 340171 675819 340174
rect 676254 340172 676260 340174
rect 676324 340172 676330 340236
rect 35574 339829 35634 340068
rect 35525 339824 35634 339829
rect 35801 339826 35867 339829
rect 35525 339768 35530 339824
rect 35586 339768 35634 339824
rect 35525 339766 35634 339768
rect 35758 339824 35867 339826
rect 35758 339768 35806 339824
rect 35862 339768 35867 339824
rect 35525 339763 35591 339766
rect 35758 339763 35867 339768
rect 39849 339826 39915 339829
rect 44214 339826 44220 339828
rect 39849 339824 44220 339826
rect 39849 339768 39854 339824
rect 39910 339768 44220 339824
rect 39849 339766 44220 339768
rect 39849 339763 39915 339766
rect 44214 339764 44220 339766
rect 44284 339764 44290 339828
rect 35758 339660 35818 339763
rect 675477 339420 675543 339421
rect 675477 339416 675524 339420
rect 675588 339418 675594 339420
rect 675477 339360 675482 339416
rect 675477 339356 675524 339360
rect 675588 339358 675634 339418
rect 675588 339356 675594 339358
rect 675477 339355 675543 339356
rect 44398 339282 44404 339284
rect 41492 339222 44404 339282
rect 44398 339220 44404 339222
rect 44468 339220 44474 339284
rect 35206 338605 35266 338844
rect 653581 338738 653647 338741
rect 675109 338738 675175 338741
rect 653581 338736 675175 338738
rect 653581 338680 653586 338736
rect 653642 338680 675114 338736
rect 675170 338680 675175 338736
rect 653581 338678 675175 338680
rect 653581 338675 653647 338678
rect 675109 338675 675175 338678
rect 35157 338600 35266 338605
rect 35157 338544 35162 338600
rect 35218 338544 35266 338600
rect 35157 338542 35266 338544
rect 35157 338539 35223 338542
rect 46565 338466 46631 338469
rect 41492 338464 46631 338466
rect 41492 338408 46570 338464
rect 46626 338408 46631 338464
rect 41492 338406 46631 338408
rect 46565 338403 46631 338406
rect 45369 338058 45435 338061
rect 41492 338056 45435 338058
rect 41492 338000 45374 338056
rect 45430 338000 45435 338056
rect 41492 337998 45435 338000
rect 45369 337995 45435 337998
rect 674281 338058 674347 338061
rect 675109 338058 675175 338061
rect 674281 338056 675175 338058
rect 674281 338000 674286 338056
rect 674342 338000 675114 338056
rect 675170 338000 675175 338056
rect 674281 337998 675175 338000
rect 674281 337995 674347 337998
rect 675109 337995 675175 337998
rect 675753 337922 675819 337925
rect 676070 337922 676076 337924
rect 675753 337920 676076 337922
rect 675753 337864 675758 337920
rect 675814 337864 676076 337920
rect 675753 337862 676076 337864
rect 675753 337859 675819 337862
rect 676070 337860 676076 337862
rect 676140 337860 676146 337924
rect 672165 337786 672231 337789
rect 675293 337786 675359 337789
rect 672165 337784 675359 337786
rect 672165 337728 672170 337784
rect 672226 337728 675298 337784
rect 675354 337728 675359 337784
rect 672165 337726 675359 337728
rect 672165 337723 672231 337726
rect 675293 337723 675359 337726
rect 46381 337650 46447 337653
rect 41492 337648 46447 337650
rect 41492 337592 46386 337648
rect 46442 337592 46447 337648
rect 41492 337590 46447 337592
rect 46381 337587 46447 337590
rect 40542 336972 40602 337212
rect 40534 336908 40540 336972
rect 40604 336908 40610 336972
rect 40726 336564 40786 336804
rect 40718 336500 40724 336564
rect 40788 336500 40794 336564
rect 675753 336562 675819 336565
rect 676438 336562 676444 336564
rect 675753 336560 676444 336562
rect 675753 336504 675758 336560
rect 675814 336504 676444 336560
rect 675753 336502 676444 336504
rect 675753 336499 675819 336502
rect 676438 336500 676444 336502
rect 676508 336500 676514 336564
rect 40910 336156 40970 336396
rect 40902 336092 40908 336156
rect 40972 336092 40978 336156
rect 35758 335749 35818 335988
rect 673361 335882 673427 335885
rect 674925 335882 674991 335885
rect 673361 335880 674991 335882
rect 673361 335824 673366 335880
rect 673422 335824 674930 335880
rect 674986 335824 674991 335880
rect 673361 335822 674991 335824
rect 673361 335819 673427 335822
rect 674925 335819 674991 335822
rect 35758 335744 35867 335749
rect 35758 335688 35806 335744
rect 35862 335688 35867 335744
rect 35758 335686 35867 335688
rect 35801 335683 35867 335686
rect 38929 335746 38995 335749
rect 42190 335746 42196 335748
rect 38929 335744 42196 335746
rect 38929 335688 38934 335744
rect 38990 335688 42196 335744
rect 38929 335686 42196 335688
rect 38929 335683 38995 335686
rect 42190 335684 42196 335686
rect 42260 335684 42266 335748
rect 672993 335610 673059 335613
rect 675109 335610 675175 335613
rect 672993 335608 675175 335610
rect 41462 335474 41522 335580
rect 672993 335552 672998 335608
rect 673054 335552 675114 335608
rect 675170 335552 675175 335608
rect 672993 335550 675175 335552
rect 672993 335547 673059 335550
rect 675109 335547 675175 335550
rect 44582 335474 44588 335476
rect 41462 335414 44588 335474
rect 44582 335412 44588 335414
rect 44652 335412 44658 335476
rect 35758 334933 35818 335172
rect 35758 334928 35867 334933
rect 35758 334872 35806 334928
rect 35862 334872 35867 334928
rect 35758 334870 35867 334872
rect 35801 334867 35867 334870
rect 41270 334868 41276 334932
rect 41340 334930 41346 334932
rect 41340 334870 44650 334930
rect 41340 334868 41346 334870
rect 41270 334460 41276 334524
rect 41340 334460 41346 334524
rect 41462 334522 41522 334764
rect 42057 334660 42123 334661
rect 42006 334658 42012 334660
rect 41966 334598 42012 334658
rect 42076 334656 42123 334660
rect 43805 334660 43871 334661
rect 43805 334658 43852 334660
rect 42118 334600 42123 334656
rect 42006 334596 42012 334598
rect 42076 334596 42123 334600
rect 43760 334656 43852 334658
rect 43760 334600 43810 334656
rect 43760 334598 43852 334600
rect 42057 334595 42123 334596
rect 43805 334596 43852 334598
rect 43916 334596 43922 334660
rect 44590 334658 44650 334870
rect 45093 334658 45159 334661
rect 44590 334656 45159 334658
rect 44590 334600 45098 334656
rect 45154 334600 45159 334656
rect 44590 334598 45159 334600
rect 43805 334595 43871 334596
rect 45093 334595 45159 334598
rect 43989 334524 44055 334525
rect 41462 334462 41890 334522
rect 41278 334356 41338 334460
rect 41830 334386 41890 334462
rect 43989 334520 44036 334524
rect 44100 334522 44106 334524
rect 43989 334464 43994 334520
rect 43989 334460 44036 334464
rect 44100 334462 44146 334522
rect 44100 334460 44106 334462
rect 43989 334459 44055 334460
rect 44357 334386 44423 334389
rect 44582 334386 44588 334388
rect 41830 334326 43178 334386
rect 43118 334250 43178 334326
rect 44357 334384 44588 334386
rect 44357 334328 44362 334384
rect 44418 334328 44588 334384
rect 44357 334326 44588 334328
rect 44357 334323 44423 334326
rect 44582 334324 44588 334326
rect 44652 334324 44658 334388
rect 44173 334250 44239 334253
rect 43118 334248 44239 334250
rect 43118 334192 44178 334248
rect 44234 334192 44239 334248
rect 43118 334190 44239 334192
rect 44173 334187 44239 334190
rect 40217 334114 40283 334117
rect 42977 334114 43043 334117
rect 40217 334112 43043 334114
rect 40217 334056 40222 334112
rect 40278 334056 42982 334112
rect 43038 334056 43043 334112
rect 40217 334054 43043 334056
rect 40217 334051 40283 334054
rect 42977 334051 43043 334054
rect 673729 333978 673795 333981
rect 675109 333978 675175 333981
rect 673729 333976 675175 333978
rect 41462 333298 41522 333948
rect 673729 333920 673734 333976
rect 673790 333920 675114 333976
rect 675170 333920 675175 333976
rect 673729 333918 675175 333920
rect 673729 333915 673795 333918
rect 675109 333915 675175 333918
rect 41462 333238 51090 333298
rect 37917 332890 37983 332893
rect 41822 332890 41828 332892
rect 37917 332888 41828 332890
rect 37917 332832 37922 332888
rect 37978 332832 41828 332888
rect 37917 332830 41828 332832
rect 37917 332827 37983 332830
rect 41822 332828 41828 332830
rect 41892 332828 41898 332892
rect 51030 332618 51090 333238
rect 673545 332754 673611 332757
rect 675109 332754 675175 332757
rect 673545 332752 675175 332754
rect 673545 332696 673550 332752
rect 673606 332696 675114 332752
rect 675170 332696 675175 332752
rect 673545 332694 675175 332696
rect 673545 332691 673611 332694
rect 675109 332691 675175 332694
rect 62481 332618 62547 332621
rect 51030 332616 62547 332618
rect 51030 332560 62486 332616
rect 62542 332560 62547 332616
rect 51030 332558 62547 332560
rect 62481 332555 62547 332558
rect 39757 332482 39823 332485
rect 42793 332482 42859 332485
rect 39757 332480 42859 332482
rect 39757 332424 39762 332480
rect 39818 332424 42798 332480
rect 42854 332424 42859 332480
rect 39757 332422 42859 332424
rect 39757 332419 39823 332422
rect 42793 332419 42859 332422
rect 35157 331802 35223 331805
rect 41638 331802 41644 331804
rect 35157 331800 41644 331802
rect 35157 331744 35162 331800
rect 35218 331744 41644 331800
rect 35157 331742 41644 331744
rect 35157 331739 35223 331742
rect 41638 331740 41644 331742
rect 41708 331740 41714 331804
rect 671705 331258 671771 331261
rect 675109 331258 675175 331261
rect 671705 331256 675175 331258
rect 671705 331200 671710 331256
rect 671766 331200 675114 331256
rect 675170 331200 675175 331256
rect 671705 331198 675175 331200
rect 671705 331195 671771 331198
rect 675109 331195 675175 331198
rect 652569 329762 652635 329765
rect 649950 329760 652635 329762
rect 649950 329704 652574 329760
rect 652630 329704 652635 329760
rect 649950 329702 652635 329704
rect 649950 329234 650010 329702
rect 652569 329699 652635 329702
rect 651465 328130 651531 328133
rect 649950 328128 651531 328130
rect 649950 328072 651470 328128
rect 651526 328072 651531 328128
rect 649950 328070 651531 328072
rect 649950 328052 650010 328070
rect 651465 328067 651531 328070
rect 675017 327994 675083 327997
rect 675385 327996 675451 327997
rect 675334 327994 675340 327996
rect 675017 327992 675340 327994
rect 675404 327994 675451 327996
rect 675404 327992 675496 327994
rect 675017 327936 675022 327992
rect 675078 327936 675340 327992
rect 675446 327936 675496 327992
rect 675017 327934 675340 327936
rect 675017 327931 675083 327934
rect 675334 327932 675340 327934
rect 675404 327934 675496 327936
rect 675404 327932 675451 327934
rect 675385 327931 675451 327932
rect 42057 327722 42123 327725
rect 62246 327722 62252 327724
rect 42057 327720 62252 327722
rect 42057 327664 42062 327720
rect 42118 327664 62252 327720
rect 42057 327662 62252 327664
rect 42057 327659 42123 327662
rect 62246 327660 62252 327662
rect 62316 327660 62322 327724
rect 42425 327042 42491 327045
rect 45277 327042 45343 327045
rect 42425 327040 45343 327042
rect 42425 326984 42430 327040
rect 42486 326984 45282 327040
rect 45338 326984 45343 327040
rect 42425 326982 45343 326984
rect 42425 326979 42491 326982
rect 45277 326979 45343 326982
rect 652201 326906 652267 326909
rect 650502 326904 652267 326906
rect 650502 326900 652206 326904
rect 649980 326848 652206 326900
rect 652262 326848 652267 326904
rect 649980 326846 652267 326848
rect 649980 326840 650562 326846
rect 652201 326843 652267 326846
rect 674649 326906 674715 326909
rect 675385 326906 675451 326909
rect 674649 326904 675451 326906
rect 674649 326848 674654 326904
rect 674710 326848 675390 326904
rect 675446 326848 675451 326904
rect 674649 326846 675451 326848
rect 674649 326843 674715 326846
rect 675385 326843 675451 326846
rect 649950 325682 650010 325710
rect 651741 325682 651807 325685
rect 649950 325680 651807 325682
rect 649950 325624 651746 325680
rect 651802 325624 651807 325680
rect 649950 325622 651807 325624
rect 651741 325619 651807 325622
rect 675201 325682 675267 325685
rect 676622 325682 676628 325684
rect 675201 325680 676628 325682
rect 675201 325624 675206 325680
rect 675262 325624 676628 325680
rect 675201 325622 676628 325624
rect 675201 325619 675267 325622
rect 676622 325620 676628 325622
rect 676692 325620 676698 325684
rect 672901 325002 672967 325005
rect 675017 325002 675083 325005
rect 672901 325000 675083 325002
rect 672901 324944 672906 325000
rect 672962 324944 675022 325000
rect 675078 324944 675083 325000
rect 672901 324942 675083 324944
rect 672901 324939 672967 324942
rect 675017 324939 675083 324942
rect 41781 324868 41847 324869
rect 41781 324864 41828 324868
rect 41892 324866 41898 324868
rect 41781 324808 41786 324864
rect 41781 324804 41828 324808
rect 41892 324806 41938 324866
rect 41892 324804 41898 324806
rect 41781 324803 41847 324804
rect 40902 322764 40908 322828
rect 40972 322826 40978 322828
rect 41781 322826 41847 322829
rect 40972 322824 41847 322826
rect 40972 322768 41786 322824
rect 41842 322768 41847 322824
rect 40972 322766 41847 322768
rect 40972 322764 40978 322766
rect 41781 322763 41847 322766
rect 42057 321602 42123 321605
rect 44173 321602 44239 321605
rect 42057 321600 44239 321602
rect 42057 321544 42062 321600
rect 42118 321544 44178 321600
rect 44234 321544 44239 321600
rect 42057 321542 44239 321544
rect 42057 321539 42123 321542
rect 44173 321539 44239 321542
rect 42057 321194 42123 321197
rect 42977 321194 43043 321197
rect 42057 321192 43043 321194
rect 42057 321136 42062 321192
rect 42118 321136 42982 321192
rect 43038 321136 43043 321192
rect 42057 321134 43043 321136
rect 42057 321131 42123 321134
rect 42977 321131 43043 321134
rect 42425 320786 42491 320789
rect 53833 320786 53899 320789
rect 42425 320784 53899 320786
rect 42425 320728 42430 320784
rect 42486 320728 53838 320784
rect 53894 320728 53899 320784
rect 42425 320726 53899 320728
rect 42425 320723 42491 320726
rect 53833 320723 53899 320726
rect 42609 319426 42675 319429
rect 61561 319426 61627 319429
rect 42609 319424 61627 319426
rect 42609 319368 42614 319424
rect 42670 319368 61566 319424
rect 61622 319368 61627 319424
rect 42609 319366 61627 319368
rect 42609 319363 42675 319366
rect 61561 319363 61627 319366
rect 42425 319018 42491 319021
rect 46565 319018 46631 319021
rect 42425 319016 46631 319018
rect 42425 318960 42430 319016
rect 42486 318960 46570 319016
rect 46626 318960 46631 319016
rect 42425 318958 46631 318960
rect 42425 318955 42491 318958
rect 46565 318955 46631 318958
rect 40718 317460 40724 317524
rect 40788 317522 40794 317524
rect 42241 317522 42307 317525
rect 40788 317520 42307 317522
rect 40788 317464 42246 317520
rect 42302 317464 42307 317520
rect 40788 317462 42307 317464
rect 40788 317460 40794 317462
rect 42241 317459 42307 317462
rect 62113 317386 62179 317389
rect 62113 317384 64706 317386
rect 62113 317328 62118 317384
rect 62174 317328 64706 317384
rect 62113 317326 64706 317328
rect 62113 317323 62179 317326
rect 42057 317250 42123 317253
rect 44357 317250 44423 317253
rect 42057 317248 44423 317250
rect 42057 317192 42062 317248
rect 42118 317192 44362 317248
rect 44418 317192 44423 317248
rect 42057 317190 44423 317192
rect 42057 317187 42123 317190
rect 44357 317187 44423 317190
rect 64646 317106 64706 317326
rect 40534 315964 40540 316028
rect 40604 316026 40610 316028
rect 41781 316026 41847 316029
rect 40604 316024 41847 316026
rect 40604 315968 41786 316024
rect 41842 315968 41847 316024
rect 40604 315966 41847 315968
rect 40604 315964 40610 315966
rect 41781 315963 41847 315966
rect 61561 316026 61627 316029
rect 61561 316024 64706 316026
rect 61561 315968 61566 316024
rect 61622 315968 64706 316024
rect 61561 315966 64706 315968
rect 61561 315963 61627 315966
rect 64646 315924 64706 315966
rect 41781 315620 41847 315621
rect 41781 315616 41828 315620
rect 41892 315618 41898 315620
rect 41781 315560 41786 315616
rect 41781 315556 41828 315560
rect 41892 315558 41938 315618
rect 41892 315556 41898 315558
rect 41781 315555 41847 315556
rect 62113 314802 62179 314805
rect 62113 314800 64706 314802
rect 62113 314744 62118 314800
rect 62174 314744 64706 314800
rect 62113 314742 64706 314744
rect 62113 314739 62179 314742
rect 62389 314122 62455 314125
rect 62389 314120 64706 314122
rect 62389 314064 62394 314120
rect 62450 314064 64706 314120
rect 62389 314062 64706 314064
rect 62389 314059 62455 314062
rect 42149 313716 42215 313717
rect 42149 313714 42196 313716
rect 42104 313712 42196 313714
rect 42104 313656 42154 313712
rect 42104 313654 42196 313656
rect 42149 313652 42196 313654
rect 42260 313652 42266 313716
rect 42149 313651 42215 313652
rect 64646 313560 64706 314062
rect 676213 313986 676279 313989
rect 676213 313984 676322 313986
rect 676213 313928 676218 313984
rect 676274 313928 676322 313984
rect 676213 313923 676322 313928
rect 676262 313684 676322 313923
rect 653397 313306 653463 313309
rect 653397 313304 676292 313306
rect 653397 313248 653402 313304
rect 653458 313248 676292 313304
rect 653397 313246 676292 313248
rect 653397 313243 653463 313246
rect 42425 313170 42491 313173
rect 46381 313170 46447 313173
rect 42425 313168 46447 313170
rect 42425 313112 42430 313168
rect 42486 313112 46386 313168
rect 46442 313112 46447 313168
rect 42425 313110 46447 313112
rect 42425 313107 42491 313110
rect 46381 313107 46447 313110
rect 63217 313034 63283 313037
rect 63217 313032 64706 313034
rect 63217 312976 63222 313032
rect 63278 312976 64706 313032
rect 63217 312974 64706 312976
rect 63217 312971 63283 312974
rect 42241 312490 42307 312493
rect 53833 312490 53899 312493
rect 42241 312488 53899 312490
rect 42241 312432 42246 312488
rect 42302 312432 53838 312488
rect 53894 312432 53899 312488
rect 42241 312430 53899 312432
rect 42241 312427 42307 312430
rect 53833 312427 53899 312430
rect 64646 312378 64706 312974
rect 674833 312898 674899 312901
rect 674833 312896 676292 312898
rect 674833 312840 674838 312896
rect 674894 312840 676292 312896
rect 674833 312838 676292 312840
rect 674833 312835 674899 312838
rect 672349 312490 672415 312493
rect 672349 312488 676292 312490
rect 672349 312432 672354 312488
rect 672410 312432 676292 312488
rect 672349 312430 676292 312432
rect 672349 312427 672415 312430
rect 675477 312082 675543 312085
rect 675477 312080 676292 312082
rect 675477 312024 675482 312080
rect 675538 312024 676292 312080
rect 675477 312022 676292 312024
rect 675477 312019 675543 312022
rect 42057 311946 42123 311949
rect 44398 311946 44404 311948
rect 42057 311944 44404 311946
rect 42057 311888 42062 311944
rect 42118 311888 44404 311944
rect 42057 311886 44404 311888
rect 42057 311883 42123 311886
rect 44398 311884 44404 311886
rect 44468 311884 44474 311948
rect 658917 311946 658983 311949
rect 674833 311946 674899 311949
rect 658917 311944 674899 311946
rect 658917 311888 658922 311944
rect 658978 311888 674838 311944
rect 674894 311888 674899 311944
rect 658917 311886 674899 311888
rect 658917 311883 658983 311886
rect 674833 311883 674899 311886
rect 62757 311810 62823 311813
rect 62757 311808 64706 311810
rect 62757 311752 62762 311808
rect 62818 311752 64706 311808
rect 62757 311750 64706 311752
rect 62757 311747 62823 311750
rect 44265 311268 44331 311269
rect 44214 311266 44220 311268
rect 44174 311206 44220 311266
rect 44284 311264 44331 311268
rect 44326 311208 44331 311264
rect 44214 311204 44220 311206
rect 44284 311204 44331 311208
rect 44265 311203 44331 311204
rect 64646 311196 64706 311750
rect 672533 311674 672599 311677
rect 672533 311672 676292 311674
rect 672533 311616 672538 311672
rect 672594 311616 676292 311672
rect 672533 311614 676292 311616
rect 672533 311611 672599 311614
rect 674741 311266 674807 311269
rect 674741 311264 676292 311266
rect 674741 311208 674746 311264
rect 674802 311208 676292 311264
rect 674741 311206 676292 311208
rect 674741 311203 674807 311206
rect 673177 310858 673243 310861
rect 673177 310856 676292 310858
rect 673177 310800 673182 310856
rect 673238 310800 676292 310856
rect 673177 310798 676292 310800
rect 673177 310795 673243 310798
rect 674557 310450 674623 310453
rect 674557 310448 676292 310450
rect 674557 310392 674562 310448
rect 674618 310392 676292 310448
rect 674557 310390 676292 310392
rect 674557 310387 674623 310390
rect 673913 310042 673979 310045
rect 673913 310040 676292 310042
rect 673913 309984 673918 310040
rect 673974 309984 676292 310040
rect 673913 309982 676292 309984
rect 673913 309979 673979 309982
rect 652477 309906 652543 309909
rect 652477 309904 663810 309906
rect 652477 309848 652482 309904
rect 652538 309848 663810 309904
rect 652477 309846 663810 309848
rect 652477 309843 652543 309846
rect 663750 309770 663810 309846
rect 675937 309770 676003 309773
rect 663750 309768 676003 309770
rect 663750 309712 675942 309768
rect 675998 309712 676003 309768
rect 663750 309710 676003 309712
rect 675937 309707 676003 309710
rect 676170 309574 676292 309634
rect 673269 309498 673335 309501
rect 676170 309498 676230 309574
rect 673269 309496 676230 309498
rect 673269 309440 673274 309496
rect 673330 309440 676230 309496
rect 673269 309438 676230 309440
rect 673269 309435 673335 309438
rect 675334 309164 675340 309228
rect 675404 309226 675410 309228
rect 675404 309166 676292 309226
rect 675404 309164 675410 309166
rect 675886 308756 675892 308820
rect 675956 308818 675962 308820
rect 675956 308758 676292 308818
rect 675956 308756 675962 308758
rect 675109 308410 675175 308413
rect 675109 308408 676292 308410
rect 675109 308352 675114 308408
rect 675170 308352 676292 308408
rect 675109 308350 676292 308352
rect 675109 308347 675175 308350
rect 675293 308002 675359 308005
rect 675293 308000 676292 308002
rect 675293 307944 675298 308000
rect 675354 307944 676292 308000
rect 675293 307942 676292 307944
rect 675293 307939 675359 307942
rect 676029 307594 676095 307597
rect 676029 307592 676292 307594
rect 676029 307536 676034 307592
rect 676090 307536 676292 307592
rect 676029 307534 676292 307536
rect 676029 307531 676095 307534
rect 676029 307186 676095 307189
rect 676029 307184 676292 307186
rect 676029 307128 676034 307184
rect 676090 307128 676292 307184
rect 676029 307126 676292 307128
rect 676029 307123 676095 307126
rect 678237 306778 678303 306781
rect 678237 306776 678316 306778
rect 678237 306720 678242 306776
rect 678298 306720 678316 306776
rect 678237 306718 678316 306720
rect 678237 306715 678303 306718
rect 674925 306370 674991 306373
rect 674925 306368 676292 306370
rect 674925 306312 674930 306368
rect 674986 306312 676292 306368
rect 674925 306310 676292 306312
rect 674925 306307 674991 306310
rect 673821 305962 673887 305965
rect 673821 305960 676292 305962
rect 673821 305904 673826 305960
rect 673882 305904 676292 305960
rect 673821 305902 676292 305904
rect 673821 305899 673887 305902
rect 672533 305554 672599 305557
rect 672533 305552 676292 305554
rect 672533 305496 672538 305552
rect 672594 305496 676292 305552
rect 672533 305494 676292 305496
rect 672533 305491 672599 305494
rect 675894 305086 676292 305146
rect 675894 304602 675954 305086
rect 676581 304738 676647 304741
rect 676581 304736 676660 304738
rect 676581 304680 676586 304736
rect 676642 304680 676660 304736
rect 676581 304678 676660 304680
rect 676581 304675 676647 304678
rect 676070 304602 676076 304604
rect 675894 304542 676076 304602
rect 676070 304540 676076 304542
rect 676140 304540 676146 304604
rect 673085 304330 673151 304333
rect 673085 304328 676292 304330
rect 673085 304272 673090 304328
rect 673146 304272 676292 304328
rect 673085 304270 676292 304272
rect 673085 304267 673151 304270
rect 674373 303922 674439 303925
rect 674373 303920 676292 303922
rect 674373 303864 674378 303920
rect 674434 303864 676292 303920
rect 674373 303862 676292 303864
rect 674373 303859 674439 303862
rect 676029 303514 676095 303517
rect 676029 303512 676292 303514
rect 676029 303456 676034 303512
rect 676090 303456 676292 303512
rect 676029 303454 676292 303456
rect 676029 303451 676095 303454
rect 651373 303378 651439 303381
rect 649950 303376 651439 303378
rect 649950 303320 651378 303376
rect 651434 303320 651439 303376
rect 649950 303318 651439 303320
rect 649950 302776 650010 303318
rect 651373 303315 651439 303318
rect 675886 302636 675892 302700
rect 675956 302698 675962 302700
rect 676262 302698 676322 303076
rect 675956 302668 676322 302698
rect 675956 302638 676292 302668
rect 675956 302636 675962 302638
rect 671521 302290 671587 302293
rect 671521 302288 676292 302290
rect 671521 302232 671526 302288
rect 671582 302232 676292 302288
rect 671521 302230 676292 302232
rect 671521 302227 671587 302230
rect 652477 302154 652543 302157
rect 649950 302152 652543 302154
rect 649950 302096 652482 302152
rect 652538 302096 652543 302152
rect 649950 302094 652543 302096
rect 649950 301594 650010 302094
rect 652477 302091 652543 302094
rect 669865 302018 669931 302021
rect 676029 302018 676095 302021
rect 669865 302016 676095 302018
rect 669865 301960 669870 302016
rect 669926 301960 676034 302016
rect 676090 301960 676095 302016
rect 669865 301958 676095 301960
rect 669865 301955 669931 301958
rect 676029 301955 676095 301958
rect 676581 301612 676647 301613
rect 676581 301608 676628 301612
rect 676692 301610 676698 301612
rect 676581 301552 676586 301608
rect 676581 301548 676628 301552
rect 676692 301550 676738 301610
rect 676692 301548 676698 301550
rect 676581 301547 676647 301548
rect 51717 301338 51783 301341
rect 41492 301336 51783 301338
rect 41492 301280 51722 301336
rect 51778 301280 51783 301336
rect 41492 301278 51783 301280
rect 51717 301275 51783 301278
rect 41137 300930 41203 300933
rect 41124 300928 41203 300930
rect 41124 300872 41142 300928
rect 41198 300872 41203 300928
rect 41124 300870 41203 300872
rect 41137 300867 41203 300870
rect 651465 300658 651531 300661
rect 649950 300656 651531 300658
rect 649950 300600 651470 300656
rect 651526 300600 651531 300656
rect 649950 300598 651531 300600
rect 54477 300522 54543 300525
rect 41492 300520 54543 300522
rect 41492 300464 54482 300520
rect 54538 300464 54543 300520
rect 41492 300462 54543 300464
rect 54477 300459 54543 300462
rect 649950 300412 650010 300598
rect 651465 300595 651531 300598
rect 45553 300114 45619 300117
rect 41492 300112 45619 300114
rect 41492 300056 45558 300112
rect 45614 300056 45619 300112
rect 41492 300054 45619 300056
rect 45553 300051 45619 300054
rect 44633 299706 44699 299709
rect 41492 299704 44699 299706
rect 41492 299648 44638 299704
rect 44694 299648 44699 299704
rect 41492 299646 44699 299648
rect 44633 299643 44699 299646
rect 45737 299298 45803 299301
rect 41492 299296 45803 299298
rect 41492 299240 45742 299296
rect 45798 299240 45803 299296
rect 41492 299238 45803 299240
rect 45737 299235 45803 299238
rect 42793 299026 42859 299029
rect 41784 299024 42859 299026
rect 41784 298968 42798 299024
rect 42854 298968 42859 299024
rect 41784 298966 42859 298968
rect 41784 298890 41844 298966
rect 42793 298963 42859 298966
rect 41492 298830 41844 298890
rect 41965 298754 42031 298757
rect 63125 298754 63191 298757
rect 41965 298752 63191 298754
rect 41965 298696 41970 298752
rect 42026 298696 63130 298752
rect 63186 298696 63191 298752
rect 41965 298694 63191 298696
rect 649950 298754 650010 299230
rect 651465 298754 651531 298757
rect 649950 298752 651531 298754
rect 649950 298696 651470 298752
rect 651526 298696 651531 298752
rect 649950 298694 651531 298696
rect 41965 298691 42031 298694
rect 63125 298691 63191 298694
rect 651465 298691 651531 298694
rect 46013 298482 46079 298485
rect 41492 298480 46079 298482
rect 41492 298424 46018 298480
rect 46074 298424 46079 298480
rect 41492 298422 46079 298424
rect 46013 298419 46079 298422
rect 675150 298148 675156 298212
rect 675220 298210 675226 298212
rect 675477 298210 675543 298213
rect 675220 298208 675543 298210
rect 675220 298152 675482 298208
rect 675538 298152 675543 298208
rect 675220 298150 675543 298152
rect 675220 298148 675226 298150
rect 675477 298147 675543 298150
rect 44265 298074 44331 298077
rect 41492 298072 44331 298074
rect 41492 298016 44270 298072
rect 44326 298016 44331 298072
rect 41492 298014 44331 298016
rect 44265 298011 44331 298014
rect 44449 297666 44515 297669
rect 41492 297664 44515 297666
rect 41492 297608 44454 297664
rect 44510 297608 44515 297664
rect 41492 297606 44515 297608
rect 44449 297603 44515 297606
rect 649950 297530 650010 298048
rect 675017 297666 675083 297669
rect 675518 297666 675524 297668
rect 675017 297664 675524 297666
rect 675017 297608 675022 297664
rect 675078 297608 675524 297664
rect 675017 297606 675524 297608
rect 675017 297603 675083 297606
rect 675518 297604 675524 297606
rect 675588 297604 675594 297668
rect 652293 297530 652359 297533
rect 649950 297528 652359 297530
rect 649950 297472 652298 297528
rect 652354 297472 652359 297528
rect 649950 297470 652359 297472
rect 652293 297467 652359 297470
rect 675702 297332 675708 297396
rect 675772 297394 675778 297396
rect 676857 297394 676923 297397
rect 675772 297392 676923 297394
rect 675772 297336 676862 297392
rect 676918 297336 676923 297392
rect 675772 297334 676923 297336
rect 675772 297332 675778 297334
rect 676857 297331 676923 297334
rect 43161 297258 43227 297261
rect 41492 297256 43227 297258
rect 41492 297200 43166 297256
rect 43222 297200 43227 297256
rect 41492 297198 43227 297200
rect 43161 297195 43227 297198
rect 46933 296850 46999 296853
rect 41492 296848 46999 296850
rect 41492 296792 46938 296848
rect 46994 296792 46999 296848
rect 41492 296790 46999 296792
rect 649950 296850 650010 296866
rect 651649 296850 651715 296853
rect 649950 296848 651715 296850
rect 649950 296792 651654 296848
rect 651710 296792 651715 296848
rect 649950 296790 651715 296792
rect 46933 296787 46999 296790
rect 651649 296787 651715 296790
rect 41321 296442 41387 296445
rect 41308 296440 41387 296442
rect 41308 296384 41326 296440
rect 41382 296384 41387 296440
rect 41308 296382 41387 296384
rect 41321 296379 41387 296382
rect 39297 296034 39363 296037
rect 39284 296032 39363 296034
rect 39284 295976 39302 296032
rect 39358 295976 39363 296032
rect 39284 295974 39363 295976
rect 39297 295971 39363 295974
rect 670969 295898 671035 295901
rect 675385 295898 675451 295901
rect 670969 295896 675451 295898
rect 670969 295840 670974 295896
rect 671030 295840 675390 295896
rect 675446 295840 675451 295896
rect 670969 295838 675451 295840
rect 670969 295835 671035 295838
rect 675385 295835 675451 295838
rect 675569 295764 675635 295765
rect 675518 295700 675524 295764
rect 675588 295762 675635 295764
rect 675588 295760 675680 295762
rect 675630 295704 675680 295760
rect 675588 295702 675680 295704
rect 675588 295700 675635 295702
rect 675569 295699 675635 295700
rect 41822 295626 41828 295628
rect 41492 295566 41828 295626
rect 41822 295564 41828 295566
rect 41892 295564 41898 295628
rect 62297 295354 62363 295357
rect 64646 295354 64706 295684
rect 62297 295352 64706 295354
rect 62297 295296 62302 295352
rect 62358 295296 64706 295352
rect 62297 295294 64706 295296
rect 649950 295354 650010 295684
rect 651925 295354 651991 295357
rect 649950 295352 651991 295354
rect 649950 295296 651930 295352
rect 651986 295296 651991 295352
rect 649950 295294 651991 295296
rect 62297 295291 62363 295294
rect 651925 295291 651991 295294
rect 42333 295218 42399 295221
rect 41492 295216 42399 295218
rect 41492 295160 42338 295216
rect 42394 295160 42399 295216
rect 41492 295158 42399 295160
rect 42333 295155 42399 295158
rect 33041 294810 33107 294813
rect 33028 294808 33107 294810
rect 33028 294752 33046 294808
rect 33102 294752 33107 294808
rect 33028 294750 33107 294752
rect 33041 294747 33107 294750
rect 675753 294674 675819 294677
rect 676438 294674 676444 294676
rect 675753 294672 676444 294674
rect 675753 294616 675758 294672
rect 675814 294616 676444 294672
rect 675753 294614 676444 294616
rect 675753 294611 675819 294614
rect 676438 294612 676444 294614
rect 676508 294612 676514 294676
rect 33777 294402 33843 294405
rect 33764 294400 33843 294402
rect 33764 294344 33782 294400
rect 33838 294344 33843 294400
rect 33764 294342 33843 294344
rect 33777 294339 33843 294342
rect 62113 294130 62179 294133
rect 64646 294130 64706 294502
rect 649950 294266 650010 294502
rect 651465 294266 651531 294269
rect 649950 294264 651531 294266
rect 649950 294208 651470 294264
rect 651526 294208 651531 294264
rect 649950 294206 651531 294208
rect 651465 294203 651531 294206
rect 62113 294128 64706 294130
rect 62113 294072 62118 294128
rect 62174 294072 64706 294128
rect 62113 294070 64706 294072
rect 62113 294067 62179 294070
rect 41781 293994 41847 293997
rect 41492 293992 41847 293994
rect 41492 293936 41786 293992
rect 41842 293936 41847 293992
rect 41492 293934 41847 293936
rect 41781 293931 41847 293934
rect 660573 293858 660639 293861
rect 670969 293858 671035 293861
rect 660573 293856 671035 293858
rect 660573 293800 660578 293856
rect 660634 293800 670974 293856
rect 671030 293800 671035 293856
rect 660573 293798 671035 293800
rect 660573 293795 660639 293798
rect 670969 293795 671035 293798
rect 42977 293586 43043 293589
rect 41492 293584 43043 293586
rect 41492 293528 42982 293584
rect 43038 293528 43043 293584
rect 41492 293526 43043 293528
rect 42977 293523 43043 293526
rect 44449 293178 44515 293181
rect 41492 293176 44515 293178
rect 41492 293120 44454 293176
rect 44510 293120 44515 293176
rect 41492 293118 44515 293120
rect 44449 293115 44515 293118
rect 45277 292770 45343 292773
rect 41492 292768 45343 292770
rect 41492 292712 45282 292768
rect 45338 292712 45343 292768
rect 41492 292710 45343 292712
rect 45277 292707 45343 292710
rect 62757 292770 62823 292773
rect 64646 292770 64706 293320
rect 649950 293042 650010 293320
rect 651465 293042 651531 293045
rect 649950 293040 651531 293042
rect 649950 292984 651470 293040
rect 651526 292984 651531 293040
rect 649950 292982 651531 292984
rect 651465 292979 651531 292982
rect 62757 292768 64706 292770
rect 62757 292712 62762 292768
rect 62818 292712 64706 292768
rect 62757 292710 64706 292712
rect 62757 292707 62823 292710
rect 40585 292592 40651 292593
rect 40534 292590 40540 292592
rect 40494 292530 40540 292590
rect 40604 292588 40651 292592
rect 40646 292532 40651 292588
rect 40534 292528 40540 292530
rect 40604 292528 40651 292532
rect 41362 292528 41368 292592
rect 41432 292528 41438 292592
rect 40585 292527 40651 292528
rect 41370 292362 41430 292528
rect 62113 292498 62179 292501
rect 674833 292498 674899 292501
rect 675150 292498 675156 292500
rect 62113 292496 64706 292498
rect 62113 292440 62118 292496
rect 62174 292440 64706 292496
rect 62113 292438 64706 292440
rect 62113 292435 62179 292438
rect 41370 292302 41492 292362
rect 64646 292138 64706 292438
rect 674833 292496 675156 292498
rect 674833 292440 674838 292496
rect 674894 292440 675156 292496
rect 674833 292438 675156 292440
rect 674833 292435 674899 292438
rect 675150 292436 675156 292438
rect 675220 292436 675226 292500
rect 35801 291954 35867 291957
rect 35788 291952 35867 291954
rect 35788 291896 35806 291952
rect 35862 291896 35867 291952
rect 35788 291894 35867 291896
rect 35801 291891 35867 291894
rect 45461 291546 45527 291549
rect 41492 291544 45527 291546
rect 41492 291488 45466 291544
rect 45522 291488 45527 291544
rect 41492 291486 45527 291488
rect 649950 291546 650010 292138
rect 651925 291818 651991 291821
rect 674005 291818 674071 291821
rect 651925 291816 674071 291818
rect 651925 291760 651930 291816
rect 651986 291760 674010 291816
rect 674066 291760 674071 291816
rect 651925 291758 674071 291760
rect 651925 291755 651991 291758
rect 674005 291755 674071 291758
rect 652109 291546 652175 291549
rect 649950 291544 652175 291546
rect 649950 291488 652114 291544
rect 652170 291488 652175 291544
rect 649950 291486 652175 291488
rect 45461 291483 45527 291486
rect 652109 291483 652175 291486
rect 673821 291546 673887 291549
rect 675385 291546 675451 291549
rect 673821 291544 675451 291546
rect 673821 291488 673826 291544
rect 673882 291488 675390 291544
rect 675446 291488 675451 291544
rect 673821 291486 675451 291488
rect 673821 291483 673887 291486
rect 675385 291483 675451 291486
rect 49141 291138 49207 291141
rect 41492 291136 49207 291138
rect 41492 291080 49146 291136
rect 49202 291080 49207 291136
rect 41492 291078 49207 291080
rect 49141 291075 49207 291078
rect 62113 291002 62179 291005
rect 675753 291002 675819 291005
rect 676622 291002 676628 291004
rect 62113 291000 64154 291002
rect 62113 290944 62118 291000
rect 62174 290986 64154 291000
rect 675753 291000 676628 291002
rect 62174 290944 64676 290986
rect 62113 290942 64676 290944
rect 62113 290939 62179 290942
rect 64094 290926 64676 290942
rect 47577 290730 47643 290733
rect 41492 290728 47643 290730
rect 41492 290672 47582 290728
rect 47638 290672 47643 290728
rect 41492 290670 47643 290672
rect 47577 290667 47643 290670
rect 41781 290458 41847 290461
rect 43345 290458 43411 290461
rect 41781 290456 43411 290458
rect 41781 290400 41786 290456
rect 41842 290400 43350 290456
rect 43406 290400 43411 290456
rect 41781 290398 43411 290400
rect 649950 290458 650010 290956
rect 675753 290944 675758 291000
rect 675814 290944 676628 291000
rect 675753 290942 676628 290944
rect 675753 290939 675819 290942
rect 676622 290940 676628 290942
rect 676692 290940 676698 291004
rect 651465 290458 651531 290461
rect 649950 290456 651531 290458
rect 649950 290400 651470 290456
rect 651526 290400 651531 290456
rect 649950 290398 651531 290400
rect 41781 290395 41847 290398
rect 43345 290395 43411 290398
rect 651465 290395 651531 290398
rect 35157 290322 35223 290325
rect 35157 290320 35236 290322
rect 35157 290264 35162 290320
rect 35218 290264 35236 290320
rect 35157 290262 35236 290264
rect 35157 290259 35223 290262
rect 63125 289778 63191 289781
rect 63125 289776 64706 289778
rect 63125 289720 63130 289776
rect 63186 289720 64706 289776
rect 63125 289718 64706 289720
rect 63125 289715 63191 289718
rect 649950 289234 650010 289774
rect 651649 289234 651715 289237
rect 649950 289232 651715 289234
rect 649950 289176 651654 289232
rect 651710 289176 651715 289232
rect 649950 289174 651715 289176
rect 651649 289171 651715 289174
rect 651465 288690 651531 288693
rect 649950 288688 651531 288690
rect 649950 288632 651470 288688
rect 651526 288632 651531 288688
rect 649950 288630 651531 288632
rect 649950 288592 650010 288630
rect 651465 288627 651531 288630
rect 62113 288554 62179 288557
rect 64646 288554 64706 288592
rect 62113 288552 64706 288554
rect 62113 288496 62118 288552
rect 62174 288496 64706 288552
rect 62113 288494 64706 288496
rect 62113 288491 62179 288494
rect 673085 287874 673151 287877
rect 675109 287874 675175 287877
rect 673085 287872 675175 287874
rect 673085 287816 673090 287872
rect 673146 287816 675114 287872
rect 675170 287816 675175 287872
rect 673085 287814 675175 287816
rect 673085 287811 673151 287814
rect 675109 287811 675175 287814
rect 651649 287738 651715 287741
rect 651649 287736 663810 287738
rect 651649 287680 651654 287736
rect 651710 287680 663810 287736
rect 651649 287678 663810 287680
rect 651649 287675 651715 287678
rect 663750 287602 663810 287678
rect 673453 287602 673519 287605
rect 663750 287600 673519 287602
rect 663750 287544 673458 287600
rect 673514 287544 673519 287600
rect 663750 287542 673519 287544
rect 673453 287539 673519 287542
rect 651465 287466 651531 287469
rect 649766 287464 651531 287466
rect 62757 287194 62823 287197
rect 64646 287194 64706 287410
rect 649766 287408 651470 287464
rect 651526 287408 651531 287464
rect 649766 287406 651531 287408
rect 651465 287403 651531 287406
rect 62757 287192 64706 287194
rect 62757 287136 62762 287192
rect 62818 287136 64706 287192
rect 62757 287134 64706 287136
rect 62757 287131 62823 287134
rect 675753 287058 675819 287061
rect 676254 287058 676260 287060
rect 675753 287056 676260 287058
rect 675753 287000 675758 287056
rect 675814 287000 676260 287056
rect 675753 286998 676260 287000
rect 675753 286995 675819 286998
rect 676254 286996 676260 286998
rect 676324 286996 676330 287060
rect 62113 285970 62179 285973
rect 64646 285970 64706 286228
rect 62113 285968 64706 285970
rect 62113 285912 62118 285968
rect 62174 285912 64706 285968
rect 62113 285910 64706 285912
rect 649950 285970 650010 286228
rect 651465 285970 651531 285973
rect 649950 285968 651531 285970
rect 649950 285912 651470 285968
rect 651526 285912 651531 285968
rect 649950 285910 651531 285912
rect 62113 285907 62179 285910
rect 651465 285907 651531 285910
rect 672533 285562 672599 285565
rect 675109 285562 675175 285565
rect 672533 285560 675175 285562
rect 672533 285504 672538 285560
rect 672594 285504 675114 285560
rect 675170 285504 675175 285560
rect 672533 285502 675175 285504
rect 672533 285499 672599 285502
rect 675109 285499 675175 285502
rect 33777 284882 33843 284885
rect 41822 284882 41828 284884
rect 33777 284880 41828 284882
rect 33777 284824 33782 284880
rect 33838 284824 41828 284880
rect 33777 284822 41828 284824
rect 33777 284819 33843 284822
rect 41822 284820 41828 284822
rect 41892 284820 41898 284884
rect 62941 284610 63007 284613
rect 64646 284610 64706 285046
rect 649950 284746 650010 285046
rect 651465 284746 651531 284749
rect 649950 284744 651531 284746
rect 649950 284688 651470 284744
rect 651526 284688 651531 284744
rect 649950 284686 651531 284688
rect 651465 284683 651531 284686
rect 62941 284608 64706 284610
rect 62941 284552 62946 284608
rect 63002 284552 64706 284608
rect 62941 284550 64706 284552
rect 62941 284547 63007 284550
rect 39297 284338 39363 284341
rect 42006 284338 42012 284340
rect 39297 284336 42012 284338
rect 39297 284280 39302 284336
rect 39358 284280 42012 284336
rect 39297 284278 42012 284280
rect 39297 284275 39363 284278
rect 42006 284276 42012 284278
rect 42076 284276 42082 284340
rect 44817 284338 44883 284341
rect 45553 284338 45619 284341
rect 44817 284336 45619 284338
rect 44817 284280 44822 284336
rect 44878 284280 45558 284336
rect 45614 284280 45619 284336
rect 44817 284278 45619 284280
rect 44817 284275 44883 284278
rect 45553 284275 45619 284278
rect 63125 283250 63191 283253
rect 64646 283250 64706 283864
rect 649950 283386 650010 283864
rect 675753 283658 675819 283661
rect 676070 283658 676076 283660
rect 675753 283656 676076 283658
rect 675753 283600 675758 283656
rect 675814 283600 676076 283656
rect 675753 283598 676076 283600
rect 675753 283595 675819 283598
rect 676070 283596 676076 283598
rect 676140 283596 676146 283660
rect 651465 283386 651531 283389
rect 649950 283384 651531 283386
rect 649950 283328 651470 283384
rect 651526 283328 651531 283384
rect 649950 283326 651531 283328
rect 651465 283323 651531 283326
rect 63125 283248 64706 283250
rect 63125 283192 63130 283248
rect 63186 283192 64706 283248
rect 63125 283190 64706 283192
rect 63125 283187 63191 283190
rect 675753 282706 675819 282709
rect 676070 282706 676076 282708
rect 675753 282704 676076 282706
rect 62481 282162 62547 282165
rect 64646 282162 64706 282682
rect 62481 282160 64706 282162
rect 62481 282104 62486 282160
rect 62542 282104 64706 282160
rect 62481 282102 64706 282104
rect 649950 282162 650010 282682
rect 675753 282648 675758 282704
rect 675814 282648 676076 282704
rect 675753 282646 676076 282648
rect 675753 282643 675819 282646
rect 676070 282644 676076 282646
rect 676140 282644 676146 282708
rect 652017 282162 652083 282165
rect 649950 282160 652083 282162
rect 649950 282104 652022 282160
rect 652078 282104 652083 282160
rect 649950 282102 652083 282104
rect 62481 282099 62547 282102
rect 652017 282099 652083 282102
rect 675661 281620 675727 281621
rect 675661 281616 675708 281620
rect 675772 281618 675778 281620
rect 675661 281560 675666 281616
rect 675661 281556 675708 281560
rect 675772 281558 675818 281618
rect 675772 281556 675778 281558
rect 675661 281555 675727 281556
rect 62297 280938 62363 280941
rect 64646 280938 64706 281500
rect 62297 280936 64706 280938
rect 62297 280880 62302 280936
rect 62358 280880 64706 280936
rect 62297 280878 64706 280880
rect 649950 280938 650010 281500
rect 651465 280938 651531 280941
rect 649950 280936 651531 280938
rect 649950 280880 651470 280936
rect 651526 280880 651531 280936
rect 649950 280878 651531 280880
rect 62297 280875 62363 280878
rect 651465 280875 651531 280878
rect 62113 280394 62179 280397
rect 652385 280394 652451 280397
rect 62113 280392 64706 280394
rect 62113 280336 62118 280392
rect 62174 280336 64706 280392
rect 62113 280334 64706 280336
rect 62113 280331 62179 280334
rect 64646 280318 64706 280334
rect 649950 280392 652451 280394
rect 649950 280336 652390 280392
rect 652446 280336 652451 280392
rect 649950 280334 652451 280336
rect 649950 280318 650010 280334
rect 652385 280331 652451 280334
rect 62246 280060 62252 280124
rect 62316 280122 62322 280124
rect 62941 280122 63007 280125
rect 62316 280120 63007 280122
rect 62316 280064 62946 280120
rect 63002 280064 63007 280120
rect 62316 280062 63007 280064
rect 62316 280060 62322 280062
rect 62941 280059 63007 280062
rect 42149 279850 42215 279853
rect 44449 279850 44515 279853
rect 42149 279848 44515 279850
rect 42149 279792 42154 279848
rect 42210 279792 44454 279848
rect 44510 279792 44515 279848
rect 42149 279790 44515 279792
rect 42149 279787 42215 279790
rect 44449 279787 44515 279790
rect 42425 279442 42491 279445
rect 61929 279442 61995 279445
rect 42425 279440 61995 279442
rect 42425 279384 42430 279440
rect 42486 279384 61934 279440
rect 61990 279384 61995 279440
rect 42425 279382 61995 279384
rect 42425 279379 42491 279382
rect 61929 279379 61995 279382
rect 652569 279442 652635 279445
rect 676857 279442 676923 279445
rect 652569 279440 676923 279442
rect 652569 279384 652574 279440
rect 652630 279384 676862 279440
rect 676918 279384 676923 279440
rect 652569 279382 676923 279384
rect 652569 279379 652635 279382
rect 676857 279379 676923 279382
rect 45369 279034 45435 279037
rect 42198 279032 45435 279034
rect 42198 278976 45374 279032
rect 45430 278976 45435 279032
rect 42198 278974 45435 278976
rect 41965 278490 42031 278493
rect 42198 278490 42258 278974
rect 45369 278971 45435 278974
rect 43989 278762 44055 278765
rect 45461 278762 45527 278765
rect 43989 278760 45527 278762
rect 43989 278704 43994 278760
rect 44050 278704 45466 278760
rect 45522 278704 45527 278760
rect 43989 278702 45527 278704
rect 43989 278699 44055 278702
rect 45461 278699 45527 278702
rect 63401 278762 63467 278765
rect 675293 278762 675359 278765
rect 63401 278760 675359 278762
rect 63401 278704 63406 278760
rect 63462 278704 675298 278760
rect 675354 278704 675359 278760
rect 63401 278702 675359 278704
rect 63401 278699 63467 278702
rect 675293 278699 675359 278702
rect 41965 278488 42258 278490
rect 41965 278432 41970 278488
rect 42026 278432 42258 278488
rect 41965 278430 42258 278432
rect 671705 278490 671771 278493
rect 672809 278490 672875 278493
rect 671705 278488 672875 278490
rect 671705 278432 671710 278488
rect 671766 278432 672814 278488
rect 672870 278432 672875 278488
rect 671705 278430 672875 278432
rect 41965 278427 42031 278430
rect 671705 278427 671771 278430
rect 672809 278427 672875 278430
rect 43805 278354 43871 278357
rect 636193 278354 636259 278357
rect 43805 278352 636259 278354
rect 43805 278296 43810 278352
rect 43866 278296 636198 278352
rect 636254 278296 636259 278352
rect 43805 278294 636259 278296
rect 43805 278291 43871 278294
rect 636193 278291 636259 278294
rect 62062 278020 62068 278084
rect 62132 278082 62138 278084
rect 63401 278082 63467 278085
rect 62132 278080 63467 278082
rect 62132 278024 63406 278080
rect 63462 278024 63467 278080
rect 62132 278022 63467 278024
rect 62132 278020 62138 278022
rect 63401 278019 63467 278022
rect 63585 278082 63651 278085
rect 675477 278082 675543 278085
rect 63585 278080 675543 278082
rect 63585 278024 63590 278080
rect 63646 278024 675482 278080
rect 675538 278024 675543 278080
rect 63585 278022 675543 278024
rect 63585 278019 63651 278022
rect 675477 278019 675543 278022
rect 635089 277810 635155 277813
rect 51030 277808 635155 277810
rect 51030 277752 635094 277808
rect 635150 277752 635155 277808
rect 51030 277750 635155 277752
rect 43662 277612 43668 277676
rect 43732 277674 43738 277676
rect 51030 277674 51090 277750
rect 635089 277747 635155 277750
rect 43732 277614 51090 277674
rect 43732 277612 43738 277614
rect 55857 277538 55923 277541
rect 63585 277538 63651 277541
rect 55857 277536 63651 277538
rect 55857 277480 55862 277536
rect 55918 277480 63590 277536
rect 63646 277480 63651 277536
rect 55857 277478 63651 277480
rect 55857 277475 55923 277478
rect 63585 277475 63651 277478
rect 42057 277266 42123 277269
rect 45369 277266 45435 277269
rect 42057 277264 45435 277266
rect 42057 277208 42062 277264
rect 42118 277208 45374 277264
rect 45430 277208 45435 277264
rect 42057 277206 45435 277208
rect 42057 277203 42123 277206
rect 45369 277203 45435 277206
rect 42517 275906 42583 275909
rect 57421 275906 57487 275909
rect 42517 275904 57487 275906
rect 42517 275848 42522 275904
rect 42578 275848 57426 275904
rect 57482 275848 57487 275904
rect 42517 275846 57487 275848
rect 42517 275843 42583 275846
rect 57421 275843 57487 275846
rect 40718 274212 40724 274276
rect 40788 274274 40794 274276
rect 41781 274274 41847 274277
rect 40788 274272 41847 274274
rect 40788 274216 41786 274272
rect 41842 274216 41847 274272
rect 40788 274214 41847 274216
rect 40788 274212 40794 274214
rect 41781 274211 41847 274214
rect 539317 274002 539383 274005
rect 545941 274002 546007 274005
rect 539317 274000 546007 274002
rect 539317 273944 539322 274000
rect 539378 273944 545946 274000
rect 546002 273944 546007 274000
rect 539317 273942 546007 273944
rect 539317 273939 539383 273942
rect 545941 273939 546007 273942
rect 43345 273866 43411 273869
rect 62297 273866 62363 273869
rect 43345 273864 62363 273866
rect 43345 273808 43350 273864
rect 43406 273808 62302 273864
rect 62358 273808 62363 273864
rect 43345 273806 62363 273808
rect 43345 273803 43411 273806
rect 62297 273803 62363 273806
rect 40534 272988 40540 273052
rect 40604 273050 40610 273052
rect 41781 273050 41847 273053
rect 40604 273048 41847 273050
rect 40604 272992 41786 273048
rect 41842 272992 41847 273048
rect 40604 272990 41847 272992
rect 40604 272988 40610 272990
rect 41781 272987 41847 272990
rect 464797 272506 464863 272509
rect 470685 272506 470751 272509
rect 464797 272504 470751 272506
rect 464797 272448 464802 272504
rect 464858 272448 470690 272504
rect 470746 272448 470751 272504
rect 464797 272446 470751 272448
rect 464797 272443 464863 272446
rect 470685 272443 470751 272446
rect 536557 272506 536623 272509
rect 547689 272506 547755 272509
rect 536557 272504 547755 272506
rect 536557 272448 536562 272504
rect 536618 272448 547694 272504
rect 547750 272448 547755 272504
rect 536557 272446 547755 272448
rect 536557 272443 536623 272446
rect 547689 272443 547755 272446
rect 460933 272370 460999 272373
rect 463693 272370 463759 272373
rect 460933 272368 463759 272370
rect 460933 272312 460938 272368
rect 460994 272312 463698 272368
rect 463754 272312 463759 272368
rect 460933 272310 463759 272312
rect 460933 272307 460999 272310
rect 463693 272307 463759 272310
rect 41454 272172 41460 272236
rect 41524 272234 41530 272236
rect 41781 272234 41847 272237
rect 41524 272232 41847 272234
rect 41524 272176 41786 272232
rect 41842 272176 41847 272232
rect 41524 272174 41847 272176
rect 41524 272172 41530 272174
rect 41781 272171 41847 272174
rect 547505 272098 547571 272101
rect 547873 272098 547939 272101
rect 547505 272096 547939 272098
rect 547505 272040 547510 272096
rect 547566 272040 547878 272096
rect 547934 272040 547939 272096
rect 547505 272038 547939 272040
rect 547505 272035 547571 272038
rect 547873 272035 547939 272038
rect 470593 271962 470659 271965
rect 478045 271962 478111 271965
rect 470593 271960 478111 271962
rect 470593 271904 470598 271960
rect 470654 271904 478050 271960
rect 478106 271904 478111 271960
rect 470593 271902 478111 271904
rect 470593 271899 470659 271902
rect 478045 271899 478111 271902
rect 479517 271962 479583 271965
rect 480529 271962 480595 271965
rect 479517 271960 480595 271962
rect 479517 271904 479522 271960
rect 479578 271904 480534 271960
rect 480590 271904 480595 271960
rect 479517 271902 480595 271904
rect 479517 271899 479583 271902
rect 480529 271899 480595 271902
rect 501597 271962 501663 271965
rect 504541 271962 504607 271965
rect 501597 271960 504607 271962
rect 501597 271904 501602 271960
rect 501658 271904 504546 271960
rect 504602 271904 504607 271960
rect 501597 271902 504607 271904
rect 501597 271899 501663 271902
rect 504541 271899 504607 271902
rect 532233 270194 532299 270197
rect 534073 270194 534139 270197
rect 532233 270192 534139 270194
rect 532233 270136 532238 270192
rect 532294 270136 534078 270192
rect 534134 270136 534139 270192
rect 532233 270134 534139 270136
rect 532233 270131 532299 270134
rect 534073 270131 534139 270134
rect 41781 270060 41847 270061
rect 41781 270056 41828 270060
rect 41892 270058 41898 270060
rect 41781 270000 41786 270056
rect 41781 269996 41828 270000
rect 41892 269998 41938 270058
rect 41892 269996 41898 269998
rect 41781 269995 41847 269996
rect 509233 269922 509299 269925
rect 516409 269922 516475 269925
rect 509233 269920 516475 269922
rect 509233 269864 509238 269920
rect 509294 269864 516414 269920
rect 516470 269864 516475 269920
rect 509233 269862 516475 269864
rect 509233 269859 509299 269862
rect 516409 269859 516475 269862
rect 43621 269786 43687 269789
rect 62481 269786 62547 269789
rect 43621 269784 62547 269786
rect 43621 269728 43626 269784
rect 43682 269728 62486 269784
rect 62542 269728 62547 269784
rect 43621 269726 62547 269728
rect 43621 269723 43687 269726
rect 62481 269723 62547 269726
rect 538029 269786 538095 269789
rect 542445 269786 542511 269789
rect 538029 269784 542511 269786
rect 538029 269728 538034 269784
rect 538090 269728 542450 269784
rect 542506 269728 542511 269784
rect 538029 269726 542511 269728
rect 538029 269723 538095 269726
rect 542445 269723 542511 269726
rect 509141 269514 509207 269517
rect 509877 269514 509943 269517
rect 509141 269512 509943 269514
rect 509141 269456 509146 269512
rect 509202 269456 509882 269512
rect 509938 269456 509943 269512
rect 509141 269454 509943 269456
rect 509141 269451 509207 269454
rect 509877 269451 509943 269454
rect 41965 269108 42031 269109
rect 41965 269104 42012 269108
rect 42076 269106 42082 269108
rect 41965 269048 41970 269104
rect 41965 269044 42012 269048
rect 42076 269046 42122 269106
rect 42076 269044 42082 269046
rect 41965 269043 42031 269044
rect 676262 268562 676322 268668
rect 676857 268562 676923 268565
rect 663750 268502 676322 268562
rect 676814 268560 676923 268562
rect 676814 268504 676862 268560
rect 676918 268504 676923 268560
rect 658917 268154 658983 268157
rect 663750 268154 663810 268502
rect 676814 268499 676923 268504
rect 676814 268260 676874 268499
rect 658917 268152 663810 268154
rect 658917 268096 658922 268152
rect 658978 268096 663810 268152
rect 658917 268094 663810 268096
rect 674005 268154 674071 268157
rect 676213 268154 676279 268157
rect 674005 268152 676279 268154
rect 674005 268096 674010 268152
rect 674066 268096 676218 268152
rect 676274 268096 676279 268152
rect 674005 268094 676279 268096
rect 658917 268091 658983 268094
rect 674005 268091 674071 268094
rect 676213 268091 676279 268094
rect 676262 267749 676322 267852
rect 42425 267746 42491 267749
rect 46933 267746 46999 267749
rect 42425 267744 46999 267746
rect 42425 267688 42430 267744
rect 42486 267688 46938 267744
rect 46994 267688 46999 267744
rect 42425 267686 46999 267688
rect 42425 267683 42491 267686
rect 46933 267683 46999 267686
rect 676213 267744 676322 267749
rect 676213 267688 676218 267744
rect 676274 267688 676322 267744
rect 676213 267686 676322 267688
rect 676213 267683 676279 267686
rect 674373 267474 674439 267477
rect 674373 267472 676292 267474
rect 674373 267416 674378 267472
rect 674434 267416 676292 267472
rect 674373 267414 676292 267416
rect 674373 267411 674439 267414
rect 673913 267066 673979 267069
rect 673913 267064 676292 267066
rect 673913 267008 673918 267064
rect 673974 267008 676292 267064
rect 673913 267006 676292 267008
rect 673913 267003 673979 267006
rect 674741 266658 674807 266661
rect 674741 266656 676292 266658
rect 674741 266600 674746 266656
rect 674802 266600 676292 266656
rect 674741 266598 676292 266600
rect 674741 266595 674807 266598
rect 42149 266250 42215 266253
rect 56041 266250 56107 266253
rect 42149 266248 56107 266250
rect 42149 266192 42154 266248
rect 42210 266192 56046 266248
rect 56102 266192 56107 266248
rect 42149 266190 56107 266192
rect 42149 266187 42215 266190
rect 56041 266187 56107 266190
rect 673085 266114 673151 266117
rect 676262 266114 676322 266220
rect 673085 266112 676322 266114
rect 673085 266056 673090 266112
rect 673146 266056 676322 266112
rect 673085 266054 676322 266056
rect 673085 266051 673151 266054
rect 674557 265842 674623 265845
rect 674557 265840 676292 265842
rect 674557 265784 674562 265840
rect 674618 265784 676292 265840
rect 674557 265782 676292 265784
rect 674557 265779 674623 265782
rect 62849 265570 62915 265573
rect 665214 265570 665220 265572
rect 62849 265568 665220 265570
rect 62849 265512 62854 265568
rect 62910 265512 665220 265568
rect 62849 265510 665220 265512
rect 62849 265507 62915 265510
rect 665214 265508 665220 265510
rect 665284 265508 665290 265572
rect 672533 265298 672599 265301
rect 676262 265298 676322 265404
rect 672533 265296 676322 265298
rect 672533 265240 672538 265296
rect 672594 265240 676322 265296
rect 672533 265238 676322 265240
rect 672533 265235 672599 265238
rect 673269 265026 673335 265029
rect 673269 265024 676292 265026
rect 673269 264968 673274 265024
rect 673330 264968 676292 265024
rect 673269 264966 676292 264968
rect 673269 264963 673335 264966
rect 673729 264618 673795 264621
rect 673729 264616 676292 264618
rect 673729 264560 673734 264616
rect 673790 264560 676292 264616
rect 673729 264558 676292 264560
rect 673729 264555 673795 264558
rect 61377 264210 61443 264213
rect 674782 264210 674788 264212
rect 61377 264208 674788 264210
rect 61377 264152 61382 264208
rect 61438 264152 674788 264208
rect 61377 264150 674788 264152
rect 61377 264147 61443 264150
rect 674782 264148 674788 264150
rect 674852 264148 674858 264212
rect 676446 264077 676506 264180
rect 676397 264072 676506 264077
rect 676397 264016 676402 264072
rect 676458 264016 676506 264072
rect 676397 264014 676506 264016
rect 676397 264011 676463 264014
rect 679574 263669 679634 263772
rect 679574 263664 679683 263669
rect 679574 263608 679622 263664
rect 679678 263608 679683 263664
rect 679574 263606 679683 263608
rect 679617 263603 679683 263606
rect 673085 263394 673151 263397
rect 673085 263392 676292 263394
rect 673085 263336 673090 263392
rect 673146 263336 676292 263392
rect 673085 263334 676292 263336
rect 673085 263331 673151 263334
rect 43253 263258 43319 263261
rect 43621 263258 43687 263261
rect 43253 263256 43687 263258
rect 43253 263200 43258 263256
rect 43314 263200 43626 263256
rect 43682 263200 43687 263256
rect 43253 263198 43687 263200
rect 43253 263195 43319 263198
rect 43621 263195 43687 263198
rect 676262 262853 676322 262956
rect 676213 262848 676322 262853
rect 676213 262792 676218 262848
rect 676274 262792 676322 262848
rect 676213 262790 676322 262792
rect 676213 262787 676279 262790
rect 674649 262578 674715 262581
rect 674649 262576 676292 262578
rect 674649 262520 674654 262576
rect 674710 262520 676292 262576
rect 674649 262518 676292 262520
rect 674649 262515 674715 262518
rect 554405 262170 554471 262173
rect 552460 262168 554471 262170
rect 552460 262112 554410 262168
rect 554466 262112 554471 262168
rect 552460 262110 554471 262112
rect 554405 262107 554471 262110
rect 670325 262170 670391 262173
rect 670325 262168 676292 262170
rect 670325 262112 670330 262168
rect 670386 262112 676292 262168
rect 670325 262110 676292 262112
rect 670325 262107 670391 262110
rect 676998 261628 677058 261732
rect 676990 261564 676996 261628
rect 677060 261564 677066 261628
rect 676814 261220 676874 261324
rect 676806 261156 676812 261220
rect 676876 261156 676882 261220
rect 674097 260946 674163 260949
rect 674097 260944 676292 260946
rect 674097 260888 674102 260944
rect 674158 260888 676292 260944
rect 674097 260886 676292 260888
rect 674097 260883 674163 260886
rect 671337 260538 671403 260541
rect 671337 260536 676292 260538
rect 671337 260480 671342 260536
rect 671398 260480 676292 260536
rect 671337 260478 676292 260480
rect 671337 260475 671403 260478
rect 674281 260130 674347 260133
rect 674281 260128 676292 260130
rect 674281 260072 674286 260128
rect 674342 260072 676292 260128
rect 674281 260070 676292 260072
rect 674281 260067 674347 260070
rect 554313 259994 554379 259997
rect 552460 259992 554379 259994
rect 552460 259936 554318 259992
rect 554374 259936 554379 259992
rect 552460 259934 554379 259936
rect 554313 259931 554379 259934
rect 671705 259722 671771 259725
rect 671705 259720 676292 259722
rect 671705 259664 671710 259720
rect 671766 259664 676292 259720
rect 671705 259662 676292 259664
rect 671705 259659 671771 259662
rect 672901 259314 672967 259317
rect 672901 259312 676292 259314
rect 672901 259256 672906 259312
rect 672962 259256 676292 259312
rect 672901 259254 676292 259256
rect 672901 259251 672967 259254
rect 674465 258906 674531 258909
rect 674465 258904 676292 258906
rect 674465 258848 674470 258904
rect 674526 258848 676292 258904
rect 674465 258846 676292 258848
rect 674465 258843 674531 258846
rect 670141 258498 670207 258501
rect 670141 258496 676292 258498
rect 670141 258440 670146 258496
rect 670202 258440 676292 258496
rect 670141 258438 676292 258440
rect 670141 258435 670207 258438
rect 46381 258090 46447 258093
rect 675477 258092 675543 258093
rect 675477 258090 675524 258092
rect 41492 258088 46447 258090
rect 41492 258032 46386 258088
rect 46442 258032 46447 258088
rect 41492 258030 46447 258032
rect 675396 258088 675524 258090
rect 675588 258090 675594 258092
rect 675396 258032 675482 258088
rect 675588 258060 676292 258090
rect 675396 258030 675524 258032
rect 46381 258027 46447 258030
rect 675477 258028 675524 258030
rect 675588 258030 676322 258060
rect 675588 258028 675594 258030
rect 675477 258027 675543 258028
rect 553945 257818 554011 257821
rect 552460 257816 554011 257818
rect 552460 257760 553950 257816
rect 554006 257760 554011 257816
rect 552460 257758 554011 257760
rect 553945 257755 554011 257758
rect 44725 257682 44791 257685
rect 41492 257680 44791 257682
rect 41492 257624 44730 257680
rect 44786 257624 44791 257680
rect 676262 257652 676322 258030
rect 41492 257622 44791 257624
rect 44725 257619 44791 257622
rect 670693 257274 670759 257277
rect 670693 257272 676292 257274
rect 35758 257141 35818 257244
rect 670693 257216 670698 257272
rect 670754 257216 676292 257272
rect 670693 257214 676292 257216
rect 670693 257211 670759 257214
rect 35758 257136 35867 257141
rect 35758 257080 35806 257136
rect 35862 257080 35867 257136
rect 35758 257078 35867 257080
rect 35801 257075 35867 257078
rect 39573 257138 39639 257141
rect 43253 257138 43319 257141
rect 39573 257136 43319 257138
rect 39573 257080 39578 257136
rect 39634 257080 43258 257136
rect 43314 257080 43319 257136
rect 39573 257078 43319 257080
rect 39573 257075 39639 257078
rect 43253 257075 43319 257078
rect 44541 256866 44607 256869
rect 41492 256864 44607 256866
rect 41492 256808 44546 256864
rect 44602 256808 44607 256864
rect 41492 256806 44607 256808
rect 44541 256803 44607 256806
rect 44909 256458 44975 256461
rect 41492 256456 44975 256458
rect 41492 256400 44914 256456
rect 44970 256400 44975 256456
rect 41492 256398 44975 256400
rect 44909 256395 44975 256398
rect 35574 255917 35634 256020
rect 35574 255912 35683 255917
rect 35574 255856 35622 255912
rect 35678 255856 35683 255912
rect 35574 255854 35683 255856
rect 35617 255851 35683 255854
rect 39941 255914 40007 255917
rect 43069 255914 43135 255917
rect 39941 255912 43135 255914
rect 39941 255856 39946 255912
rect 40002 255856 43074 255912
rect 43130 255856 43135 255912
rect 39941 255854 43135 255856
rect 39941 255851 40007 255854
rect 43069 255851 43135 255854
rect 554497 255642 554563 255645
rect 552460 255640 554563 255642
rect 35758 255509 35818 255612
rect 552460 255584 554502 255640
rect 554558 255584 554563 255640
rect 552460 255582 554563 255584
rect 554497 255579 554563 255582
rect 35758 255504 35867 255509
rect 35758 255448 35806 255504
rect 35862 255448 35867 255504
rect 35758 255446 35867 255448
rect 35801 255443 35867 255446
rect 44265 255234 44331 255237
rect 41492 255232 44331 255234
rect 41492 255176 44270 255232
rect 44326 255176 44331 255232
rect 41492 255174 44331 255176
rect 44265 255171 44331 255174
rect 35758 254693 35818 254796
rect 35758 254688 35867 254693
rect 35758 254632 35806 254688
rect 35862 254632 35867 254688
rect 35758 254630 35867 254632
rect 35801 254627 35867 254630
rect 40493 254690 40559 254693
rect 43805 254690 43871 254693
rect 40493 254688 43871 254690
rect 40493 254632 40498 254688
rect 40554 254632 43810 254688
rect 43866 254632 43871 254688
rect 40493 254630 43871 254632
rect 40493 254627 40559 254630
rect 43805 254627 43871 254630
rect 35574 254285 35634 254388
rect 35574 254280 35683 254285
rect 35574 254224 35622 254280
rect 35678 254224 35683 254280
rect 35574 254222 35683 254224
rect 35617 254219 35683 254222
rect 35758 253877 35818 253980
rect 35758 253872 35867 253877
rect 35758 253816 35806 253872
rect 35862 253816 35867 253872
rect 35758 253814 35867 253816
rect 35801 253811 35867 253814
rect 41505 253874 41571 253877
rect 43621 253874 43687 253877
rect 41505 253872 43687 253874
rect 41505 253816 41510 253872
rect 41566 253816 43626 253872
rect 43682 253816 43687 253872
rect 41505 253814 43687 253816
rect 41505 253811 41571 253814
rect 43621 253811 43687 253814
rect 35574 253469 35634 253572
rect 35574 253464 35683 253469
rect 554405 253466 554471 253469
rect 35574 253408 35622 253464
rect 35678 253408 35683 253464
rect 35574 253406 35683 253408
rect 552460 253464 554471 253466
rect 552460 253408 554410 253464
rect 554466 253408 554471 253464
rect 552460 253406 554471 253408
rect 35617 253403 35683 253406
rect 554405 253403 554471 253406
rect 674925 253194 674991 253197
rect 675845 253194 675911 253197
rect 674925 253192 675911 253194
rect 35758 253061 35818 253164
rect 674925 253136 674930 253192
rect 674986 253136 675850 253192
rect 675906 253136 675911 253192
rect 674925 253134 675911 253136
rect 674925 253131 674991 253134
rect 675845 253131 675911 253134
rect 35758 253056 35867 253061
rect 35758 253000 35806 253056
rect 35862 253000 35867 253056
rect 35758 252998 35867 253000
rect 35801 252995 35867 252998
rect 40677 253058 40743 253061
rect 42885 253058 42951 253061
rect 40677 253056 42951 253058
rect 40677 253000 40682 253056
rect 40738 253000 42890 253056
rect 42946 253000 42951 253056
rect 40677 252998 42951 253000
rect 40677 252995 40743 252998
rect 42885 252995 42951 252998
rect 46933 252786 46999 252789
rect 41492 252784 46999 252786
rect 41492 252728 46938 252784
rect 46994 252728 46999 252784
rect 41492 252726 46999 252728
rect 46933 252723 46999 252726
rect 35758 252245 35818 252348
rect 35758 252240 35867 252245
rect 35758 252184 35806 252240
rect 35862 252184 35867 252240
rect 35758 252182 35867 252184
rect 35801 252179 35867 252182
rect 47117 251970 47183 251973
rect 41492 251968 47183 251970
rect 41492 251912 47122 251968
rect 47178 251912 47183 251968
rect 41492 251910 47183 251912
rect 47117 251907 47183 251910
rect 44449 251562 44515 251565
rect 41492 251560 44515 251562
rect 41492 251504 44454 251560
rect 44510 251504 44515 251560
rect 41492 251502 44515 251504
rect 44449 251499 44515 251502
rect 554129 251290 554195 251293
rect 552460 251288 554195 251290
rect 552460 251232 554134 251288
rect 554190 251232 554195 251288
rect 552460 251230 554195 251232
rect 554129 251227 554195 251230
rect 44633 251154 44699 251157
rect 41492 251152 44699 251154
rect 41492 251096 44638 251152
rect 44694 251096 44699 251152
rect 41492 251094 44699 251096
rect 44633 251091 44699 251094
rect 673085 250746 673151 250749
rect 675477 250746 675543 250749
rect 673085 250744 675543 250746
rect 35758 250613 35818 250716
rect 673085 250688 673090 250744
rect 673146 250688 675482 250744
rect 675538 250688 675543 250744
rect 673085 250686 675543 250688
rect 673085 250683 673151 250686
rect 675477 250683 675543 250686
rect 35758 250608 35867 250613
rect 35758 250552 35806 250608
rect 35862 250552 35867 250608
rect 35758 250550 35867 250552
rect 35801 250547 35867 250550
rect 44173 250338 44239 250341
rect 41492 250336 44239 250338
rect 41492 250280 44178 250336
rect 44234 250280 44239 250336
rect 41492 250278 44239 250280
rect 44173 250275 44239 250278
rect 675753 250338 675819 250341
rect 676990 250338 676996 250340
rect 675753 250336 676996 250338
rect 675753 250280 675758 250336
rect 675814 250280 676996 250336
rect 675753 250278 676996 250280
rect 675753 250275 675819 250278
rect 676990 250276 676996 250278
rect 677060 250276 677066 250340
rect 40542 249796 40602 249900
rect 40534 249732 40540 249796
rect 40604 249732 40610 249796
rect 673085 249658 673151 249661
rect 674782 249658 674788 249660
rect 673085 249656 674788 249658
rect 673085 249600 673090 249656
rect 673146 249600 674788 249656
rect 673085 249598 674788 249600
rect 673085 249595 673151 249598
rect 674782 249596 674788 249598
rect 674852 249596 674858 249660
rect 675518 249658 675524 249660
rect 674974 249598 675524 249658
rect 40726 249388 40786 249492
rect 40718 249324 40724 249388
rect 40788 249324 40794 249388
rect 45553 249114 45619 249117
rect 554037 249114 554103 249117
rect 41492 249112 45619 249114
rect 41492 249056 45558 249112
rect 45614 249056 45619 249112
rect 41492 249054 45619 249056
rect 552460 249112 554103 249114
rect 552460 249056 554042 249112
rect 554098 249056 554103 249112
rect 552460 249054 554103 249056
rect 45553 249051 45619 249054
rect 554037 249051 554103 249054
rect 674974 248845 675034 249598
rect 675518 249596 675524 249598
rect 675588 249596 675594 249660
rect 674925 248840 675034 248845
rect 674925 248784 674930 248840
rect 674986 248784 675034 248840
rect 674925 248782 675034 248784
rect 674925 248779 674991 248782
rect 45921 248706 45987 248709
rect 41492 248704 45987 248706
rect 41492 248648 45926 248704
rect 45982 248648 45987 248704
rect 41492 248646 45987 248648
rect 45921 248643 45987 248646
rect 45737 248298 45803 248301
rect 41492 248296 45803 248298
rect 41492 248240 45742 248296
rect 45798 248240 45803 248296
rect 41492 248238 45803 248240
rect 45737 248235 45803 248238
rect 664437 248298 664503 248301
rect 675385 248298 675451 248301
rect 664437 248296 675451 248298
rect 664437 248240 664442 248296
rect 664498 248240 675390 248296
rect 675446 248240 675451 248296
rect 664437 248238 675451 248240
rect 664437 248235 664503 248238
rect 675385 248235 675451 248238
rect 50521 247890 50587 247893
rect 41492 247888 50587 247890
rect 41492 247832 50526 247888
rect 50582 247832 50587 247888
rect 41492 247830 50587 247832
rect 50521 247827 50587 247830
rect 47761 247482 47827 247485
rect 41492 247480 47827 247482
rect 41492 247424 47766 247480
rect 47822 247424 47827 247480
rect 41492 247422 47827 247424
rect 47761 247419 47827 247422
rect 46105 247074 46171 247077
rect 41492 247072 46171 247074
rect 41492 247016 46110 247072
rect 46166 247016 46171 247072
rect 41492 247014 46171 247016
rect 46105 247011 46171 247014
rect 553853 246938 553919 246941
rect 552460 246936 553919 246938
rect 552460 246880 553858 246936
rect 553914 246880 553919 246936
rect 552460 246878 553919 246880
rect 553853 246875 553919 246878
rect 674097 246666 674163 246669
rect 675293 246666 675359 246669
rect 674097 246664 675359 246666
rect 674097 246608 674102 246664
rect 674158 246608 675298 246664
rect 675354 246608 675359 246664
rect 674097 246606 675359 246608
rect 674097 246603 674163 246606
rect 675293 246603 675359 246606
rect 675753 246666 675819 246669
rect 676806 246666 676812 246668
rect 675753 246664 676812 246666
rect 675753 246608 675758 246664
rect 675814 246608 676812 246664
rect 675753 246606 676812 246608
rect 675753 246603 675819 246606
rect 676806 246604 676812 246606
rect 676876 246604 676882 246668
rect 673453 246258 673519 246261
rect 674598 246258 674604 246260
rect 673453 246256 674604 246258
rect 673453 246200 673458 246256
rect 673514 246200 674604 246256
rect 673453 246198 674604 246200
rect 673453 246195 673519 246198
rect 674598 246196 674604 246198
rect 674668 246196 674674 246260
rect 672165 246122 672231 246125
rect 673310 246122 673316 246124
rect 672165 246120 673316 246122
rect 672165 246064 672170 246120
rect 672226 246064 673316 246120
rect 672165 246062 673316 246064
rect 672165 246059 672231 246062
rect 673310 246060 673316 246062
rect 673380 246060 673386 246124
rect 673085 245850 673151 245853
rect 675334 245850 675340 245852
rect 673085 245848 675340 245850
rect 673085 245792 673090 245848
rect 673146 245792 675340 245848
rect 673085 245790 675340 245792
rect 673085 245787 673151 245790
rect 675334 245788 675340 245790
rect 675404 245788 675410 245852
rect 40309 245714 40375 245717
rect 43069 245714 43135 245717
rect 40309 245712 43135 245714
rect 40309 245656 40314 245712
rect 40370 245656 43074 245712
rect 43130 245656 43135 245712
rect 40309 245654 43135 245656
rect 40309 245651 40375 245654
rect 43069 245651 43135 245654
rect 671705 245578 671771 245581
rect 675201 245578 675267 245581
rect 671705 245576 675267 245578
rect 671705 245520 671710 245576
rect 671766 245520 675206 245576
rect 675262 245520 675267 245576
rect 671705 245518 675267 245520
rect 671705 245515 671771 245518
rect 675201 245515 675267 245518
rect 553485 244762 553551 244765
rect 552460 244760 553551 244762
rect 552460 244704 553490 244760
rect 553546 244704 553551 244760
rect 552460 244702 553551 244704
rect 553485 244699 553551 244702
rect 672901 242722 672967 242725
rect 675385 242722 675451 242725
rect 672901 242720 675451 242722
rect 672901 242664 672906 242720
rect 672962 242664 675390 242720
rect 675446 242664 675451 242720
rect 672901 242662 675451 242664
rect 672901 242659 672967 242662
rect 675385 242659 675451 242662
rect 553669 242586 553735 242589
rect 552460 242584 553735 242586
rect 552460 242528 553674 242584
rect 553730 242528 553735 242584
rect 552460 242526 553735 242528
rect 553669 242523 553735 242526
rect 674281 242314 674347 242317
rect 675385 242314 675451 242317
rect 674281 242312 675451 242314
rect 674281 242256 674286 242312
rect 674342 242256 675390 242312
rect 675446 242256 675451 242312
rect 674281 242254 675451 242256
rect 674281 242251 674347 242254
rect 675385 242251 675451 242254
rect 673729 242042 673795 242045
rect 676806 242042 676812 242044
rect 673729 242040 676812 242042
rect 673729 241984 673734 242040
rect 673790 241984 676812 242040
rect 673729 241982 676812 241984
rect 673729 241979 673795 241982
rect 676806 241980 676812 241982
rect 676876 241980 676882 242044
rect 673269 241770 673335 241773
rect 674833 241770 674899 241773
rect 673269 241768 674899 241770
rect 673269 241712 673274 241768
rect 673330 241712 674838 241768
rect 674894 241712 674899 241768
rect 673269 241710 674899 241712
rect 673269 241707 673335 241710
rect 674833 241707 674899 241710
rect 674465 241498 674531 241501
rect 675385 241498 675451 241501
rect 674465 241496 675451 241498
rect 674465 241440 674470 241496
rect 674526 241440 675390 241496
rect 675446 241440 675451 241496
rect 674465 241438 675451 241440
rect 674465 241435 674531 241438
rect 675385 241435 675451 241438
rect 554497 240410 554563 240413
rect 552460 240408 554563 240410
rect 552460 240352 554502 240408
rect 554558 240352 554563 240408
rect 552460 240350 554563 240352
rect 554497 240347 554563 240350
rect 671337 240274 671403 240277
rect 675385 240274 675451 240277
rect 671337 240272 675451 240274
rect 671337 240216 671342 240272
rect 671398 240216 675390 240272
rect 675446 240216 675451 240272
rect 671337 240214 675451 240216
rect 671337 240211 671403 240214
rect 675385 240211 675451 240214
rect 42241 240138 42307 240141
rect 44449 240138 44515 240141
rect 42241 240136 44515 240138
rect 42241 240080 42246 240136
rect 42302 240080 44454 240136
rect 44510 240080 44515 240136
rect 42241 240078 44515 240080
rect 42241 240075 42307 240078
rect 44449 240075 44515 240078
rect 42241 238506 42307 238509
rect 46105 238506 46171 238509
rect 42241 238504 46171 238506
rect 42241 238448 42246 238504
rect 42302 238448 46110 238504
rect 46166 238448 46171 238504
rect 42241 238446 46171 238448
rect 42241 238443 42307 238446
rect 46105 238443 46171 238446
rect 554313 238234 554379 238237
rect 552460 238232 554379 238234
rect 552460 238176 554318 238232
rect 554374 238176 554379 238232
rect 552460 238174 554379 238176
rect 554313 238171 554379 238174
rect 42006 237356 42012 237420
rect 42076 237418 42082 237420
rect 42701 237418 42767 237421
rect 42076 237416 42767 237418
rect 42076 237360 42706 237416
rect 42762 237360 42767 237416
rect 42076 237358 42767 237360
rect 42076 237356 42082 237358
rect 42701 237355 42767 237358
rect 670325 237282 670391 237285
rect 675109 237282 675175 237285
rect 670325 237280 675175 237282
rect 670325 237224 670330 237280
rect 670386 237224 675114 237280
rect 675170 237224 675175 237280
rect 670325 237222 675175 237224
rect 670325 237219 670391 237222
rect 675109 237219 675175 237222
rect 670734 236676 670740 236740
rect 670804 236738 670810 236740
rect 671797 236738 671863 236741
rect 670804 236736 671863 236738
rect 670804 236680 671802 236736
rect 671858 236680 671863 236736
rect 670804 236678 671863 236680
rect 670804 236676 670810 236678
rect 671797 236675 671863 236678
rect 672947 236738 673013 236741
rect 674189 236738 674255 236741
rect 672947 236736 674255 236738
rect 672947 236680 672952 236736
rect 673008 236680 674194 236736
rect 674250 236680 674255 236736
rect 672947 236678 674255 236680
rect 672947 236675 673013 236678
rect 674189 236675 674255 236678
rect 40534 236540 40540 236604
rect 40604 236602 40610 236604
rect 41781 236602 41847 236605
rect 40604 236600 41847 236602
rect 40604 236544 41786 236600
rect 41842 236544 41847 236600
rect 40604 236542 41847 236544
rect 40604 236540 40610 236542
rect 41781 236539 41847 236542
rect 553761 236058 553827 236061
rect 552460 236056 553827 236058
rect 552460 236000 553766 236056
rect 553822 236000 553827 236056
rect 552460 235998 553827 236000
rect 553761 235995 553827 235998
rect 42333 235922 42399 235925
rect 45737 235922 45803 235925
rect 42333 235920 45803 235922
rect 42333 235864 42338 235920
rect 42394 235864 45742 235920
rect 45798 235864 45803 235920
rect 42333 235862 45803 235864
rect 42333 235859 42399 235862
rect 45737 235859 45803 235862
rect 675334 235180 675340 235244
rect 675404 235242 675410 235244
rect 676029 235242 676095 235245
rect 675404 235240 676095 235242
rect 675404 235184 676034 235240
rect 676090 235184 676095 235240
rect 675404 235182 676095 235184
rect 675404 235180 675410 235182
rect 676029 235179 676095 235182
rect 40718 234636 40724 234700
rect 40788 234698 40794 234700
rect 41781 234698 41847 234701
rect 40788 234696 41847 234698
rect 40788 234640 41786 234696
rect 41842 234640 41847 234696
rect 40788 234638 41847 234640
rect 40788 234636 40794 234638
rect 41781 234635 41847 234638
rect 554405 233882 554471 233885
rect 552460 233880 554471 233882
rect 552460 233824 554410 233880
rect 554466 233824 554471 233880
rect 552460 233822 554471 233824
rect 554405 233819 554471 233822
rect 668761 232930 668827 232933
rect 672809 232930 672875 232933
rect 668761 232928 672875 232930
rect 668761 232872 668766 232928
rect 668822 232872 672814 232928
rect 672870 232872 672875 232928
rect 668761 232870 672875 232872
rect 668761 232867 668827 232870
rect 672809 232867 672875 232870
rect 42701 232250 42767 232253
rect 45921 232250 45987 232253
rect 42701 232248 45987 232250
rect 42701 232192 42706 232248
rect 42762 232192 45926 232248
rect 45982 232192 45987 232248
rect 42701 232190 45987 232192
rect 42701 232187 42767 232190
rect 45921 232187 45987 232190
rect 42333 231978 42399 231981
rect 47117 231978 47183 231981
rect 42333 231976 47183 231978
rect 42333 231920 42338 231976
rect 42394 231920 47122 231976
rect 47178 231920 47183 231976
rect 42333 231918 47183 231920
rect 42333 231915 42399 231918
rect 47117 231915 47183 231918
rect 42333 231298 42399 231301
rect 45553 231298 45619 231301
rect 42333 231296 45619 231298
rect 42333 231240 42338 231296
rect 42394 231240 45558 231296
rect 45614 231240 45619 231296
rect 42333 231238 45619 231240
rect 42333 231235 42399 231238
rect 45553 231235 45619 231238
rect 64137 231162 64203 231165
rect 667054 231162 667060 231164
rect 64137 231160 667060 231162
rect 64137 231104 64142 231160
rect 64198 231104 667060 231160
rect 64137 231102 667060 231104
rect 64137 231099 64203 231102
rect 667054 231100 667060 231102
rect 667124 231100 667130 231164
rect 664897 230482 664963 230485
rect 674669 230482 674735 230485
rect 664897 230480 674735 230482
rect 664897 230424 664902 230480
rect 664958 230424 674674 230480
rect 674730 230424 674735 230480
rect 664897 230422 674735 230424
rect 664897 230419 664963 230422
rect 674669 230419 674735 230422
rect 674833 230482 674899 230485
rect 675150 230482 675156 230484
rect 674833 230480 675156 230482
rect 674833 230424 674838 230480
rect 674894 230424 675156 230480
rect 674833 230422 675156 230424
rect 674833 230419 674899 230422
rect 675150 230420 675156 230422
rect 675220 230420 675226 230484
rect 42149 230346 42215 230349
rect 44173 230346 44239 230349
rect 42149 230344 44239 230346
rect 42149 230288 42154 230344
rect 42210 230288 44178 230344
rect 44234 230288 44239 230344
rect 42149 230286 44239 230288
rect 42149 230283 42215 230286
rect 44173 230283 44239 230286
rect 142153 230210 142219 230213
rect 150525 230210 150591 230213
rect 157425 230210 157491 230213
rect 142153 230208 150591 230210
rect 142153 230152 142158 230208
rect 142214 230152 150530 230208
rect 150586 230152 150591 230208
rect 142153 230150 150591 230152
rect 142153 230147 142219 230150
rect 150525 230147 150591 230150
rect 157382 230208 157491 230210
rect 157382 230152 157430 230208
rect 157486 230152 157491 230208
rect 157382 230147 157491 230152
rect 157793 230210 157859 230213
rect 161289 230210 161355 230213
rect 157793 230208 161355 230210
rect 157793 230152 157798 230208
rect 157854 230152 161294 230208
rect 161350 230152 161355 230208
rect 157793 230150 161355 230152
rect 157793 230147 157859 230150
rect 161289 230147 161355 230150
rect 673867 230210 673933 230213
rect 676765 230210 676831 230213
rect 673867 230208 676831 230210
rect 673867 230152 673872 230208
rect 673928 230152 676770 230208
rect 676826 230152 676831 230208
rect 673867 230150 676831 230152
rect 673867 230147 673933 230150
rect 676765 230147 676831 230150
rect 157149 230074 157215 230077
rect 157382 230074 157442 230147
rect 157149 230072 157442 230074
rect 157149 230016 157154 230072
rect 157210 230016 157442 230072
rect 157149 230014 157442 230016
rect 157149 230011 157215 230014
rect 141969 229938 142035 229941
rect 142613 229938 142679 229941
rect 141969 229936 142679 229938
rect 141969 229880 141974 229936
rect 142030 229880 142618 229936
rect 142674 229880 142679 229936
rect 141969 229878 142679 229880
rect 141969 229875 142035 229878
rect 142613 229875 142679 229878
rect 195053 229938 195119 229941
rect 196893 229938 196959 229941
rect 195053 229936 196959 229938
rect 195053 229880 195058 229936
rect 195114 229880 196898 229936
rect 196954 229880 196959 229936
rect 195053 229878 196959 229880
rect 195053 229875 195119 229878
rect 196893 229875 196959 229878
rect 157609 229666 157675 229669
rect 158713 229666 158779 229669
rect 157609 229664 158779 229666
rect 157609 229608 157614 229664
rect 157670 229608 158718 229664
rect 158774 229608 158779 229664
rect 157609 229606 158779 229608
rect 157609 229603 157675 229606
rect 158713 229603 158779 229606
rect 144637 229394 144703 229397
rect 148317 229394 148383 229397
rect 144637 229392 148383 229394
rect 144637 229336 144642 229392
rect 144698 229336 148322 229392
rect 148378 229336 148383 229392
rect 144637 229334 148383 229336
rect 144637 229331 144703 229334
rect 148317 229331 148383 229334
rect 167361 229258 167427 229261
rect 174353 229258 174419 229261
rect 167361 229256 174419 229258
rect 167361 229200 167366 229256
rect 167422 229200 174358 229256
rect 174414 229200 174419 229256
rect 167361 229198 174419 229200
rect 167361 229195 167427 229198
rect 174353 229195 174419 229198
rect 140037 229122 140103 229125
rect 143533 229122 143599 229125
rect 140037 229120 143599 229122
rect 140037 229064 140042 229120
rect 140098 229064 143538 229120
rect 143594 229064 143599 229120
rect 140037 229062 143599 229064
rect 140037 229059 140103 229062
rect 143533 229059 143599 229062
rect 150341 229122 150407 229125
rect 157149 229122 157215 229125
rect 150341 229120 157215 229122
rect 150341 229064 150346 229120
rect 150402 229064 157154 229120
rect 157210 229064 157215 229120
rect 150341 229062 157215 229064
rect 150341 229059 150407 229062
rect 157149 229059 157215 229062
rect 663701 229122 663767 229125
rect 673269 229122 673335 229125
rect 663701 229120 673335 229122
rect 663701 229064 663706 229120
rect 663762 229064 673274 229120
rect 673330 229064 673335 229120
rect 663701 229062 673335 229064
rect 663701 229059 663767 229062
rect 673269 229059 673335 229062
rect 193029 228986 193095 228989
rect 195605 228986 195671 228989
rect 193029 228984 195671 228986
rect 193029 228928 193034 228984
rect 193090 228928 195610 228984
rect 195666 228928 195671 228984
rect 193029 228926 195671 228928
rect 193029 228923 193095 228926
rect 195605 228923 195671 228926
rect 166349 228850 166415 228853
rect 167545 228850 167611 228853
rect 166349 228848 167611 228850
rect 166349 228792 166354 228848
rect 166410 228792 167550 228848
rect 167606 228792 167611 228848
rect 166349 228790 167611 228792
rect 166349 228787 166415 228790
rect 167545 228787 167611 228790
rect 673867 228714 673933 228717
rect 673867 228712 675218 228714
rect 673867 228656 673872 228712
rect 673928 228656 675218 228712
rect 673867 228654 675218 228656
rect 673867 228651 673933 228654
rect 160001 228578 160067 228581
rect 166809 228578 166875 228581
rect 160001 228576 166875 228578
rect 160001 228520 160006 228576
rect 160062 228520 166814 228576
rect 166870 228520 166875 228576
rect 160001 228518 166875 228520
rect 160001 228515 160067 228518
rect 166809 228515 166875 228518
rect 662137 228578 662203 228581
rect 673085 228578 673151 228581
rect 662137 228576 673151 228578
rect 662137 228520 662142 228576
rect 662198 228520 673090 228576
rect 673146 228520 673151 228576
rect 662137 228518 673151 228520
rect 675158 228578 675218 228654
rect 676397 228578 676463 228581
rect 675158 228576 676463 228578
rect 675158 228520 676402 228576
rect 676458 228520 676463 228576
rect 675158 228518 676463 228520
rect 662137 228515 662203 228518
rect 673085 228515 673151 228518
rect 676397 228515 676463 228518
rect 145925 228034 145991 228037
rect 147121 228034 147187 228037
rect 145925 228032 147187 228034
rect 145925 227976 145930 228032
rect 145986 227976 147126 228032
rect 147182 227976 147187 228032
rect 145925 227974 147187 227976
rect 145925 227971 145991 227974
rect 147121 227971 147187 227974
rect 136633 227898 136699 227901
rect 141509 227898 141575 227901
rect 136633 227896 141575 227898
rect 136633 227840 136638 227896
rect 136694 227840 141514 227896
rect 141570 227840 141575 227896
rect 136633 227838 141575 227840
rect 136633 227835 136699 227838
rect 141509 227835 141575 227838
rect 204805 227626 204871 227629
rect 205633 227626 205699 227629
rect 204805 227624 205699 227626
rect 204805 227568 204810 227624
rect 204866 227568 205638 227624
rect 205694 227568 205699 227624
rect 204805 227566 205699 227568
rect 204805 227563 204871 227566
rect 205633 227563 205699 227566
rect 157333 227490 157399 227493
rect 166533 227490 166599 227493
rect 157333 227488 166599 227490
rect 157333 227432 157338 227488
rect 157394 227432 166538 227488
rect 166594 227432 166599 227488
rect 157333 227430 166599 227432
rect 157333 227427 157399 227430
rect 166533 227427 166599 227430
rect 41965 227356 42031 227357
rect 41965 227352 42012 227356
rect 42076 227354 42082 227356
rect 169385 227354 169451 227357
rect 171685 227354 171751 227357
rect 41965 227296 41970 227352
rect 41965 227292 42012 227296
rect 42076 227294 42122 227354
rect 169385 227352 171751 227354
rect 169385 227296 169390 227352
rect 169446 227296 171690 227352
rect 171746 227296 171751 227352
rect 169385 227294 171751 227296
rect 42076 227292 42082 227294
rect 41965 227291 42031 227292
rect 169385 227291 169451 227294
rect 171685 227291 171751 227294
rect 157425 227218 157491 227221
rect 157382 227216 157491 227218
rect 157382 227160 157430 227216
rect 157486 227160 157491 227216
rect 157382 227155 157491 227160
rect 155861 227082 155927 227085
rect 157382 227082 157442 227155
rect 155861 227080 157442 227082
rect 155861 227024 155866 227080
rect 155922 227024 157442 227080
rect 155861 227022 157442 227024
rect 672349 227082 672415 227085
rect 672574 227082 672580 227084
rect 672349 227080 672580 227082
rect 672349 227024 672354 227080
rect 672410 227024 672580 227080
rect 672349 227022 672580 227024
rect 155861 227019 155927 227022
rect 672349 227019 672415 227022
rect 672574 227020 672580 227022
rect 672644 227020 672650 227084
rect 673453 227082 673519 227085
rect 677317 227082 677383 227085
rect 673453 227080 677383 227082
rect 673453 227024 673458 227080
rect 673514 227024 677322 227080
rect 677378 227024 677383 227080
rect 673453 227022 677383 227024
rect 673453 227019 673519 227022
rect 677317 227019 677383 227022
rect 652385 226946 652451 226949
rect 652385 226944 663810 226946
rect 652385 226888 652390 226944
rect 652446 226888 663810 226944
rect 652385 226886 663810 226888
rect 652385 226883 652451 226886
rect 663750 226810 663810 226886
rect 674046 226810 674052 226812
rect 663750 226750 674052 226810
rect 674046 226748 674052 226750
rect 674116 226748 674122 226812
rect 42149 226674 42215 226677
rect 44633 226674 44699 226677
rect 42149 226672 44699 226674
rect 42149 226616 42154 226672
rect 42210 226616 44638 226672
rect 44694 226616 44699 226672
rect 42149 226614 44699 226616
rect 42149 226611 42215 226614
rect 44633 226611 44699 226614
rect 141785 226538 141851 226541
rect 142245 226538 142311 226541
rect 141785 226536 142311 226538
rect 141785 226480 141790 226536
rect 141846 226480 142250 226536
rect 142306 226480 142311 226536
rect 141785 226478 142311 226480
rect 141785 226475 141851 226478
rect 142245 226475 142311 226478
rect 658917 226402 658983 226405
rect 672717 226402 672783 226405
rect 658917 226400 672783 226402
rect 658917 226344 658922 226400
rect 658978 226344 672722 226400
rect 672778 226344 672783 226400
rect 658917 226342 672783 226344
rect 658917 226339 658983 226342
rect 672717 226339 672783 226342
rect 151353 226266 151419 226269
rect 157149 226266 157215 226269
rect 151353 226264 157215 226266
rect 151353 226208 151358 226264
rect 151414 226208 157154 226264
rect 157210 226208 157215 226264
rect 151353 226206 157215 226208
rect 151353 226203 151419 226206
rect 157149 226203 157215 226206
rect 672597 226130 672663 226133
rect 674833 226130 674899 226133
rect 672597 226128 674899 226130
rect 672597 226072 672602 226128
rect 672658 226072 674838 226128
rect 674894 226072 674899 226128
rect 672597 226070 674899 226072
rect 672597 226067 672663 226070
rect 674833 226067 674899 226070
rect 142613 225994 142679 225997
rect 149789 225994 149855 225997
rect 142613 225992 149855 225994
rect 142613 225936 142618 225992
rect 142674 225936 149794 225992
rect 149850 225936 149855 225992
rect 142613 225934 149855 225936
rect 142613 225931 142679 225934
rect 149789 225931 149855 225934
rect 667013 225994 667079 225997
rect 672487 225994 672553 225997
rect 667013 225992 672553 225994
rect 667013 225936 667018 225992
rect 667074 225936 672492 225992
rect 672548 225936 672553 225992
rect 667013 225934 672553 225936
rect 667013 225931 667079 225934
rect 672487 225931 672553 225934
rect 156597 225858 156663 225861
rect 157793 225858 157859 225861
rect 156597 225856 157859 225858
rect 156597 225800 156602 225856
rect 156658 225800 157798 225856
rect 157854 225800 157859 225856
rect 156597 225798 157859 225800
rect 156597 225795 156663 225798
rect 157793 225795 157859 225798
rect 652753 225722 652819 225725
rect 671981 225722 672047 225725
rect 652753 225720 672047 225722
rect 652753 225664 652758 225720
rect 652814 225664 671986 225720
rect 672042 225664 672047 225720
rect 652753 225662 672047 225664
rect 652753 225659 652819 225662
rect 671981 225659 672047 225662
rect 672165 225722 672231 225725
rect 675201 225722 675267 225725
rect 672165 225720 675267 225722
rect 672165 225664 672170 225720
rect 672226 225664 675206 225720
rect 675262 225664 675267 225720
rect 672165 225662 675267 225664
rect 672165 225659 672231 225662
rect 675201 225659 675267 225662
rect 148869 225450 148935 225453
rect 157149 225450 157215 225453
rect 148869 225448 157215 225450
rect 148869 225392 148874 225448
rect 148930 225392 157154 225448
rect 157210 225392 157215 225448
rect 148869 225390 157215 225392
rect 148869 225387 148935 225390
rect 157149 225387 157215 225390
rect 656157 225314 656223 225317
rect 667013 225314 667079 225317
rect 672257 225314 672323 225317
rect 656157 225312 667079 225314
rect 656157 225256 656162 225312
rect 656218 225256 667018 225312
rect 667074 225256 667079 225312
rect 656157 225254 667079 225256
rect 656157 225251 656223 225254
rect 667013 225251 667079 225254
rect 667982 225312 672323 225314
rect 667982 225256 672262 225312
rect 672318 225256 672323 225312
rect 667982 225254 672323 225256
rect 650637 225042 650703 225045
rect 667982 225042 668042 225254
rect 672257 225251 672323 225254
rect 650637 225040 668042 225042
rect 650637 224984 650642 225040
rect 650698 224984 668042 225040
rect 650637 224982 668042 224984
rect 672165 225042 672231 225045
rect 675661 225042 675727 225045
rect 672165 225040 675727 225042
rect 672165 224984 672170 225040
rect 672226 224984 675666 225040
rect 675722 224984 675727 225040
rect 672165 224982 675727 224984
rect 650637 224979 650703 224982
rect 672165 224979 672231 224982
rect 675661 224979 675727 224982
rect 554773 224906 554839 224909
rect 561673 224906 561739 224909
rect 554773 224904 561739 224906
rect 554773 224848 554778 224904
rect 554834 224848 561678 224904
rect 561734 224848 561739 224904
rect 554773 224846 561739 224848
rect 554773 224843 554839 224846
rect 561673 224843 561739 224846
rect 562133 224770 562199 224773
rect 563789 224770 563855 224773
rect 671613 224772 671679 224773
rect 671613 224770 671660 224772
rect 562133 224768 563855 224770
rect 562133 224712 562138 224768
rect 562194 224712 563794 224768
rect 563850 224712 563855 224768
rect 562133 224710 563855 224712
rect 671568 224768 671660 224770
rect 671568 224712 671618 224768
rect 671568 224710 671660 224712
rect 562133 224707 562199 224710
rect 563789 224707 563855 224710
rect 671613 224708 671660 224710
rect 671724 224708 671730 224772
rect 671613 224707 671679 224708
rect 549253 224498 549319 224501
rect 549897 224498 549963 224501
rect 552841 224498 552907 224501
rect 549253 224496 552907 224498
rect 549253 224440 549258 224496
rect 549314 224440 549902 224496
rect 549958 224440 552846 224496
rect 552902 224440 552907 224496
rect 549253 224438 552907 224440
rect 549253 224435 549319 224438
rect 549897 224435 549963 224438
rect 552841 224435 552907 224438
rect 670509 224500 670575 224501
rect 670509 224496 670556 224500
rect 670620 224498 670626 224500
rect 671475 224498 671541 224501
rect 672073 224498 672139 224501
rect 670509 224440 670514 224496
rect 670509 224436 670556 224440
rect 670620 224438 670666 224498
rect 671475 224496 672139 224498
rect 671475 224440 671480 224496
rect 671536 224440 672078 224496
rect 672134 224440 672139 224496
rect 671475 224438 672139 224440
rect 670620 224436 670626 224438
rect 670509 224435 670575 224436
rect 671475 224435 671541 224438
rect 672073 224435 672139 224438
rect 138013 224362 138079 224365
rect 152365 224362 152431 224365
rect 138013 224360 152431 224362
rect 138013 224304 138018 224360
rect 138074 224304 152370 224360
rect 152426 224304 152431 224360
rect 138013 224302 152431 224304
rect 138013 224299 138079 224302
rect 152365 224299 152431 224302
rect 671589 224226 671655 224229
rect 663750 224224 671655 224226
rect 663750 224168 671594 224224
rect 671650 224168 671655 224224
rect 663750 224166 671655 224168
rect 137277 224090 137343 224093
rect 138105 224090 138171 224093
rect 137277 224088 138171 224090
rect 137277 224032 137282 224088
rect 137338 224032 138110 224088
rect 138166 224032 138171 224088
rect 137277 224030 138171 224032
rect 137277 224027 137343 224030
rect 138105 224027 138171 224030
rect 654777 223954 654843 223957
rect 663750 223954 663810 224166
rect 671589 224163 671655 224166
rect 654777 223952 663810 223954
rect 654777 223896 654782 223952
rect 654838 223896 663810 223952
rect 654777 223894 663810 223896
rect 669681 223954 669747 223957
rect 671613 223956 671679 223957
rect 669998 223954 670004 223956
rect 669681 223952 670004 223954
rect 669681 223896 669686 223952
rect 669742 223896 670004 223952
rect 669681 223894 670004 223896
rect 654777 223891 654843 223894
rect 669681 223891 669747 223894
rect 669998 223892 670004 223894
rect 670068 223892 670074 223956
rect 671613 223952 671660 223956
rect 671724 223954 671730 223956
rect 671613 223896 671618 223952
rect 671613 223892 671660 223896
rect 671724 223894 671770 223954
rect 671724 223892 671730 223894
rect 671613 223891 671679 223892
rect 678237 223818 678303 223821
rect 678237 223816 678346 223818
rect 678237 223760 678242 223816
rect 678298 223760 678346 223816
rect 678237 223755 678346 223760
rect 657537 223682 657603 223685
rect 670509 223682 670575 223685
rect 657537 223680 670575 223682
rect 657537 223624 657542 223680
rect 657598 223624 670514 223680
rect 670570 223624 670575 223680
rect 657537 223622 670575 223624
rect 657537 223619 657603 223622
rect 670509 223619 670575 223622
rect 42425 223546 42491 223549
rect 46933 223546 46999 223549
rect 51717 223546 51783 223549
rect 42425 223544 46999 223546
rect 42425 223488 42430 223544
rect 42486 223488 46938 223544
rect 46994 223488 46999 223544
rect 42425 223486 46999 223488
rect 42425 223483 42491 223486
rect 46933 223483 46999 223486
rect 51030 223544 51783 223546
rect 51030 223488 51722 223544
rect 51778 223488 51783 223544
rect 51030 223486 51783 223488
rect 42149 223274 42215 223277
rect 51030 223274 51090 223486
rect 51717 223483 51783 223486
rect 63401 223546 63467 223549
rect 591982 223546 591988 223548
rect 63401 223544 591988 223546
rect 63401 223488 63406 223544
rect 63462 223488 591988 223544
rect 63401 223486 591988 223488
rect 63401 223483 63467 223486
rect 591982 223484 591988 223486
rect 592052 223484 592058 223548
rect 678286 223516 678346 223755
rect 42149 223272 51090 223274
rect 42149 223216 42154 223272
rect 42210 223216 51090 223272
rect 42149 223214 51090 223216
rect 42149 223211 42215 223214
rect 142521 223138 142587 223141
rect 143625 223138 143691 223141
rect 683297 223138 683363 223141
rect 142521 223136 143691 223138
rect 142521 223080 142526 223136
rect 142582 223080 143630 223136
rect 143686 223080 143691 223136
rect 142521 223078 143691 223080
rect 683284 223136 683363 223138
rect 683284 223080 683302 223136
rect 683358 223080 683363 223136
rect 683284 223078 683363 223080
rect 142521 223075 142587 223078
rect 143625 223075 143691 223078
rect 683297 223075 683363 223078
rect 649574 222940 649580 223004
rect 649644 223002 649650 223004
rect 651966 223002 651972 223004
rect 649644 222942 651972 223002
rect 649644 222940 649650 222942
rect 651966 222940 651972 222942
rect 652036 222940 652042 223004
rect 139853 222866 139919 222869
rect 143809 222866 143875 222869
rect 139853 222864 143875 222866
rect 139853 222808 139858 222864
rect 139914 222808 143814 222864
rect 143870 222808 143875 222864
rect 139853 222806 143875 222808
rect 139853 222803 139919 222806
rect 143809 222803 143875 222806
rect 653397 222866 653463 222869
rect 665817 222866 665883 222869
rect 670509 222866 670575 222869
rect 653397 222864 663810 222866
rect 653397 222808 653402 222864
rect 653458 222808 663810 222864
rect 653397 222806 663810 222808
rect 653397 222803 653463 222806
rect 663750 222594 663810 222806
rect 665817 222864 670575 222866
rect 665817 222808 665822 222864
rect 665878 222808 670514 222864
rect 670570 222808 670575 222864
rect 665817 222806 670575 222808
rect 665817 222803 665883 222806
rect 670509 222803 670575 222806
rect 683113 222730 683179 222733
rect 683100 222728 683179 222730
rect 683100 222672 683118 222728
rect 683174 222672 683179 222728
rect 683100 222670 683179 222672
rect 683113 222667 683179 222670
rect 673269 222594 673335 222597
rect 663750 222592 673335 222594
rect 663750 222536 673274 222592
rect 673330 222536 673335 222592
rect 663750 222534 673335 222536
rect 673269 222531 673335 222534
rect 669773 222322 669839 222325
rect 669998 222322 670004 222324
rect 669773 222320 670004 222322
rect 669773 222264 669778 222320
rect 669834 222264 670004 222320
rect 669773 222262 670004 222264
rect 669773 222259 669839 222262
rect 669998 222260 670004 222262
rect 670068 222260 670074 222324
rect 674557 222322 674623 222325
rect 674557 222320 676292 222322
rect 674557 222264 674562 222320
rect 674618 222264 676292 222320
rect 674557 222262 676292 222264
rect 674557 222259 674623 222262
rect 535729 222050 535795 222053
rect 539777 222050 539843 222053
rect 535729 222048 539843 222050
rect 535729 221992 535734 222048
rect 535790 221992 539782 222048
rect 539838 221992 539843 222048
rect 535729 221990 539843 221992
rect 535729 221987 535795 221990
rect 539777 221987 539843 221990
rect 173341 221914 173407 221917
rect 177389 221914 177455 221917
rect 173341 221912 177455 221914
rect 173341 221856 173346 221912
rect 173402 221856 177394 221912
rect 177450 221856 177455 221912
rect 173341 221854 177455 221856
rect 173341 221851 173407 221854
rect 177389 221851 177455 221854
rect 553945 221914 554011 221917
rect 558545 221914 558611 221917
rect 553945 221912 558611 221914
rect 553945 221856 553950 221912
rect 554006 221856 558550 221912
rect 558606 221856 558611 221912
rect 553945 221854 558611 221856
rect 553945 221851 554011 221854
rect 558545 221851 558611 221854
rect 559373 221914 559439 221917
rect 561489 221914 561555 221917
rect 559373 221912 561555 221914
rect 559373 221856 559378 221912
rect 559434 221856 561494 221912
rect 561550 221856 561555 221912
rect 559373 221854 561555 221856
rect 559373 221851 559439 221854
rect 561489 221851 561555 221854
rect 676029 221914 676095 221917
rect 676029 221912 676292 221914
rect 676029 221856 676034 221912
rect 676090 221856 676292 221912
rect 676029 221854 676292 221856
rect 676029 221851 676095 221854
rect 161427 221778 161493 221781
rect 167637 221778 167703 221781
rect 161427 221776 167703 221778
rect 161427 221720 161432 221776
rect 161488 221720 167642 221776
rect 167698 221720 167703 221776
rect 161427 221718 167703 221720
rect 161427 221715 161493 221718
rect 167637 221715 167703 221718
rect 547827 221778 547893 221781
rect 549253 221778 549319 221781
rect 547827 221776 549319 221778
rect 547827 221720 547832 221776
rect 547888 221720 549258 221776
rect 549314 221720 549319 221776
rect 547827 221718 549319 221720
rect 547827 221715 547893 221718
rect 549253 221715 549319 221718
rect 563789 221778 563855 221781
rect 572621 221778 572687 221781
rect 563789 221776 572687 221778
rect 563789 221720 563794 221776
rect 563850 221720 572626 221776
rect 572682 221720 572687 221776
rect 563789 221718 572687 221720
rect 563789 221715 563855 221718
rect 572621 221715 572687 221718
rect 660757 221778 660823 221781
rect 674833 221778 674899 221781
rect 660757 221776 674899 221778
rect 660757 221720 660762 221776
rect 660818 221720 674838 221776
rect 674894 221720 674899 221776
rect 660757 221718 674899 221720
rect 660757 221715 660823 221718
rect 674833 221715 674899 221718
rect 138473 221642 138539 221645
rect 141509 221642 141575 221645
rect 138473 221640 141575 221642
rect 138473 221584 138478 221640
rect 138534 221584 141514 221640
rect 141570 221584 141575 221640
rect 138473 221582 141575 221584
rect 138473 221579 138539 221582
rect 141509 221579 141575 221582
rect 142061 221642 142127 221645
rect 147581 221642 147647 221645
rect 142061 221640 147647 221642
rect 142061 221584 142066 221640
rect 142122 221584 147586 221640
rect 147642 221584 147647 221640
rect 142061 221582 147647 221584
rect 142061 221579 142127 221582
rect 147581 221579 147647 221582
rect 513557 221506 513623 221509
rect 599485 221506 599551 221509
rect 513557 221504 599551 221506
rect 513557 221448 513562 221504
rect 513618 221448 599490 221504
rect 599546 221448 599551 221504
rect 513557 221446 599551 221448
rect 513557 221443 513623 221446
rect 599485 221443 599551 221446
rect 651465 221506 651531 221509
rect 668577 221506 668643 221509
rect 651465 221504 668643 221506
rect 651465 221448 651470 221504
rect 651526 221448 668582 221504
rect 668638 221448 668643 221504
rect 651465 221446 668643 221448
rect 651465 221443 651531 221446
rect 668577 221443 668643 221446
rect 675017 221506 675083 221509
rect 675017 221504 676292 221506
rect 675017 221448 675022 221504
rect 675078 221448 676292 221504
rect 675017 221446 676292 221448
rect 675017 221443 675083 221446
rect 515765 221234 515831 221237
rect 600681 221234 600747 221237
rect 515765 221232 600747 221234
rect 515765 221176 515770 221232
rect 515826 221176 600686 221232
rect 600742 221176 600747 221232
rect 515765 221174 600747 221176
rect 515765 221171 515831 221174
rect 600681 221171 600747 221174
rect 673269 221098 673335 221101
rect 673269 221096 676292 221098
rect 673269 221040 673274 221096
rect 673330 221040 676292 221096
rect 673269 221038 676292 221040
rect 673269 221035 673335 221038
rect 158345 220962 158411 220965
rect 161565 220962 161631 220965
rect 158345 220960 161631 220962
rect 158345 220904 158350 220960
rect 158406 220904 161570 220960
rect 161626 220904 161631 220960
rect 158345 220902 161631 220904
rect 158345 220899 158411 220902
rect 161565 220899 161631 220902
rect 180793 220962 180859 220965
rect 185117 220962 185183 220965
rect 180793 220960 185183 220962
rect 180793 220904 180798 220960
rect 180854 220904 185122 220960
rect 185178 220904 185183 220960
rect 180793 220902 185183 220904
rect 180793 220899 180859 220902
rect 185117 220899 185183 220902
rect 522573 220962 522639 220965
rect 618253 220962 618319 220965
rect 522573 220960 618319 220962
rect 522573 220904 522578 220960
rect 522634 220904 618258 220960
rect 618314 220904 618319 220960
rect 522573 220902 618319 220904
rect 522573 220899 522639 220902
rect 618253 220899 618319 220902
rect 147213 220826 147279 220829
rect 151169 220826 151235 220829
rect 147213 220824 151235 220826
rect 147213 220768 147218 220824
rect 147274 220768 151174 220824
rect 151230 220768 151235 220824
rect 147213 220766 151235 220768
rect 147213 220763 147279 220766
rect 151169 220763 151235 220766
rect 185945 220826 186011 220829
rect 190545 220826 190611 220829
rect 185945 220824 190611 220826
rect 185945 220768 185950 220824
rect 186006 220768 190550 220824
rect 190606 220768 190611 220824
rect 185945 220766 190611 220768
rect 185945 220763 186011 220766
rect 190545 220763 190611 220766
rect 176285 220690 176351 220693
rect 180885 220690 180951 220693
rect 176285 220688 180951 220690
rect 176285 220632 176290 220688
rect 176346 220632 180890 220688
rect 180946 220632 180951 220688
rect 176285 220630 180951 220632
rect 176285 220627 176351 220630
rect 180885 220627 180951 220630
rect 565629 220690 565695 220693
rect 569953 220690 570019 220693
rect 565629 220688 570019 220690
rect 565629 220632 565634 220688
rect 565690 220632 569958 220688
rect 570014 220632 570019 220688
rect 565629 220630 570019 220632
rect 565629 220627 565695 220630
rect 569953 220627 570019 220630
rect 673085 220690 673151 220693
rect 673085 220688 676292 220690
rect 673085 220632 673090 220688
rect 673146 220632 676292 220688
rect 673085 220630 676292 220632
rect 673085 220627 673151 220630
rect 150709 220554 150775 220557
rect 151905 220554 151971 220557
rect 150709 220552 151971 220554
rect 150709 220496 150714 220552
rect 150770 220496 151910 220552
rect 151966 220496 151971 220552
rect 150709 220494 151971 220496
rect 150709 220491 150775 220494
rect 151905 220491 151971 220494
rect 557993 220554 558059 220557
rect 558729 220554 558795 220557
rect 557993 220552 558795 220554
rect 557993 220496 557998 220552
rect 558054 220496 558734 220552
rect 558790 220496 558795 220552
rect 557993 220494 558795 220496
rect 557993 220491 558059 220494
rect 558729 220491 558795 220494
rect 562869 220554 562935 220557
rect 563329 220554 563395 220557
rect 562869 220552 563395 220554
rect 562869 220496 562874 220552
rect 562930 220496 563334 220552
rect 563390 220496 563395 220552
rect 562869 220494 563395 220496
rect 562869 220491 562935 220494
rect 563329 220491 563395 220494
rect 572253 220556 572319 220557
rect 572253 220552 572300 220556
rect 572364 220554 572370 220556
rect 572253 220496 572258 220552
rect 572253 220492 572300 220496
rect 572364 220494 572410 220554
rect 572364 220492 572370 220494
rect 572253 220491 572319 220492
rect 147213 220418 147279 220421
rect 148317 220418 148383 220421
rect 147213 220416 148383 220418
rect 147213 220360 147218 220416
rect 147274 220360 148322 220416
rect 148378 220360 148383 220416
rect 147213 220358 148383 220360
rect 147213 220355 147279 220358
rect 148317 220355 148383 220358
rect 654133 220418 654199 220421
rect 669221 220418 669287 220421
rect 654133 220416 669287 220418
rect 654133 220360 654138 220416
rect 654194 220360 669226 220416
rect 669282 220360 669287 220416
rect 654133 220358 669287 220360
rect 654133 220355 654199 220358
rect 669221 220355 669287 220358
rect 151721 220282 151787 220285
rect 154389 220282 154455 220285
rect 151721 220280 154455 220282
rect 151721 220224 151726 220280
rect 151782 220224 154394 220280
rect 154450 220224 154455 220280
rect 151721 220222 154455 220224
rect 151721 220219 151787 220222
rect 154389 220219 154455 220222
rect 486969 220282 487035 220285
rect 611629 220282 611695 220285
rect 486969 220280 611695 220282
rect 486969 220224 486974 220280
rect 487030 220224 611634 220280
rect 611690 220224 611695 220280
rect 486969 220222 611695 220224
rect 486969 220219 487035 220222
rect 611629 220219 611695 220222
rect 672533 220282 672599 220285
rect 672533 220280 676292 220282
rect 672533 220224 672538 220280
rect 672594 220224 676292 220280
rect 672533 220222 676292 220224
rect 672533 220219 672599 220222
rect 669313 220148 669379 220149
rect 669262 220084 669268 220148
rect 669332 220146 669379 220148
rect 669332 220144 669424 220146
rect 669374 220088 669424 220144
rect 669332 220086 669424 220088
rect 669332 220084 669379 220086
rect 669313 220083 669379 220084
rect 515121 220010 515187 220013
rect 617149 220010 617215 220013
rect 515121 220008 617215 220010
rect 515121 219952 515126 220008
rect 515182 219952 617154 220008
rect 617210 219952 617215 220008
rect 515121 219950 617215 219952
rect 515121 219947 515187 219950
rect 617149 219947 617215 219950
rect 645853 219874 645919 219877
rect 675201 219874 675267 219877
rect 645853 219872 675267 219874
rect 645853 219816 645858 219872
rect 645914 219816 675206 219872
rect 675262 219816 675267 219872
rect 645853 219814 675267 219816
rect 645853 219811 645919 219814
rect 675201 219811 675267 219814
rect 676024 219812 676030 219876
rect 676094 219874 676100 219876
rect 676094 219814 676292 219874
rect 676094 219812 676100 219814
rect 492949 219738 493015 219741
rect 493685 219738 493751 219741
rect 612917 219738 612983 219741
rect 492949 219736 612983 219738
rect 492949 219680 492954 219736
rect 493010 219680 493690 219736
rect 493746 219680 612922 219736
rect 612978 219680 612983 219736
rect 492949 219678 612983 219680
rect 492949 219675 493015 219678
rect 493685 219675 493751 219678
rect 612917 219675 612983 219678
rect 520181 219466 520247 219469
rect 618437 219466 618503 219469
rect 520181 219464 618503 219466
rect 520181 219408 520186 219464
rect 520242 219408 618442 219464
rect 618498 219408 618503 219464
rect 520181 219406 618503 219408
rect 520181 219403 520247 219406
rect 618437 219403 618503 219406
rect 666645 219466 666711 219469
rect 666645 219464 676292 219466
rect 666645 219408 666650 219464
rect 666706 219408 676292 219464
rect 666645 219406 676292 219408
rect 666645 219403 666711 219406
rect 136173 219330 136239 219333
rect 137277 219330 137343 219333
rect 136173 219328 137343 219330
rect 136173 219272 136178 219328
rect 136234 219272 137282 219328
rect 137338 219272 137343 219328
rect 136173 219270 137343 219272
rect 136173 219267 136239 219270
rect 137277 219267 137343 219270
rect 170949 219330 171015 219333
rect 171777 219330 171843 219333
rect 170949 219328 171843 219330
rect 170949 219272 170954 219328
rect 171010 219272 171782 219328
rect 171838 219272 171843 219328
rect 170949 219270 171843 219272
rect 170949 219267 171015 219270
rect 171777 219267 171843 219270
rect 562869 219194 562935 219197
rect 563513 219194 563579 219197
rect 562869 219192 563579 219194
rect 562869 219136 562874 219192
rect 562930 219136 563518 219192
rect 563574 219136 563579 219192
rect 562869 219134 563579 219136
rect 562869 219131 562935 219134
rect 563513 219131 563579 219134
rect 572069 219194 572135 219197
rect 574553 219194 574619 219197
rect 572069 219192 574619 219194
rect 572069 219136 572074 219192
rect 572130 219136 574558 219192
rect 574614 219136 574619 219192
rect 572069 219134 574619 219136
rect 572069 219131 572135 219134
rect 574553 219131 574619 219134
rect 674833 219058 674899 219061
rect 674833 219056 676292 219058
rect 674833 219000 674838 219056
rect 674894 219000 676292 219056
rect 674833 218998 676292 219000
rect 674833 218995 674899 218998
rect 563421 218922 563487 218925
rect 564157 218922 564223 218925
rect 563421 218920 564223 218922
rect 563421 218864 563426 218920
rect 563482 218864 564162 218920
rect 564218 218864 564223 218920
rect 563421 218862 564223 218864
rect 563421 218859 563487 218862
rect 564157 218859 564223 218862
rect 564801 218922 564867 218925
rect 574737 218922 574803 218925
rect 564801 218920 574803 218922
rect 564801 218864 564806 218920
rect 564862 218864 574742 218920
rect 574798 218864 574803 218920
rect 564801 218862 574803 218864
rect 564801 218859 564867 218862
rect 574737 218859 574803 218862
rect 656801 218922 656867 218925
rect 670509 218922 670575 218925
rect 656801 218920 670575 218922
rect 656801 218864 656806 218920
rect 656862 218864 670514 218920
rect 670570 218864 670575 218920
rect 656801 218862 670575 218864
rect 656801 218859 656867 218862
rect 670509 218859 670575 218862
rect 675477 218786 675543 218789
rect 672168 218784 675543 218786
rect 672168 218728 675482 218784
rect 675538 218728 675543 218784
rect 672168 218726 675543 218728
rect 154481 218650 154547 218653
rect 160185 218650 160251 218653
rect 154481 218648 160251 218650
rect 154481 218592 154486 218648
rect 154542 218592 160190 218648
rect 160246 218592 160251 218648
rect 154481 218590 160251 218592
rect 154481 218587 154547 218590
rect 160185 218587 160251 218590
rect 563053 218650 563119 218653
rect 574737 218650 574803 218653
rect 563053 218648 574803 218650
rect 563053 218592 563058 218648
rect 563114 218592 574742 218648
rect 574798 218592 574803 218648
rect 563053 218590 574803 218592
rect 563053 218587 563119 218590
rect 574737 218587 574803 218590
rect 648429 218650 648495 218653
rect 672168 218650 672228 218726
rect 675477 218723 675543 218726
rect 648429 218648 672228 218650
rect 648429 218592 648434 218648
rect 648490 218592 672228 218648
rect 648429 218590 672228 218592
rect 648429 218587 648495 218590
rect 675702 218588 675708 218652
rect 675772 218650 675778 218652
rect 675772 218590 676292 218650
rect 675772 218588 675778 218590
rect 494697 218378 494763 218381
rect 630673 218378 630739 218381
rect 494697 218376 630739 218378
rect 494697 218320 494702 218376
rect 494758 218320 630678 218376
rect 630734 218320 630739 218376
rect 494697 218318 630739 218320
rect 494697 218315 494763 218318
rect 630673 218315 630739 218318
rect 669313 218242 669379 218245
rect 669630 218242 669636 218244
rect 669313 218240 669636 218242
rect 669313 218184 669318 218240
rect 669374 218184 669636 218240
rect 669313 218182 669636 218184
rect 669313 218179 669379 218182
rect 669630 218180 669636 218182
rect 669700 218180 669706 218244
rect 675569 218242 675635 218245
rect 675569 218240 676292 218242
rect 675569 218184 675574 218240
rect 675630 218184 676292 218240
rect 675569 218182 676292 218184
rect 675569 218179 675635 218182
rect 487797 218106 487863 218109
rect 623957 218106 624023 218109
rect 487797 218104 624023 218106
rect 487797 218048 487802 218104
rect 487858 218048 623962 218104
rect 624018 218048 624023 218104
rect 487797 218046 624023 218048
rect 487797 218043 487863 218046
rect 623957 218043 624023 218046
rect 35801 217970 35867 217973
rect 54477 217970 54543 217973
rect 670550 217970 670556 217972
rect 35801 217968 54543 217970
rect 35801 217912 35806 217968
rect 35862 217912 54482 217968
rect 54538 217912 54543 217968
rect 35801 217910 54543 217912
rect 35801 217907 35867 217910
rect 54477 217907 54543 217910
rect 663750 217910 670556 217970
rect 562869 217834 562935 217837
rect 568297 217834 568363 217837
rect 562869 217832 568363 217834
rect 562869 217776 562874 217832
rect 562930 217776 568302 217832
rect 568358 217776 568363 217832
rect 562869 217774 568363 217776
rect 562869 217771 562935 217774
rect 568297 217771 568363 217774
rect 572069 217834 572135 217837
rect 574921 217834 574987 217837
rect 572069 217832 574987 217834
rect 572069 217776 572074 217832
rect 572130 217776 574926 217832
rect 574982 217776 574987 217832
rect 572069 217774 574987 217776
rect 572069 217771 572135 217774
rect 574921 217771 574987 217774
rect 651097 217834 651163 217837
rect 663750 217834 663810 217910
rect 670550 217908 670556 217910
rect 670620 217908 670626 217972
rect 675886 217908 675892 217972
rect 675956 217970 675962 217972
rect 675956 217910 676230 217970
rect 675956 217908 675962 217910
rect 651097 217832 663810 217834
rect 651097 217776 651102 217832
rect 651158 217776 663810 217832
rect 651097 217774 663810 217776
rect 676170 217834 676230 217910
rect 676170 217774 676292 217834
rect 651097 217771 651163 217774
rect 673913 217698 673979 217701
rect 676029 217698 676095 217701
rect 673913 217696 676095 217698
rect 673913 217640 673918 217696
rect 673974 217640 676034 217696
rect 676090 217640 676095 217696
rect 673913 217638 676095 217640
rect 673913 217635 673979 217638
rect 676029 217635 676095 217638
rect 510981 217564 511047 217565
rect 519997 217564 520063 217565
rect 510981 217562 511028 217564
rect 510936 217560 511028 217562
rect 510936 217504 510986 217560
rect 510936 217502 511028 217504
rect 510981 217500 511028 217502
rect 511092 217500 511098 217564
rect 519997 217562 520044 217564
rect 519952 217560 520044 217562
rect 519952 217504 520002 217560
rect 519952 217502 520044 217504
rect 519997 217500 520044 217502
rect 520108 217500 520114 217564
rect 531497 217562 531563 217565
rect 532509 217564 532575 217565
rect 532509 217562 532556 217564
rect 531497 217560 532556 217562
rect 531497 217504 531502 217560
rect 531558 217504 532514 217560
rect 531497 217502 532556 217504
rect 510981 217499 511047 217500
rect 519997 217499 520063 217500
rect 531497 217499 531563 217502
rect 532509 217500 532556 217502
rect 532620 217500 532626 217564
rect 560753 217562 560819 217565
rect 563145 217562 563211 217565
rect 572253 217564 572319 217565
rect 572253 217562 572300 217564
rect 560753 217560 563211 217562
rect 560753 217504 560758 217560
rect 560814 217504 563150 217560
rect 563206 217504 563211 217560
rect 560753 217502 563211 217504
rect 572208 217560 572300 217562
rect 572208 217504 572258 217560
rect 572208 217502 572300 217504
rect 532509 217499 532575 217500
rect 560753 217499 560819 217502
rect 563145 217499 563211 217502
rect 572253 217500 572300 217502
rect 572364 217500 572370 217564
rect 572897 217562 572963 217565
rect 574185 217562 574251 217565
rect 572897 217560 574251 217562
rect 572897 217504 572902 217560
rect 572958 217504 574190 217560
rect 574246 217504 574251 217560
rect 572897 217502 574251 217504
rect 572253 217499 572319 217500
rect 572897 217499 572963 217502
rect 574185 217499 574251 217502
rect 653765 217562 653831 217565
rect 672073 217562 672139 217565
rect 653765 217560 672139 217562
rect 653765 217504 653770 217560
rect 653826 217504 672078 217560
rect 672134 217504 672139 217560
rect 653765 217502 672139 217504
rect 653765 217499 653831 217502
rect 672073 217499 672139 217502
rect 676170 217366 676292 217426
rect 502241 217290 502307 217293
rect 595161 217290 595227 217293
rect 502241 217288 595227 217290
rect 502241 217232 502246 217288
rect 502302 217232 595166 217288
rect 595222 217232 595227 217288
rect 502241 217230 595227 217232
rect 502241 217227 502307 217230
rect 595161 217227 595227 217230
rect 671981 217290 672047 217293
rect 676170 217290 676230 217366
rect 671981 217288 676230 217290
rect 671981 217232 671986 217288
rect 672042 217232 676230 217288
rect 671981 217230 676230 217232
rect 671981 217227 672047 217230
rect 488809 217154 488875 217157
rect 495157 217154 495223 217157
rect 488809 217152 491034 217154
rect 488809 217096 488814 217152
rect 488870 217096 491034 217152
rect 488809 217094 491034 217096
rect 488809 217091 488875 217094
rect 490974 216746 491034 217094
rect 495157 217152 499590 217154
rect 495157 217096 495162 217152
rect 495218 217096 499590 217152
rect 495157 217094 499590 217096
rect 495157 217091 495223 217094
rect 499530 217018 499590 217094
rect 595713 217018 595779 217021
rect 499530 217016 595779 217018
rect 499530 216960 595718 217016
rect 595774 216960 595779 217016
rect 499530 216958 595779 216960
rect 595713 216955 595779 216958
rect 669221 217018 669287 217021
rect 669221 217016 676292 217018
rect 669221 216960 669226 217016
rect 669282 216960 676292 217016
rect 669221 216958 676292 216960
rect 669221 216955 669287 216958
rect 575473 216746 575539 216749
rect 490974 216744 575539 216746
rect 490974 216688 575478 216744
rect 575534 216688 575539 216744
rect 490974 216686 575539 216688
rect 575473 216683 575539 216686
rect 670509 216746 670575 216749
rect 671981 216746 672047 216749
rect 670509 216744 672047 216746
rect 670509 216688 670514 216744
rect 670570 216688 671986 216744
rect 672042 216688 672047 216744
rect 670509 216686 672047 216688
rect 670509 216683 670575 216686
rect 671981 216683 672047 216686
rect 672533 216746 672599 216749
rect 676029 216746 676095 216749
rect 672533 216744 676095 216746
rect 672533 216688 672538 216744
rect 672594 216688 676034 216744
rect 676090 216688 676095 216744
rect 672533 216686 676095 216688
rect 672533 216683 672599 216686
rect 676029 216683 676095 216686
rect 676170 216550 676292 216610
rect 673453 216474 673519 216477
rect 676170 216474 676230 216550
rect 673453 216472 676230 216474
rect 673453 216416 673458 216472
rect 673514 216416 676230 216472
rect 673453 216414 676230 216416
rect 673453 216411 673519 216414
rect 673085 216202 673151 216205
rect 673085 216200 676292 216202
rect 673085 216144 673090 216200
rect 673146 216144 676292 216200
rect 673085 216142 676292 216144
rect 673085 216139 673151 216142
rect 672073 216066 672139 216069
rect 669270 216064 672139 216066
rect 669270 216008 672078 216064
rect 672134 216008 672139 216064
rect 669270 216006 672139 216008
rect 520038 215868 520044 215932
rect 520108 215930 520114 215932
rect 617793 215930 617859 215933
rect 669270 215930 669330 216006
rect 672073 216003 672139 216006
rect 520108 215928 617859 215930
rect 520108 215872 617798 215928
rect 617854 215872 617859 215928
rect 520108 215870 617859 215872
rect 520108 215868 520114 215870
rect 617793 215867 617859 215870
rect 663750 215870 669330 215930
rect 511022 215596 511028 215660
rect 511092 215658 511098 215660
rect 599025 215658 599091 215661
rect 511092 215656 599091 215658
rect 511092 215600 599030 215656
rect 599086 215600 599091 215656
rect 511092 215598 599091 215600
rect 511092 215596 511098 215598
rect 599025 215595 599091 215598
rect 532550 215324 532556 215388
rect 532620 215386 532626 215388
rect 621105 215386 621171 215389
rect 532620 215384 621171 215386
rect 532620 215328 621110 215384
rect 621166 215328 621171 215384
rect 532620 215326 621171 215328
rect 532620 215324 532626 215326
rect 621105 215323 621171 215326
rect 659561 215386 659627 215389
rect 663750 215386 663810 215870
rect 669822 215734 676292 215794
rect 664621 215658 664687 215661
rect 668393 215658 668459 215661
rect 664621 215656 668459 215658
rect 664621 215600 664626 215656
rect 664682 215600 668398 215656
rect 668454 215600 668459 215656
rect 664621 215598 668459 215600
rect 664621 215595 664687 215598
rect 668393 215595 668459 215598
rect 659561 215384 663810 215386
rect 659561 215328 659566 215384
rect 659622 215328 663810 215384
rect 659561 215326 663810 215328
rect 666829 215386 666895 215389
rect 669822 215386 669882 215734
rect 675886 215460 675892 215524
rect 675956 215522 675962 215524
rect 675956 215462 676230 215522
rect 675956 215460 675962 215462
rect 666829 215384 669146 215386
rect 666829 215328 666834 215384
rect 666890 215328 669146 215384
rect 666829 215326 669146 215328
rect 659561 215323 659627 215326
rect 666829 215323 666895 215326
rect 53281 215114 53347 215117
rect 41462 215112 53347 215114
rect 41462 215056 53286 215112
rect 53342 215056 53347 215112
rect 41462 215054 53347 215056
rect 669086 215114 669146 215326
rect 669638 215326 669882 215386
rect 672073 215386 672139 215389
rect 675753 215386 675819 215389
rect 672073 215384 675819 215386
rect 672073 215328 672078 215384
rect 672134 215328 675758 215384
rect 675814 215328 675819 215384
rect 672073 215326 675819 215328
rect 676170 215386 676230 215462
rect 676170 215326 676292 215386
rect 669638 215114 669698 215326
rect 672073 215323 672139 215326
rect 675753 215323 675819 215326
rect 669086 215054 669698 215114
rect 41462 214948 41522 215054
rect 53281 215051 53347 215054
rect 674465 214978 674531 214981
rect 674465 214976 676292 214978
rect 674465 214920 674470 214976
rect 674526 214920 676292 214976
rect 674465 214918 676292 214920
rect 674465 214915 674531 214918
rect 35801 214706 35867 214709
rect 675845 214706 675911 214709
rect 35758 214704 35867 214706
rect 35758 214648 35806 214704
rect 35862 214648 35867 214704
rect 35758 214643 35867 214648
rect 663750 214704 675911 214706
rect 663750 214648 675850 214704
rect 675906 214648 675911 214704
rect 663750 214646 675911 214648
rect 35758 214540 35818 214643
rect 660389 214570 660455 214573
rect 663750 214570 663810 214646
rect 675845 214643 675911 214646
rect 660389 214568 663810 214570
rect 660389 214512 660394 214568
rect 660450 214512 663810 214568
rect 660389 214510 663810 214512
rect 676029 214570 676095 214573
rect 676029 214568 676292 214570
rect 676029 214512 676034 214568
rect 676090 214512 676292 214568
rect 676029 214510 676292 214512
rect 660389 214507 660455 214510
rect 676029 214507 676095 214510
rect 35801 214298 35867 214301
rect 35758 214296 35867 214298
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 35758 214235 35867 214240
rect 39757 214298 39823 214301
rect 43437 214298 43503 214301
rect 39757 214296 43503 214298
rect 39757 214240 39762 214296
rect 39818 214240 43442 214296
rect 43498 214240 43503 214296
rect 39757 214238 43503 214240
rect 39757 214235 39823 214238
rect 43437 214235 43503 214238
rect 35758 214132 35818 214235
rect 575982 214026 576042 214404
rect 672073 214162 672139 214165
rect 672073 214160 676292 214162
rect 672073 214104 672078 214160
rect 672134 214104 676292 214160
rect 672073 214102 676292 214104
rect 672073 214099 672139 214102
rect 578877 214026 578943 214029
rect 575982 214024 578943 214026
rect 575982 213968 578882 214024
rect 578938 213968 578943 214024
rect 575982 213966 578943 213968
rect 578877 213963 578943 213966
rect 669589 213890 669655 213893
rect 673453 213890 673519 213893
rect 669589 213888 673519 213890
rect 669589 213832 669594 213888
rect 669650 213832 673458 213888
rect 673514 213832 673519 213888
rect 669589 213830 673519 213832
rect 669589 213827 669655 213830
rect 673453 213827 673519 213830
rect 44909 213754 44975 213757
rect 41492 213752 44975 213754
rect 41492 213696 44914 213752
rect 44970 213696 44975 213752
rect 41492 213694 44975 213696
rect 44909 213691 44975 213694
rect 674649 213754 674715 213757
rect 674649 213752 676292 213754
rect 674649 213696 674654 213752
rect 674710 213696 676292 213752
rect 674649 213694 676292 213696
rect 674649 213691 674715 213694
rect 672717 213618 672783 213621
rect 663750 213616 672783 213618
rect 663750 213560 672722 213616
rect 672778 213560 672783 213616
rect 663750 213558 672783 213560
rect 661493 213482 661559 213485
rect 663750 213482 663810 213558
rect 672717 213555 672783 213558
rect 661493 213480 663810 213482
rect 661493 213424 661498 213480
rect 661554 213424 663810 213480
rect 661493 213422 663810 213424
rect 661493 213419 661559 213422
rect 672809 213346 672875 213349
rect 672809 213344 676292 213346
rect 672809 213288 672814 213344
rect 672870 213288 676292 213344
rect 672809 213286 676292 213288
rect 672809 213283 672875 213286
rect 658733 213210 658799 213213
rect 672533 213210 672599 213213
rect 658733 213208 672599 213210
rect 658733 213152 658738 213208
rect 658794 213152 672538 213208
rect 672594 213152 672599 213208
rect 658733 213150 672599 213152
rect 658733 213147 658799 213150
rect 672533 213147 672599 213150
rect 39849 213074 39915 213077
rect 43805 213074 43871 213077
rect 39849 213072 43871 213074
rect 39849 213016 39854 213072
rect 39910 213016 43810 213072
rect 43866 213016 43871 213072
rect 39849 213014 43871 213016
rect 39849 213011 39915 213014
rect 43805 213011 43871 213014
rect 35758 212669 35818 212908
rect 35758 212664 35867 212669
rect 35758 212608 35806 212664
rect 35862 212608 35867 212664
rect 35758 212606 35867 212608
rect 35801 212603 35867 212606
rect 675385 212530 675451 212533
rect 675886 212530 675892 212532
rect 675385 212528 675892 212530
rect 675385 212472 675390 212528
rect 675446 212472 675892 212528
rect 675385 212470 675892 212472
rect 675385 212467 675451 212470
rect 675886 212468 675892 212470
rect 675956 212530 675962 212532
rect 683070 212530 683130 212908
rect 675956 212500 683130 212530
rect 675956 212470 683100 212500
rect 675956 212468 675962 212470
rect 40769 212258 40835 212261
rect 42885 212258 42951 212261
rect 40769 212256 42951 212258
rect 40769 212200 40774 212256
rect 40830 212200 42890 212256
rect 42946 212200 42951 212256
rect 40769 212198 42951 212200
rect 40769 212195 40835 212198
rect 42885 212195 42951 212198
rect 35574 211853 35634 212092
rect 35574 211848 35683 211853
rect 35574 211792 35622 211848
rect 35678 211792 35683 211848
rect 35574 211790 35683 211792
rect 35617 211787 35683 211790
rect 40125 211850 40191 211853
rect 43621 211850 43687 211853
rect 40125 211848 43687 211850
rect 40125 211792 40130 211848
rect 40186 211792 43626 211848
rect 43682 211792 43687 211848
rect 40125 211790 43687 211792
rect 40125 211787 40191 211790
rect 43621 211787 43687 211790
rect 575982 211714 576042 212228
rect 672625 212122 672691 212125
rect 672625 212120 676292 212122
rect 672625 212064 672630 212120
rect 672686 212064 676292 212120
rect 672625 212062 676292 212064
rect 672625 212059 672691 212062
rect 578509 211714 578575 211717
rect 575982 211712 578575 211714
rect 575982 211656 578514 211712
rect 578570 211656 578575 211712
rect 575982 211654 578575 211656
rect 578509 211651 578575 211654
rect 35801 211442 35867 211445
rect 35758 211440 35867 211442
rect 35758 211384 35806 211440
rect 35862 211384 35867 211440
rect 35758 211379 35867 211384
rect 676029 211442 676095 211445
rect 676622 211442 676628 211444
rect 676029 211440 676628 211442
rect 676029 211384 676034 211440
rect 676090 211384 676628 211440
rect 676029 211382 676628 211384
rect 676029 211379 676095 211382
rect 676622 211380 676628 211382
rect 676692 211380 676698 211444
rect 35758 211276 35818 211379
rect 35758 210221 35818 210460
rect 35758 210216 35867 210221
rect 35758 210160 35806 210216
rect 35862 210160 35867 210216
rect 35758 210158 35867 210160
rect 35801 210155 35867 210158
rect 41462 209812 41522 210052
rect 41454 209748 41460 209812
rect 41524 209748 41530 209812
rect 575982 209810 576042 210052
rect 579521 209810 579587 209813
rect 575982 209808 579587 209810
rect 575982 209752 579526 209808
rect 579582 209752 579587 209808
rect 575982 209750 579587 209752
rect 579521 209747 579587 209750
rect 35574 209405 35634 209644
rect 35574 209400 35683 209405
rect 35574 209344 35622 209400
rect 35678 209344 35683 209400
rect 35574 209342 35683 209344
rect 35617 209339 35683 209342
rect 41462 208994 41522 209236
rect 41638 208994 41644 208996
rect 41462 208934 41644 208994
rect 41638 208932 41644 208934
rect 41708 208932 41714 208996
rect 41278 208586 41338 208828
rect 44449 208586 44515 208589
rect 41278 208584 44515 208586
rect 41278 208528 44454 208584
rect 44510 208528 44515 208584
rect 41278 208526 44515 208528
rect 44449 208523 44515 208526
rect 35758 208181 35818 208420
rect 35758 208176 35867 208181
rect 35758 208120 35806 208176
rect 35862 208120 35867 208176
rect 35758 208118 35867 208120
rect 35801 208115 35867 208118
rect 44173 208042 44239 208045
rect 41492 208040 44239 208042
rect 41492 207984 44178 208040
rect 44234 207984 44239 208040
rect 41492 207982 44239 207984
rect 44173 207979 44239 207982
rect 589457 208042 589523 208045
rect 589457 208040 592572 208042
rect 589457 207984 589462 208040
rect 589518 207984 592572 208040
rect 589457 207982 592572 207984
rect 589457 207979 589523 207982
rect 40953 207770 41019 207773
rect 43253 207770 43319 207773
rect 40953 207768 43319 207770
rect 40953 207712 40958 207768
rect 41014 207712 43258 207768
rect 43314 207712 43319 207768
rect 40953 207710 43319 207712
rect 40953 207707 41019 207710
rect 43253 207707 43319 207710
rect 35801 207362 35867 207365
rect 40726 207364 40786 207604
rect 575982 207498 576042 207876
rect 579521 207498 579587 207501
rect 575982 207496 579587 207498
rect 575982 207440 579526 207496
rect 579582 207440 579587 207496
rect 575982 207438 579587 207440
rect 579521 207435 579587 207438
rect 35758 207360 35867 207362
rect 35758 207304 35806 207360
rect 35862 207304 35867 207360
rect 35758 207299 35867 207304
rect 40718 207300 40724 207364
rect 40788 207300 40794 207364
rect 40953 207362 41019 207365
rect 43069 207362 43135 207365
rect 40953 207360 43135 207362
rect 40953 207304 40958 207360
rect 41014 207304 43074 207360
rect 43130 207304 43135 207360
rect 40953 207302 43135 207304
rect 40953 207299 41019 207302
rect 43069 207299 43135 207302
rect 35758 207196 35818 207299
rect 39205 206954 39271 206957
rect 42885 206954 42951 206957
rect 39205 206952 42951 206954
rect 39205 206896 39210 206952
rect 39266 206896 42890 206952
rect 42946 206896 42951 206952
rect 39205 206894 42951 206896
rect 39205 206891 39271 206894
rect 42885 206891 42951 206894
rect 674598 206892 674604 206956
rect 674668 206954 674674 206956
rect 675477 206954 675543 206957
rect 674668 206952 675543 206954
rect 674668 206896 675482 206952
rect 675538 206896 675543 206952
rect 674668 206894 675543 206896
rect 674668 206892 674674 206894
rect 675477 206891 675543 206894
rect 40910 206548 40970 206788
rect 40902 206484 40908 206548
rect 40972 206484 40978 206548
rect 589457 206410 589523 206413
rect 589457 206408 592572 206410
rect 35801 206138 35867 206141
rect 40542 206140 40602 206380
rect 589457 206352 589462 206408
rect 589518 206352 592572 206408
rect 589457 206350 592572 206352
rect 589457 206347 589523 206350
rect 35758 206136 35867 206138
rect 35758 206080 35806 206136
rect 35862 206080 35867 206136
rect 35758 206075 35867 206080
rect 40534 206076 40540 206140
rect 40604 206076 40610 206140
rect 35758 205972 35818 206075
rect 579521 205866 579587 205869
rect 575798 205864 579587 205866
rect 575798 205808 579526 205864
rect 579582 205808 579587 205864
rect 575798 205806 579587 205808
rect 575798 205700 575858 205806
rect 579521 205803 579587 205806
rect 669262 205668 669268 205732
rect 669332 205730 669338 205732
rect 669630 205730 669636 205732
rect 669332 205670 669636 205730
rect 669332 205668 669338 205670
rect 669630 205668 669636 205670
rect 669700 205668 669706 205732
rect 44633 205594 44699 205597
rect 41492 205592 44699 205594
rect 41492 205536 44638 205592
rect 44694 205536 44699 205592
rect 41492 205534 44699 205536
rect 44633 205531 44699 205534
rect 669262 205396 669268 205460
rect 669332 205458 669338 205460
rect 669630 205458 669636 205460
rect 669332 205398 669636 205458
rect 669332 205396 669338 205398
rect 669630 205396 669636 205398
rect 669700 205396 669706 205460
rect 39941 205322 40007 205325
rect 43437 205322 43503 205325
rect 39941 205320 43503 205322
rect 39941 205264 39946 205320
rect 40002 205264 43442 205320
rect 43498 205264 43503 205320
rect 39941 205262 43503 205264
rect 39941 205259 40007 205262
rect 43437 205259 43503 205262
rect 35758 204917 35818 205156
rect 35758 204912 35867 204917
rect 35758 204856 35806 204912
rect 35862 204856 35867 204912
rect 35758 204854 35867 204856
rect 35801 204851 35867 204854
rect 41505 204914 41571 204917
rect 46197 204914 46263 204917
rect 41505 204912 46263 204914
rect 41505 204856 41510 204912
rect 41566 204856 46202 204912
rect 46258 204856 46263 204912
rect 41505 204854 46263 204856
rect 41505 204851 41571 204854
rect 46197 204851 46263 204854
rect 589457 204778 589523 204781
rect 589457 204776 592572 204778
rect 35758 204509 35818 204748
rect 589457 204720 589462 204776
rect 589518 204720 592572 204776
rect 589457 204718 592572 204720
rect 589457 204715 589523 204718
rect 35758 204504 35867 204509
rect 41505 204506 41571 204509
rect 35758 204448 35806 204504
rect 35862 204448 35867 204504
rect 35758 204446 35867 204448
rect 35801 204443 35867 204446
rect 41462 204504 41571 204506
rect 41462 204448 41510 204504
rect 41566 204448 41571 204504
rect 41462 204443 41571 204448
rect 41689 204506 41755 204509
rect 43805 204506 43871 204509
rect 41689 204504 43871 204506
rect 41689 204448 41694 204504
rect 41750 204448 43810 204504
rect 43866 204448 43871 204504
rect 41689 204446 43871 204448
rect 41689 204443 41755 204446
rect 43805 204443 43871 204446
rect 41462 204340 41522 204443
rect 666502 204172 666508 204236
rect 666572 204234 666578 204236
rect 674925 204234 674991 204237
rect 675385 204234 675451 204237
rect 666572 204174 666754 204234
rect 666572 204172 666578 204174
rect 39389 204098 39455 204101
rect 42701 204098 42767 204101
rect 39389 204096 42767 204098
rect 39389 204040 39394 204096
rect 39450 204040 42706 204096
rect 42762 204040 42767 204096
rect 39389 204038 42767 204040
rect 39389 204035 39455 204038
rect 42701 204035 42767 204038
rect 666694 204030 666754 204174
rect 674925 204232 675451 204234
rect 674925 204176 674930 204232
rect 674986 204176 675390 204232
rect 675446 204176 675451 204232
rect 674925 204174 675451 204176
rect 674925 204171 674991 204174
rect 675385 204171 675451 204174
rect 666356 203970 666754 204030
rect 35758 203693 35818 203932
rect 35758 203688 35867 203693
rect 35758 203632 35806 203688
rect 35862 203632 35867 203688
rect 35758 203630 35867 203632
rect 35801 203627 35867 203630
rect 575982 203282 576042 203524
rect 578325 203282 578391 203285
rect 575982 203280 578391 203282
rect 575982 203224 578330 203280
rect 578386 203224 578391 203280
rect 575982 203222 578391 203224
rect 578325 203219 578391 203222
rect 589457 203146 589523 203149
rect 589457 203144 592572 203146
rect 589457 203088 589462 203144
rect 589518 203088 592572 203144
rect 589457 203086 592572 203088
rect 589457 203083 589523 203086
rect 669589 202874 669655 202877
rect 674925 202874 674991 202877
rect 669589 202872 674991 202874
rect 669589 202816 669594 202872
rect 669650 202816 674930 202872
rect 674986 202816 674991 202872
rect 669589 202814 674991 202816
rect 669589 202811 669655 202814
rect 674925 202811 674991 202814
rect 675753 202738 675819 202741
rect 676438 202738 676444 202740
rect 675753 202736 676444 202738
rect 675753 202680 675758 202736
rect 675814 202680 676444 202736
rect 675753 202678 676444 202680
rect 675753 202675 675819 202678
rect 676438 202676 676444 202678
rect 676508 202676 676514 202740
rect 589457 201514 589523 201517
rect 589457 201512 592572 201514
rect 589457 201456 589462 201512
rect 589518 201456 592572 201512
rect 589457 201454 592572 201456
rect 589457 201451 589523 201454
rect 42425 201378 42491 201381
rect 43437 201378 43503 201381
rect 42425 201376 43503 201378
rect 42425 201320 42430 201376
rect 42486 201320 43442 201376
rect 43498 201320 43503 201376
rect 672993 201378 673059 201381
rect 675477 201378 675543 201381
rect 672993 201376 675543 201378
rect 42425 201318 43503 201320
rect 42425 201315 42491 201318
rect 43437 201315 43503 201318
rect 575982 200834 576042 201348
rect 672993 201320 672998 201376
rect 673054 201320 675482 201376
rect 675538 201320 675543 201376
rect 672993 201318 675543 201320
rect 672993 201315 673059 201318
rect 675477 201315 675543 201318
rect 578785 200834 578851 200837
rect 575982 200832 578851 200834
rect 575982 200776 578790 200832
rect 578846 200776 578851 200832
rect 575982 200774 578851 200776
rect 578785 200771 578851 200774
rect 672574 200772 672580 200836
rect 672644 200834 672650 200836
rect 673085 200834 673151 200837
rect 672644 200832 673151 200834
rect 672644 200776 673090 200832
rect 673146 200776 673151 200832
rect 672644 200774 673151 200776
rect 672644 200772 672650 200774
rect 673085 200771 673151 200774
rect 675753 200018 675819 200021
rect 676622 200018 676628 200020
rect 675753 200016 676628 200018
rect 675753 199960 675758 200016
rect 675814 199960 676628 200016
rect 675753 199958 676628 199960
rect 675753 199955 675819 199958
rect 676622 199956 676628 199958
rect 676692 199956 676698 200020
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 672073 199746 672139 199749
rect 674925 199746 674991 199749
rect 672073 199744 674991 199746
rect 672073 199688 672078 199744
rect 672134 199688 674930 199744
rect 674986 199688 674991 199744
rect 672073 199686 674991 199688
rect 672073 199683 672139 199686
rect 674925 199683 674991 199686
rect 668025 199202 668091 199205
rect 666694 199200 668091 199202
rect 575982 198930 576042 199172
rect 666694 199144 668030 199200
rect 668086 199144 668091 199200
rect 666694 199142 668091 199144
rect 666694 199134 666754 199142
rect 668025 199139 668091 199142
rect 666356 199074 666754 199134
rect 579521 198930 579587 198933
rect 575982 198928 579587 198930
rect 575982 198872 579526 198928
rect 579582 198872 579587 198928
rect 575982 198870 579587 198872
rect 579521 198867 579587 198870
rect 668393 198794 668459 198797
rect 670734 198794 670740 198796
rect 668393 198792 670740 198794
rect 668393 198736 668398 198792
rect 668454 198736 670740 198792
rect 668393 198734 670740 198736
rect 668393 198731 668459 198734
rect 670734 198732 670740 198734
rect 670804 198732 670810 198796
rect 666829 198522 666895 198525
rect 675109 198522 675175 198525
rect 666829 198520 675175 198522
rect 666829 198464 666834 198520
rect 666890 198464 675114 198520
rect 675170 198464 675175 198520
rect 666829 198462 675175 198464
rect 666829 198459 666895 198462
rect 675109 198459 675175 198462
rect 590377 198250 590443 198253
rect 670509 198250 670575 198253
rect 675477 198250 675543 198253
rect 590377 198248 592572 198250
rect 590377 198192 590382 198248
rect 590438 198192 592572 198248
rect 590377 198190 592572 198192
rect 670509 198248 675543 198250
rect 670509 198192 670514 198248
rect 670570 198192 675482 198248
rect 675538 198192 675543 198248
rect 670509 198190 675543 198192
rect 590377 198187 590443 198190
rect 670509 198187 670575 198190
rect 675477 198187 675543 198190
rect 673269 197978 673335 197981
rect 676806 197978 676812 197980
rect 673269 197976 676812 197978
rect 673269 197920 673274 197976
rect 673330 197920 676812 197976
rect 673269 197918 676812 197920
rect 673269 197915 673335 197918
rect 676806 197916 676812 197918
rect 676876 197916 676882 197980
rect 39297 197842 39363 197845
rect 41822 197842 41828 197844
rect 39297 197840 41828 197842
rect 39297 197784 39302 197840
rect 39358 197784 41828 197840
rect 39297 197782 41828 197784
rect 39297 197779 39363 197782
rect 41822 197780 41828 197782
rect 41892 197780 41898 197844
rect 674465 197162 674531 197165
rect 675385 197162 675451 197165
rect 674465 197160 675451 197162
rect 674465 197104 674470 197160
rect 674526 197104 675390 197160
rect 675446 197104 675451 197160
rect 674465 197102 675451 197104
rect 674465 197099 674531 197102
rect 675385 197099 675451 197102
rect 575982 196482 576042 196996
rect 589457 196618 589523 196621
rect 589457 196616 592572 196618
rect 589457 196560 589462 196616
rect 589518 196560 592572 196616
rect 589457 196558 592572 196560
rect 589457 196555 589523 196558
rect 578509 196482 578575 196485
rect 575982 196480 578575 196482
rect 575982 196424 578514 196480
rect 578570 196424 578575 196480
rect 575982 196422 578575 196424
rect 578509 196419 578575 196422
rect 669262 196148 669268 196212
rect 669332 196210 669338 196212
rect 669630 196210 669636 196212
rect 669332 196150 669636 196210
rect 669332 196148 669338 196150
rect 669630 196148 669636 196150
rect 669700 196148 669706 196212
rect 669262 195876 669268 195940
rect 669332 195938 669338 195940
rect 669630 195938 669636 195940
rect 669332 195878 669636 195938
rect 669332 195876 669338 195878
rect 669630 195876 669636 195878
rect 669700 195876 669706 195940
rect 41873 195804 41939 195805
rect 41822 195802 41828 195804
rect 41782 195742 41828 195802
rect 41892 195800 41939 195804
rect 41934 195744 41939 195800
rect 41822 195740 41828 195742
rect 41892 195740 41939 195744
rect 41873 195739 41939 195740
rect 41638 195468 41644 195532
rect 41708 195530 41714 195532
rect 42333 195530 42399 195533
rect 41708 195528 42399 195530
rect 41708 195472 42338 195528
rect 42394 195472 42399 195528
rect 41708 195470 42399 195472
rect 41708 195468 41714 195470
rect 42333 195467 42399 195470
rect 41454 195196 41460 195260
rect 41524 195258 41530 195260
rect 41781 195258 41847 195261
rect 41524 195256 41847 195258
rect 41524 195200 41786 195256
rect 41842 195200 41847 195256
rect 41524 195198 41847 195200
rect 41524 195196 41530 195198
rect 41781 195195 41847 195198
rect 40718 194924 40724 194988
rect 40788 194986 40794 194988
rect 42190 194986 42196 194988
rect 40788 194926 42196 194986
rect 40788 194924 40794 194926
rect 42190 194924 42196 194926
rect 42260 194924 42266 194988
rect 579521 194986 579587 194989
rect 575798 194984 579587 194986
rect 575798 194928 579526 194984
rect 579582 194928 579587 194984
rect 575798 194926 579587 194928
rect 575798 194820 575858 194926
rect 579521 194923 579587 194926
rect 589273 194986 589339 194989
rect 589273 194984 592572 194986
rect 589273 194928 589278 194984
rect 589334 194928 592572 194984
rect 589273 194926 592572 194928
rect 589273 194923 589339 194926
rect 675753 194578 675819 194581
rect 676254 194578 676260 194580
rect 675753 194576 676260 194578
rect 675753 194520 675758 194576
rect 675814 194520 676260 194576
rect 675753 194518 676260 194520
rect 675753 194515 675819 194518
rect 676254 194516 676260 194518
rect 676324 194516 676330 194580
rect 669313 194306 669379 194309
rect 666694 194304 669379 194306
rect 666694 194248 669318 194304
rect 669374 194248 669379 194304
rect 666694 194246 669379 194248
rect 666694 194238 666754 194246
rect 669313 194243 669379 194246
rect 666356 194178 666754 194238
rect 40902 193428 40908 193492
rect 40972 193490 40978 193492
rect 41781 193490 41847 193493
rect 40972 193488 41847 193490
rect 40972 193432 41786 193488
rect 41842 193432 41847 193488
rect 40972 193430 41847 193432
rect 40972 193428 40978 193430
rect 41781 193427 41847 193430
rect 589457 193354 589523 193357
rect 589457 193352 592572 193354
rect 589457 193296 589462 193352
rect 589518 193296 592572 193352
rect 589457 193294 592572 193296
rect 589457 193291 589523 193294
rect 42333 193220 42399 193221
rect 42333 193218 42380 193220
rect 42288 193216 42380 193218
rect 42288 193160 42338 193216
rect 42288 193158 42380 193160
rect 42333 193156 42380 193158
rect 42444 193156 42450 193220
rect 675753 193218 675819 193221
rect 676070 193218 676076 193220
rect 675753 193216 676076 193218
rect 675753 193160 675758 193216
rect 675814 193160 676076 193216
rect 675753 193158 676076 193160
rect 42333 193155 42399 193156
rect 675753 193155 675819 193158
rect 676070 193156 676076 193158
rect 676140 193156 676146 193220
rect 40534 192748 40540 192812
rect 40604 192810 40610 192812
rect 42241 192810 42307 192813
rect 40604 192808 42307 192810
rect 40604 192752 42246 192808
rect 42302 192752 42307 192808
rect 40604 192750 42307 192752
rect 40604 192748 40610 192750
rect 42241 192747 42307 192750
rect 675661 192810 675727 192813
rect 675886 192810 675892 192812
rect 675661 192808 675892 192810
rect 675661 192752 675666 192808
rect 675722 192752 675892 192808
rect 675661 192750 675892 192752
rect 675661 192747 675727 192750
rect 675886 192748 675892 192750
rect 675956 192748 675962 192812
rect 575982 192266 576042 192644
rect 579521 192266 579587 192269
rect 575982 192264 579587 192266
rect 575982 192208 579526 192264
rect 579582 192208 579587 192264
rect 575982 192206 579587 192208
rect 579521 192203 579587 192206
rect 589457 191722 589523 191725
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 589457 191659 589523 191662
rect 42057 191586 42123 191589
rect 43805 191586 43871 191589
rect 42057 191584 43871 191586
rect 42057 191528 42062 191584
rect 42118 191528 43810 191584
rect 43866 191528 43871 191584
rect 42057 191526 43871 191528
rect 42057 191523 42123 191526
rect 43805 191523 43871 191526
rect 669129 191586 669195 191589
rect 675385 191586 675451 191589
rect 669129 191584 675451 191586
rect 669129 191528 669134 191584
rect 669190 191528 675390 191584
rect 675446 191528 675451 191584
rect 669129 191526 675451 191528
rect 669129 191523 669195 191526
rect 675385 191523 675451 191526
rect 579521 190770 579587 190773
rect 575798 190768 579587 190770
rect 575798 190712 579526 190768
rect 579582 190712 579587 190768
rect 575798 190710 579587 190712
rect 42425 190498 42491 190501
rect 44633 190498 44699 190501
rect 42425 190496 44699 190498
rect 42425 190440 42430 190496
rect 42486 190440 44638 190496
rect 44694 190440 44699 190496
rect 575798 190468 575858 190710
rect 579521 190707 579587 190710
rect 42425 190438 44699 190440
rect 42425 190435 42491 190438
rect 44633 190435 44699 190438
rect 590561 190090 590627 190093
rect 590561 190088 592572 190090
rect 590561 190032 590566 190088
rect 590622 190032 592572 190088
rect 590561 190030 592572 190032
rect 590561 190027 590627 190030
rect 675150 190028 675156 190092
rect 675220 190090 675226 190092
rect 676029 190090 676095 190093
rect 675220 190088 676095 190090
rect 675220 190032 676034 190088
rect 676090 190032 676095 190088
rect 675220 190030 676095 190032
rect 675220 190028 675226 190030
rect 676029 190027 676095 190030
rect 42425 189954 42491 189957
rect 44449 189954 44515 189957
rect 42425 189952 44515 189954
rect 42425 189896 42430 189952
rect 42486 189896 44454 189952
rect 44510 189896 44515 189952
rect 42425 189894 44515 189896
rect 42425 189891 42491 189894
rect 44449 189891 44515 189894
rect 668945 189410 669011 189413
rect 666694 189408 669011 189410
rect 666694 189352 668950 189408
rect 669006 189352 669011 189408
rect 666694 189350 669011 189352
rect 666694 189342 666754 189350
rect 668945 189347 669011 189350
rect 666356 189282 666754 189342
rect 589641 188458 589707 188461
rect 669129 188458 669195 188461
rect 669446 188458 669452 188460
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 669129 188456 669452 188458
rect 669129 188400 669134 188456
rect 669190 188400 669452 188456
rect 669129 188398 669452 188400
rect 589641 188395 589707 188398
rect 669129 188395 669195 188398
rect 669446 188396 669452 188398
rect 669516 188396 669522 188460
rect 575982 188050 576042 188292
rect 579521 188050 579587 188053
rect 575982 188048 579587 188050
rect 575982 187992 579526 188048
rect 579582 187992 579587 188048
rect 575982 187990 579587 187992
rect 579521 187987 579587 187990
rect 42425 187642 42491 187645
rect 43621 187642 43687 187645
rect 42425 187640 43687 187642
rect 42425 187584 42430 187640
rect 42486 187584 43626 187640
rect 43682 187584 43687 187640
rect 42425 187582 43687 187584
rect 42425 187579 42491 187582
rect 43621 187579 43687 187582
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 42333 186284 42399 186285
rect 42333 186282 42380 186284
rect 42288 186280 42380 186282
rect 42288 186224 42338 186280
rect 42288 186222 42380 186224
rect 42333 186220 42380 186222
rect 42444 186220 42450 186284
rect 579521 186282 579587 186285
rect 575798 186280 579587 186282
rect 575798 186224 579526 186280
rect 579582 186224 579587 186280
rect 575798 186222 579587 186224
rect 42333 186219 42399 186220
rect 575798 186116 575858 186222
rect 579521 186219 579587 186222
rect 42149 186012 42215 186013
rect 42149 186010 42196 186012
rect 42104 186008 42196 186010
rect 42104 185952 42154 186008
rect 42104 185950 42196 185952
rect 42149 185948 42196 185950
rect 42260 185948 42266 186012
rect 42149 185947 42215 185948
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 668209 184514 668275 184517
rect 666694 184512 668275 184514
rect 666694 184456 668214 184512
rect 668270 184456 668275 184512
rect 666694 184454 668275 184456
rect 666694 184446 666754 184454
rect 668209 184451 668275 184454
rect 666356 184386 666754 184446
rect 579521 184378 579587 184381
rect 575798 184376 579587 184378
rect 575798 184320 579526 184376
rect 579582 184320 579587 184376
rect 575798 184318 579587 184320
rect 575798 183940 575858 184318
rect 579521 184315 579587 184318
rect 589457 183562 589523 183565
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 589457 183499 589523 183502
rect 42425 183154 42491 183157
rect 44173 183154 44239 183157
rect 42425 183152 44239 183154
rect 42425 183096 42430 183152
rect 42486 183096 44178 183152
rect 44234 183096 44239 183152
rect 42425 183094 44239 183096
rect 42425 183091 42491 183094
rect 44173 183091 44239 183094
rect 579521 181930 579587 181933
rect 575798 181928 579587 181930
rect 575798 181872 579526 181928
rect 579582 181872 579587 181928
rect 575798 181870 579587 181872
rect 575798 181764 575858 181870
rect 579521 181867 579587 181870
rect 590561 181930 590627 181933
rect 590561 181928 592572 181930
rect 590561 181872 590566 181928
rect 590622 181872 592572 181928
rect 590561 181870 592572 181872
rect 590561 181867 590627 181870
rect 673085 181524 673151 181525
rect 673085 181522 673132 181524
rect 673040 181520 673132 181522
rect 673040 181464 673090 181520
rect 673040 181462 673132 181464
rect 673085 181460 673132 181462
rect 673196 181460 673202 181524
rect 673085 181459 673151 181460
rect 667749 181386 667815 181389
rect 667749 181384 669330 181386
rect 667749 181328 667754 181384
rect 667810 181328 669330 181384
rect 667749 181326 669330 181328
rect 667749 181323 667815 181326
rect 669270 181250 669330 181326
rect 676213 181250 676279 181253
rect 669270 181248 676279 181250
rect 669270 181192 676218 181248
rect 676274 181192 676279 181248
rect 669270 181190 676279 181192
rect 676213 181187 676279 181190
rect 589641 180298 589707 180301
rect 667565 180298 667631 180301
rect 675845 180298 675911 180301
rect 589641 180296 592572 180298
rect 589641 180240 589646 180296
rect 589702 180240 592572 180296
rect 589641 180238 592572 180240
rect 667565 180296 675911 180298
rect 667565 180240 667570 180296
rect 667626 180240 675850 180296
rect 675906 180240 675911 180296
rect 667565 180238 675911 180240
rect 589641 180235 589707 180238
rect 667565 180235 667631 180238
rect 675845 180235 675911 180238
rect 578785 180162 578851 180165
rect 575798 180160 578851 180162
rect 575798 180104 578790 180160
rect 578846 180104 578851 180160
rect 575798 180102 578851 180104
rect 575798 179588 575858 180102
rect 578785 180099 578851 180102
rect 667974 179618 667980 179620
rect 666694 179558 667980 179618
rect 666694 179550 666754 179558
rect 667974 179556 667980 179558
rect 668044 179556 668050 179620
rect 666356 179490 666754 179550
rect 42057 179346 42123 179349
rect 51901 179346 51967 179349
rect 42057 179344 51967 179346
rect 42057 179288 42062 179344
rect 42118 179288 51906 179344
rect 51962 179288 51967 179344
rect 42057 179286 51967 179288
rect 42057 179283 42123 179286
rect 51901 179283 51967 179286
rect 676213 178938 676279 178941
rect 676213 178936 676322 178938
rect 676213 178880 676218 178936
rect 676274 178880 676322 178936
rect 676213 178875 676322 178880
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 676262 178500 676322 178875
rect 673310 178060 673316 178124
rect 673380 178122 673386 178124
rect 673380 178062 676292 178122
rect 673380 178060 673386 178062
rect 668209 177986 668275 177989
rect 666694 177984 668275 177986
rect 666694 177928 668214 177984
rect 668270 177928 668275 177984
rect 666694 177926 668275 177928
rect 666694 177918 666754 177926
rect 668209 177923 668275 177926
rect 670785 177986 670851 177989
rect 671337 177986 671403 177989
rect 670785 177984 671403 177986
rect 670785 177928 670790 177984
rect 670846 177928 671342 177984
rect 671398 177928 671403 177984
rect 670785 177926 671403 177928
rect 670785 177923 670851 177926
rect 671337 177923 671403 177926
rect 666356 177858 666754 177918
rect 579521 177714 579587 177717
rect 575798 177712 579587 177714
rect 575798 177656 579526 177712
rect 579582 177656 579587 177712
rect 575798 177654 579587 177656
rect 575798 177412 575858 177654
rect 579521 177651 579587 177654
rect 675845 177714 675911 177717
rect 675845 177712 676292 177714
rect 675845 177656 675850 177712
rect 675906 177656 676292 177712
rect 675845 177654 676292 177656
rect 675845 177651 675911 177654
rect 673913 177306 673979 177309
rect 673913 177304 676292 177306
rect 673913 177248 673918 177304
rect 673974 177248 676292 177304
rect 673913 177246 676292 177248
rect 673913 177243 673979 177246
rect 589641 177034 589707 177037
rect 589641 177032 592572 177034
rect 589641 176976 589646 177032
rect 589702 176976 592572 177032
rect 589641 176974 592572 176976
rect 589641 176971 589707 176974
rect 673177 176898 673243 176901
rect 673177 176896 676292 176898
rect 673177 176840 673182 176896
rect 673238 176840 676292 176896
rect 673177 176838 676292 176840
rect 673177 176835 673243 176838
rect 676806 176608 676812 176672
rect 676876 176608 676882 176672
rect 676814 176460 676874 176608
rect 674465 176082 674531 176085
rect 674465 176080 676292 176082
rect 674465 176024 674470 176080
rect 674526 176024 676292 176080
rect 674465 176022 676292 176024
rect 674465 176019 674531 176022
rect 672441 175674 672507 175677
rect 672441 175672 676292 175674
rect 672441 175616 672446 175672
rect 672502 175616 676292 175672
rect 672441 175614 676292 175616
rect 672441 175611 672507 175614
rect 589457 175402 589523 175405
rect 589457 175400 592572 175402
rect 589457 175344 589462 175400
rect 589518 175344 592572 175400
rect 589457 175342 592572 175344
rect 589457 175339 589523 175342
rect 674649 175266 674715 175269
rect 674649 175264 676292 175266
rect 575982 175130 576042 175236
rect 674649 175208 674654 175264
rect 674710 175208 676292 175264
rect 674649 175206 676292 175208
rect 674649 175203 674715 175206
rect 578785 175130 578851 175133
rect 575982 175128 578851 175130
rect 575982 175072 578790 175128
rect 578846 175072 578851 175128
rect 575982 175070 578851 175072
rect 578785 175067 578851 175070
rect 666737 174994 666803 174997
rect 666737 174992 669330 174994
rect 666737 174936 666742 174992
rect 666798 174936 669330 174992
rect 666737 174934 669330 174936
rect 666737 174931 666803 174934
rect 669270 174858 669330 174934
rect 669270 174798 676292 174858
rect 668025 174722 668091 174725
rect 666694 174720 668091 174722
rect 666694 174664 668030 174720
rect 668086 174664 668091 174720
rect 666694 174662 668091 174664
rect 666694 174654 666754 174662
rect 668025 174659 668091 174662
rect 666356 174594 666754 174654
rect 673913 174450 673979 174453
rect 673913 174448 676292 174450
rect 673913 174392 673918 174448
rect 673974 174392 676292 174448
rect 673913 174390 676292 174392
rect 673913 174387 673979 174390
rect 674833 174042 674899 174045
rect 674833 174040 676292 174042
rect 674833 173984 674838 174040
rect 674894 173984 676292 174040
rect 674833 173982 676292 173984
rect 674833 173979 674899 173982
rect 589457 173770 589523 173773
rect 589457 173768 592572 173770
rect 589457 173712 589462 173768
rect 589518 173712 592572 173768
rect 589457 173710 592572 173712
rect 589457 173707 589523 173710
rect 680997 173634 681063 173637
rect 680997 173632 681076 173634
rect 680997 173576 681002 173632
rect 681058 173576 681076 173632
rect 680997 173574 681076 173576
rect 680997 173571 681063 173574
rect 578417 173498 578483 173501
rect 575798 173496 578483 173498
rect 575798 173440 578422 173496
rect 578478 173440 578483 173496
rect 575798 173438 578483 173440
rect 575798 173060 575858 173438
rect 578417 173435 578483 173438
rect 676029 173226 676095 173229
rect 676029 173224 676292 173226
rect 676029 173168 676034 173224
rect 676090 173168 676292 173224
rect 676029 173166 676292 173168
rect 676029 173163 676095 173166
rect 666356 172962 666938 173022
rect 666878 172954 666938 172962
rect 674097 172954 674163 172957
rect 666878 172952 674163 172954
rect 666878 172896 674102 172952
rect 674158 172896 674163 172952
rect 666878 172894 674163 172896
rect 674097 172891 674163 172894
rect 675886 172756 675892 172820
rect 675956 172818 675962 172820
rect 675956 172758 676292 172818
rect 675956 172756 675962 172758
rect 669497 172410 669563 172413
rect 669497 172408 676292 172410
rect 669497 172352 669502 172408
rect 669558 172352 676292 172408
rect 669497 172350 676292 172352
rect 669497 172347 669563 172350
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 671981 172002 672047 172005
rect 671981 172000 676292 172002
rect 671981 171944 671986 172000
rect 672042 171944 676292 172000
rect 671981 171942 676292 171944
rect 671981 171939 672047 171942
rect 682377 171594 682443 171597
rect 682364 171592 682443 171594
rect 682364 171536 682382 171592
rect 682438 171536 682443 171592
rect 682364 171534 682443 171536
rect 682377 171531 682443 171534
rect 670417 171186 670483 171189
rect 670417 171184 676292 171186
rect 670417 171128 670422 171184
rect 670478 171128 676292 171184
rect 670417 171126 676292 171128
rect 670417 171123 670483 171126
rect 578233 171050 578299 171053
rect 575798 171048 578299 171050
rect 575798 170992 578238 171048
rect 578294 170992 578299 171048
rect 575798 170990 578299 170992
rect 575798 170884 575858 170990
rect 578233 170987 578299 170990
rect 673453 170778 673519 170781
rect 673453 170776 676292 170778
rect 673453 170720 673458 170776
rect 673514 170720 676292 170776
rect 673453 170718 676292 170720
rect 673453 170715 673519 170718
rect 589641 170506 589707 170509
rect 589641 170504 592572 170506
rect 589641 170448 589646 170504
rect 589702 170448 592572 170504
rect 589641 170446 592572 170448
rect 589641 170443 589707 170446
rect 674606 170310 676292 170370
rect 670601 170234 670667 170237
rect 674606 170234 674666 170310
rect 670601 170232 674666 170234
rect 670601 170176 670606 170232
rect 670662 170176 674666 170232
rect 670601 170174 674666 170176
rect 670601 170171 670667 170174
rect 676581 169962 676647 169965
rect 676581 169960 676660 169962
rect 676581 169904 676586 169960
rect 676642 169904 676660 169960
rect 676581 169902 676660 169904
rect 676581 169899 676647 169902
rect 666356 169698 666754 169758
rect 666694 169690 666754 169698
rect 667933 169690 667999 169693
rect 666694 169688 667999 169690
rect 666694 169632 667938 169688
rect 667994 169632 667999 169688
rect 666694 169630 667999 169632
rect 667933 169627 667999 169630
rect 676170 169494 676292 169554
rect 675886 169356 675892 169420
rect 675956 169418 675962 169420
rect 676170 169418 676230 169494
rect 675956 169358 676230 169418
rect 675956 169356 675962 169358
rect 578693 169282 578759 169285
rect 575798 169280 578759 169282
rect 575798 169224 578698 169280
rect 578754 169224 578759 169280
rect 575798 169222 578759 169224
rect 575798 168708 575858 169222
rect 578693 169219 578759 169222
rect 672993 169146 673059 169149
rect 672993 169144 676292 169146
rect 672993 169088 672998 169144
rect 673054 169088 676292 169144
rect 672993 169086 676292 169088
rect 672993 169083 673059 169086
rect 589457 168874 589523 168877
rect 589457 168872 592572 168874
rect 589457 168816 589462 168872
rect 589518 168816 592572 168872
rect 589457 168814 592572 168816
rect 589457 168811 589523 168814
rect 673085 168738 673151 168741
rect 673085 168736 676292 168738
rect 673085 168680 673090 168736
rect 673146 168680 676292 168736
rect 673085 168678 676292 168680
rect 673085 168675 673151 168678
rect 672349 168330 672415 168333
rect 672349 168328 676292 168330
rect 672349 168272 672354 168328
rect 672410 168272 676292 168328
rect 672349 168270 676292 168272
rect 672349 168267 672415 168270
rect 666356 168066 666754 168126
rect 666694 168058 666754 168066
rect 672165 168058 672231 168061
rect 666694 168056 672231 168058
rect 666694 168000 672170 168056
rect 672226 168000 672231 168056
rect 666694 167998 672231 168000
rect 672165 167995 672231 167998
rect 683113 167922 683179 167925
rect 683100 167920 683179 167922
rect 683100 167864 683118 167920
rect 683174 167864 683179 167920
rect 683100 167862 683179 167864
rect 683113 167859 683179 167862
rect 675334 167452 675340 167516
rect 675404 167514 675410 167516
rect 675661 167514 675727 167517
rect 675404 167512 676292 167514
rect 675404 167456 675666 167512
rect 675722 167456 676292 167512
rect 675404 167454 676292 167456
rect 675404 167452 675410 167454
rect 675661 167451 675727 167454
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 676170 167046 676292 167106
rect 578233 166970 578299 166973
rect 575798 166968 578299 166970
rect 575798 166912 578238 166968
rect 578294 166912 578299 166968
rect 575798 166910 578299 166912
rect 575798 166532 575858 166910
rect 578233 166907 578299 166910
rect 672349 166970 672415 166973
rect 676170 166970 676230 167046
rect 672349 166968 676230 166970
rect 672349 166912 672354 166968
rect 672410 166912 676230 166968
rect 672349 166910 676230 166912
rect 672349 166907 672415 166910
rect 676581 166428 676647 166429
rect 676581 166424 676628 166428
rect 676692 166426 676698 166428
rect 676581 166368 676586 166424
rect 676581 166364 676628 166368
rect 676692 166366 676738 166426
rect 676692 166364 676698 166366
rect 676581 166363 676647 166364
rect 589457 165610 589523 165613
rect 589457 165608 592572 165610
rect 589457 165552 589462 165608
rect 589518 165552 592572 165608
rect 589457 165550 592572 165552
rect 589457 165547 589523 165550
rect 667933 164930 667999 164933
rect 666694 164928 667999 164930
rect 666694 164872 667938 164928
rect 667994 164872 667999 164928
rect 666694 164870 667999 164872
rect 666694 164862 666754 164870
rect 667933 164867 667999 164870
rect 666356 164802 666754 164862
rect 579521 164522 579587 164525
rect 575798 164520 579587 164522
rect 575798 164464 579526 164520
rect 579582 164464 579587 164520
rect 575798 164462 579587 164464
rect 575798 164356 575858 164462
rect 579521 164459 579587 164462
rect 589457 163978 589523 163981
rect 589457 163976 592572 163978
rect 589457 163920 589462 163976
rect 589518 163920 592572 163976
rect 589457 163918 592572 163920
rect 589457 163915 589523 163918
rect 668761 163298 668827 163301
rect 666694 163296 668827 163298
rect 666694 163240 668766 163296
rect 668822 163240 668827 163296
rect 666694 163238 668827 163240
rect 666694 163230 666754 163238
rect 668761 163235 668827 163238
rect 666356 163170 666754 163230
rect 669313 162890 669379 162893
rect 673821 162890 673887 162893
rect 669313 162888 673887 162890
rect 669313 162832 669318 162888
rect 669374 162832 673826 162888
rect 673882 162832 673887 162888
rect 669313 162830 673887 162832
rect 669313 162827 669379 162830
rect 673821 162827 673887 162830
rect 579337 162754 579403 162757
rect 575798 162752 579403 162754
rect 575798 162696 579342 162752
rect 579398 162696 579403 162752
rect 575798 162694 579403 162696
rect 575798 162180 575858 162694
rect 579337 162691 579403 162694
rect 676070 162692 676076 162756
rect 676140 162754 676146 162756
rect 680997 162754 681063 162757
rect 676140 162752 681063 162754
rect 676140 162696 681002 162752
rect 681058 162696 681063 162752
rect 676140 162694 681063 162696
rect 676140 162692 676146 162694
rect 680997 162691 681063 162694
rect 589457 162346 589523 162349
rect 675201 162346 675267 162349
rect 675845 162346 675911 162349
rect 589457 162344 592572 162346
rect 589457 162288 589462 162344
rect 589518 162288 592572 162344
rect 589457 162286 592572 162288
rect 675201 162344 675911 162346
rect 675201 162288 675206 162344
rect 675262 162288 675850 162344
rect 675906 162288 675911 162344
rect 675201 162286 675911 162288
rect 589457 162283 589523 162286
rect 675201 162283 675267 162286
rect 675845 162283 675911 162286
rect 674097 162074 674163 162077
rect 683113 162074 683179 162077
rect 674097 162072 683179 162074
rect 674097 162016 674102 162072
rect 674158 162016 683118 162072
rect 683174 162016 683179 162072
rect 674097 162014 683179 162016
rect 674097 162011 674163 162014
rect 683113 162011 683179 162014
rect 673126 161468 673132 161532
rect 673196 161530 673202 161532
rect 675477 161530 675543 161533
rect 673196 161528 675543 161530
rect 673196 161472 675482 161528
rect 675538 161472 675543 161528
rect 673196 161470 675543 161472
rect 673196 161468 673202 161470
rect 675477 161467 675543 161470
rect 589457 160714 589523 160717
rect 589457 160712 592572 160714
rect 589457 160656 589462 160712
rect 589518 160656 592572 160712
rect 589457 160654 592572 160656
rect 589457 160651 589523 160654
rect 668209 160034 668275 160037
rect 666694 160032 668275 160034
rect 575982 159898 576042 160004
rect 666694 159976 668214 160032
rect 668270 159976 668275 160032
rect 666694 159974 668275 159976
rect 666694 159966 666754 159974
rect 668209 159971 668275 159974
rect 666356 159906 666754 159966
rect 578233 159898 578299 159901
rect 575982 159896 578299 159898
rect 575982 159840 578238 159896
rect 578294 159840 578299 159896
rect 575982 159838 578299 159840
rect 578233 159835 578299 159838
rect 589457 159082 589523 159085
rect 589457 159080 592572 159082
rect 589457 159024 589462 159080
rect 589518 159024 592572 159080
rect 589457 159022 592572 159024
rect 589457 159019 589523 159022
rect 578417 158402 578483 158405
rect 669313 158402 669379 158405
rect 575798 158400 578483 158402
rect 575798 158344 578422 158400
rect 578478 158344 578483 158400
rect 575798 158342 578483 158344
rect 575798 157828 575858 158342
rect 578417 158339 578483 158342
rect 666694 158400 669379 158402
rect 666694 158344 669318 158400
rect 669374 158344 669379 158400
rect 666694 158342 669379 158344
rect 666694 158334 666754 158342
rect 669313 158339 669379 158342
rect 666356 158274 666754 158334
rect 589273 157450 589339 157453
rect 589273 157448 592572 157450
rect 589273 157392 589278 157448
rect 589334 157392 592572 157448
rect 589273 157390 592572 157392
rect 589273 157387 589339 157390
rect 675753 157042 675819 157045
rect 676438 157042 676444 157044
rect 675753 157040 676444 157042
rect 675753 156984 675758 157040
rect 675814 156984 676444 157040
rect 675753 156982 676444 156984
rect 675753 156979 675819 156982
rect 676438 156980 676444 156982
rect 676508 156980 676514 157044
rect 673545 156498 673611 156501
rect 675293 156498 675359 156501
rect 673545 156496 675359 156498
rect 673545 156440 673550 156496
rect 673606 156440 675298 156496
rect 675354 156440 675359 156496
rect 673545 156438 675359 156440
rect 673545 156435 673611 156438
rect 675293 156435 675359 156438
rect 668761 156226 668827 156229
rect 673545 156226 673611 156229
rect 668761 156224 673611 156226
rect 668761 156168 668766 156224
rect 668822 156168 673550 156224
rect 673606 156168 673611 156224
rect 668761 156166 673611 156168
rect 668761 156163 668827 156166
rect 673545 156163 673611 156166
rect 578877 155954 578943 155957
rect 575798 155952 578943 155954
rect 575798 155896 578882 155952
rect 578938 155896 578943 155952
rect 575798 155894 578943 155896
rect 575798 155652 575858 155894
rect 578877 155891 578943 155894
rect 670417 155954 670483 155957
rect 675109 155954 675175 155957
rect 670417 155952 675175 155954
rect 670417 155896 670422 155952
rect 670478 155896 675114 155952
rect 675170 155896 675175 155952
rect 670417 155894 675175 155896
rect 670417 155891 670483 155894
rect 675109 155891 675175 155894
rect 589457 155818 589523 155821
rect 675753 155818 675819 155821
rect 676254 155818 676260 155820
rect 589457 155816 592572 155818
rect 589457 155760 589462 155816
rect 589518 155760 592572 155816
rect 589457 155758 592572 155760
rect 675753 155816 676260 155818
rect 675753 155760 675758 155816
rect 675814 155760 676260 155816
rect 675753 155758 676260 155760
rect 589457 155755 589523 155758
rect 675753 155755 675819 155758
rect 676254 155756 676260 155758
rect 676324 155756 676330 155820
rect 668209 155138 668275 155141
rect 666694 155136 668275 155138
rect 666694 155080 668214 155136
rect 668270 155080 668275 155136
rect 666694 155078 668275 155080
rect 666694 155070 666754 155078
rect 668209 155075 668275 155078
rect 666356 155010 666754 155070
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 578325 154050 578391 154053
rect 575798 154048 578391 154050
rect 575798 153992 578330 154048
rect 578386 153992 578391 154048
rect 575798 153990 578391 153992
rect 575798 153476 575858 153990
rect 578325 153987 578391 153990
rect 666356 153378 666938 153438
rect 666878 153370 666938 153378
rect 666878 153310 673470 153370
rect 673410 153234 673470 153310
rect 674281 153234 674347 153237
rect 673410 153232 674347 153234
rect 673410 153176 674286 153232
rect 674342 153176 674347 153232
rect 673410 153174 674347 153176
rect 674281 153171 674347 153174
rect 673085 152690 673151 152693
rect 675109 152690 675175 152693
rect 673085 152688 675175 152690
rect 673085 152632 673090 152688
rect 673146 152632 675114 152688
rect 675170 152632 675175 152688
rect 673085 152630 675175 152632
rect 673085 152627 673151 152630
rect 675109 152627 675175 152630
rect 589457 152554 589523 152557
rect 589457 152552 592572 152554
rect 589457 152496 589462 152552
rect 589518 152496 592572 152552
rect 589457 152494 592572 152496
rect 589457 152491 589523 152494
rect 578233 151738 578299 151741
rect 575798 151736 578299 151738
rect 575798 151680 578238 151736
rect 578294 151680 578299 151736
rect 575798 151678 578299 151680
rect 575798 151300 575858 151678
rect 578233 151675 578299 151678
rect 675753 151466 675819 151469
rect 676622 151466 676628 151468
rect 675753 151464 676628 151466
rect 675753 151408 675758 151464
rect 675814 151408 676628 151464
rect 675753 151406 676628 151408
rect 675753 151403 675819 151406
rect 676622 151404 676628 151406
rect 676692 151404 676698 151468
rect 673177 151330 673243 151333
rect 675109 151330 675175 151333
rect 673177 151328 675175 151330
rect 673177 151272 673182 151328
rect 673238 151272 675114 151328
rect 675170 151272 675175 151328
rect 673177 151270 675175 151272
rect 673177 151267 673243 151270
rect 675109 151267 675175 151270
rect 590009 150922 590075 150925
rect 590009 150920 592572 150922
rect 590009 150864 590014 150920
rect 590070 150864 592572 150920
rect 590009 150862 592572 150864
rect 590009 150859 590075 150862
rect 669589 150378 669655 150381
rect 674925 150378 674991 150381
rect 669589 150376 674991 150378
rect 669589 150320 669594 150376
rect 669650 150320 674930 150376
rect 674986 150320 674991 150376
rect 669589 150318 674991 150320
rect 669589 150315 669655 150318
rect 674925 150315 674991 150318
rect 666356 150114 666754 150174
rect 666694 150106 666754 150114
rect 671705 150106 671771 150109
rect 666694 150104 671771 150106
rect 666694 150048 671710 150104
rect 671766 150048 671771 150104
rect 666694 150046 671771 150048
rect 671705 150043 671771 150046
rect 578877 149698 578943 149701
rect 575798 149696 578943 149698
rect 575798 149640 578882 149696
rect 578938 149640 578943 149696
rect 575798 149638 578943 149640
rect 575798 149124 575858 149638
rect 578877 149635 578943 149638
rect 589457 149290 589523 149293
rect 589457 149288 592572 149290
rect 589457 149232 589462 149288
rect 589518 149232 592572 149288
rect 589457 149230 592572 149232
rect 589457 149227 589523 149230
rect 668761 148610 668827 148613
rect 666694 148608 668827 148610
rect 666694 148552 668766 148608
rect 668822 148552 668827 148608
rect 666694 148550 668827 148552
rect 666694 148542 666754 148550
rect 668761 148547 668827 148550
rect 666356 148482 666754 148542
rect 675753 148474 675819 148477
rect 676070 148474 676076 148476
rect 675753 148472 676076 148474
rect 675753 148416 675758 148472
rect 675814 148416 676076 148472
rect 675753 148414 676076 148416
rect 675753 148411 675819 148414
rect 676070 148412 676076 148414
rect 676140 148412 676146 148476
rect 588537 147658 588603 147661
rect 670601 147658 670667 147661
rect 675109 147658 675175 147661
rect 675385 147660 675451 147661
rect 588537 147656 592572 147658
rect 588537 147600 588542 147656
rect 588598 147600 592572 147656
rect 588537 147598 592572 147600
rect 670601 147656 675175 147658
rect 670601 147600 670606 147656
rect 670662 147600 675114 147656
rect 675170 147600 675175 147656
rect 670601 147598 675175 147600
rect 588537 147595 588603 147598
rect 670601 147595 670667 147598
rect 675109 147595 675175 147598
rect 675334 147596 675340 147660
rect 675404 147658 675451 147660
rect 675404 147656 675496 147658
rect 675446 147600 675496 147656
rect 675404 147598 675496 147600
rect 675404 147596 675451 147598
rect 675385 147595 675451 147596
rect 579521 147522 579587 147525
rect 575798 147520 579587 147522
rect 575798 147464 579526 147520
rect 579582 147464 579587 147520
rect 575798 147462 579587 147464
rect 575798 146948 575858 147462
rect 579521 147459 579587 147462
rect 589457 146026 589523 146029
rect 589457 146024 592572 146026
rect 589457 145968 589462 146024
rect 589518 145968 592572 146024
rect 589457 145966 592572 145968
rect 589457 145963 589523 145966
rect 668761 145346 668827 145349
rect 666694 145344 668827 145346
rect 666694 145288 668766 145344
rect 668822 145288 668827 145344
rect 666694 145286 668827 145288
rect 666694 145278 666754 145286
rect 668761 145283 668827 145286
rect 666356 145218 666754 145278
rect 671981 144938 672047 144941
rect 675109 144938 675175 144941
rect 671981 144936 675175 144938
rect 671981 144880 671986 144936
rect 672042 144880 675114 144936
rect 675170 144880 675175 144936
rect 671981 144878 675175 144880
rect 671981 144875 672047 144878
rect 675109 144875 675175 144878
rect 575982 144666 576042 144772
rect 579245 144666 579311 144669
rect 575982 144664 579311 144666
rect 575982 144608 579250 144664
rect 579306 144608 579311 144664
rect 575982 144606 579311 144608
rect 579245 144603 579311 144606
rect 589457 144394 589523 144397
rect 589457 144392 592572 144394
rect 589457 144336 589462 144392
rect 589518 144336 592572 144392
rect 589457 144334 592572 144336
rect 589457 144331 589523 144334
rect 668393 143714 668459 143717
rect 666694 143712 668459 143714
rect 666694 143656 668398 143712
rect 668454 143656 668459 143712
rect 666694 143654 668459 143656
rect 666694 143646 666754 143654
rect 668393 143651 668459 143654
rect 666356 143586 666754 143646
rect 579521 143034 579587 143037
rect 575798 143032 579587 143034
rect 575798 142976 579526 143032
rect 579582 142976 579587 143032
rect 575798 142974 579587 142976
rect 575798 142596 575858 142974
rect 579521 142971 579587 142974
rect 589825 142762 589891 142765
rect 589825 142760 592572 142762
rect 589825 142704 589830 142760
rect 589886 142704 592572 142760
rect 589825 142702 592572 142704
rect 589825 142699 589891 142702
rect 589457 141130 589523 141133
rect 589457 141128 592572 141130
rect 589457 141072 589462 141128
rect 589518 141072 592572 141128
rect 589457 141070 592572 141072
rect 589457 141067 589523 141070
rect 578601 140586 578667 140589
rect 575798 140584 578667 140586
rect 575798 140528 578606 140584
rect 578662 140528 578667 140584
rect 575798 140526 578667 140528
rect 575798 140420 575858 140526
rect 578601 140523 578667 140526
rect 669262 140450 669268 140452
rect 666694 140390 669268 140450
rect 666694 140382 666754 140390
rect 669262 140388 669268 140390
rect 669332 140388 669338 140452
rect 666356 140322 666754 140382
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 578601 138818 578667 138821
rect 668577 138818 668643 138821
rect 575798 138816 578667 138818
rect 575798 138760 578606 138816
rect 578662 138760 578667 138816
rect 575798 138758 578667 138760
rect 575798 138244 575858 138758
rect 578601 138755 578667 138758
rect 666694 138816 668643 138818
rect 666694 138760 668582 138816
rect 668638 138760 668643 138816
rect 666694 138758 668643 138760
rect 666694 138750 666754 138758
rect 668577 138755 668643 138758
rect 666356 138690 666754 138750
rect 589457 137866 589523 137869
rect 589457 137864 592572 137866
rect 589457 137808 589462 137864
rect 589518 137808 592572 137864
rect 589457 137806 592572 137808
rect 589457 137803 589523 137806
rect 578877 136642 578943 136645
rect 575798 136640 578943 136642
rect 575798 136584 578882 136640
rect 578938 136584 578943 136640
rect 575798 136582 578943 136584
rect 575798 136068 575858 136582
rect 578877 136579 578943 136582
rect 589457 136234 589523 136237
rect 589457 136232 592572 136234
rect 589457 136176 589462 136232
rect 589518 136176 592572 136232
rect 589457 136174 592572 136176
rect 589457 136171 589523 136174
rect 669129 135554 669195 135557
rect 666694 135552 669195 135554
rect 666694 135496 669134 135552
rect 669190 135496 669195 135552
rect 666694 135494 669195 135496
rect 666694 135486 666754 135494
rect 669129 135491 669195 135494
rect 666356 135426 666754 135486
rect 668761 135146 668827 135149
rect 672165 135146 672231 135149
rect 668761 135144 672231 135146
rect 668761 135088 668766 135144
rect 668822 135088 672170 135144
rect 672226 135088 672231 135144
rect 668761 135086 672231 135088
rect 668761 135083 668827 135086
rect 672165 135083 672231 135086
rect 590377 134602 590443 134605
rect 667197 134602 667263 134605
rect 675845 134602 675911 134605
rect 590377 134600 592572 134602
rect 590377 134544 590382 134600
rect 590438 134544 592572 134600
rect 590377 134542 592572 134544
rect 667197 134600 675911 134602
rect 667197 134544 667202 134600
rect 667258 134544 675850 134600
rect 675906 134544 675911 134600
rect 667197 134542 675911 134544
rect 590377 134539 590443 134542
rect 667197 134539 667263 134542
rect 675845 134539 675911 134542
rect 579521 134466 579587 134469
rect 575798 134464 579587 134466
rect 575798 134408 579526 134464
rect 579582 134408 579587 134464
rect 575798 134406 579587 134408
rect 575798 133892 575858 134406
rect 579521 134403 579587 134406
rect 666356 133794 666754 133854
rect 666694 133786 666754 133794
rect 667933 133786 667999 133789
rect 666694 133784 667999 133786
rect 666694 133728 667938 133784
rect 667994 133728 667999 133784
rect 666694 133726 667999 133728
rect 667933 133723 667999 133726
rect 667381 133514 667447 133517
rect 672993 133514 673059 133517
rect 667381 133512 673059 133514
rect 667381 133456 667386 133512
rect 667442 133456 672998 133512
rect 673054 133456 673059 133512
rect 667381 133454 673059 133456
rect 667381 133451 667447 133454
rect 672993 133451 673059 133454
rect 676262 133106 676322 133348
rect 676489 133106 676555 133109
rect 669270 133046 676322 133106
rect 676446 133104 676555 133106
rect 676446 133048 676494 133104
rect 676550 133048 676555 133104
rect 589457 132970 589523 132973
rect 589457 132968 592572 132970
rect 589457 132912 589462 132968
rect 589518 132912 592572 132968
rect 589457 132910 592572 132912
rect 589457 132907 589523 132910
rect 667013 132698 667079 132701
rect 669270 132698 669330 133046
rect 676446 133043 676555 133048
rect 676446 132940 676506 133043
rect 667013 132696 669330 132698
rect 667013 132640 667018 132696
rect 667074 132640 669330 132696
rect 667013 132638 669330 132640
rect 672993 132698 673059 132701
rect 672993 132696 676322 132698
rect 672993 132640 672998 132696
rect 673054 132640 676322 132696
rect 672993 132638 676322 132640
rect 667013 132635 667079 132638
rect 672993 132635 673059 132638
rect 676262 132532 676322 132638
rect 579061 132290 579127 132293
rect 575798 132288 579127 132290
rect 575798 132232 579066 132288
rect 579122 132232 579127 132288
rect 575798 132230 579127 132232
rect 575798 131716 575858 132230
rect 579061 132227 579127 132230
rect 673361 132154 673427 132157
rect 673361 132152 676292 132154
rect 673361 132096 673366 132152
rect 673422 132096 676292 132152
rect 673361 132094 676292 132096
rect 673361 132091 673427 132094
rect 671337 131746 671403 131749
rect 671337 131744 676292 131746
rect 671337 131688 671342 131744
rect 671398 131688 676292 131744
rect 671337 131686 676292 131688
rect 671337 131683 671403 131686
rect 589457 131338 589523 131341
rect 674465 131338 674531 131341
rect 589457 131336 592572 131338
rect 589457 131280 589462 131336
rect 589518 131280 592572 131336
rect 589457 131278 592572 131280
rect 674465 131336 676292 131338
rect 674465 131280 674470 131336
rect 674526 131280 676292 131336
rect 674465 131278 676292 131280
rect 589457 131275 589523 131278
rect 674465 131275 674531 131278
rect 669957 130930 670023 130933
rect 669957 130928 676292 130930
rect 669957 130872 669962 130928
rect 670018 130872 676292 130928
rect 669957 130870 676292 130872
rect 669957 130867 670023 130870
rect 668577 130658 668643 130661
rect 666694 130656 668643 130658
rect 666694 130600 668582 130656
rect 668638 130600 668643 130656
rect 666694 130598 668643 130600
rect 666694 130590 666754 130598
rect 668577 130595 668643 130598
rect 666356 130530 666754 130590
rect 674649 130522 674715 130525
rect 674649 130520 676292 130522
rect 674649 130464 674654 130520
rect 674710 130464 676292 130520
rect 674649 130462 676292 130464
rect 674649 130459 674715 130462
rect 676213 130250 676279 130253
rect 676213 130248 676322 130250
rect 676213 130192 676218 130248
rect 676274 130192 676322 130248
rect 676213 130187 676322 130192
rect 676262 130084 676322 130187
rect 578877 129706 578943 129709
rect 575798 129704 578943 129706
rect 575798 129648 578882 129704
rect 578938 129648 578943 129704
rect 575798 129646 578943 129648
rect 575798 129540 575858 129646
rect 578877 129643 578943 129646
rect 588537 129706 588603 129709
rect 673913 129706 673979 129709
rect 588537 129704 592572 129706
rect 588537 129648 588542 129704
rect 588598 129648 592572 129704
rect 588537 129646 592572 129648
rect 673913 129704 676292 129706
rect 673913 129648 673918 129704
rect 673974 129648 676292 129704
rect 673913 129646 676292 129648
rect 588537 129643 588603 129646
rect 673913 129643 673979 129646
rect 671521 129298 671587 129301
rect 671521 129296 676292 129298
rect 671521 129240 671526 129296
rect 671582 129240 676292 129296
rect 671521 129238 676292 129240
rect 671521 129235 671587 129238
rect 668025 129026 668091 129029
rect 666694 129024 668091 129026
rect 666694 128968 668030 129024
rect 668086 128968 668091 129024
rect 666694 128966 668091 128968
rect 666694 128958 666754 128966
rect 668025 128963 668091 128966
rect 666356 128898 666754 128958
rect 674925 128890 674991 128893
rect 674925 128888 676292 128890
rect 674925 128832 674930 128888
rect 674986 128832 676292 128888
rect 674925 128830 676292 128832
rect 674925 128827 674991 128830
rect 674557 128482 674623 128485
rect 674557 128480 676292 128482
rect 674557 128424 674562 128480
rect 674618 128424 676292 128480
rect 674557 128422 676292 128424
rect 674557 128419 674623 128422
rect 589457 128074 589523 128077
rect 589457 128072 592572 128074
rect 589457 128016 589462 128072
rect 589518 128016 592572 128072
rect 589457 128014 592572 128016
rect 589457 128011 589523 128014
rect 579521 127938 579587 127941
rect 575798 127936 579587 127938
rect 575798 127880 579526 127936
rect 579582 127880 579587 127936
rect 575798 127878 579587 127880
rect 575798 127364 575858 127878
rect 579521 127875 579587 127878
rect 676446 127805 676506 128044
rect 668577 127802 668643 127805
rect 676213 127802 676279 127805
rect 668577 127800 676279 127802
rect 668577 127744 668582 127800
rect 668638 127744 676218 127800
rect 676274 127744 676279 127800
rect 668577 127742 676279 127744
rect 668577 127739 668643 127742
rect 676213 127739 676279 127742
rect 676397 127800 676506 127805
rect 676397 127744 676402 127800
rect 676458 127744 676506 127800
rect 676397 127742 676506 127744
rect 676397 127739 676463 127742
rect 676630 127396 676690 127636
rect 676622 127332 676628 127396
rect 676692 127332 676698 127396
rect 676070 126924 676076 126988
rect 676140 126986 676146 126988
rect 676262 126986 676322 127228
rect 676140 126926 676322 126986
rect 676140 126924 676146 126926
rect 673361 126578 673427 126581
rect 676262 126578 676322 126820
rect 673361 126576 676322 126578
rect 673361 126520 673366 126576
rect 673422 126520 676322 126576
rect 673361 126518 676322 126520
rect 673361 126515 673427 126518
rect 589917 126442 589983 126445
rect 589917 126440 592572 126442
rect 589917 126384 589922 126440
rect 589978 126384 592572 126440
rect 589917 126382 592572 126384
rect 589917 126379 589983 126382
rect 679574 126173 679634 126412
rect 679574 126168 679683 126173
rect 679574 126112 679622 126168
rect 679678 126112 679683 126168
rect 679574 126110 679683 126112
rect 679617 126107 679683 126110
rect 668945 125762 669011 125765
rect 676262 125764 676322 126004
rect 666694 125760 669011 125762
rect 666694 125704 668950 125760
rect 669006 125704 669011 125760
rect 666694 125702 669011 125704
rect 666694 125694 666754 125702
rect 668945 125699 669011 125702
rect 676254 125700 676260 125764
rect 676324 125700 676330 125764
rect 666356 125634 666754 125694
rect 682334 125357 682394 125596
rect 578325 125354 578391 125357
rect 575798 125352 578391 125354
rect 575798 125296 578330 125352
rect 578386 125296 578391 125352
rect 575798 125294 578391 125296
rect 682334 125352 682443 125357
rect 682334 125296 682382 125352
rect 682438 125296 682443 125352
rect 682334 125294 682443 125296
rect 575798 125188 575858 125294
rect 578325 125291 578391 125294
rect 682377 125291 682443 125294
rect 672165 124946 672231 124949
rect 676262 124946 676322 125188
rect 672165 124944 676322 124946
rect 672165 124888 672170 124944
rect 672226 124888 676322 124944
rect 672165 124886 676322 124888
rect 672165 124883 672231 124886
rect 589457 124810 589523 124813
rect 589457 124808 592572 124810
rect 589457 124752 589462 124808
rect 589518 124752 592572 124808
rect 589457 124750 592572 124752
rect 589457 124747 589523 124750
rect 673913 124538 673979 124541
rect 676262 124538 676322 124780
rect 673913 124536 676322 124538
rect 673913 124480 673918 124536
rect 673974 124480 676322 124536
rect 673913 124478 676322 124480
rect 673913 124475 673979 124478
rect 672809 124130 672875 124133
rect 676446 124132 676506 124372
rect 666694 124128 672875 124130
rect 666694 124072 672814 124128
rect 672870 124072 672875 124128
rect 666694 124070 672875 124072
rect 666694 124062 666754 124070
rect 672809 124067 672875 124070
rect 676438 124068 676444 124132
rect 676508 124068 676514 124132
rect 666356 124002 666754 124062
rect 674373 123722 674439 123725
rect 676262 123722 676322 123964
rect 674373 123720 676322 123722
rect 674373 123664 674378 123720
rect 674434 123664 676322 123720
rect 674373 123662 676322 123664
rect 674373 123659 674439 123662
rect 578417 123586 578483 123589
rect 575798 123584 578483 123586
rect 575798 123528 578422 123584
rect 578478 123528 578483 123584
rect 575798 123526 578483 123528
rect 575798 123012 575858 123526
rect 578417 123523 578483 123526
rect 676446 123317 676506 123556
rect 672993 123314 673059 123317
rect 672993 123312 676322 123314
rect 672993 123256 672998 123312
rect 673054 123256 676322 123312
rect 672993 123254 676322 123256
rect 676446 123312 676555 123317
rect 676446 123256 676494 123312
rect 676550 123256 676555 123312
rect 676446 123254 676555 123256
rect 672993 123251 673059 123254
rect 589457 123178 589523 123181
rect 589457 123176 592572 123178
rect 589457 123120 589462 123176
rect 589518 123120 592572 123176
rect 676262 123148 676322 123254
rect 676489 123251 676555 123254
rect 589457 123118 592572 123120
rect 589457 123115 589523 123118
rect 673177 123042 673243 123045
rect 674373 123042 674439 123045
rect 673177 123040 674439 123042
rect 673177 122984 673182 123040
rect 673238 122984 674378 123040
rect 674434 122984 674439 123040
rect 673177 122982 674439 122984
rect 673177 122979 673243 122982
rect 674373 122979 674439 122982
rect 674741 123042 674807 123045
rect 674741 123040 674850 123042
rect 674741 122984 674746 123040
rect 674802 122984 674850 123040
rect 674741 122979 674850 122984
rect 674790 122906 674850 122979
rect 676489 122906 676555 122909
rect 674790 122904 676555 122906
rect 674790 122848 676494 122904
rect 676550 122848 676555 122904
rect 674790 122846 676555 122848
rect 676489 122843 676555 122846
rect 675017 122498 675083 122501
rect 676262 122498 676322 122740
rect 675017 122496 676322 122498
rect 675017 122440 675022 122496
rect 675078 122440 676322 122496
rect 675017 122438 676322 122440
rect 675017 122435 675083 122438
rect 667054 122028 667060 122092
rect 667124 122090 667130 122092
rect 675334 122090 675340 122092
rect 667124 122030 675340 122090
rect 667124 122028 667130 122030
rect 675334 122028 675340 122030
rect 675404 122090 675410 122092
rect 676262 122090 676322 122332
rect 675404 122030 676322 122090
rect 675404 122028 675410 122030
rect 670417 121682 670483 121685
rect 675017 121682 675083 121685
rect 676262 121682 676322 121924
rect 670417 121680 675083 121682
rect 670417 121624 670422 121680
rect 670478 121624 675022 121680
rect 675078 121624 675083 121680
rect 670417 121622 675083 121624
rect 670417 121619 670483 121622
rect 675017 121619 675083 121622
rect 676032 121622 676322 121682
rect 590009 121546 590075 121549
rect 590009 121544 592572 121546
rect 590009 121488 590014 121544
rect 590070 121488 592572 121544
rect 590009 121486 592572 121488
rect 590009 121483 590075 121486
rect 578877 121410 578943 121413
rect 575798 121408 578943 121410
rect 575798 121352 578882 121408
rect 578938 121352 578943 121408
rect 575798 121350 578943 121352
rect 575798 120836 575858 121350
rect 578877 121347 578943 121350
rect 672533 120866 672599 120869
rect 666694 120864 672599 120866
rect 666694 120808 672538 120864
rect 672594 120808 672599 120864
rect 666694 120806 672599 120808
rect 666694 120798 666754 120806
rect 672533 120803 672599 120806
rect 666356 120738 666754 120798
rect 672993 120730 673059 120733
rect 676032 120730 676092 121622
rect 672993 120728 676092 120730
rect 672993 120672 672998 120728
rect 673054 120672 676092 120728
rect 672993 120670 676092 120672
rect 672993 120667 673059 120670
rect 589641 119914 589707 119917
rect 589641 119912 592572 119914
rect 589641 119856 589646 119912
rect 589702 119856 592572 119912
rect 589641 119854 592572 119856
rect 589641 119851 589707 119854
rect 668761 119234 668827 119237
rect 666694 119232 668827 119234
rect 666694 119176 668766 119232
rect 668822 119176 668827 119232
rect 666694 119174 668827 119176
rect 666694 119166 666754 119174
rect 668761 119171 668827 119174
rect 666356 119106 666754 119166
rect 669221 118826 669287 118829
rect 672809 118826 672875 118829
rect 669221 118824 672875 118826
rect 669221 118768 669226 118824
rect 669282 118768 672814 118824
rect 672870 118768 672875 118824
rect 669221 118766 672875 118768
rect 669221 118763 669287 118766
rect 672809 118763 672875 118766
rect 575982 118418 576042 118660
rect 578509 118418 578575 118421
rect 575982 118416 578575 118418
rect 575982 118360 578514 118416
rect 578570 118360 578575 118416
rect 575982 118358 578575 118360
rect 578509 118355 578575 118358
rect 590101 118282 590167 118285
rect 590101 118280 592572 118282
rect 590101 118224 590106 118280
rect 590162 118224 592572 118280
rect 590101 118222 592572 118224
rect 590101 118219 590167 118222
rect 666356 117474 666938 117534
rect 666878 117466 666938 117474
rect 674097 117466 674163 117469
rect 666878 117464 674163 117466
rect 666878 117408 674102 117464
rect 674158 117408 674163 117464
rect 666878 117406 674163 117408
rect 674097 117403 674163 117406
rect 675702 117268 675708 117332
rect 675772 117330 675778 117332
rect 682377 117330 682443 117333
rect 675772 117328 682443 117330
rect 675772 117272 682382 117328
rect 682438 117272 682443 117328
rect 675772 117270 682443 117272
rect 675772 117268 675778 117270
rect 682377 117267 682443 117270
rect 675201 117058 675267 117061
rect 675937 117058 676003 117061
rect 675201 117056 676003 117058
rect 675201 117000 675206 117056
rect 675262 117000 675942 117056
rect 675998 117000 676003 117056
rect 675201 116998 676003 117000
rect 675201 116995 675267 116998
rect 675937 116995 676003 116998
rect 579521 116922 579587 116925
rect 575798 116920 579587 116922
rect 575798 116864 579526 116920
rect 579582 116864 579587 116920
rect 575798 116862 579587 116864
rect 575798 116484 575858 116862
rect 579521 116859 579587 116862
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 666356 115842 666754 115902
rect 666694 115834 666754 115842
rect 672349 115834 672415 115837
rect 666694 115832 672415 115834
rect 666694 115776 672354 115832
rect 672410 115776 672415 115832
rect 666694 115774 672415 115776
rect 672349 115771 672415 115774
rect 674046 115772 674052 115836
rect 674116 115834 674122 115836
rect 675477 115834 675543 115837
rect 674116 115832 675543 115834
rect 674116 115776 675482 115832
rect 675538 115776 675543 115832
rect 674116 115774 675543 115776
rect 674116 115772 674122 115774
rect 675477 115771 675543 115774
rect 590285 115018 590351 115021
rect 590285 115016 592572 115018
rect 590285 114960 590290 115016
rect 590346 114960 592572 115016
rect 590285 114958 592572 114960
rect 590285 114955 590351 114958
rect 579245 114474 579311 114477
rect 575798 114472 579311 114474
rect 575798 114416 579250 114472
rect 579306 114416 579311 114472
rect 575798 114414 579311 114416
rect 575798 114308 575858 114414
rect 579245 114411 579311 114414
rect 669221 114338 669287 114341
rect 666694 114336 669287 114338
rect 666694 114280 669226 114336
rect 669282 114280 669287 114336
rect 666694 114278 669287 114280
rect 666694 114270 666754 114278
rect 669221 114275 669287 114278
rect 666356 114210 666754 114270
rect 589457 113386 589523 113389
rect 589457 113384 592572 113386
rect 589457 113328 589462 113384
rect 589518 113328 592572 113384
rect 589457 113326 592572 113328
rect 589457 113323 589523 113326
rect 668761 112706 668827 112709
rect 666694 112704 668827 112706
rect 666694 112648 668766 112704
rect 668822 112648 668827 112704
rect 666694 112646 668827 112648
rect 666694 112638 666754 112646
rect 668761 112643 668827 112646
rect 666356 112578 666754 112638
rect 579521 112570 579587 112573
rect 575798 112568 579587 112570
rect 575798 112512 579526 112568
rect 579582 112512 579587 112568
rect 575798 112510 579587 112512
rect 575798 112132 575858 112510
rect 579521 112507 579587 112510
rect 675753 112434 675819 112437
rect 676622 112434 676628 112436
rect 675753 112432 676628 112434
rect 675753 112376 675758 112432
rect 675814 112376 676628 112432
rect 675753 112374 676628 112376
rect 675753 112371 675819 112374
rect 676622 112372 676628 112374
rect 676692 112372 676698 112436
rect 589457 111754 589523 111757
rect 675753 111754 675819 111757
rect 676254 111754 676260 111756
rect 589457 111752 592572 111754
rect 589457 111696 589462 111752
rect 589518 111696 592572 111752
rect 589457 111694 592572 111696
rect 675753 111752 676260 111754
rect 675753 111696 675758 111752
rect 675814 111696 676260 111752
rect 675753 111694 676260 111696
rect 589457 111691 589523 111694
rect 675753 111691 675819 111694
rect 676254 111692 676260 111694
rect 676324 111692 676330 111756
rect 675753 111348 675819 111349
rect 675702 111284 675708 111348
rect 675772 111346 675819 111348
rect 675772 111344 675864 111346
rect 675814 111288 675864 111344
rect 675772 111286 675864 111288
rect 675772 111284 675819 111286
rect 675753 111283 675819 111284
rect 672993 111074 673059 111077
rect 666694 111072 673059 111074
rect 666694 111016 672998 111072
rect 673054 111016 673059 111072
rect 666694 111014 673059 111016
rect 666694 111006 666754 111014
rect 672993 111011 673059 111014
rect 666356 110946 666754 111006
rect 675753 110394 675819 110397
rect 676438 110394 676444 110396
rect 675753 110392 676444 110394
rect 675753 110336 675758 110392
rect 675814 110336 676444 110392
rect 675753 110334 676444 110336
rect 675753 110331 675819 110334
rect 676438 110332 676444 110334
rect 676508 110332 676514 110396
rect 579337 110122 579403 110125
rect 575798 110120 579403 110122
rect 575798 110064 579342 110120
rect 579398 110064 579403 110120
rect 575798 110062 579403 110064
rect 575798 109956 575858 110062
rect 579337 110059 579403 110062
rect 589273 110122 589339 110125
rect 589273 110120 592572 110122
rect 589273 110064 589278 110120
rect 589334 110064 592572 110120
rect 589273 110062 592572 110064
rect 589273 110059 589339 110062
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 578325 108354 578391 108357
rect 575798 108352 578391 108354
rect 575798 108296 578330 108352
rect 578386 108296 578391 108352
rect 575798 108294 578391 108296
rect 575798 107780 575858 108294
rect 578325 108291 578391 108294
rect 675753 108218 675819 108221
rect 676070 108218 676076 108220
rect 675753 108216 676076 108218
rect 675753 108160 675758 108216
rect 675814 108160 676076 108216
rect 675753 108158 676076 108160
rect 675753 108155 675819 108158
rect 676070 108156 676076 108158
rect 676140 108156 676146 108220
rect 667933 107810 667999 107813
rect 666694 107808 667999 107810
rect 666694 107752 667938 107808
rect 667994 107752 667999 107808
rect 666694 107750 667999 107752
rect 666694 107742 666754 107750
rect 667933 107747 667999 107750
rect 666356 107682 666754 107742
rect 673913 106994 673979 106997
rect 675385 106994 675451 106997
rect 673913 106992 675451 106994
rect 673913 106936 673918 106992
rect 673974 106936 675390 106992
rect 675446 106936 675451 106992
rect 673913 106934 675451 106936
rect 673913 106931 673979 106934
rect 675385 106931 675451 106934
rect 589825 106858 589891 106861
rect 589825 106856 592572 106858
rect 589825 106800 589830 106856
rect 589886 106800 592572 106856
rect 589825 106798 592572 106800
rect 589825 106795 589891 106798
rect 673177 106314 673243 106317
rect 675109 106314 675175 106317
rect 673177 106312 675175 106314
rect 673177 106256 673182 106312
rect 673238 106256 675114 106312
rect 675170 106256 675175 106312
rect 673177 106254 675175 106256
rect 673177 106251 673243 106254
rect 675109 106251 675175 106254
rect 668393 106178 668459 106181
rect 666694 106176 668459 106178
rect 666694 106120 668398 106176
rect 668454 106120 668459 106176
rect 666694 106118 668459 106120
rect 666694 106110 666754 106118
rect 668393 106115 668459 106118
rect 666356 106050 666754 106110
rect 579061 105906 579127 105909
rect 575798 105904 579127 105906
rect 575798 105848 579066 105904
rect 579122 105848 579127 105904
rect 575798 105846 579127 105848
rect 575798 105604 575858 105846
rect 579061 105843 579127 105846
rect 589457 105226 589523 105229
rect 589457 105224 592572 105226
rect 589457 105168 589462 105224
rect 589518 105168 592572 105224
rect 589457 105166 592572 105168
rect 589457 105163 589523 105166
rect 672165 104682 672231 104685
rect 675109 104682 675175 104685
rect 672165 104680 675175 104682
rect 672165 104624 672170 104680
rect 672226 104624 675114 104680
rect 675170 104624 675175 104680
rect 672165 104622 675175 104624
rect 672165 104619 672231 104622
rect 675109 104619 675175 104622
rect 668761 104546 668827 104549
rect 666694 104544 668827 104546
rect 666694 104488 668766 104544
rect 668822 104488 668827 104544
rect 666694 104486 668827 104488
rect 666694 104478 666754 104486
rect 668761 104483 668827 104486
rect 666356 104418 666754 104478
rect 588721 103594 588787 103597
rect 588721 103592 592572 103594
rect 588721 103536 588726 103592
rect 588782 103536 592572 103592
rect 588721 103534 592572 103536
rect 588721 103531 588787 103534
rect 575982 103322 576042 103428
rect 579521 103322 579587 103325
rect 575982 103320 579587 103322
rect 575982 103264 579526 103320
rect 579582 103264 579587 103320
rect 575982 103262 579587 103264
rect 579521 103259 579587 103262
rect 668577 102914 668643 102917
rect 666694 102912 668643 102914
rect 666694 102856 668582 102912
rect 668638 102856 668643 102912
rect 666694 102854 668643 102856
rect 666694 102846 666754 102854
rect 668577 102851 668643 102854
rect 666356 102786 666754 102846
rect 675385 102644 675451 102645
rect 675334 102642 675340 102644
rect 675294 102582 675340 102642
rect 675404 102640 675451 102644
rect 675446 102584 675451 102640
rect 675334 102580 675340 102582
rect 675404 102580 675451 102584
rect 675385 102579 675451 102580
rect 589457 101962 589523 101965
rect 589457 101960 592572 101962
rect 589457 101904 589462 101960
rect 589518 101904 592572 101960
rect 589457 101902 592572 101904
rect 589457 101899 589523 101902
rect 579521 101690 579587 101693
rect 575798 101688 579587 101690
rect 575798 101632 579526 101688
rect 579582 101632 579587 101688
rect 575798 101630 579587 101632
rect 575798 101252 575858 101630
rect 579521 101627 579587 101630
rect 673361 101010 673427 101013
rect 675109 101010 675175 101013
rect 673361 101008 675175 101010
rect 673361 100952 673366 101008
rect 673422 100952 675114 101008
rect 675170 100952 675175 101008
rect 673361 100950 675175 100952
rect 673361 100947 673427 100950
rect 675109 100947 675175 100950
rect 578601 99242 578667 99245
rect 575798 99240 578667 99242
rect 575798 99184 578606 99240
rect 578662 99184 578667 99240
rect 575798 99182 578667 99184
rect 575798 99076 575858 99182
rect 578601 99179 578667 99182
rect 578325 97474 578391 97477
rect 575798 97472 578391 97474
rect 575798 97416 578330 97472
rect 578386 97416 578391 97472
rect 575798 97414 578391 97416
rect 575798 96900 575858 97414
rect 578325 97411 578391 97414
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 641989 96522 642055 96525
rect 647182 96522 647188 96524
rect 641989 96520 647188 96522
rect 641989 96464 641994 96520
rect 642050 96464 647188 96520
rect 641989 96462 647188 96464
rect 641989 96459 642055 96462
rect 647182 96460 647188 96462
rect 647252 96460 647258 96524
rect 633934 95372 633940 95436
rect 634004 95434 634010 95436
rect 635733 95434 635799 95437
rect 634004 95432 635799 95434
rect 634004 95376 635738 95432
rect 635794 95376 635799 95432
rect 634004 95374 635799 95376
rect 634004 95372 634010 95374
rect 635733 95371 635799 95374
rect 579521 95026 579587 95029
rect 575798 95024 579587 95026
rect 575798 94968 579526 95024
rect 579582 94968 579587 95024
rect 575798 94966 579587 94968
rect 575798 94724 575858 94966
rect 579521 94963 579587 94966
rect 647141 95026 647207 95029
rect 647141 95024 647434 95026
rect 647141 94968 647146 95024
rect 647202 94968 647434 95024
rect 647141 94966 647434 94968
rect 647141 94963 647207 94966
rect 626441 94482 626507 94485
rect 626441 94480 628268 94482
rect 626441 94424 626446 94480
rect 626502 94424 628268 94480
rect 647374 94452 647434 94966
rect 626441 94422 628268 94424
rect 626441 94419 626507 94422
rect 654593 94210 654659 94213
rect 654593 94208 656788 94210
rect 654593 94152 654598 94208
rect 654654 94152 656788 94208
rect 654593 94150 656788 94152
rect 654593 94147 654659 94150
rect 626257 93666 626323 93669
rect 626257 93664 628268 93666
rect 626257 93608 626262 93664
rect 626318 93608 628268 93664
rect 626257 93606 628268 93608
rect 626257 93603 626323 93606
rect 655421 93394 655487 93397
rect 665541 93394 665607 93397
rect 655421 93392 656788 93394
rect 655421 93336 655426 93392
rect 655482 93336 656788 93392
rect 655421 93334 656788 93336
rect 663596 93392 665607 93394
rect 663596 93336 665546 93392
rect 665602 93336 665607 93392
rect 663596 93334 665607 93336
rect 655421 93331 655487 93334
rect 665541 93331 665607 93334
rect 578509 93122 578575 93125
rect 575798 93120 578575 93122
rect 575798 93064 578514 93120
rect 578570 93064 578575 93120
rect 575798 93062 578575 93064
rect 575798 92548 575858 93062
rect 578509 93059 578575 93062
rect 650310 93060 650316 93124
rect 650380 93122 650386 93124
rect 663793 93122 663859 93125
rect 650380 93062 656818 93122
rect 650380 93060 650386 93062
rect 626441 92850 626507 92853
rect 626441 92848 628268 92850
rect 626441 92792 626446 92848
rect 626502 92792 628268 92848
rect 626441 92790 628268 92792
rect 626441 92787 626507 92790
rect 656758 92548 656818 93062
rect 663566 93120 663859 93122
rect 663566 93064 663798 93120
rect 663854 93064 663859 93120
rect 663566 93062 663859 93064
rect 663566 92548 663626 93062
rect 663793 93059 663859 93062
rect 647509 92442 647575 92445
rect 647509 92440 647618 92442
rect 647509 92384 647514 92440
rect 647570 92384 647618 92440
rect 647509 92379 647618 92384
rect 625797 92034 625863 92037
rect 625797 92032 628268 92034
rect 625797 91976 625802 92032
rect 625858 91976 628268 92032
rect 647558 92004 647618 92379
rect 625797 91974 628268 91976
rect 625797 91971 625863 91974
rect 665173 91762 665239 91765
rect 663596 91760 665239 91762
rect 663596 91704 665178 91760
rect 665234 91704 665239 91760
rect 663596 91702 665239 91704
rect 665173 91699 665239 91702
rect 654317 91490 654383 91493
rect 654317 91488 656788 91490
rect 654317 91432 654322 91488
rect 654378 91432 656788 91488
rect 654317 91430 656788 91432
rect 654317 91427 654383 91430
rect 626441 91218 626507 91221
rect 626441 91216 628268 91218
rect 626441 91160 626446 91216
rect 626502 91160 628268 91216
rect 626441 91158 628268 91160
rect 626441 91155 626507 91158
rect 579061 90946 579127 90949
rect 575798 90944 579127 90946
rect 575798 90888 579066 90944
rect 579122 90888 579127 90944
rect 575798 90886 579127 90888
rect 575798 90372 575858 90886
rect 579061 90883 579127 90886
rect 655421 90674 655487 90677
rect 665357 90674 665423 90677
rect 655421 90672 656788 90674
rect 655421 90616 655426 90672
rect 655482 90616 656788 90672
rect 655421 90614 656788 90616
rect 663596 90672 665423 90674
rect 663596 90616 665362 90672
rect 665418 90616 665423 90672
rect 663596 90614 665423 90616
rect 655421 90611 655487 90614
rect 665357 90611 665423 90614
rect 626441 90402 626507 90405
rect 626441 90400 628268 90402
rect 626441 90344 626446 90400
rect 626502 90344 628268 90400
rect 626441 90342 628268 90344
rect 626441 90339 626507 90342
rect 655789 89858 655855 89861
rect 664345 89858 664411 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 655789 89798 656788 89800
rect 663596 89856 664411 89858
rect 663596 89800 664350 89856
rect 664406 89800 664411 89856
rect 663596 89798 664411 89800
rect 655789 89795 655855 89798
rect 664345 89795 664411 89798
rect 626441 89586 626507 89589
rect 648245 89586 648311 89589
rect 626441 89584 628268 89586
rect 626441 89528 626446 89584
rect 626502 89528 628268 89584
rect 626441 89526 628268 89528
rect 648140 89584 648311 89586
rect 648140 89528 648250 89584
rect 648306 89528 648311 89584
rect 648140 89526 648311 89528
rect 626441 89523 626507 89526
rect 648245 89523 648311 89526
rect 663977 89042 664043 89045
rect 663596 89040 664043 89042
rect 663596 88984 663982 89040
rect 664038 88984 664043 89040
rect 663596 88982 664043 88984
rect 663977 88979 664043 88982
rect 626398 88710 628268 88770
rect 624969 88634 625035 88637
rect 626398 88634 626458 88710
rect 624969 88632 626458 88634
rect 624969 88576 624974 88632
rect 625030 88576 626458 88632
rect 624969 88574 626458 88576
rect 624969 88571 625035 88574
rect 575982 88090 576042 88196
rect 579521 88090 579587 88093
rect 575982 88088 579587 88090
rect 575982 88032 579526 88088
rect 579582 88032 579587 88088
rect 575982 88030 579587 88032
rect 579521 88027 579587 88030
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 626257 87138 626323 87141
rect 649993 87138 650059 87141
rect 626257 87136 628268 87138
rect 626257 87080 626262 87136
rect 626318 87080 628268 87136
rect 626257 87078 628268 87080
rect 648140 87136 650059 87138
rect 648140 87080 649998 87136
rect 650054 87080 650059 87136
rect 648140 87078 650059 87080
rect 626257 87075 626323 87078
rect 649993 87075 650059 87078
rect 579337 86458 579403 86461
rect 575798 86456 579403 86458
rect 575798 86400 579342 86456
rect 579398 86400 579403 86456
rect 575798 86398 579403 86400
rect 575798 86020 575858 86398
rect 579337 86395 579403 86398
rect 626441 86322 626507 86325
rect 626441 86320 628268 86322
rect 626441 86264 626446 86320
rect 626502 86264 628268 86320
rect 626441 86262 628268 86264
rect 626441 86259 626507 86262
rect 626441 85506 626507 85509
rect 626441 85504 628268 85506
rect 626441 85448 626446 85504
rect 626502 85448 628268 85504
rect 626441 85446 628268 85448
rect 626441 85443 626507 85446
rect 625245 84690 625311 84693
rect 650545 84690 650611 84693
rect 625245 84688 628268 84690
rect 625245 84632 625250 84688
rect 625306 84632 628268 84688
rect 625245 84630 628268 84632
rect 648140 84688 650611 84690
rect 648140 84632 650550 84688
rect 650606 84632 650611 84688
rect 648140 84630 650611 84632
rect 625245 84627 625311 84630
rect 650545 84627 650611 84630
rect 579153 84010 579219 84013
rect 575798 84008 579219 84010
rect 575798 83952 579158 84008
rect 579214 83952 579219 84008
rect 575798 83950 579219 83952
rect 575798 83844 575858 83950
rect 579153 83947 579219 83950
rect 625797 83874 625863 83877
rect 625797 83872 628268 83874
rect 625797 83816 625802 83872
rect 625858 83816 628268 83872
rect 625797 83814 628268 83816
rect 625797 83811 625863 83814
rect 628741 83330 628807 83333
rect 628741 83328 628850 83330
rect 628741 83272 628746 83328
rect 628802 83272 628850 83328
rect 628741 83267 628850 83272
rect 628790 83028 628850 83267
rect 579061 82242 579127 82245
rect 650361 82242 650427 82245
rect 575798 82240 579127 82242
rect 575798 82184 579066 82240
rect 579122 82184 579127 82240
rect 648140 82240 650427 82242
rect 575798 82182 579127 82184
rect 575798 81668 575858 82182
rect 579061 82179 579127 82182
rect 628790 81698 628850 82212
rect 648140 82184 650366 82240
rect 650422 82184 650427 82240
rect 648140 82182 650427 82184
rect 650361 82179 650427 82182
rect 629201 81698 629267 81701
rect 628790 81696 629267 81698
rect 628790 81640 629206 81696
rect 629262 81640 629267 81696
rect 628790 81638 629267 81640
rect 629201 81635 629267 81638
rect 578877 80066 578943 80069
rect 575798 80064 578943 80066
rect 575798 80008 578882 80064
rect 578938 80008 578943 80064
rect 575798 80006 578943 80008
rect 575798 79492 575858 80006
rect 578877 80003 578943 80006
rect 633893 78572 633959 78573
rect 633893 78570 633940 78572
rect 633848 78568 633940 78570
rect 633848 78512 633898 78568
rect 633848 78510 633940 78512
rect 633893 78508 633940 78510
rect 634004 78508 634010 78572
rect 633893 78507 633959 78508
rect 637062 78162 637068 78164
rect 625110 78102 637068 78162
rect 579521 77890 579587 77893
rect 575798 77888 579587 77890
rect 575798 77832 579526 77888
rect 579582 77832 579587 77888
rect 575798 77830 579587 77832
rect 575798 77316 575858 77830
rect 579521 77827 579587 77830
rect 581637 77890 581703 77893
rect 625110 77890 625170 78102
rect 637062 78100 637068 78102
rect 637132 78162 637138 78164
rect 639597 78162 639663 78165
rect 637132 78160 639663 78162
rect 637132 78104 639602 78160
rect 639658 78104 639663 78160
rect 637132 78102 639663 78104
rect 637132 78100 637138 78102
rect 639597 78099 639663 78102
rect 581637 77888 625170 77890
rect 581637 77832 581642 77888
rect 581698 77832 625170 77888
rect 581637 77830 625170 77832
rect 581637 77827 581703 77830
rect 624417 77346 624483 77349
rect 633893 77346 633959 77349
rect 624417 77344 633959 77346
rect 624417 77288 624422 77344
rect 624478 77288 633898 77344
rect 633954 77288 633959 77344
rect 624417 77286 633959 77288
rect 624417 77283 624483 77286
rect 633893 77283 633959 77286
rect 578233 75578 578299 75581
rect 575798 75576 578299 75578
rect 575798 75520 578238 75576
rect 578294 75520 578299 75576
rect 575798 75518 578299 75520
rect 575798 75140 575858 75518
rect 578233 75515 578299 75518
rect 646221 74218 646287 74221
rect 646221 74216 646330 74218
rect 646221 74160 646226 74216
rect 646282 74160 646330 74216
rect 646221 74155 646330 74160
rect 646270 73848 646330 74155
rect 579061 73130 579127 73133
rect 575798 73128 579127 73130
rect 575798 73072 579066 73128
rect 579122 73072 579127 73128
rect 575798 73070 579127 73072
rect 575798 72964 575858 73070
rect 579061 73067 579127 73070
rect 646681 71770 646747 71773
rect 646638 71768 646747 71770
rect 646638 71712 646686 71768
rect 646742 71712 646747 71768
rect 646638 71707 646747 71712
rect 646638 71400 646698 71707
rect 579061 71226 579127 71229
rect 575798 71224 579127 71226
rect 575798 71168 579066 71224
rect 579122 71168 579127 71224
rect 575798 71166 579127 71168
rect 575798 70788 575858 71166
rect 579061 71163 579127 71166
rect 646638 68914 646698 68952
rect 647233 68914 647299 68917
rect 646638 68912 647299 68914
rect 646638 68856 647238 68912
rect 647294 68856 647299 68912
rect 646638 68854 647299 68856
rect 647233 68851 647299 68854
rect 646221 67146 646287 67149
rect 646221 67144 646330 67146
rect 646221 67088 646226 67144
rect 646282 67088 646330 67144
rect 646221 67083 646330 67088
rect 646270 66504 646330 67083
rect 646497 64426 646563 64429
rect 646454 64424 646563 64426
rect 646454 64368 646502 64424
rect 646558 64368 646563 64424
rect 646454 64363 646563 64368
rect 646454 64056 646514 64363
rect 648613 62114 648679 62117
rect 646638 62112 648679 62114
rect 646638 62056 648618 62112
rect 648674 62056 648679 62112
rect 646638 62054 648679 62056
rect 646638 61608 646698 62054
rect 648613 62051 648679 62054
rect 647233 59258 647299 59261
rect 646638 59256 647299 59258
rect 646638 59200 647238 59256
rect 647294 59200 647299 59256
rect 646638 59198 647299 59200
rect 646638 59160 646698 59198
rect 647233 59195 647299 59198
rect 648797 57354 648863 57357
rect 646638 57352 648863 57354
rect 646638 57296 648802 57352
rect 648858 57296 648863 57352
rect 646638 57294 648863 57296
rect 646638 56712 646698 57294
rect 648797 57291 648863 57294
rect 460790 54980 460796 55044
rect 460860 55042 460866 55044
rect 576117 55042 576183 55045
rect 460860 55040 576183 55042
rect 460860 54984 576122 55040
rect 576178 54984 576183 55040
rect 460860 54982 576183 54984
rect 460860 54980 460866 54982
rect 576117 54979 576183 54982
rect 462630 54708 462636 54772
rect 462700 54770 462706 54772
rect 580257 54770 580323 54773
rect 462700 54768 580323 54770
rect 462700 54712 580262 54768
rect 580318 54712 580323 54768
rect 462700 54710 580323 54712
rect 462700 54708 462706 54710
rect 580257 54707 580323 54710
rect 578877 54498 578943 54501
rect 466410 54496 578943 54498
rect 466410 54440 578882 54496
rect 578938 54440 578943 54496
rect 466410 54438 578943 54440
rect 466410 54226 466470 54438
rect 578877 54435 578943 54438
rect 577497 54226 577563 54229
rect 459878 54166 466470 54226
rect 469170 54224 577563 54226
rect 469170 54168 577502 54224
rect 577558 54168 577563 54224
rect 469170 54166 577563 54168
rect 459878 53685 459938 54166
rect 460790 53892 460796 53956
rect 460860 53892 460866 53956
rect 469170 53954 469230 54166
rect 577497 54163 577563 54166
rect 461718 53894 469230 53954
rect 460798 53685 460858 53892
rect 461718 53685 461778 53894
rect 459829 53680 459938 53685
rect 459829 53624 459834 53680
rect 459890 53624 459938 53680
rect 459829 53622 459938 53624
rect 460749 53680 460858 53685
rect 460749 53624 460754 53680
rect 460810 53624 460858 53680
rect 460749 53622 460858 53624
rect 461669 53680 461778 53685
rect 462589 53684 462655 53685
rect 462589 53682 462636 53684
rect 461669 53624 461674 53680
rect 461730 53624 461778 53680
rect 461669 53622 461778 53624
rect 462544 53680 462636 53682
rect 462544 53624 462594 53680
rect 462544 53622 462636 53624
rect 459829 53619 459895 53622
rect 460749 53619 460815 53622
rect 461669 53619 461735 53622
rect 462589 53620 462636 53622
rect 462700 53620 462706 53684
rect 463233 53682 463299 53685
rect 464245 53682 464311 53685
rect 463233 53680 464311 53682
rect 463233 53624 463238 53680
rect 463294 53624 464250 53680
rect 464306 53624 464311 53680
rect 463233 53622 464311 53624
rect 462589 53619 462655 53620
rect 463233 53619 463299 53622
rect 464245 53619 464311 53622
rect 476021 53682 476087 53685
rect 476573 53682 476639 53685
rect 476021 53680 476639 53682
rect 476021 53624 476026 53680
rect 476082 53624 476578 53680
rect 476634 53624 476639 53680
rect 476021 53622 476639 53624
rect 476021 53619 476087 53622
rect 476573 53619 476639 53622
rect 476205 53410 476271 53413
rect 477033 53410 477099 53413
rect 476205 53408 477099 53410
rect 476205 53352 476210 53408
rect 476266 53352 477038 53408
rect 477094 53352 477099 53408
rect 476205 53350 477099 53352
rect 476205 53347 476271 53350
rect 477033 53347 477099 53350
rect 464061 53274 464127 53277
rect 464429 53274 464495 53277
rect 464061 53272 464495 53274
rect 464061 53216 464066 53272
rect 464122 53216 464434 53272
rect 464490 53216 464495 53272
rect 464061 53214 464495 53216
rect 464061 53211 464127 53214
rect 464429 53211 464495 53214
rect 518750 48860 518756 48924
rect 518820 48922 518826 48924
rect 549989 48922 550055 48925
rect 518820 48920 550055 48922
rect 518820 48864 549994 48920
rect 550050 48864 550055 48920
rect 518820 48862 550055 48864
rect 518820 48860 518826 48862
rect 549989 48859 550055 48862
rect 661585 48512 661651 48515
rect 661480 48510 661651 48512
rect 661480 48454 661590 48510
rect 661646 48454 661651 48510
rect 661480 48452 661651 48454
rect 661585 48449 661651 48452
rect 529606 48044 529612 48108
rect 529676 48106 529682 48108
rect 553669 48106 553735 48109
rect 529676 48104 553735 48106
rect 529676 48048 553674 48104
rect 553730 48048 553735 48104
rect 529676 48046 553735 48048
rect 529676 48044 529682 48046
rect 553669 48043 553735 48046
rect 515438 47772 515444 47836
rect 515508 47834 515514 47836
rect 522941 47834 523007 47837
rect 515508 47832 523007 47834
rect 515508 47776 522946 47832
rect 523002 47776 523007 47832
rect 515508 47774 523007 47776
rect 515508 47772 515514 47774
rect 522941 47771 523007 47774
rect 526478 47772 526484 47836
rect 526548 47834 526554 47836
rect 552013 47834 552079 47837
rect 526548 47832 552079 47834
rect 526548 47776 552018 47832
rect 552074 47776 552079 47832
rect 526548 47774 552079 47776
rect 526548 47772 526554 47774
rect 552013 47771 552079 47774
rect 520958 47500 520964 47564
rect 521028 47562 521034 47564
rect 547873 47562 547939 47565
rect 521028 47560 547939 47562
rect 521028 47504 547878 47560
rect 547934 47504 547939 47560
rect 521028 47502 547939 47504
rect 521028 47500 521034 47502
rect 547873 47499 547939 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 522062 47228 522068 47292
rect 522132 47290 522138 47292
rect 545665 47290 545731 47293
rect 522132 47288 545731 47290
rect 522132 47232 545670 47288
rect 545726 47232 545731 47288
rect 522132 47230 545731 47232
rect 522132 47228 522138 47230
rect 545665 47227 545731 47230
rect 458173 47018 458239 47021
rect 465073 47018 465139 47021
rect 458173 47016 465139 47018
rect 458173 46960 458178 47016
rect 458234 46960 465078 47016
rect 465134 46960 465139 47016
rect 458173 46958 465139 46960
rect 458173 46955 458239 46958
rect 465073 46955 465139 46958
rect 458357 46746 458423 46749
rect 465257 46746 465323 46749
rect 458357 46744 465323 46746
rect 458357 46688 458362 46744
rect 458418 46688 465262 46744
rect 465318 46688 465323 46744
rect 458357 46686 465323 46688
rect 458357 46683 458423 46686
rect 465257 46683 465323 46686
rect 461025 44436 461091 44437
rect 460974 44434 460980 44436
rect 460934 44374 460980 44434
rect 461044 44432 461091 44436
rect 461086 44376 461091 44432
rect 460974 44372 460980 44374
rect 461044 44372 461091 44376
rect 462262 44372 462268 44436
rect 462332 44434 462338 44436
rect 462865 44434 462931 44437
rect 463785 44436 463851 44437
rect 463734 44434 463740 44436
rect 462332 44432 462931 44434
rect 462332 44376 462870 44432
rect 462926 44376 462931 44432
rect 462332 44374 462931 44376
rect 463694 44374 463740 44434
rect 463804 44432 463851 44436
rect 463846 44376 463851 44432
rect 462332 44372 462338 44374
rect 461025 44371 461091 44372
rect 462865 44371 462931 44374
rect 463734 44372 463740 44374
rect 463804 44372 463851 44376
rect 463785 44371 463851 44372
rect 130837 44298 130903 44301
rect 132769 44298 132835 44301
rect 142613 44298 142679 44301
rect 130837 44296 132835 44298
rect 130837 44240 130842 44296
rect 130898 44240 132774 44296
rect 132830 44240 132835 44296
rect 130837 44238 132835 44240
rect 130837 44235 130903 44238
rect 132769 44235 132835 44238
rect 142110 44296 142679 44298
rect 142110 44240 142618 44296
rect 142674 44240 142679 44296
rect 142110 44238 142679 44240
rect 141734 43964 141740 44028
rect 141804 44026 141810 44028
rect 142110 44026 142170 44238
rect 142613 44235 142679 44238
rect 255865 44162 255931 44165
rect 460105 44162 460171 44165
rect 464337 44162 464403 44165
rect 255865 44160 460171 44162
rect 255865 44104 255870 44160
rect 255926 44104 460110 44160
rect 460166 44104 460171 44160
rect 255865 44102 460171 44104
rect 255865 44099 255931 44102
rect 460105 44099 460171 44102
rect 460890 44160 464403 44162
rect 460890 44104 464342 44160
rect 464398 44104 464403 44160
rect 460890 44102 464403 44104
rect 141804 43966 142170 44026
rect 141804 43964 141810 43966
rect 361757 43890 361823 43893
rect 440233 43890 440299 43893
rect 361757 43888 440299 43890
rect 361757 43832 361762 43888
rect 361818 43832 440238 43888
rect 440294 43832 440299 43888
rect 361757 43830 440299 43832
rect 361757 43827 361823 43830
rect 440233 43827 440299 43830
rect 441061 43890 441127 43893
rect 460890 43890 460950 44102
rect 464337 44099 464403 44102
rect 441061 43888 460950 43890
rect 441061 43832 441066 43888
rect 441122 43832 460950 43888
rect 441061 43830 460950 43832
rect 441061 43827 441127 43830
rect 460841 43482 460907 43485
rect 471053 43482 471119 43485
rect 460841 43480 471119 43482
rect 460841 43424 460846 43480
rect 460902 43424 471058 43480
rect 471114 43424 471119 43480
rect 460841 43422 471119 43424
rect 460841 43419 460907 43422
rect 471053 43419 471119 43422
rect 462681 43210 462747 43213
rect 465809 43210 465875 43213
rect 462681 43208 465875 43210
rect 462681 43152 462686 43208
rect 462742 43152 465814 43208
rect 465870 43152 465875 43208
rect 462681 43150 465875 43152
rect 462681 43147 462747 43150
rect 465809 43147 465875 43150
rect 461761 42938 461827 42941
rect 463969 42938 464035 42941
rect 461761 42936 464035 42938
rect 461761 42880 461766 42936
rect 461822 42880 463974 42936
rect 464030 42880 464035 42936
rect 461761 42878 464035 42880
rect 461761 42875 461827 42878
rect 463969 42875 464035 42878
rect 518801 42804 518867 42805
rect 518750 42802 518756 42804
rect 518710 42742 518756 42802
rect 518820 42800 518867 42804
rect 518862 42744 518867 42800
rect 518750 42740 518756 42742
rect 518820 42740 518867 42744
rect 518801 42739 518867 42740
rect 415577 42394 415643 42397
rect 415577 42392 422310 42394
rect 415577 42336 415582 42392
rect 415638 42336 422310 42392
rect 415577 42334 422310 42336
rect 415577 42331 415643 42334
rect 422250 42258 422310 42334
rect 446213 42258 446279 42261
rect 461945 42258 462011 42261
rect 422250 42198 427830 42258
rect 419206 42060 419212 42124
rect 419276 42122 419282 42124
rect 419276 42062 420194 42122
rect 419276 42060 419282 42062
rect 420134 41986 420194 42062
rect 420134 41926 424978 41986
rect 365069 41852 365135 41853
rect 416681 41852 416747 41853
rect 365069 41848 365116 41852
rect 365180 41850 365186 41852
rect 416630 41850 416636 41852
rect 365069 41792 365074 41848
rect 365069 41788 365116 41792
rect 365180 41790 365226 41850
rect 416590 41790 416636 41850
rect 416700 41848 416747 41852
rect 416742 41792 416747 41848
rect 365180 41788 365186 41790
rect 416630 41788 416636 41790
rect 416700 41788 416747 41792
rect 365069 41787 365135 41788
rect 416681 41787 416747 41788
rect 419901 41852 419967 41853
rect 419901 41848 419948 41852
rect 420012 41850 420018 41852
rect 424918 41850 424978 41926
rect 425094 41850 425100 41852
rect 419901 41792 419906 41848
rect 419901 41788 419948 41792
rect 420012 41790 420058 41850
rect 424918 41790 425100 41850
rect 420012 41788 420018 41790
rect 425094 41788 425100 41790
rect 425164 41788 425170 41852
rect 419901 41787 419967 41788
rect 427770 41578 427830 42198
rect 446213 42256 462011 42258
rect 446213 42200 446218 42256
rect 446274 42200 461950 42256
rect 462006 42200 462011 42256
rect 446213 42198 462011 42200
rect 446213 42195 446279 42198
rect 461945 42195 462011 42198
rect 515397 42124 515463 42125
rect 520917 42124 520983 42125
rect 522021 42124 522087 42125
rect 526437 42124 526503 42125
rect 529565 42124 529631 42125
rect 515397 42122 515444 42124
rect 515352 42120 515444 42122
rect 515352 42064 515402 42120
rect 515352 42062 515444 42064
rect 515397 42060 515444 42062
rect 515508 42060 515514 42124
rect 520917 42122 520964 42124
rect 520872 42120 520964 42122
rect 520872 42064 520922 42120
rect 520872 42062 520964 42064
rect 520917 42060 520964 42062
rect 521028 42060 521034 42124
rect 522021 42122 522068 42124
rect 521976 42120 522068 42122
rect 521976 42064 522026 42120
rect 521976 42062 522068 42064
rect 522021 42060 522068 42062
rect 522132 42060 522138 42124
rect 526437 42122 526484 42124
rect 526392 42120 526484 42122
rect 526392 42064 526442 42120
rect 526392 42062 526484 42064
rect 526437 42060 526484 42062
rect 526548 42060 526554 42124
rect 529565 42122 529612 42124
rect 529520 42120 529612 42122
rect 529520 42064 529570 42120
rect 529520 42062 529612 42064
rect 529565 42060 529612 42062
rect 529676 42060 529682 42124
rect 515397 42059 515463 42060
rect 520917 42059 520983 42060
rect 522021 42059 522087 42060
rect 526437 42059 526503 42060
rect 529565 42059 529631 42060
rect 441838 41788 441844 41852
rect 441908 41850 441914 41852
rect 451958 41850 451964 41852
rect 441908 41790 451964 41850
rect 441908 41788 441914 41790
rect 451958 41788 451964 41790
rect 452028 41788 452034 41852
rect 446213 41578 446279 41581
rect 427770 41576 446279 41578
rect 427770 41520 446218 41576
rect 446274 41520 446279 41576
rect 427770 41518 446279 41520
rect 446213 41515 446279 41518
rect 141693 40356 141759 40357
rect 141693 40352 141740 40356
rect 141804 40354 141810 40356
rect 141693 40296 141698 40352
rect 141693 40292 141740 40296
rect 141804 40294 141850 40354
rect 141804 40292 141810 40294
rect 141693 40291 141759 40292
<< via3 >>
rect 233004 997384 233068 997388
rect 233004 997328 233018 997384
rect 233018 997328 233068 997384
rect 233004 997324 233068 997328
rect 285444 997384 285508 997388
rect 285444 997328 285458 997384
rect 285458 997328 285508 997384
rect 285444 997324 285508 997328
rect 387564 997384 387628 997388
rect 387564 997328 387578 997384
rect 387578 997328 387628 997384
rect 387564 997324 387628 997328
rect 233004 990932 233068 990996
rect 387564 990932 387628 990996
rect 285444 987940 285508 988004
rect 675892 892196 675956 892260
rect 675892 887708 675956 887772
rect 675708 885804 675772 885868
rect 675524 880636 675588 880700
rect 676260 880364 676324 880428
rect 675340 878460 675404 878524
rect 675340 874108 675404 874172
rect 676444 873020 676508 873084
rect 676260 872748 676324 872812
rect 675708 865676 675772 865740
rect 676076 865404 676140 865468
rect 675892 864860 675956 864924
rect 41828 813180 41892 813244
rect 41828 809976 41892 809980
rect 41828 809920 41842 809976
rect 41842 809920 41892 809976
rect 41828 809916 41892 809920
rect 41828 807876 41892 807940
rect 40540 805564 40604 805628
rect 40724 805156 40788 805220
rect 40908 804748 40972 804812
rect 41828 804748 41892 804812
rect 41828 802436 41892 802500
rect 42196 798144 42260 798148
rect 42196 798088 42210 798144
rect 42210 798088 42260 798144
rect 42196 798084 42260 798088
rect 40908 794820 40972 794884
rect 42196 794472 42260 794476
rect 42196 794416 42210 794472
rect 42210 794416 42260 794472
rect 42196 794412 42260 794416
rect 41644 791964 41708 792028
rect 40724 790604 40788 790668
rect 40540 789244 40604 789308
rect 41460 788292 41524 788356
rect 41828 788020 41892 788084
rect 676076 788020 676140 788084
rect 674420 786660 674484 786724
rect 675340 786720 675404 786724
rect 675340 786664 675390 786720
rect 675390 786664 675404 786720
rect 675340 786660 675404 786664
rect 41644 769796 41708 769860
rect 41460 768980 41524 769044
rect 40540 766532 40604 766596
rect 40724 765308 40788 765372
rect 40908 764900 40972 764964
rect 41828 757692 41892 757756
rect 40724 753884 40788 753948
rect 40908 750484 40972 750548
rect 40540 746676 40604 746740
rect 41644 745588 41708 745652
rect 41460 745044 41524 745108
rect 41828 743064 41892 743068
rect 41828 743008 41878 743064
rect 41878 743008 41892 743064
rect 41828 743004 41892 743008
rect 674236 742460 674300 742524
rect 674604 738108 674668 738172
rect 675340 730144 675404 730148
rect 675340 730088 675354 730144
rect 675354 730088 675404 730144
rect 675340 730084 675404 730088
rect 676812 729812 676876 729876
rect 676076 726548 676140 726612
rect 674420 726276 674484 726340
rect 41828 725868 41892 725932
rect 41828 725656 41892 725660
rect 41828 725600 41842 725656
rect 41842 725600 41892 725656
rect 41828 725596 41892 725600
rect 675156 723148 675220 723212
rect 40724 721708 40788 721772
rect 40540 718524 40604 718588
rect 41828 716892 41892 716956
rect 42012 714444 42076 714508
rect 42012 709880 42076 709884
rect 42012 709824 42062 709880
rect 42062 709824 42076 709880
rect 42012 709820 42076 709824
rect 673868 709336 673932 709340
rect 673868 709280 673882 709336
rect 673882 709280 673932 709336
rect 673868 709276 673932 709280
rect 40540 707916 40604 707980
rect 42196 707916 42260 707980
rect 40724 707372 40788 707436
rect 673868 707024 673932 707028
rect 673868 706968 673882 707024
rect 673882 706968 673932 707024
rect 673868 706964 673932 706968
rect 42196 706208 42260 706212
rect 42196 706152 42246 706208
rect 42246 706152 42260 706208
rect 42196 706148 42260 706152
rect 41644 702748 41708 702812
rect 41460 702068 41524 702132
rect 41828 701796 41892 701860
rect 675524 696824 675588 696828
rect 675524 696768 675538 696824
rect 675538 696768 675588 696824
rect 675524 696764 675588 696768
rect 674420 694588 674484 694652
rect 675524 683980 675588 684044
rect 675340 683768 675404 683772
rect 675340 683712 675354 683768
rect 675354 683712 675404 683768
rect 675340 683708 675404 683712
rect 41828 683572 41892 683636
rect 674236 682348 674300 682412
rect 41828 681728 41892 681732
rect 41828 681672 41842 681728
rect 41842 681672 41892 681728
rect 41828 681668 41892 681672
rect 40540 678928 40604 678992
rect 40724 677750 40788 677754
rect 40724 677694 40774 677750
rect 40774 677694 40788 677750
rect 40724 677690 40788 677694
rect 676076 676364 676140 676428
rect 42196 673100 42260 673164
rect 41828 672692 41892 672756
rect 40356 670924 40420 670988
rect 42196 668476 42260 668540
rect 40356 667388 40420 667452
rect 676812 665756 676876 665820
rect 40724 665212 40788 665276
rect 40540 664124 40604 664188
rect 674604 662356 674668 662420
rect 41644 658548 41708 658612
rect 41828 658336 41892 658340
rect 41828 658280 41842 658336
rect 41842 658280 41892 658336
rect 41828 658276 41892 658280
rect 41460 657188 41524 657252
rect 674236 652836 674300 652900
rect 41460 640596 41524 640660
rect 676076 637468 676140 637532
rect 40540 635292 40604 635356
rect 40724 634884 40788 634948
rect 675156 631348 675220 631412
rect 676076 631348 676140 631412
rect 41644 629852 41708 629916
rect 41828 629172 41892 629236
rect 42196 625908 42260 625972
rect 40724 623732 40788 623796
rect 40540 620876 40604 620940
rect 42196 620196 42260 620260
rect 674420 618700 674484 618764
rect 676260 617068 676324 617132
rect 41644 616796 41708 616860
rect 41460 616388 41524 616452
rect 673868 616116 673932 616180
rect 41828 615436 41892 615500
rect 40540 612308 40604 612372
rect 674420 602924 674484 602988
rect 40540 601972 40604 602036
rect 42932 598436 42996 598500
rect 40356 596974 40420 597038
rect 42932 597000 42996 597004
rect 42932 596944 42946 597000
rect 42946 596944 42996 597000
rect 42932 596940 42996 596944
rect 42012 596396 42076 596460
rect 41782 593948 41846 594012
rect 675156 593132 675220 593196
rect 41782 592724 41846 592788
rect 676076 591636 676140 591700
rect 674236 591228 674300 591292
rect 40908 589052 40972 589116
rect 40356 588780 40420 588844
rect 41460 588780 41524 588844
rect 676076 586196 676140 586260
rect 41828 585924 41892 585988
rect 62068 585652 62132 585716
rect 40356 584564 40420 584628
rect 42196 582448 42260 582452
rect 42196 582392 42246 582448
rect 42246 582392 42260 582448
rect 42196 582388 42260 582392
rect 40356 580212 40420 580276
rect 42196 580272 42260 580276
rect 42196 580216 42246 580272
rect 42246 580216 42260 580272
rect 42196 580212 42260 580216
rect 42012 579320 42076 579324
rect 42012 579264 42062 579320
rect 42062 579264 42076 579320
rect 42012 579260 42076 579264
rect 40908 577764 40972 577828
rect 676812 576812 676876 576876
rect 40540 575724 40604 575788
rect 40724 574636 40788 574700
rect 41460 572868 41524 572932
rect 42012 572656 42076 572660
rect 42012 572600 42062 572656
rect 42062 572600 42076 572656
rect 42012 572596 42076 572600
rect 41644 571508 41708 571572
rect 41828 570208 41892 570212
rect 41828 570152 41842 570208
rect 41842 570152 41892 570208
rect 41828 570148 41892 570152
rect 675340 561912 675404 561916
rect 675340 561856 675390 561912
rect 675390 561856 675404 561912
rect 675340 561852 675404 561856
rect 41092 558724 41156 558788
rect 41092 557488 41156 557552
rect 676260 557500 676324 557564
rect 41828 553964 41892 554028
rect 676812 553828 676876 553892
rect 673684 553480 673748 553484
rect 673684 553424 673698 553480
rect 673698 553424 673748 553480
rect 673684 553420 673748 553424
rect 41828 552740 41892 552804
rect 673684 551516 673748 551580
rect 42012 549476 42076 549540
rect 674972 548796 675036 548860
rect 676996 548252 677060 548316
rect 674972 547844 675036 547908
rect 676260 547572 676324 547636
rect 674420 547028 674484 547092
rect 676076 546756 676140 546820
rect 675340 545804 675404 545868
rect 40724 545592 40788 545596
rect 40724 545536 40738 545592
rect 40738 545536 40788 545592
rect 40724 545532 40788 545536
rect 40540 545260 40604 545324
rect 42012 545260 42076 545324
rect 41828 542268 41892 542332
rect 40724 539548 40788 539612
rect 673500 535060 673564 535124
rect 673500 534244 673564 534308
rect 40540 533292 40604 533356
rect 41644 531660 41708 531724
rect 41460 530164 41524 530228
rect 41828 528940 41892 529004
rect 676996 503644 677060 503708
rect 676812 500924 676876 500988
rect 675892 488820 675956 488884
rect 675892 487868 675956 487932
rect 673868 455228 673932 455292
rect 41460 426566 41524 426630
rect 40908 422248 40972 422312
rect 41828 421500 41892 421564
rect 40724 418644 40788 418708
rect 40540 418372 40604 418436
rect 41828 418372 41892 418436
rect 41644 415244 41708 415308
rect 42012 414564 42076 414628
rect 40908 406948 40972 407012
rect 40540 406676 40604 406740
rect 40724 404500 40788 404564
rect 677180 401236 677244 401300
rect 676812 400420 676876 400484
rect 41460 400012 41524 400076
rect 42012 399392 42076 399396
rect 42012 399336 42026 399392
rect 42026 399336 42076 399392
rect 42012 399332 42076 399336
rect 41828 398848 41892 398852
rect 41828 398792 41842 398848
rect 41842 398792 41892 398848
rect 41828 398788 41892 398792
rect 676076 398788 676140 398852
rect 676260 396748 676324 396812
rect 676444 396340 676508 396404
rect 676628 395116 676692 395180
rect 675892 392804 675956 392868
rect 675708 387636 675772 387700
rect 676260 384916 676324 384980
rect 676444 382196 676508 382260
rect 41460 381788 41524 381852
rect 41828 379340 41892 379404
rect 40724 378932 40788 378996
rect 675708 378720 675772 378724
rect 675708 378664 675758 378720
rect 675758 378664 675772 378720
rect 675708 378660 675772 378664
rect 40540 378524 40604 378588
rect 40908 377708 40972 377772
rect 676628 377300 676692 377364
rect 41644 374580 41708 374644
rect 676076 373628 676140 373692
rect 675340 372464 675404 372468
rect 675340 372408 675390 372464
rect 675390 372408 675404 372464
rect 675340 372404 675404 372408
rect 41828 365740 41892 365804
rect 675340 365604 675404 365668
rect 40908 364788 40972 364852
rect 40724 364108 40788 364172
rect 40540 360028 40604 360092
rect 41828 358728 41892 358732
rect 41828 358672 41878 358728
rect 41878 358672 41892 358728
rect 41828 358668 41892 358672
rect 41460 356900 41524 356964
rect 43668 354588 43732 354652
rect 675524 354180 675588 354244
rect 44772 353636 44836 353700
rect 675892 353772 675956 353836
rect 675708 352956 675772 353020
rect 44036 352140 44100 352204
rect 42012 351868 42076 351932
rect 675892 351732 675956 351796
rect 675340 347652 675404 347716
rect 676444 346564 676508 346628
rect 50108 342076 50172 342140
rect 50476 341668 50540 341732
rect 676260 340172 676324 340236
rect 44220 339764 44284 339828
rect 675524 339416 675588 339420
rect 675524 339360 675538 339416
rect 675538 339360 675588 339416
rect 675524 339356 675588 339360
rect 44404 339220 44468 339284
rect 676076 337860 676140 337924
rect 40540 336908 40604 336972
rect 40724 336500 40788 336564
rect 676444 336500 676508 336564
rect 40908 336092 40972 336156
rect 42196 335684 42260 335748
rect 44588 335412 44652 335476
rect 41276 334868 41340 334932
rect 41276 334460 41340 334524
rect 42012 334656 42076 334660
rect 42012 334600 42062 334656
rect 42062 334600 42076 334656
rect 42012 334596 42076 334600
rect 43852 334656 43916 334660
rect 43852 334600 43866 334656
rect 43866 334600 43916 334656
rect 43852 334596 43916 334600
rect 44036 334520 44100 334524
rect 44036 334464 44050 334520
rect 44050 334464 44100 334520
rect 44036 334460 44100 334464
rect 44588 334324 44652 334388
rect 41828 332828 41892 332892
rect 41644 331740 41708 331804
rect 675340 327992 675404 327996
rect 675340 327936 675390 327992
rect 675390 327936 675404 327992
rect 675340 327932 675404 327936
rect 62252 327660 62316 327724
rect 676628 325620 676692 325684
rect 41828 324864 41892 324868
rect 41828 324808 41842 324864
rect 41842 324808 41892 324864
rect 41828 324804 41892 324808
rect 40908 322764 40972 322828
rect 40724 317460 40788 317524
rect 40540 315964 40604 316028
rect 41828 315616 41892 315620
rect 41828 315560 41842 315616
rect 41842 315560 41892 315616
rect 41828 315556 41892 315560
rect 42196 313712 42260 313716
rect 42196 313656 42210 313712
rect 42210 313656 42260 313712
rect 42196 313652 42260 313656
rect 44404 311884 44468 311948
rect 44220 311264 44284 311268
rect 44220 311208 44270 311264
rect 44270 311208 44284 311264
rect 44220 311204 44284 311208
rect 675340 309164 675404 309228
rect 675892 308756 675956 308820
rect 676076 304540 676140 304604
rect 675892 302636 675956 302700
rect 676628 301608 676692 301612
rect 676628 301552 676642 301608
rect 676642 301552 676692 301608
rect 676628 301548 676692 301552
rect 675156 298148 675220 298212
rect 675524 297604 675588 297668
rect 675708 297332 675772 297396
rect 675524 295760 675588 295764
rect 675524 295704 675574 295760
rect 675574 295704 675588 295760
rect 675524 295700 675588 295704
rect 41828 295564 41892 295628
rect 676444 294612 676508 294676
rect 40540 292588 40604 292592
rect 40540 292532 40590 292588
rect 40590 292532 40604 292588
rect 40540 292528 40604 292532
rect 41368 292528 41432 292592
rect 675156 292436 675220 292500
rect 676628 290940 676692 291004
rect 676260 286996 676324 287060
rect 41828 284820 41892 284884
rect 42012 284276 42076 284340
rect 676076 283596 676140 283660
rect 676076 282644 676140 282708
rect 675708 281616 675772 281620
rect 675708 281560 675722 281616
rect 675722 281560 675772 281616
rect 675708 281556 675772 281560
rect 62252 280060 62316 280124
rect 62068 278020 62132 278084
rect 43668 277612 43732 277676
rect 40724 274212 40788 274276
rect 40540 272988 40604 273052
rect 41460 272172 41524 272236
rect 41828 270056 41892 270060
rect 41828 270000 41842 270056
rect 41842 270000 41892 270056
rect 41828 269996 41892 270000
rect 42012 269104 42076 269108
rect 42012 269048 42026 269104
rect 42026 269048 42076 269104
rect 42012 269044 42076 269048
rect 665220 265508 665284 265572
rect 674788 264148 674852 264212
rect 676996 261564 677060 261628
rect 676812 261156 676876 261220
rect 675524 258088 675588 258092
rect 675524 258032 675538 258088
rect 675538 258032 675588 258088
rect 675524 258028 675588 258032
rect 676996 250276 677060 250340
rect 40540 249732 40604 249796
rect 674788 249596 674852 249660
rect 40724 249324 40788 249388
rect 675524 249596 675588 249660
rect 676812 246604 676876 246668
rect 674604 246196 674668 246260
rect 673316 246060 673380 246124
rect 675340 245788 675404 245852
rect 676812 241980 676876 242044
rect 42012 237356 42076 237420
rect 670740 236676 670804 236740
rect 40540 236540 40604 236604
rect 675340 235180 675404 235244
rect 40724 234636 40788 234700
rect 667060 231100 667124 231164
rect 675156 230420 675220 230484
rect 42012 227352 42076 227356
rect 42012 227296 42026 227352
rect 42026 227296 42076 227352
rect 42012 227292 42076 227296
rect 672580 227020 672644 227084
rect 674052 226748 674116 226812
rect 671660 224768 671724 224772
rect 671660 224712 671674 224768
rect 671674 224712 671724 224768
rect 671660 224708 671724 224712
rect 670556 224496 670620 224500
rect 670556 224440 670570 224496
rect 670570 224440 670620 224496
rect 670556 224436 670620 224440
rect 670004 223892 670068 223956
rect 671660 223952 671724 223956
rect 671660 223896 671674 223952
rect 671674 223896 671724 223952
rect 671660 223892 671724 223896
rect 591988 223484 592052 223548
rect 649580 222940 649644 223004
rect 651972 222940 652036 223004
rect 670004 222260 670068 222324
rect 572300 220552 572364 220556
rect 572300 220496 572314 220552
rect 572314 220496 572364 220552
rect 572300 220492 572364 220496
rect 669268 220144 669332 220148
rect 669268 220088 669318 220144
rect 669318 220088 669332 220144
rect 669268 220084 669332 220088
rect 676030 219812 676094 219876
rect 675708 218588 675772 218652
rect 669636 218180 669700 218244
rect 670556 217908 670620 217972
rect 675892 217908 675956 217972
rect 511028 217560 511092 217564
rect 511028 217504 511042 217560
rect 511042 217504 511092 217560
rect 511028 217500 511092 217504
rect 520044 217560 520108 217564
rect 520044 217504 520058 217560
rect 520058 217504 520108 217560
rect 520044 217500 520108 217504
rect 532556 217560 532620 217564
rect 532556 217504 532570 217560
rect 532570 217504 532620 217560
rect 532556 217500 532620 217504
rect 572300 217560 572364 217564
rect 572300 217504 572314 217560
rect 572314 217504 572364 217560
rect 572300 217500 572364 217504
rect 520044 215868 520108 215932
rect 511028 215596 511092 215660
rect 532556 215324 532620 215388
rect 675892 215460 675956 215524
rect 675892 212468 675956 212532
rect 676628 211380 676692 211444
rect 41460 209748 41524 209812
rect 41644 208932 41708 208996
rect 40724 207300 40788 207364
rect 674604 206892 674668 206956
rect 40908 206484 40972 206548
rect 40540 206076 40604 206140
rect 669268 205668 669332 205732
rect 669636 205668 669700 205732
rect 669268 205396 669332 205460
rect 669636 205396 669700 205460
rect 666508 204172 666572 204236
rect 676444 202676 676508 202740
rect 672580 200772 672644 200836
rect 676628 199956 676692 200020
rect 670740 198732 670804 198796
rect 676812 197916 676876 197980
rect 41828 197780 41892 197844
rect 669268 196148 669332 196212
rect 669636 196148 669700 196212
rect 669268 195876 669332 195940
rect 669636 195876 669700 195940
rect 41828 195800 41892 195804
rect 41828 195744 41878 195800
rect 41878 195744 41892 195800
rect 41828 195740 41892 195744
rect 41644 195468 41708 195532
rect 41460 195196 41524 195260
rect 40724 194924 40788 194988
rect 42196 194924 42260 194988
rect 676260 194516 676324 194580
rect 40908 193428 40972 193492
rect 42380 193216 42444 193220
rect 42380 193160 42394 193216
rect 42394 193160 42444 193216
rect 42380 193156 42444 193160
rect 676076 193156 676140 193220
rect 40540 192748 40604 192812
rect 675892 192748 675956 192812
rect 675156 190028 675220 190092
rect 669452 188396 669516 188460
rect 42380 186280 42444 186284
rect 42380 186224 42394 186280
rect 42394 186224 42444 186280
rect 42380 186220 42444 186224
rect 42196 186008 42260 186012
rect 42196 185952 42210 186008
rect 42210 185952 42260 186008
rect 42196 185948 42260 185952
rect 673132 181520 673196 181524
rect 673132 181464 673146 181520
rect 673146 181464 673196 181520
rect 673132 181460 673196 181464
rect 667980 179556 668044 179620
rect 673316 178060 673380 178124
rect 676812 176608 676876 176672
rect 675892 172756 675956 172820
rect 675892 169356 675956 169420
rect 675340 167452 675404 167516
rect 676628 166424 676692 166428
rect 676628 166368 676642 166424
rect 676642 166368 676692 166424
rect 676628 166364 676692 166368
rect 676076 162692 676140 162756
rect 673132 161468 673196 161532
rect 676444 156980 676508 157044
rect 676260 155756 676324 155820
rect 676628 151404 676692 151468
rect 676076 148412 676140 148476
rect 675340 147656 675404 147660
rect 675340 147600 675390 147656
rect 675390 147600 675404 147656
rect 675340 147596 675404 147600
rect 669268 140388 669332 140452
rect 676628 127332 676692 127396
rect 676076 126924 676140 126988
rect 676260 125700 676324 125764
rect 676444 124068 676508 124132
rect 667060 122028 667124 122092
rect 675340 122028 675404 122092
rect 675708 117268 675772 117332
rect 674052 115772 674116 115836
rect 676628 112372 676692 112436
rect 676260 111692 676324 111756
rect 675708 111344 675772 111348
rect 675708 111288 675758 111344
rect 675758 111288 675772 111344
rect 675708 111284 675772 111288
rect 676444 110332 676508 110396
rect 676076 108156 676140 108220
rect 675340 102640 675404 102644
rect 675340 102584 675390 102640
rect 675390 102584 675404 102640
rect 675340 102580 675404 102584
rect 637252 96868 637316 96932
rect 647188 96460 647252 96524
rect 633940 95372 634004 95436
rect 650316 93060 650380 93124
rect 633940 78568 634004 78572
rect 633940 78512 633954 78568
rect 633954 78512 634004 78568
rect 633940 78508 634004 78512
rect 637068 78100 637132 78164
rect 460796 54980 460860 55044
rect 462636 54708 462700 54772
rect 460796 53892 460860 53956
rect 462636 53680 462700 53684
rect 462636 53624 462650 53680
rect 462650 53624 462700 53680
rect 462636 53620 462700 53624
rect 518756 48860 518820 48924
rect 529612 48044 529676 48108
rect 515444 47772 515508 47836
rect 526484 47772 526548 47836
rect 520964 47500 521028 47564
rect 522068 47228 522132 47292
rect 460980 44432 461044 44436
rect 460980 44376 461030 44432
rect 461030 44376 461044 44432
rect 460980 44372 461044 44376
rect 462268 44372 462332 44436
rect 463740 44432 463804 44436
rect 463740 44376 463790 44432
rect 463790 44376 463804 44432
rect 463740 44372 463804 44376
rect 141740 43964 141804 44028
rect 518756 42800 518820 42804
rect 518756 42744 518806 42800
rect 518806 42744 518820 42800
rect 518756 42740 518820 42744
rect 419212 42060 419276 42124
rect 365116 41848 365180 41852
rect 365116 41792 365130 41848
rect 365130 41792 365180 41848
rect 365116 41788 365180 41792
rect 416636 41848 416700 41852
rect 416636 41792 416686 41848
rect 416686 41792 416700 41848
rect 416636 41788 416700 41792
rect 419948 41848 420012 41852
rect 419948 41792 419962 41848
rect 419962 41792 420012 41848
rect 419948 41788 420012 41792
rect 425100 41788 425164 41852
rect 515444 42120 515508 42124
rect 515444 42064 515458 42120
rect 515458 42064 515508 42120
rect 515444 42060 515508 42064
rect 520964 42120 521028 42124
rect 520964 42064 520978 42120
rect 520978 42064 521028 42120
rect 520964 42060 521028 42064
rect 522068 42120 522132 42124
rect 522068 42064 522082 42120
rect 522082 42064 522132 42120
rect 522068 42060 522132 42064
rect 526484 42120 526548 42124
rect 526484 42064 526498 42120
rect 526498 42064 526548 42120
rect 526484 42060 526548 42064
rect 529612 42120 529676 42124
rect 529612 42064 529626 42120
rect 529626 42064 529676 42120
rect 529612 42060 529676 42064
rect 441844 41788 441908 41852
rect 451964 41788 452028 41852
rect 141740 40352 141804 40356
rect 141740 40296 141754 40352
rect 141754 40296 141804 40352
rect 141740 40292 141804 40296
<< metal4 >>
rect 233003 997388 233069 997389
rect 233003 997324 233004 997388
rect 233068 997324 233069 997388
rect 233003 997323 233069 997324
rect 285443 997388 285509 997389
rect 285443 997324 285444 997388
rect 285508 997324 285509 997388
rect 285443 997323 285509 997324
rect 387563 997388 387629 997389
rect 387563 997324 387564 997388
rect 387628 997324 387629 997388
rect 387563 997323 387629 997324
rect 233006 990997 233066 997323
rect 233003 990996 233069 990997
rect 233003 990932 233004 990996
rect 233068 990932 233069 990996
rect 233003 990931 233069 990932
rect 285446 988005 285506 997323
rect 387566 990997 387626 997323
rect 387563 990996 387629 990997
rect 387563 990932 387564 990996
rect 387628 990932 387629 990996
rect 387563 990931 387629 990932
rect 285443 988004 285509 988005
rect 285443 987940 285444 988004
rect 285508 987940 285509 988004
rect 285443 987939 285509 987940
rect 675891 892260 675957 892261
rect 675891 892196 675892 892260
rect 675956 892196 675957 892260
rect 675891 892195 675957 892196
rect 675894 891510 675954 892195
rect 675710 891450 675954 891510
rect 675710 887090 675770 891450
rect 675891 887772 675957 887773
rect 675891 887708 675892 887772
rect 675956 887770 675957 887772
rect 675956 887710 676322 887770
rect 675956 887708 675957 887710
rect 675891 887707 675957 887708
rect 675710 887030 675954 887090
rect 675707 885868 675773 885869
rect 675707 885804 675708 885868
rect 675772 885804 675773 885868
rect 675707 885803 675773 885804
rect 675523 880700 675589 880701
rect 675523 880636 675524 880700
rect 675588 880636 675589 880700
rect 675523 880635 675589 880636
rect 675339 878524 675405 878525
rect 675339 878460 675340 878524
rect 675404 878460 675405 878524
rect 675339 878459 675405 878460
rect 675342 874173 675402 878459
rect 675339 874172 675405 874173
rect 675339 874108 675340 874172
rect 675404 874108 675405 874172
rect 675339 874107 675405 874108
rect 675526 872190 675586 880635
rect 675710 876890 675770 885803
rect 675894 881850 675954 887030
rect 676262 881850 676322 887710
rect 675894 881790 676138 881850
rect 676262 881790 676506 881850
rect 675710 876830 675954 876890
rect 675526 872130 675770 872190
rect 675710 865741 675770 872130
rect 675707 865740 675773 865741
rect 675707 865676 675708 865740
rect 675772 865676 675773 865740
rect 675707 865675 675773 865676
rect 675894 864925 675954 876830
rect 676078 865469 676138 881790
rect 676259 880428 676325 880429
rect 676259 880364 676260 880428
rect 676324 880364 676325 880428
rect 676259 880363 676325 880364
rect 676262 872813 676322 880363
rect 676446 873085 676506 881790
rect 676443 873084 676509 873085
rect 676443 873020 676444 873084
rect 676508 873020 676509 873084
rect 676443 873019 676509 873020
rect 676259 872812 676325 872813
rect 676259 872748 676260 872812
rect 676324 872748 676325 872812
rect 676259 872747 676325 872748
rect 676075 865468 676141 865469
rect 676075 865404 676076 865468
rect 676140 865404 676141 865468
rect 676075 865403 676141 865404
rect 675891 864924 675957 864925
rect 675891 864860 675892 864924
rect 675956 864860 675957 864924
rect 675891 864859 675957 864860
rect 41827 813244 41893 813245
rect 41827 813180 41828 813244
rect 41892 813180 41893 813244
rect 41827 813179 41893 813180
rect 41830 812970 41890 813179
rect 41462 812910 41890 812970
rect 40539 805628 40605 805629
rect 40539 805564 40540 805628
rect 40604 805564 40605 805628
rect 40539 805563 40605 805564
rect 40542 789309 40602 805563
rect 40723 805220 40789 805221
rect 40723 805156 40724 805220
rect 40788 805156 40789 805220
rect 40723 805155 40789 805156
rect 40726 790669 40786 805155
rect 40907 804812 40973 804813
rect 40907 804748 40908 804812
rect 40972 804748 40973 804812
rect 40907 804747 40973 804748
rect 40910 794885 40970 804747
rect 40907 794884 40973 794885
rect 40907 794820 40908 794884
rect 40972 794820 40973 794884
rect 40907 794819 40973 794820
rect 40723 790668 40789 790669
rect 40723 790604 40724 790668
rect 40788 790604 40789 790668
rect 40723 790603 40789 790604
rect 40539 789308 40605 789309
rect 40539 789244 40540 789308
rect 40604 789244 40605 789308
rect 40539 789243 40605 789244
rect 41462 788357 41522 812910
rect 41827 809980 41893 809981
rect 41827 809916 41828 809980
rect 41892 809916 41893 809980
rect 41827 809915 41893 809916
rect 41830 808710 41890 809915
rect 41646 808650 41890 808710
rect 41646 792029 41706 808650
rect 41827 807940 41893 807941
rect 41827 807876 41828 807940
rect 41892 807876 41893 807940
rect 41827 807875 41893 807876
rect 41830 804813 41890 807875
rect 41827 804812 41893 804813
rect 41827 804748 41828 804812
rect 41892 804748 41893 804812
rect 41827 804747 41893 804748
rect 41827 802500 41893 802501
rect 41827 802436 41828 802500
rect 41892 802436 41893 802500
rect 41827 802435 41893 802436
rect 41643 792028 41709 792029
rect 41643 791964 41644 792028
rect 41708 791964 41709 792028
rect 41643 791963 41709 791964
rect 41459 788356 41525 788357
rect 41459 788292 41460 788356
rect 41524 788292 41525 788356
rect 41459 788291 41525 788292
rect 41830 788085 41890 802435
rect 42195 798148 42261 798149
rect 42195 798084 42196 798148
rect 42260 798084 42261 798148
rect 42195 798083 42261 798084
rect 42198 794477 42258 798083
rect 42195 794476 42261 794477
rect 42195 794412 42196 794476
rect 42260 794412 42261 794476
rect 42195 794411 42261 794412
rect 41827 788084 41893 788085
rect 41827 788020 41828 788084
rect 41892 788020 41893 788084
rect 41827 788019 41893 788020
rect 676075 788084 676141 788085
rect 676075 788020 676076 788084
rect 676140 788020 676141 788084
rect 676075 788019 676141 788020
rect 674419 786724 674485 786725
rect 674419 786660 674420 786724
rect 674484 786660 674485 786724
rect 674419 786659 674485 786660
rect 675339 786724 675405 786725
rect 675339 786660 675340 786724
rect 675404 786660 675405 786724
rect 675339 786659 675405 786660
rect 41643 769860 41709 769861
rect 41643 769796 41644 769860
rect 41708 769796 41709 769860
rect 41643 769795 41709 769796
rect 41459 769044 41525 769045
rect 41459 768980 41460 769044
rect 41524 768980 41525 769044
rect 41459 768979 41525 768980
rect 40539 766596 40605 766597
rect 40539 766532 40540 766596
rect 40604 766532 40605 766596
rect 40539 766531 40605 766532
rect 40542 746741 40602 766531
rect 40723 765372 40789 765373
rect 40723 765308 40724 765372
rect 40788 765308 40789 765372
rect 40723 765307 40789 765308
rect 40726 753949 40786 765307
rect 40907 764964 40973 764965
rect 40907 764900 40908 764964
rect 40972 764900 40973 764964
rect 40907 764899 40973 764900
rect 40723 753948 40789 753949
rect 40723 753884 40724 753948
rect 40788 753884 40789 753948
rect 40723 753883 40789 753884
rect 40910 750549 40970 764899
rect 40907 750548 40973 750549
rect 40907 750484 40908 750548
rect 40972 750484 40973 750548
rect 40907 750483 40973 750484
rect 40539 746740 40605 746741
rect 40539 746676 40540 746740
rect 40604 746676 40605 746740
rect 40539 746675 40605 746676
rect 41462 745109 41522 768979
rect 41646 745653 41706 769795
rect 41827 757756 41893 757757
rect 41827 757692 41828 757756
rect 41892 757692 41893 757756
rect 41827 757691 41893 757692
rect 41643 745652 41709 745653
rect 41643 745588 41644 745652
rect 41708 745588 41709 745652
rect 41643 745587 41709 745588
rect 41459 745108 41525 745109
rect 41459 745044 41460 745108
rect 41524 745044 41525 745108
rect 41459 745043 41525 745044
rect 41830 743069 41890 757691
rect 41827 743068 41893 743069
rect 41827 743004 41828 743068
rect 41892 743004 41893 743068
rect 41827 743003 41893 743004
rect 674235 742524 674301 742525
rect 674235 742460 674236 742524
rect 674300 742460 674301 742524
rect 674235 742459 674301 742460
rect 41827 725932 41893 725933
rect 41827 725930 41828 725932
rect 41646 725870 41828 725930
rect 41646 724530 41706 725870
rect 41827 725868 41828 725870
rect 41892 725868 41893 725932
rect 41827 725867 41893 725868
rect 41827 725660 41893 725661
rect 41827 725596 41828 725660
rect 41892 725596 41893 725660
rect 41827 725595 41893 725596
rect 41462 724470 41706 724530
rect 40723 721772 40789 721773
rect 40723 721708 40724 721772
rect 40788 721708 40789 721772
rect 40723 721707 40789 721708
rect 40539 718588 40605 718589
rect 40539 718524 40540 718588
rect 40604 718524 40605 718588
rect 40539 718523 40605 718524
rect 40542 707981 40602 718523
rect 40539 707980 40605 707981
rect 40539 707916 40540 707980
rect 40604 707916 40605 707980
rect 40539 707915 40605 707916
rect 40726 707437 40786 721707
rect 40723 707436 40789 707437
rect 40723 707372 40724 707436
rect 40788 707372 40789 707436
rect 40723 707371 40789 707372
rect 41462 702133 41522 724470
rect 41830 717630 41890 725595
rect 41646 717570 41890 717630
rect 41646 702813 41706 717570
rect 41827 716956 41893 716957
rect 41827 716892 41828 716956
rect 41892 716892 41893 716956
rect 41827 716891 41893 716892
rect 41643 702812 41709 702813
rect 41643 702748 41644 702812
rect 41708 702748 41709 702812
rect 41643 702747 41709 702748
rect 41459 702132 41525 702133
rect 41459 702068 41460 702132
rect 41524 702068 41525 702132
rect 41459 702067 41525 702068
rect 41830 701861 41890 716891
rect 42011 714508 42077 714509
rect 42011 714444 42012 714508
rect 42076 714444 42077 714508
rect 42011 714443 42077 714444
rect 42014 709885 42074 714443
rect 42011 709884 42077 709885
rect 42011 709820 42012 709884
rect 42076 709820 42077 709884
rect 42011 709819 42077 709820
rect 673867 709340 673933 709341
rect 673867 709276 673868 709340
rect 673932 709276 673933 709340
rect 673867 709275 673933 709276
rect 42195 707980 42261 707981
rect 42195 707916 42196 707980
rect 42260 707916 42261 707980
rect 42195 707915 42261 707916
rect 42198 706213 42258 707915
rect 673870 707029 673930 709275
rect 673867 707028 673933 707029
rect 673867 706964 673868 707028
rect 673932 706964 673933 707028
rect 673867 706963 673933 706964
rect 42195 706212 42261 706213
rect 42195 706148 42196 706212
rect 42260 706148 42261 706212
rect 42195 706147 42261 706148
rect 41827 701860 41893 701861
rect 41827 701796 41828 701860
rect 41892 701796 41893 701860
rect 41827 701795 41893 701796
rect 41827 683636 41893 683637
rect 41827 683572 41828 683636
rect 41892 683572 41893 683636
rect 41827 683571 41893 683572
rect 41830 683090 41890 683571
rect 41462 683030 41890 683090
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40355 670988 40421 670989
rect 40355 670924 40356 670988
rect 40420 670924 40421 670988
rect 40355 670923 40421 670924
rect 40358 667453 40418 670923
rect 40355 667452 40421 667453
rect 40355 667388 40356 667452
rect 40420 667388 40421 667452
rect 40355 667387 40421 667388
rect 40542 664189 40602 678927
rect 40723 677754 40789 677755
rect 40723 677690 40724 677754
rect 40788 677690 40789 677754
rect 40723 677689 40789 677690
rect 40726 665277 40786 677689
rect 40723 665276 40789 665277
rect 40723 665212 40724 665276
rect 40788 665212 40789 665276
rect 40723 665211 40789 665212
rect 40539 664188 40605 664189
rect 40539 664124 40540 664188
rect 40604 664124 40605 664188
rect 40539 664123 40605 664124
rect 41462 657253 41522 683030
rect 674238 682413 674298 742459
rect 674422 726341 674482 786659
rect 674603 738172 674669 738173
rect 674603 738108 674604 738172
rect 674668 738108 674669 738172
rect 674603 738107 674669 738108
rect 674419 726340 674485 726341
rect 674419 726276 674420 726340
rect 674484 726276 674485 726340
rect 674419 726275 674485 726276
rect 674419 694652 674485 694653
rect 674419 694588 674420 694652
rect 674484 694588 674485 694652
rect 674419 694587 674485 694588
rect 674235 682412 674301 682413
rect 674235 682348 674236 682412
rect 674300 682348 674301 682412
rect 674235 682347 674301 682348
rect 41827 681732 41893 681733
rect 41827 681730 41828 681732
rect 41646 681670 41828 681730
rect 41646 658613 41706 681670
rect 41827 681668 41828 681670
rect 41892 681668 41893 681732
rect 41827 681667 41893 681668
rect 42195 673164 42261 673165
rect 42195 673100 42196 673164
rect 42260 673100 42261 673164
rect 42195 673099 42261 673100
rect 41827 672756 41893 672757
rect 41827 672692 41828 672756
rect 41892 672692 41893 672756
rect 41827 672691 41893 672692
rect 41643 658612 41709 658613
rect 41643 658548 41644 658612
rect 41708 658548 41709 658612
rect 41643 658547 41709 658548
rect 41830 658341 41890 672691
rect 42198 668541 42258 673099
rect 42195 668540 42261 668541
rect 42195 668476 42196 668540
rect 42260 668476 42261 668540
rect 42195 668475 42261 668476
rect 41827 658340 41893 658341
rect 41827 658276 41828 658340
rect 41892 658276 41893 658340
rect 41827 658275 41893 658276
rect 41459 657252 41525 657253
rect 41459 657188 41460 657252
rect 41524 657188 41525 657252
rect 41459 657187 41525 657188
rect 674235 652900 674301 652901
rect 674235 652836 674236 652900
rect 674300 652836 674301 652900
rect 674235 652835 674301 652836
rect 41459 640660 41525 640661
rect 41459 640596 41460 640660
rect 41524 640596 41525 640660
rect 41459 640595 41525 640596
rect 40539 635356 40605 635357
rect 40539 635292 40540 635356
rect 40604 635292 40605 635356
rect 40539 635291 40605 635292
rect 40542 620941 40602 635291
rect 40723 634948 40789 634949
rect 40723 634884 40724 634948
rect 40788 634884 40789 634948
rect 40723 634883 40789 634884
rect 40726 623797 40786 634883
rect 40723 623796 40789 623797
rect 40723 623732 40724 623796
rect 40788 623732 40789 623796
rect 40723 623731 40789 623732
rect 40539 620940 40605 620941
rect 40539 620876 40540 620940
rect 40604 620876 40605 620940
rect 40539 620875 40605 620876
rect 41462 616453 41522 640595
rect 41643 629916 41709 629917
rect 41643 629852 41644 629916
rect 41708 629852 41709 629916
rect 41643 629851 41709 629852
rect 41646 616861 41706 629851
rect 41827 629236 41893 629237
rect 41827 629172 41828 629236
rect 41892 629172 41893 629236
rect 41827 629171 41893 629172
rect 41643 616860 41709 616861
rect 41643 616796 41644 616860
rect 41708 616796 41709 616860
rect 41643 616795 41709 616796
rect 41459 616452 41525 616453
rect 41459 616388 41460 616452
rect 41524 616388 41525 616452
rect 41459 616387 41525 616388
rect 41830 615501 41890 629171
rect 42195 625972 42261 625973
rect 42195 625908 42196 625972
rect 42260 625908 42261 625972
rect 42195 625907 42261 625908
rect 42198 620261 42258 625907
rect 42195 620260 42261 620261
rect 42195 620196 42196 620260
rect 42260 620196 42261 620260
rect 42195 620195 42261 620196
rect 673867 616180 673933 616181
rect 673867 616116 673868 616180
rect 673932 616116 673933 616180
rect 673867 616115 673933 616116
rect 41827 615500 41893 615501
rect 41827 615436 41828 615500
rect 41892 615436 41893 615500
rect 41827 615435 41893 615436
rect 40539 612372 40605 612373
rect 40539 612308 40540 612372
rect 40604 612308 40605 612372
rect 40539 612307 40605 612308
rect 40542 602037 40602 612307
rect 40539 602036 40605 602037
rect 40539 601972 40540 602036
rect 40604 601972 40605 602036
rect 40539 601971 40605 601972
rect 42931 598500 42997 598501
rect 42931 598436 42932 598500
rect 42996 598436 42997 598500
rect 42931 598435 42997 598436
rect 40355 597038 40421 597039
rect 40355 596974 40356 597038
rect 40420 596974 40421 597038
rect 42934 597005 42994 598435
rect 40355 596973 40421 596974
rect 42931 597004 42997 597005
rect 40358 588845 40418 596973
rect 42931 596940 42932 597004
rect 42996 596940 42997 597004
rect 42931 596939 42997 596940
rect 42011 596460 42077 596461
rect 42011 596396 42012 596460
rect 42076 596396 42077 596460
rect 42011 596395 42077 596396
rect 41781 594012 41847 594013
rect 41781 594010 41782 594012
rect 40542 593950 41782 594010
rect 40355 588844 40421 588845
rect 40355 588780 40356 588844
rect 40420 588780 40421 588844
rect 40355 588779 40421 588780
rect 40355 584628 40421 584629
rect 40355 584564 40356 584628
rect 40420 584564 40421 584628
rect 40355 584563 40421 584564
rect 40358 580277 40418 584563
rect 40355 580276 40421 580277
rect 40355 580212 40356 580276
rect 40420 580212 40421 580276
rect 40355 580211 40421 580212
rect 40542 575789 40602 593950
rect 41781 593948 41782 593950
rect 41846 593948 41847 594012
rect 41781 593947 41847 593948
rect 41781 592788 41847 592789
rect 41781 592724 41782 592788
rect 41846 592724 41847 592788
rect 41781 592723 41847 592724
rect 41784 592514 41844 592723
rect 40726 592454 41844 592514
rect 40539 575788 40605 575789
rect 40539 575724 40540 575788
rect 40604 575724 40605 575788
rect 40539 575723 40605 575724
rect 40726 574701 40786 592454
rect 40907 589116 40973 589117
rect 40907 589052 40908 589116
rect 40972 589052 40973 589116
rect 40907 589051 40973 589052
rect 40910 577829 40970 589051
rect 41459 588844 41525 588845
rect 41459 588780 41460 588844
rect 41524 588780 41525 588844
rect 41459 588779 41525 588780
rect 40907 577828 40973 577829
rect 40907 577764 40908 577828
rect 40972 577764 40973 577828
rect 40907 577763 40973 577764
rect 40723 574700 40789 574701
rect 40723 574636 40724 574700
rect 40788 574636 40789 574700
rect 40723 574635 40789 574636
rect 41462 572933 41522 588779
rect 42014 587910 42074 596395
rect 41830 587850 42074 587910
rect 41830 587210 41890 587850
rect 41646 587150 41890 587210
rect 41459 572932 41525 572933
rect 41459 572868 41460 572932
rect 41524 572868 41525 572932
rect 41459 572867 41525 572868
rect 41646 571573 41706 587150
rect 41827 585988 41893 585989
rect 41827 585924 41828 585988
rect 41892 585924 41893 585988
rect 41827 585923 41893 585924
rect 41643 571572 41709 571573
rect 41643 571508 41644 571572
rect 41708 571508 41709 571572
rect 41643 571507 41709 571508
rect 41830 570213 41890 585923
rect 62067 585716 62133 585717
rect 62067 585652 62068 585716
rect 62132 585652 62133 585716
rect 62067 585651 62133 585652
rect 42195 582452 42261 582453
rect 42195 582388 42196 582452
rect 42260 582388 42261 582452
rect 42195 582387 42261 582388
rect 42198 580277 42258 582387
rect 42195 580276 42261 580277
rect 42195 580212 42196 580276
rect 42260 580212 42261 580276
rect 42195 580211 42261 580212
rect 42011 579324 42077 579325
rect 42011 579260 42012 579324
rect 42076 579260 42077 579324
rect 42011 579259 42077 579260
rect 42014 572661 42074 579259
rect 42011 572660 42077 572661
rect 42011 572596 42012 572660
rect 42076 572596 42077 572660
rect 42011 572595 42077 572596
rect 41827 570212 41893 570213
rect 41827 570148 41828 570212
rect 41892 570148 41893 570212
rect 41827 570147 41893 570148
rect 41091 558788 41157 558789
rect 41091 558724 41092 558788
rect 41156 558724 41157 558788
rect 41091 558723 41157 558724
rect 41094 557553 41154 558723
rect 41091 557552 41157 557553
rect 41091 557488 41092 557552
rect 41156 557488 41157 557552
rect 41091 557487 41157 557488
rect 41827 554028 41893 554029
rect 41827 553964 41828 554028
rect 41892 553964 41893 554028
rect 41827 553963 41893 553964
rect 41830 553410 41890 553963
rect 41462 553350 41890 553410
rect 40723 545596 40789 545597
rect 40723 545532 40724 545596
rect 40788 545532 40789 545596
rect 40723 545531 40789 545532
rect 40539 545324 40605 545325
rect 40539 545260 40540 545324
rect 40604 545260 40605 545324
rect 40539 545259 40605 545260
rect 40542 533357 40602 545259
rect 40726 539613 40786 545531
rect 40723 539612 40789 539613
rect 40723 539548 40724 539612
rect 40788 539548 40789 539612
rect 40723 539547 40789 539548
rect 40539 533356 40605 533357
rect 40539 533292 40540 533356
rect 40604 533292 40605 533356
rect 40539 533291 40605 533292
rect 41462 530229 41522 553350
rect 41827 552804 41893 552805
rect 41827 552740 41828 552804
rect 41892 552740 41893 552804
rect 41827 552739 41893 552740
rect 41830 543750 41890 552739
rect 42011 549540 42077 549541
rect 42011 549476 42012 549540
rect 42076 549476 42077 549540
rect 42011 549475 42077 549476
rect 42014 545325 42074 549475
rect 42011 545324 42077 545325
rect 42011 545260 42012 545324
rect 42076 545260 42077 545324
rect 42011 545259 42077 545260
rect 41646 543690 41890 543750
rect 41646 531725 41706 543690
rect 41827 542332 41893 542333
rect 41827 542268 41828 542332
rect 41892 542268 41893 542332
rect 41827 542267 41893 542268
rect 41643 531724 41709 531725
rect 41643 531660 41644 531724
rect 41708 531660 41709 531724
rect 41643 531659 41709 531660
rect 41459 530228 41525 530229
rect 41459 530164 41460 530228
rect 41524 530164 41525 530228
rect 41459 530163 41525 530164
rect 41830 529005 41890 542267
rect 41827 529004 41893 529005
rect 41827 528940 41828 529004
rect 41892 528940 41893 529004
rect 41827 528939 41893 528940
rect 41459 426630 41525 426631
rect 41459 426566 41460 426630
rect 41524 426566 41525 426630
rect 41459 426565 41525 426566
rect 40907 422312 40973 422313
rect 40907 422248 40908 422312
rect 40972 422248 40973 422312
rect 40907 422247 40973 422248
rect 40723 418708 40789 418709
rect 40723 418644 40724 418708
rect 40788 418644 40789 418708
rect 40723 418643 40789 418644
rect 40539 418436 40605 418437
rect 40539 418372 40540 418436
rect 40604 418372 40605 418436
rect 40539 418371 40605 418372
rect 40542 406741 40602 418371
rect 40539 406740 40605 406741
rect 40539 406676 40540 406740
rect 40604 406676 40605 406740
rect 40539 406675 40605 406676
rect 40726 404565 40786 418643
rect 40910 407013 40970 422247
rect 40907 407012 40973 407013
rect 40907 406948 40908 407012
rect 40972 406948 40973 407012
rect 40907 406947 40973 406948
rect 40723 404564 40789 404565
rect 40723 404500 40724 404564
rect 40788 404500 40789 404564
rect 40723 404499 40789 404500
rect 41462 400077 41522 426565
rect 41827 421564 41893 421565
rect 41827 421500 41828 421564
rect 41892 421500 41893 421564
rect 41827 421499 41893 421500
rect 41830 418437 41890 421499
rect 41827 418436 41893 418437
rect 41827 418372 41828 418436
rect 41892 418372 41893 418436
rect 41827 418371 41893 418372
rect 41643 415308 41709 415309
rect 41643 415244 41644 415308
rect 41708 415244 41709 415308
rect 41643 415243 41709 415244
rect 41646 402990 41706 415243
rect 42011 414628 42077 414629
rect 42011 414564 42012 414628
rect 42076 414564 42077 414628
rect 42011 414563 42077 414564
rect 41646 402930 41890 402990
rect 41459 400076 41525 400077
rect 41459 400012 41460 400076
rect 41524 400012 41525 400076
rect 41459 400011 41525 400012
rect 41830 398853 41890 402930
rect 42014 399397 42074 414563
rect 42011 399396 42077 399397
rect 42011 399332 42012 399396
rect 42076 399332 42077 399396
rect 42011 399331 42077 399332
rect 41827 398852 41893 398853
rect 41827 398788 41828 398852
rect 41892 398788 41893 398852
rect 41827 398787 41893 398788
rect 41459 381852 41525 381853
rect 41459 381788 41460 381852
rect 41524 381788 41525 381852
rect 41459 381787 41525 381788
rect 40723 378996 40789 378997
rect 40723 378932 40724 378996
rect 40788 378932 40789 378996
rect 40723 378931 40789 378932
rect 40539 378588 40605 378589
rect 40539 378524 40540 378588
rect 40604 378524 40605 378588
rect 40539 378523 40605 378524
rect 40542 360093 40602 378523
rect 40726 364173 40786 378931
rect 40907 377772 40973 377773
rect 40907 377708 40908 377772
rect 40972 377708 40973 377772
rect 40907 377707 40973 377708
rect 40910 364853 40970 377707
rect 40907 364852 40973 364853
rect 40907 364788 40908 364852
rect 40972 364788 40973 364852
rect 40907 364787 40973 364788
rect 40723 364172 40789 364173
rect 40723 364108 40724 364172
rect 40788 364108 40789 364172
rect 40723 364107 40789 364108
rect 40539 360092 40605 360093
rect 40539 360028 40540 360092
rect 40604 360028 40605 360092
rect 40539 360027 40605 360028
rect 41462 356965 41522 381787
rect 41827 379404 41893 379405
rect 41827 379340 41828 379404
rect 41892 379340 41893 379404
rect 41827 379339 41893 379340
rect 41643 374644 41709 374645
rect 41643 374580 41644 374644
rect 41708 374580 41709 374644
rect 41643 374579 41709 374580
rect 41646 360210 41706 374579
rect 41830 365805 41890 379339
rect 41827 365804 41893 365805
rect 41827 365740 41828 365804
rect 41892 365740 41893 365804
rect 41827 365739 41893 365740
rect 41646 360150 41890 360210
rect 41830 358733 41890 360150
rect 41827 358732 41893 358733
rect 41827 358668 41828 358732
rect 41892 358668 41893 358732
rect 41827 358667 41893 358668
rect 41459 356964 41525 356965
rect 41459 356900 41460 356964
rect 41524 356900 41525 356964
rect 41459 356899 41525 356900
rect 43667 354652 43733 354653
rect 43667 354588 43668 354652
rect 43732 354588 43733 354652
rect 43667 354587 43733 354588
rect 42011 351932 42077 351933
rect 42011 351868 42012 351932
rect 42076 351868 42077 351932
rect 42011 351867 42077 351868
rect 40539 336972 40605 336973
rect 40539 336908 40540 336972
rect 40604 336908 40605 336972
rect 40539 336907 40605 336908
rect 40542 316029 40602 336907
rect 40723 336564 40789 336565
rect 40723 336500 40724 336564
rect 40788 336500 40789 336564
rect 40723 336499 40789 336500
rect 40726 317525 40786 336499
rect 40907 336156 40973 336157
rect 40907 336092 40908 336156
rect 40972 336092 40973 336156
rect 40907 336091 40973 336092
rect 40910 322829 40970 336091
rect 41275 334932 41341 334933
rect 41275 334868 41276 334932
rect 41340 334868 41341 334932
rect 41275 334867 41341 334868
rect 41278 334525 41338 334867
rect 42014 334661 42074 351867
rect 42195 335748 42261 335749
rect 42195 335684 42196 335748
rect 42260 335684 42261 335748
rect 42195 335683 42261 335684
rect 42011 334660 42077 334661
rect 42011 334596 42012 334660
rect 42076 334596 42077 334660
rect 42011 334595 42077 334596
rect 41275 334524 41341 334525
rect 41275 334460 41276 334524
rect 41340 334460 41341 334524
rect 41275 334459 41341 334460
rect 41827 332892 41893 332893
rect 41827 332828 41828 332892
rect 41892 332828 41893 332892
rect 41827 332827 41893 332828
rect 41643 331804 41709 331805
rect 41643 331740 41644 331804
rect 41708 331740 41709 331804
rect 41643 331739 41709 331740
rect 40907 322828 40973 322829
rect 40907 322764 40908 322828
rect 40972 322764 40973 322828
rect 40907 322763 40973 322764
rect 40723 317524 40789 317525
rect 40723 317460 40724 317524
rect 40788 317460 40789 317524
rect 40723 317459 40789 317460
rect 41646 316050 41706 331739
rect 41830 324869 41890 332827
rect 41827 324868 41893 324869
rect 41827 324804 41828 324868
rect 41892 324804 41893 324868
rect 41827 324803 41893 324804
rect 40539 316028 40605 316029
rect 40539 315964 40540 316028
rect 40604 315964 40605 316028
rect 41646 315990 41890 316050
rect 40539 315963 40605 315964
rect 41830 315621 41890 315990
rect 41827 315620 41893 315621
rect 41827 315556 41828 315620
rect 41892 315556 41893 315620
rect 41827 315555 41893 315556
rect 42198 313717 42258 335683
rect 42195 313716 42261 313717
rect 42195 313652 42196 313716
rect 42260 313652 42261 313716
rect 42195 313651 42261 313652
rect 41827 295628 41893 295629
rect 41827 295564 41828 295628
rect 41892 295564 41893 295628
rect 41827 295563 41893 295564
rect 40539 292592 40605 292593
rect 40539 292528 40540 292592
rect 40604 292528 40605 292592
rect 40539 292527 40605 292528
rect 41367 292592 41433 292593
rect 41367 292528 41368 292592
rect 41432 292528 41433 292592
rect 41830 292590 41890 295563
rect 41367 292527 41433 292528
rect 41646 292530 41890 292590
rect 40542 273053 40602 292527
rect 41370 292090 41430 292527
rect 40726 292030 41430 292090
rect 40726 274277 40786 292030
rect 40723 274276 40789 274277
rect 40723 274212 40724 274276
rect 40788 274212 40789 274276
rect 40723 274211 40789 274212
rect 41646 273270 41706 292530
rect 41827 284884 41893 284885
rect 41827 284820 41828 284884
rect 41892 284820 41893 284884
rect 41827 284819 41893 284820
rect 41462 273210 41706 273270
rect 40539 273052 40605 273053
rect 40539 272988 40540 273052
rect 40604 272988 40605 273052
rect 40539 272987 40605 272988
rect 41462 272237 41522 273210
rect 41459 272236 41525 272237
rect 41459 272172 41460 272236
rect 41524 272172 41525 272236
rect 41459 272171 41525 272172
rect 41830 270061 41890 284819
rect 42011 284340 42077 284341
rect 42011 284276 42012 284340
rect 42076 284276 42077 284340
rect 42011 284275 42077 284276
rect 41827 270060 41893 270061
rect 41827 269996 41828 270060
rect 41892 269996 41893 270060
rect 41827 269995 41893 269996
rect 42014 269109 42074 284275
rect 43670 277677 43730 354587
rect 44771 353700 44837 353701
rect 44771 353636 44772 353700
rect 44836 353636 44837 353700
rect 44771 353635 44837 353636
rect 44774 353290 44834 353635
rect 43854 353230 44834 353290
rect 43854 334661 43914 353230
rect 44035 352204 44101 352205
rect 44035 352140 44036 352204
rect 44100 352140 44101 352204
rect 44035 352139 44101 352140
rect 43851 334660 43917 334661
rect 43851 334596 43852 334660
rect 43916 334596 43917 334660
rect 43851 334595 43917 334596
rect 44038 334525 44098 352139
rect 50107 342140 50173 342141
rect 50107 342076 50108 342140
rect 50172 342076 50173 342140
rect 50107 342075 50173 342076
rect 50110 341730 50170 342075
rect 50475 341732 50541 341733
rect 50475 341730 50476 341732
rect 50110 341670 50476 341730
rect 50475 341668 50476 341670
rect 50540 341668 50541 341732
rect 50475 341667 50541 341668
rect 44219 339828 44285 339829
rect 44219 339764 44220 339828
rect 44284 339764 44285 339828
rect 44219 339763 44285 339764
rect 44035 334524 44101 334525
rect 44035 334460 44036 334524
rect 44100 334460 44101 334524
rect 44035 334459 44101 334460
rect 44222 311269 44282 339763
rect 44403 339284 44469 339285
rect 44403 339220 44404 339284
rect 44468 339220 44469 339284
rect 44403 339219 44469 339220
rect 44406 311949 44466 339219
rect 44587 335476 44653 335477
rect 44587 335412 44588 335476
rect 44652 335412 44653 335476
rect 44587 335411 44653 335412
rect 44590 334389 44650 335411
rect 44587 334388 44653 334389
rect 44587 334324 44588 334388
rect 44652 334324 44653 334388
rect 44587 334323 44653 334324
rect 44403 311948 44469 311949
rect 44403 311884 44404 311948
rect 44468 311884 44469 311948
rect 44403 311883 44469 311884
rect 44219 311268 44285 311269
rect 44219 311204 44220 311268
rect 44284 311204 44285 311268
rect 44219 311203 44285 311204
rect 62070 278085 62130 585651
rect 673683 553484 673749 553485
rect 673683 553420 673684 553484
rect 673748 553420 673749 553484
rect 673683 553419 673749 553420
rect 673686 551581 673746 553419
rect 673683 551580 673749 551581
rect 673683 551516 673684 551580
rect 673748 551516 673749 551580
rect 673683 551515 673749 551516
rect 673499 535124 673565 535125
rect 673499 535060 673500 535124
rect 673564 535060 673565 535124
rect 673499 535059 673565 535060
rect 673502 534309 673562 535059
rect 673499 534308 673565 534309
rect 673499 534244 673500 534308
rect 673564 534244 673565 534308
rect 673499 534243 673565 534244
rect 673870 455293 673930 616115
rect 674238 591293 674298 652835
rect 674422 618765 674482 694587
rect 674606 662421 674666 738107
rect 675342 730149 675402 786659
rect 675339 730148 675405 730149
rect 675339 730084 675340 730148
rect 675404 730084 675405 730148
rect 675339 730083 675405 730084
rect 676078 726613 676138 788019
rect 676811 729876 676877 729877
rect 676811 729812 676812 729876
rect 676876 729812 676877 729876
rect 676811 729811 676877 729812
rect 676075 726612 676141 726613
rect 676075 726548 676076 726612
rect 676140 726548 676141 726612
rect 676075 726547 676141 726548
rect 675155 723212 675221 723213
rect 675155 723148 675156 723212
rect 675220 723148 675221 723212
rect 675155 723147 675221 723148
rect 675158 717630 675218 723147
rect 675158 717570 675402 717630
rect 675342 683773 675402 717570
rect 675523 696828 675589 696829
rect 675523 696764 675524 696828
rect 675588 696764 675589 696828
rect 675523 696763 675589 696764
rect 675526 684045 675586 696763
rect 675523 684044 675589 684045
rect 675523 683980 675524 684044
rect 675588 683980 675589 684044
rect 675523 683979 675589 683980
rect 675339 683772 675405 683773
rect 675339 683708 675340 683772
rect 675404 683708 675405 683772
rect 675339 683707 675405 683708
rect 676075 676428 676141 676429
rect 676075 676364 676076 676428
rect 676140 676364 676141 676428
rect 676075 676363 676141 676364
rect 674603 662420 674669 662421
rect 674603 662356 674604 662420
rect 674668 662356 674669 662420
rect 674603 662355 674669 662356
rect 676078 637533 676138 676363
rect 676814 665821 676874 729811
rect 676811 665820 676877 665821
rect 676811 665756 676812 665820
rect 676876 665756 676877 665820
rect 676811 665755 676877 665756
rect 676075 637532 676141 637533
rect 676075 637468 676076 637532
rect 676140 637468 676141 637532
rect 676075 637467 676141 637468
rect 675155 631412 675221 631413
rect 675155 631348 675156 631412
rect 675220 631348 675221 631412
rect 675155 631347 675221 631348
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 674419 618764 674485 618765
rect 674419 618700 674420 618764
rect 674484 618700 674485 618764
rect 674419 618699 674485 618700
rect 674419 602988 674485 602989
rect 674419 602924 674420 602988
rect 674484 602924 674485 602988
rect 674419 602923 674485 602924
rect 674235 591292 674301 591293
rect 674235 591228 674236 591292
rect 674300 591228 674301 591292
rect 674235 591227 674301 591228
rect 674422 547093 674482 602923
rect 675158 593197 675218 631347
rect 675155 593196 675221 593197
rect 675155 593132 675156 593196
rect 675220 593132 675221 593196
rect 675155 593131 675221 593132
rect 676078 591701 676138 631347
rect 676259 617132 676325 617133
rect 676259 617068 676260 617132
rect 676324 617068 676325 617132
rect 676259 617067 676325 617068
rect 676262 615510 676322 617067
rect 676262 615450 676874 615510
rect 676075 591700 676141 591701
rect 676075 591636 676076 591700
rect 676140 591636 676141 591700
rect 676075 591635 676141 591636
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675339 561916 675405 561917
rect 675339 561852 675340 561916
rect 675404 561852 675405 561916
rect 675339 561851 675405 561852
rect 674971 548860 675037 548861
rect 674971 548796 674972 548860
rect 675036 548796 675037 548860
rect 674971 548795 675037 548796
rect 674974 547909 675034 548795
rect 674971 547908 675037 547909
rect 674971 547844 674972 547908
rect 675036 547844 675037 547908
rect 674971 547843 675037 547844
rect 674419 547092 674485 547093
rect 674419 547028 674420 547092
rect 674484 547028 674485 547092
rect 674419 547027 674485 547028
rect 675342 545869 675402 561851
rect 676078 546821 676138 586195
rect 676814 576877 676874 615450
rect 676811 576876 676877 576877
rect 676811 576812 676812 576876
rect 676876 576812 676877 576876
rect 676811 576811 676877 576812
rect 676259 557564 676325 557565
rect 676259 557500 676260 557564
rect 676324 557500 676325 557564
rect 676259 557499 676325 557500
rect 676262 547637 676322 557499
rect 676811 553892 676877 553893
rect 676811 553828 676812 553892
rect 676876 553828 676877 553892
rect 676811 553827 676877 553828
rect 676259 547636 676325 547637
rect 676259 547572 676260 547636
rect 676324 547572 676325 547636
rect 676259 547571 676325 547572
rect 676075 546820 676141 546821
rect 676075 546756 676076 546820
rect 676140 546756 676141 546820
rect 676075 546755 676141 546756
rect 675339 545868 675405 545869
rect 675339 545804 675340 545868
rect 675404 545804 675405 545868
rect 675339 545803 675405 545804
rect 676814 500989 676874 553827
rect 676995 548316 677061 548317
rect 676995 548252 676996 548316
rect 677060 548252 677061 548316
rect 676995 548251 677061 548252
rect 676998 503709 677058 548251
rect 676995 503708 677061 503709
rect 676995 503644 676996 503708
rect 677060 503644 677061 503708
rect 676995 503643 677061 503644
rect 676811 500988 676877 500989
rect 676811 500924 676812 500988
rect 676876 500924 676877 500988
rect 676811 500923 676877 500924
rect 675894 489230 676138 489290
rect 675894 488885 675954 489230
rect 675891 488884 675957 488885
rect 675891 488820 675892 488884
rect 675956 488820 675957 488884
rect 675891 488819 675957 488820
rect 676078 488610 676138 489230
rect 676078 488550 676506 488610
rect 675891 487932 675957 487933
rect 675891 487868 675892 487932
rect 675956 487930 675957 487932
rect 676446 487930 676506 488550
rect 675956 487870 676322 487930
rect 676446 487870 677058 487930
rect 675956 487868 675957 487870
rect 675891 487867 675957 487868
rect 676262 483030 676322 487870
rect 676998 483030 677058 487870
rect 676262 482970 676874 483030
rect 676998 482970 677242 483030
rect 673867 455292 673933 455293
rect 673867 455228 673868 455292
rect 673932 455228 673933 455292
rect 673867 455227 673933 455228
rect 676814 400485 676874 482970
rect 677182 401301 677242 482970
rect 677179 401300 677245 401301
rect 677179 401236 677180 401300
rect 677244 401236 677245 401300
rect 677179 401235 677245 401236
rect 676811 400484 676877 400485
rect 676811 400420 676812 400484
rect 676876 400420 676877 400484
rect 676811 400419 676877 400420
rect 676075 398852 676141 398853
rect 676075 398788 676076 398852
rect 676140 398788 676141 398852
rect 676075 398787 676141 398788
rect 675891 392868 675957 392869
rect 675891 392804 675892 392868
rect 675956 392804 675957 392868
rect 675891 392803 675957 392804
rect 675707 387700 675773 387701
rect 675707 387636 675708 387700
rect 675772 387636 675773 387700
rect 675707 387635 675773 387636
rect 675710 378725 675770 387635
rect 675707 378724 675773 378725
rect 675707 378660 675708 378724
rect 675772 378660 675773 378724
rect 675707 378659 675773 378660
rect 675894 374010 675954 392803
rect 675342 373950 675954 374010
rect 675342 372469 675402 373950
rect 676078 373693 676138 398787
rect 676259 396812 676325 396813
rect 676259 396748 676260 396812
rect 676324 396748 676325 396812
rect 676259 396747 676325 396748
rect 676262 384981 676322 396747
rect 676443 396404 676509 396405
rect 676443 396340 676444 396404
rect 676508 396340 676509 396404
rect 676443 396339 676509 396340
rect 676259 384980 676325 384981
rect 676259 384916 676260 384980
rect 676324 384916 676325 384980
rect 676259 384915 676325 384916
rect 676446 382261 676506 396339
rect 676627 395180 676693 395181
rect 676627 395116 676628 395180
rect 676692 395116 676693 395180
rect 676627 395115 676693 395116
rect 676443 382260 676509 382261
rect 676443 382196 676444 382260
rect 676508 382196 676509 382260
rect 676443 382195 676509 382196
rect 676630 377365 676690 395115
rect 676627 377364 676693 377365
rect 676627 377300 676628 377364
rect 676692 377300 676693 377364
rect 676627 377299 676693 377300
rect 676075 373692 676141 373693
rect 676075 373628 676076 373692
rect 676140 373628 676141 373692
rect 676075 373627 676141 373628
rect 675339 372468 675405 372469
rect 675339 372404 675340 372468
rect 675404 372404 675405 372468
rect 675339 372403 675405 372404
rect 675342 365669 675402 372403
rect 675339 365668 675405 365669
rect 675339 365604 675340 365668
rect 675404 365604 675405 365668
rect 675339 365603 675405 365604
rect 675523 354244 675589 354245
rect 675523 354180 675524 354244
rect 675588 354180 675589 354244
rect 675523 354179 675589 354180
rect 675339 347716 675405 347717
rect 675339 347652 675340 347716
rect 675404 347652 675405 347716
rect 675339 347651 675405 347652
rect 675342 327997 675402 347651
rect 675526 339421 675586 354179
rect 675891 353836 675957 353837
rect 675891 353772 675892 353836
rect 675956 353772 675957 353836
rect 675891 353771 675957 353772
rect 675894 353290 675954 353771
rect 675894 353230 676690 353290
rect 675707 353020 675773 353021
rect 675707 352956 675708 353020
rect 675772 352956 675773 353020
rect 675707 352955 675773 352956
rect 675710 349210 675770 352955
rect 675891 351796 675957 351797
rect 675891 351732 675892 351796
rect 675956 351732 675957 351796
rect 675891 351731 675957 351732
rect 675894 349890 675954 351731
rect 675894 349830 676322 349890
rect 675710 349150 676138 349210
rect 675523 339420 675589 339421
rect 675523 339356 675524 339420
rect 675588 339356 675589 339420
rect 675523 339355 675589 339356
rect 676078 337925 676138 349150
rect 676262 340237 676322 349830
rect 676443 346628 676509 346629
rect 676443 346564 676444 346628
rect 676508 346564 676509 346628
rect 676443 346563 676509 346564
rect 676259 340236 676325 340237
rect 676259 340172 676260 340236
rect 676324 340172 676325 340236
rect 676259 340171 676325 340172
rect 676075 337924 676141 337925
rect 676075 337860 676076 337924
rect 676140 337860 676141 337924
rect 676075 337859 676141 337860
rect 676446 336565 676506 346563
rect 676443 336564 676509 336565
rect 676443 336500 676444 336564
rect 676508 336500 676509 336564
rect 676443 336499 676509 336500
rect 675339 327996 675405 327997
rect 675339 327932 675340 327996
rect 675404 327932 675405 327996
rect 675339 327931 675405 327932
rect 62251 327724 62317 327725
rect 62251 327660 62252 327724
rect 62316 327660 62317 327724
rect 62251 327659 62317 327660
rect 62254 325710 62314 327659
rect 62254 325650 63050 325710
rect 676630 325685 676690 353230
rect 62990 296730 63050 325650
rect 676627 325684 676693 325685
rect 676627 325620 676628 325684
rect 676692 325620 676693 325684
rect 676627 325619 676693 325620
rect 675342 309710 675770 309770
rect 675342 309229 675402 309710
rect 675339 309228 675405 309229
rect 675339 309164 675340 309228
rect 675404 309164 675405 309228
rect 675339 309163 675405 309164
rect 675710 309090 675770 309710
rect 675710 309030 676506 309090
rect 675891 308820 675957 308821
rect 675891 308756 675892 308820
rect 675956 308756 675957 308820
rect 675891 308755 675957 308756
rect 675894 303650 675954 308755
rect 676075 304604 676141 304605
rect 676075 304540 676076 304604
rect 676140 304540 676141 304604
rect 676075 304539 676141 304540
rect 676078 304330 676138 304539
rect 676078 304270 676322 304330
rect 675894 303590 676138 303650
rect 675891 302700 675957 302701
rect 675891 302636 675892 302700
rect 675956 302636 675957 302700
rect 675891 302635 675957 302636
rect 675155 298212 675221 298213
rect 675155 298148 675156 298212
rect 675220 298148 675221 298212
rect 675155 298147 675221 298148
rect 62254 296670 63050 296730
rect 62254 280125 62314 296670
rect 675158 292501 675218 298147
rect 675523 297668 675589 297669
rect 675523 297604 675524 297668
rect 675588 297604 675589 297668
rect 675523 297603 675589 297604
rect 675526 295765 675586 297603
rect 675707 297396 675773 297397
rect 675707 297332 675708 297396
rect 675772 297332 675773 297396
rect 675707 297331 675773 297332
rect 675523 295764 675589 295765
rect 675523 295700 675524 295764
rect 675588 295700 675589 295764
rect 675523 295699 675589 295700
rect 675155 292500 675221 292501
rect 675155 292436 675156 292500
rect 675220 292436 675221 292500
rect 675155 292435 675221 292436
rect 675710 281621 675770 297331
rect 675894 282930 675954 302635
rect 676078 283661 676138 303590
rect 676262 287061 676322 304270
rect 676446 294677 676506 309030
rect 676627 301612 676693 301613
rect 676627 301548 676628 301612
rect 676692 301548 676693 301612
rect 676627 301547 676693 301548
rect 676443 294676 676509 294677
rect 676443 294612 676444 294676
rect 676508 294612 676509 294676
rect 676443 294611 676509 294612
rect 676630 291005 676690 301547
rect 676627 291004 676693 291005
rect 676627 290940 676628 291004
rect 676692 290940 676693 291004
rect 676627 290939 676693 290940
rect 676259 287060 676325 287061
rect 676259 286996 676260 287060
rect 676324 286996 676325 287060
rect 676259 286995 676325 286996
rect 676075 283660 676141 283661
rect 676075 283596 676076 283660
rect 676140 283596 676141 283660
rect 676075 283595 676141 283596
rect 675894 282870 676138 282930
rect 676078 282709 676138 282870
rect 676075 282708 676141 282709
rect 676075 282644 676076 282708
rect 676140 282644 676141 282708
rect 676075 282643 676141 282644
rect 675707 281620 675773 281621
rect 675707 281556 675708 281620
rect 675772 281556 675773 281620
rect 675707 281555 675773 281556
rect 62251 280124 62317 280125
rect 62251 280060 62252 280124
rect 62316 280060 62317 280124
rect 62251 280059 62317 280060
rect 62067 278084 62133 278085
rect 62067 278020 62068 278084
rect 62132 278020 62133 278084
rect 62067 278019 62133 278020
rect 43667 277676 43733 277677
rect 43667 277612 43668 277676
rect 43732 277612 43733 277676
rect 43667 277611 43733 277612
rect 42011 269108 42077 269109
rect 42011 269044 42012 269108
rect 42076 269044 42077 269108
rect 42011 269043 42077 269044
rect 665219 265572 665285 265573
rect 665219 265508 665220 265572
rect 665284 265508 665285 265572
rect 665219 265507 665285 265508
rect 40539 249796 40605 249797
rect 40539 249732 40540 249796
rect 40604 249732 40605 249796
rect 40539 249731 40605 249732
rect 40542 236605 40602 249731
rect 40723 249388 40789 249389
rect 40723 249324 40724 249388
rect 40788 249324 40789 249388
rect 40723 249323 40789 249324
rect 40539 236604 40605 236605
rect 40539 236540 40540 236604
rect 40604 236540 40605 236604
rect 40539 236539 40605 236540
rect 40726 234701 40786 249323
rect 42011 237420 42077 237421
rect 42011 237356 42012 237420
rect 42076 237356 42077 237420
rect 42011 237355 42077 237356
rect 40723 234700 40789 234701
rect 40723 234636 40724 234700
rect 40788 234636 40789 234700
rect 40723 234635 40789 234636
rect 42014 227357 42074 237355
rect 42011 227356 42077 227357
rect 42011 227292 42012 227356
rect 42076 227292 42077 227356
rect 42011 227291 42077 227292
rect 591987 223548 592053 223549
rect 591987 223484 591988 223548
rect 592052 223484 592053 223548
rect 591987 223483 592053 223484
rect 591990 222818 592050 223483
rect 649579 223004 649645 223005
rect 649579 222940 649580 223004
rect 649644 222940 649645 223004
rect 649579 222939 649645 222940
rect 651971 223004 652037 223005
rect 651971 222940 651972 223004
rect 652036 222940 652037 223004
rect 651971 222939 652037 222940
rect 649582 222818 649642 222939
rect 651974 222818 652034 222939
rect 572299 220556 572365 220557
rect 572299 220492 572300 220556
rect 572364 220492 572365 220556
rect 572299 220491 572365 220492
rect 572302 217565 572362 220491
rect 511027 217564 511093 217565
rect 511027 217500 511028 217564
rect 511092 217500 511093 217564
rect 511027 217499 511093 217500
rect 520043 217564 520109 217565
rect 520043 217500 520044 217564
rect 520108 217500 520109 217564
rect 520043 217499 520109 217500
rect 532555 217564 532621 217565
rect 532555 217500 532556 217564
rect 532620 217500 532621 217564
rect 532555 217499 532621 217500
rect 572299 217564 572365 217565
rect 572299 217500 572300 217564
rect 572364 217500 572365 217564
rect 572299 217499 572365 217500
rect 511030 215661 511090 217499
rect 520046 215933 520106 217499
rect 520043 215932 520109 215933
rect 520043 215868 520044 215932
rect 520108 215868 520109 215932
rect 520043 215867 520109 215868
rect 511027 215660 511093 215661
rect 511027 215596 511028 215660
rect 511092 215596 511093 215660
rect 511027 215595 511093 215596
rect 532558 215389 532618 217499
rect 532555 215388 532621 215389
rect 532555 215324 532556 215388
rect 532620 215324 532621 215388
rect 532555 215323 532621 215324
rect 41459 209812 41525 209813
rect 41459 209748 41460 209812
rect 41524 209748 41525 209812
rect 41459 209747 41525 209748
rect 665222 209790 665282 265507
rect 674787 264212 674853 264213
rect 674787 264148 674788 264212
rect 674852 264148 674853 264212
rect 674787 264147 674853 264148
rect 674790 249661 674850 264147
rect 676995 261628 677061 261629
rect 676995 261564 676996 261628
rect 677060 261564 677061 261628
rect 676995 261563 677061 261564
rect 676811 261220 676877 261221
rect 676811 261156 676812 261220
rect 676876 261156 676877 261220
rect 676811 261155 676877 261156
rect 675523 258092 675589 258093
rect 675523 258028 675524 258092
rect 675588 258028 675589 258092
rect 675523 258027 675589 258028
rect 675526 249661 675586 258027
rect 674787 249660 674853 249661
rect 674787 249596 674788 249660
rect 674852 249596 674853 249660
rect 674787 249595 674853 249596
rect 675523 249660 675589 249661
rect 675523 249596 675524 249660
rect 675588 249596 675589 249660
rect 675523 249595 675589 249596
rect 676814 246669 676874 261155
rect 676998 250341 677058 261563
rect 676995 250340 677061 250341
rect 676995 250276 676996 250340
rect 677060 250276 677061 250340
rect 676995 250275 677061 250276
rect 676811 246668 676877 246669
rect 676811 246604 676812 246668
rect 676876 246604 676877 246668
rect 676811 246603 676877 246604
rect 674603 246260 674669 246261
rect 674603 246196 674604 246260
rect 674668 246196 674669 246260
rect 674603 246195 674669 246196
rect 673315 246124 673381 246125
rect 673315 246060 673316 246124
rect 673380 246060 673381 246124
rect 673315 246059 673381 246060
rect 670739 236740 670805 236741
rect 670739 236676 670740 236740
rect 670804 236676 670805 236740
rect 670739 236675 670805 236676
rect 667059 231164 667125 231165
rect 667059 231100 667060 231164
rect 667124 231100 667125 231164
rect 667059 231099 667125 231100
rect 40723 207364 40789 207365
rect 40723 207300 40724 207364
rect 40788 207300 40789 207364
rect 40723 207299 40789 207300
rect 40539 206140 40605 206141
rect 40539 206076 40540 206140
rect 40604 206076 40605 206140
rect 40539 206075 40605 206076
rect 40542 192813 40602 206075
rect 40726 194989 40786 207299
rect 40907 206548 40973 206549
rect 40907 206484 40908 206548
rect 40972 206484 40973 206548
rect 40907 206483 40973 206484
rect 40723 194988 40789 194989
rect 40723 194924 40724 194988
rect 40788 194924 40789 194988
rect 40723 194923 40789 194924
rect 40910 193493 40970 206483
rect 41462 195261 41522 209747
rect 665222 209730 666570 209790
rect 41643 208996 41709 208997
rect 41643 208932 41644 208996
rect 41708 208932 41709 208996
rect 41643 208931 41709 208932
rect 41646 195533 41706 208931
rect 666510 204237 666570 209730
rect 666507 204236 666573 204237
rect 666507 204172 666508 204236
rect 666572 204172 666573 204236
rect 666507 204171 666573 204172
rect 41827 197844 41893 197845
rect 41827 197780 41828 197844
rect 41892 197780 41893 197844
rect 41827 197779 41893 197780
rect 41830 195805 41890 197779
rect 41827 195804 41893 195805
rect 41827 195740 41828 195804
rect 41892 195740 41893 195804
rect 41827 195739 41893 195740
rect 41643 195532 41709 195533
rect 41643 195468 41644 195532
rect 41708 195468 41709 195532
rect 41643 195467 41709 195468
rect 41459 195260 41525 195261
rect 41459 195196 41460 195260
rect 41524 195196 41525 195260
rect 41459 195195 41525 195196
rect 42195 194988 42261 194989
rect 42195 194924 42196 194988
rect 42260 194924 42261 194988
rect 42195 194923 42261 194924
rect 40907 193492 40973 193493
rect 40907 193428 40908 193492
rect 40972 193428 40973 193492
rect 40907 193427 40973 193428
rect 40539 192812 40605 192813
rect 40539 192748 40540 192812
rect 40604 192748 40605 192812
rect 40539 192747 40605 192748
rect 42198 186013 42258 194923
rect 42379 193220 42445 193221
rect 42379 193156 42380 193220
rect 42444 193156 42445 193220
rect 42379 193155 42445 193156
rect 42382 186285 42442 193155
rect 42379 186284 42445 186285
rect 42379 186220 42380 186284
rect 42444 186220 42445 186284
rect 42379 186219 42445 186220
rect 42195 186012 42261 186013
rect 42195 185948 42196 186012
rect 42260 185948 42261 186012
rect 42195 185947 42261 185948
rect 667062 122093 667122 231099
rect 670555 224500 670621 224501
rect 670555 224436 670556 224500
rect 670620 224436 670621 224500
rect 670555 224435 670621 224436
rect 670003 223956 670069 223957
rect 670003 223892 670004 223956
rect 670068 223892 670069 223956
rect 670003 223891 670069 223892
rect 667982 179621 668042 222582
rect 670006 222325 670066 223891
rect 670003 222324 670069 222325
rect 670003 222260 670004 222324
rect 670068 222260 670069 222324
rect 670003 222259 670069 222260
rect 669267 220148 669333 220149
rect 669267 220084 669268 220148
rect 669332 220084 669333 220148
rect 669267 220083 669333 220084
rect 669270 212550 669330 220083
rect 669635 218244 669701 218245
rect 669635 218180 669636 218244
rect 669700 218180 669701 218244
rect 669635 218179 669701 218180
rect 669270 212490 669514 212550
rect 669267 205732 669333 205733
rect 669267 205668 669268 205732
rect 669332 205668 669333 205732
rect 669267 205667 669333 205668
rect 669270 205461 669330 205667
rect 669267 205460 669333 205461
rect 669267 205396 669268 205460
rect 669332 205396 669333 205460
rect 669267 205395 669333 205396
rect 669267 196212 669333 196213
rect 669267 196148 669268 196212
rect 669332 196148 669333 196212
rect 669267 196147 669333 196148
rect 669270 195941 669330 196147
rect 669267 195940 669333 195941
rect 669267 195876 669268 195940
rect 669332 195876 669333 195940
rect 669267 195875 669333 195876
rect 669454 188461 669514 212490
rect 669638 205733 669698 218179
rect 670558 217973 670618 224435
rect 670555 217972 670621 217973
rect 670555 217908 670556 217972
rect 670620 217908 670621 217972
rect 670555 217907 670621 217908
rect 669635 205732 669701 205733
rect 669635 205668 669636 205732
rect 669700 205668 669701 205732
rect 669635 205667 669701 205668
rect 669635 205460 669701 205461
rect 669635 205396 669636 205460
rect 669700 205396 669701 205460
rect 669635 205395 669701 205396
rect 669638 196213 669698 205395
rect 670742 198797 670802 236675
rect 672579 227084 672645 227085
rect 672579 227020 672580 227084
rect 672644 227020 672645 227084
rect 672579 227019 672645 227020
rect 671659 224772 671725 224773
rect 671659 224708 671660 224772
rect 671724 224708 671725 224772
rect 671659 224707 671725 224708
rect 671662 223957 671722 224707
rect 671659 223956 671725 223957
rect 671659 223892 671660 223956
rect 671724 223892 671725 223956
rect 671659 223891 671725 223892
rect 672582 200837 672642 227019
rect 672579 200836 672645 200837
rect 672579 200772 672580 200836
rect 672644 200772 672645 200836
rect 672579 200771 672645 200772
rect 670739 198796 670805 198797
rect 670739 198732 670740 198796
rect 670804 198732 670805 198796
rect 670739 198731 670805 198732
rect 669635 196212 669701 196213
rect 669635 196148 669636 196212
rect 669700 196148 669701 196212
rect 669635 196147 669701 196148
rect 669635 195940 669701 195941
rect 669635 195876 669636 195940
rect 669700 195876 669701 195940
rect 669635 195875 669701 195876
rect 669451 188460 669517 188461
rect 669451 188396 669452 188460
rect 669516 188396 669517 188460
rect 669451 188395 669517 188396
rect 667979 179620 668045 179621
rect 667979 179556 667980 179620
rect 668044 179556 668045 179620
rect 667979 179555 668045 179556
rect 669638 176670 669698 195875
rect 673131 181524 673197 181525
rect 673131 181460 673132 181524
rect 673196 181460 673197 181524
rect 673131 181459 673197 181460
rect 669454 176610 669698 176670
rect 669454 157350 669514 176610
rect 673134 161533 673194 181459
rect 673318 178125 673378 246059
rect 674051 226812 674117 226813
rect 674051 226748 674052 226812
rect 674116 226748 674117 226812
rect 674051 226747 674117 226748
rect 673315 178124 673381 178125
rect 673315 178060 673316 178124
rect 673380 178060 673381 178124
rect 673315 178059 673381 178060
rect 673131 161532 673197 161533
rect 673131 161468 673132 161532
rect 673196 161468 673197 161532
rect 673131 161467 673197 161468
rect 669270 157290 669514 157350
rect 669270 140453 669330 157290
rect 669267 140452 669333 140453
rect 669267 140388 669268 140452
rect 669332 140388 669333 140452
rect 669267 140387 669333 140388
rect 667059 122092 667125 122093
rect 667059 122028 667060 122092
rect 667124 122028 667125 122092
rect 667059 122027 667125 122028
rect 674054 115837 674114 226747
rect 674606 206957 674666 246195
rect 675339 245852 675405 245853
rect 675339 245788 675340 245852
rect 675404 245788 675405 245852
rect 675339 245787 675405 245788
rect 675342 235245 675402 245787
rect 676811 242044 676877 242045
rect 676811 241980 676812 242044
rect 676876 241980 676877 242044
rect 676811 241979 676877 241980
rect 675339 235244 675405 235245
rect 675339 235180 675340 235244
rect 675404 235180 675405 235244
rect 675339 235179 675405 235180
rect 675155 230484 675221 230485
rect 675155 230420 675156 230484
rect 675220 230420 675221 230484
rect 675155 230419 675221 230420
rect 674603 206956 674669 206957
rect 674603 206892 674604 206956
rect 674668 206892 674669 206956
rect 674603 206891 674669 206892
rect 675158 190093 675218 230419
rect 676814 220010 676874 241979
rect 676078 219950 676874 220010
rect 676078 219877 676138 219950
rect 676029 219876 676138 219877
rect 676029 219812 676030 219876
rect 676094 219814 676138 219876
rect 676094 219812 676095 219814
rect 676029 219811 676095 219812
rect 675707 218652 675773 218653
rect 675707 218588 675708 218652
rect 675772 218588 675773 218652
rect 675707 218587 675773 218588
rect 675710 215310 675770 218587
rect 675891 217972 675957 217973
rect 675891 217908 675892 217972
rect 675956 217970 675957 217972
rect 675956 217910 676322 217970
rect 675956 217908 675957 217910
rect 675891 217907 675957 217908
rect 676262 217290 676322 217910
rect 676262 217230 676506 217290
rect 675894 215870 676322 215930
rect 675894 215525 675954 215870
rect 675891 215524 675957 215525
rect 675891 215460 675892 215524
rect 675956 215460 675957 215524
rect 675891 215459 675957 215460
rect 675710 215250 676138 215310
rect 675891 212532 675957 212533
rect 675891 212468 675892 212532
rect 675956 212468 675957 212532
rect 675891 212467 675957 212468
rect 675894 192813 675954 212467
rect 676078 193221 676138 215250
rect 676262 194581 676322 215870
rect 676446 202741 676506 217230
rect 676627 211444 676693 211445
rect 676627 211380 676628 211444
rect 676692 211380 676693 211444
rect 676627 211379 676693 211380
rect 676443 202740 676509 202741
rect 676443 202676 676444 202740
rect 676508 202676 676509 202740
rect 676443 202675 676509 202676
rect 676630 200021 676690 211379
rect 676627 200020 676693 200021
rect 676627 199956 676628 200020
rect 676692 199956 676693 200020
rect 676627 199955 676693 199956
rect 676811 197980 676877 197981
rect 676811 197916 676812 197980
rect 676876 197916 676877 197980
rect 676811 197915 676877 197916
rect 676259 194580 676325 194581
rect 676259 194516 676260 194580
rect 676324 194516 676325 194580
rect 676259 194515 676325 194516
rect 676075 193220 676141 193221
rect 676075 193156 676076 193220
rect 676140 193156 676141 193220
rect 676075 193155 676141 193156
rect 675891 192812 675957 192813
rect 675891 192748 675892 192812
rect 675956 192748 675957 192812
rect 675891 192747 675957 192748
rect 675155 190092 675221 190093
rect 675155 190028 675156 190092
rect 675220 190028 675221 190092
rect 675155 190027 675221 190028
rect 676814 176673 676874 197915
rect 676811 176672 676877 176673
rect 676811 176608 676812 176672
rect 676876 176608 676877 176672
rect 676811 176607 676877 176608
rect 675891 172820 675957 172821
rect 675891 172756 675892 172820
rect 675956 172756 675957 172820
rect 675891 172755 675957 172756
rect 675894 172410 675954 172755
rect 675894 172350 676506 172410
rect 675891 169420 675957 169421
rect 675891 169356 675892 169420
rect 675956 169356 675957 169420
rect 675891 169355 675957 169356
rect 675894 169010 675954 169355
rect 675894 168950 676322 169010
rect 675339 167516 675405 167517
rect 675339 167452 675340 167516
rect 675404 167452 675405 167516
rect 675339 167451 675405 167452
rect 675342 147661 675402 167451
rect 676075 162756 676141 162757
rect 676075 162692 676076 162756
rect 676140 162692 676141 162756
rect 676075 162691 676141 162692
rect 676078 148477 676138 162691
rect 676262 155821 676322 168950
rect 676446 157045 676506 172350
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676443 157044 676509 157045
rect 676443 156980 676444 157044
rect 676508 156980 676509 157044
rect 676443 156979 676509 156980
rect 676259 155820 676325 155821
rect 676259 155756 676260 155820
rect 676324 155756 676325 155820
rect 676259 155755 676325 155756
rect 676630 151469 676690 166363
rect 676627 151468 676693 151469
rect 676627 151404 676628 151468
rect 676692 151404 676693 151468
rect 676627 151403 676693 151404
rect 676075 148476 676141 148477
rect 676075 148412 676076 148476
rect 676140 148412 676141 148476
rect 676075 148411 676141 148412
rect 675339 147660 675405 147661
rect 675339 147596 675340 147660
rect 675404 147596 675405 147660
rect 675339 147595 675405 147596
rect 676627 127396 676693 127397
rect 676627 127332 676628 127396
rect 676692 127332 676693 127396
rect 676627 127331 676693 127332
rect 676075 126988 676141 126989
rect 676075 126924 676076 126988
rect 676140 126924 676141 126988
rect 676075 126923 676141 126924
rect 675339 122092 675405 122093
rect 675339 122028 675340 122092
rect 675404 122028 675405 122092
rect 675339 122027 675405 122028
rect 674051 115836 674117 115837
rect 674051 115772 674052 115836
rect 674116 115772 674117 115836
rect 674051 115771 674117 115772
rect 675342 102645 675402 122027
rect 675707 117332 675773 117333
rect 675707 117268 675708 117332
rect 675772 117268 675773 117332
rect 675707 117267 675773 117268
rect 675710 111349 675770 117267
rect 675707 111348 675773 111349
rect 675707 111284 675708 111348
rect 675772 111284 675773 111348
rect 675707 111283 675773 111284
rect 676078 108221 676138 126923
rect 676259 125764 676325 125765
rect 676259 125700 676260 125764
rect 676324 125700 676325 125764
rect 676259 125699 676325 125700
rect 676262 111757 676322 125699
rect 676443 124132 676509 124133
rect 676443 124068 676444 124132
rect 676508 124068 676509 124132
rect 676443 124067 676509 124068
rect 676259 111756 676325 111757
rect 676259 111692 676260 111756
rect 676324 111692 676325 111756
rect 676259 111691 676325 111692
rect 676446 110397 676506 124067
rect 676630 112437 676690 127331
rect 676627 112436 676693 112437
rect 676627 112372 676628 112436
rect 676692 112372 676693 112436
rect 676627 112371 676693 112372
rect 676443 110396 676509 110397
rect 676443 110332 676444 110396
rect 676508 110332 676509 110396
rect 676443 110331 676509 110332
rect 676075 108220 676141 108221
rect 676075 108156 676076 108220
rect 676140 108156 676141 108220
rect 676075 108155 676141 108156
rect 675339 102644 675405 102645
rect 675339 102580 675340 102644
rect 675404 102580 675405 102644
rect 675339 102579 675405 102580
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 633939 95436 634005 95437
rect 633939 95372 633940 95436
rect 634004 95372 634005 95436
rect 633939 95371 634005 95372
rect 633942 78573 634002 95371
rect 637254 84210 637314 96867
rect 647187 96524 647253 96525
rect 647187 96460 647188 96524
rect 647252 96460 647253 96524
rect 647187 96459 647253 96460
rect 647190 94298 647250 96459
rect 650318 93125 650378 93382
rect 650315 93124 650381 93125
rect 650315 93060 650316 93124
rect 650380 93060 650381 93124
rect 650315 93059 650381 93060
rect 637070 84150 637314 84210
rect 633939 78572 634005 78573
rect 633939 78508 633940 78572
rect 634004 78508 634005 78572
rect 633939 78507 634005 78508
rect 637070 78165 637130 84150
rect 637067 78164 637133 78165
rect 637067 78100 637068 78164
rect 637132 78100 637133 78164
rect 637067 78099 637133 78100
rect 460795 55044 460861 55045
rect 460795 54980 460796 55044
rect 460860 54980 460861 55044
rect 460795 54979 460861 54980
rect 460798 53957 460858 54979
rect 462635 54772 462701 54773
rect 462635 54708 462636 54772
rect 462700 54708 462701 54772
rect 462635 54707 462701 54708
rect 460795 53956 460861 53957
rect 460795 53892 460796 53956
rect 460860 53892 460861 53956
rect 460795 53891 460861 53892
rect 462638 53685 462698 54707
rect 462635 53684 462701 53685
rect 462635 53620 462636 53684
rect 462700 53620 462701 53684
rect 462635 53619 462701 53620
rect 518755 48924 518821 48925
rect 518755 48860 518756 48924
rect 518820 48860 518821 48924
rect 518755 48859 518821 48860
rect 515443 47836 515509 47837
rect 515443 47772 515444 47836
rect 515508 47772 515509 47836
rect 515443 47771 515509 47772
rect 460979 44436 461045 44437
rect 460979 44372 460980 44436
rect 461044 44372 461045 44436
rect 460979 44371 461045 44372
rect 462267 44436 462333 44437
rect 462267 44372 462268 44436
rect 462332 44372 462333 44436
rect 462267 44371 462333 44372
rect 463739 44436 463805 44437
rect 463739 44372 463740 44436
rect 463804 44372 463805 44436
rect 463739 44371 463805 44372
rect 141739 44028 141805 44029
rect 141739 43964 141740 44028
rect 141804 43964 141805 44028
rect 141739 43963 141805 43964
rect 141742 40357 141802 43963
rect 419211 42124 419277 42125
rect 419211 42060 419212 42124
rect 419276 42060 419277 42124
rect 419211 42059 419277 42060
rect 419214 41938 419274 42059
rect 416635 41852 416701 41853
rect 416635 41788 416636 41852
rect 416700 41788 416701 41852
rect 416635 41787 416701 41788
rect 416638 40578 416698 41787
rect 441843 41852 441909 41853
rect 441843 41850 441844 41852
rect 441626 41790 441844 41850
rect 441843 41788 441844 41790
rect 441908 41788 441909 41852
rect 441843 41787 441909 41788
rect 451963 41852 452029 41853
rect 451963 41788 451964 41852
rect 452028 41788 452029 41852
rect 451963 41787 452029 41788
rect 451966 41258 452026 41787
rect 458958 41170 459018 41702
rect 458958 41110 460342 41170
rect 460982 40578 461042 44371
rect 462270 41258 462330 44371
rect 463742 41938 463802 44371
rect 515446 42125 515506 47771
rect 518758 42805 518818 48859
rect 529611 48108 529677 48109
rect 529611 48044 529612 48108
rect 529676 48044 529677 48108
rect 529611 48043 529677 48044
rect 526483 47836 526549 47837
rect 526483 47772 526484 47836
rect 526548 47772 526549 47836
rect 526483 47771 526549 47772
rect 520963 47564 521029 47565
rect 520963 47500 520964 47564
rect 521028 47500 521029 47564
rect 520963 47499 521029 47500
rect 518755 42804 518821 42805
rect 518755 42740 518756 42804
rect 518820 42740 518821 42804
rect 518755 42739 518821 42740
rect 520966 42125 521026 47499
rect 522067 47292 522133 47293
rect 522067 47228 522068 47292
rect 522132 47228 522133 47292
rect 522067 47227 522133 47228
rect 522070 42125 522130 47227
rect 526486 42125 526546 47771
rect 529614 42125 529674 48043
rect 515443 42124 515509 42125
rect 515443 42060 515444 42124
rect 515508 42060 515509 42124
rect 515443 42059 515509 42060
rect 520963 42124 521029 42125
rect 520963 42060 520964 42124
rect 521028 42060 521029 42124
rect 520963 42059 521029 42060
rect 522067 42124 522133 42125
rect 522067 42060 522068 42124
rect 522132 42060 522133 42124
rect 522067 42059 522133 42060
rect 526483 42124 526549 42125
rect 526483 42060 526484 42124
rect 526548 42060 526549 42124
rect 526483 42059 526549 42060
rect 529611 42124 529677 42125
rect 529611 42060 529612 42124
rect 529676 42060 529677 42124
rect 529611 42059 529677 42060
rect 141739 40356 141805 40357
rect 141739 40292 141740 40356
rect 141804 40292 141805 40356
rect 141739 40291 141805 40292
<< via4 >>
rect 591902 222582 592138 222818
rect 649494 222582 649730 222818
rect 651886 222582 652122 222818
rect 667894 222582 668130 222818
rect 647102 94062 647338 94298
rect 650230 93382 650466 93618
rect 365030 41852 365266 41938
rect 365030 41788 365116 41852
rect 365116 41788 365180 41852
rect 365180 41788 365266 41852
rect 365030 41702 365266 41788
rect 419126 41702 419362 41938
rect 419862 41852 420098 41938
rect 419862 41788 419948 41852
rect 419948 41788 420012 41852
rect 420012 41788 420098 41852
rect 419862 41702 420098 41788
rect 425014 41852 425250 41938
rect 425014 41788 425100 41852
rect 425100 41788 425164 41852
rect 425164 41788 425250 41852
rect 425014 41702 425250 41788
rect 441390 41702 441626 41938
rect 458870 41702 459106 41938
rect 451878 41022 452114 41258
rect 460342 41022 460578 41258
rect 463654 41702 463890 41938
rect 462182 41022 462418 41258
rect 416550 40342 416786 40578
rect 460894 40342 461130 40578
<< metal5 >>
rect 78610 1018624 90778 1030789
rect 130010 1018624 142178 1030789
rect 181410 1018624 193578 1030789
rect 231810 1018624 243978 1030789
rect 284410 1018624 296578 1030789
rect 334810 1018624 346978 1030789
rect 386210 1018624 398378 1030789
rect 475210 1018624 487378 1030789
rect 526610 1018624 538778 1030789
rect 577010 1018624 589178 1030789
rect 628410 1018624 640578 1030789
rect 6811 956610 18976 968778
rect 698624 953022 710789 965190
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 591860 222818 649772 222860
rect 591860 222582 591902 222818
rect 592138 222582 649494 222818
rect 649730 222582 649772 222818
rect 591860 222540 649772 222582
rect 651844 222818 668172 222860
rect 651844 222582 651886 222818
rect 652122 222582 667894 222818
rect 668130 222582 668172 222818
rect 651844 222540 668172 222582
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 647060 94298 647748 94340
rect 647060 94062 647102 94298
rect 647338 94062 647748 94298
rect 647060 94020 647748 94062
rect 647428 93660 647748 94020
rect 647428 93618 650508 93660
rect 647428 93382 650230 93618
rect 650466 93382 650508 93618
rect 647428 93340 650508 93382
rect 6167 70054 19620 80934
rect 364988 41938 419404 41980
rect 364988 41702 365030 41938
rect 365266 41702 419126 41938
rect 419362 41702 419404 41938
rect 364988 41660 419404 41702
rect 419820 41938 424556 41980
rect 419820 41702 419862 41938
rect 420098 41702 424556 41938
rect 419820 41660 424556 41702
rect 424972 41938 441668 41980
rect 424972 41702 425014 41938
rect 425250 41702 441390 41938
rect 441626 41702 441668 41938
rect 424972 41660 441668 41702
rect 442084 41660 450684 41980
rect 424236 41300 424556 41660
rect 442084 41300 442404 41660
rect 424236 40980 442404 41300
rect 450364 41300 450684 41660
rect 451100 41938 459148 41980
rect 451100 41702 458870 41938
rect 459106 41702 459148 41938
rect 451100 41660 459148 41702
rect 459564 41938 463932 41980
rect 459564 41702 463654 41938
rect 463890 41702 463932 41938
rect 459564 41660 463932 41702
rect 451100 41300 451420 41660
rect 459564 41300 459884 41660
rect 450364 40980 451420 41300
rect 451836 41258 459884 41300
rect 451836 41022 451878 41258
rect 452114 41022 459884 41258
rect 451836 40980 459884 41022
rect 460300 41258 462460 41300
rect 460300 41022 460342 41258
rect 460578 41022 462182 41258
rect 462418 41022 462460 41258
rect 460300 40980 462460 41022
rect 416508 40578 461172 40620
rect 416508 40342 416550 40578
rect 416786 40342 460894 40578
rect 461130 40342 461172 40578
rect 416508 40300 461172 40342
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use caravan_logo  caravan_logo
timestamp 0
transform 1 0 255300 0 1 6032
box 0 0 1 1
use caravan_motto  caravan_motto
timestamp 0
transform 1 0 -54560 0 1 -52
box 0 0 1 1
use copyright_block_a  copyright_block_a
timestamp 0
transform 1 0 149582 0 1 16298
box 0 0 1 1
use open_source  open_source
timestamp 0
transform 1 0 206074 0 1 2336
box 0 0 1 1
use xres_buf  rstb_level
timestamp 1666198072
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use user_id_textblock  user_id_textblock
timestamp 0
transform 1 0 96272 0 1 6890
box 0 0 1 1
use caravel_clocking  clock_ctrl
timestamp 1666198072
transform 1 0 626764 0 1 55284
box 136 496 20000 20000
use buff_flash_clkrst  flash_clkrst_buffers
timestamp 1666198072
transform 1 0 458400 0 1 47600
box 330 0 7699 5000
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1666198072
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1666198072
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1666198072
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use digital_pll  pll
timestamp 1666198072
transform 1 0 628146 0 1 80944
box 0 0 20000 15000
use simple_por  por
timestamp 1666198072
transform 1 0 650146 0 -1 55282
box -14 11 11344 8684
use user_id_programming  user_id_value
timestamp 1666198072
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1666198072
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1666198072
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1666198072
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1666198072
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1666198072
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1666198072
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1666198072
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use spare_logic_block  spare_logic\[2\]
timestamp 1666198072
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1666198072
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1666198072
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1666198072
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use mgmt_protect  mgmt_buffers
timestamp 1666198072
transform 1 0 128180 0 1 232036
box 1066 -400 424400 32400
use spare_logic_block  spare_logic\[0\]
timestamp 1666198072
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1666198072
transform 1 0 108632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1666198072
transform 1 0 578632 0 1 232528
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1666198072
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1666198072
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1666198072
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1666198072
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1666198072
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1666198072
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1666198072
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1666198072
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1666198072
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1666198072
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1666198072
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1666198072
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1666198072
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1666198072
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1666198072
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1666198072
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1666198072
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1666198072
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1666198072
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1666198072
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1666198072
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1666198072
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1666198072
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1666198072
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1666198072
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1666198072
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1666198072
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1666198072
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1666198072
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1666198072
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1666198072
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1666198072
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1666198072
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1666198072
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1666198072
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1666198072
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1666198072
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1666198072
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1666198072
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1666198072
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1666198072
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1666198072
transform -1 0 710203 0 1 884800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1666198072
transform -1 0 709467 0 1 897800
box -38 0 6018 2224
use caravan_power_routing  caravan_power_routing
timestamp 1666198072
transform 1 0 0 0 1 0
box 6022 30806 711814 1006847
use user_analog_project_wrapper  mprj
timestamp 1666198072
transform 1 0 65308 0 1 278718
box -800 -800 584800 704800
use chip_io_alt  padframe
timestamp 1666198072
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use gpio_signal_buffering_alt  sigbuf
timestamp 1666198072
transform 1 0 0 0 1 0
box 40023 41960 677583 728321
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698624 953022 710789 965190 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 628410 1018624 640578 1030789 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 526610 1018624 538778 1030789 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 475210 1018624 487378 1030789 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 386210 1018624 398378 1030789 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 284410 1018624 296578 1030789 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 231810 1018624 243978 1030789 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 181410 1018624 193578 1030789 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 130010 1018624 142178 1030789 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 78610 1018624 90778 1030789 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6811 956610 18976 968778 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144150 18309 6 resetb
port 44 nsew signal input
rlabel metal5 s 6167 70054 19620 80934 6 vccd
port 45 nsew signal bidirectional
rlabel metal5 s 697980 909666 711433 920546 6 vccd1
port 46 nsew signal bidirectional
rlabel metal5 s 6167 914054 19620 924934 6 vccd2
port 47 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18976 6 vdda
port 48 nsew signal bidirectional
rlabel metal5 s 698624 819822 710789 831990 6 vdda1
port 49 nsew signal bidirectional
rlabel metal5 s 698624 505222 710789 517390 6 vdda1_2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 484410 18976 496578 6 vdda2
port 51 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio
port 52 nsew signal bidirectional
rlabel metal5 s 6811 871210 18976 883378 6 vddio_2
port 53 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18976 6 vssa
port 54 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1
port 55 nsew signal bidirectional
rlabel metal5 s 698624 417022 710789 429190 6 vssa1_2
port 56 nsew signal bidirectional
rlabel metal5 s 6811 829010 18976 841178 6 vssa2
port 57 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19620 6 vssd
port 58 nsew signal bidirectional
rlabel metal5 s 697980 461866 711433 472746 6 vssd1
port 59 nsew signal bidirectional
rlabel metal5 s 6167 442854 19620 453734 6 vssd2
port 60 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio
port 61 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030789 6 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
