magic
tech sky130A
magscale 1 2
timestamp 1661979173
<< checkpaint >>
rect 3127 15264 5715 15266
rect 839 15258 5715 15264
rect 425 15220 5715 15258
rect 425 12732 10890 15220
rect -378 4132 11142 12732
rect -102 372 11142 4132
rect 1738 -220 11142 372
<< isosubstrate >>
rect 1110 1538 2650 4514
<< viali >>
rect 1317 11305 1351 11339
rect 1777 11305 1811 11339
rect 5825 11305 5859 11339
rect 8493 11305 8527 11339
rect 9413 11305 9447 11339
rect 2053 11237 2087 11271
rect 2145 11237 2179 11271
rect 2881 11237 2915 11271
rect 2973 11237 3007 11271
rect 3249 11237 3283 11271
rect 6377 11237 6411 11271
rect 7757 11237 7791 11271
rect 4445 11169 4479 11203
rect 1501 11101 1535 11135
rect 1593 11101 1627 11135
rect 1869 11101 1903 11135
rect 2329 11101 2363 11135
rect 2421 11101 2455 11135
rect 2697 11101 2731 11135
rect 3157 11101 3191 11135
rect 3433 11101 3467 11135
rect 3801 11101 3835 11135
rect 4077 11101 4111 11135
rect 4721 11101 4755 11135
rect 5733 11101 5767 11135
rect 6009 11101 6043 11135
rect 6561 11101 6595 11135
rect 7481 11101 7515 11135
rect 7573 11101 7607 11135
rect 7941 11101 7975 11135
rect 8309 11101 8343 11135
rect 8861 11101 8895 11135
rect 9229 11101 9263 11135
rect 4261 11033 4295 11067
rect 6653 11033 6687 11067
rect 6837 11033 6871 11067
rect 7021 11033 7055 11067
rect 2605 10965 2639 10999
rect 3985 10965 4019 10999
rect 5365 10965 5399 10999
rect 5549 10965 5583 10999
rect 7297 10965 7331 10999
rect 8125 10965 8159 10999
rect 9045 10965 9079 10999
rect 2513 10761 2547 10795
rect 1225 10625 1259 10659
rect 2237 10625 2271 10659
rect 2329 10625 2363 10659
rect 2789 10649 2823 10683
rect 4905 10625 4939 10659
rect 4997 10625 5031 10659
rect 5549 10625 5583 10659
rect 5733 10625 5767 10659
rect 6285 10625 6319 10659
rect 8677 10625 8711 10659
rect 9229 10625 9263 10659
rect 2870 10557 2904 10591
rect 4629 10557 4663 10591
rect 5457 10557 5491 10591
rect 6837 10557 6871 10591
rect 7205 10557 7239 10591
rect 1869 10489 1903 10523
rect 5917 10489 5951 10523
rect 6745 10489 6779 10523
rect 2053 10421 2087 10455
rect 2605 10421 2639 10455
rect 3144 10421 3178 10455
rect 4721 10421 4755 10455
rect 5273 10421 5307 10455
rect 6377 10421 6411 10455
rect 9137 10421 9171 10455
rect 9413 10421 9447 10455
rect 6837 10217 6871 10251
rect 9505 10217 9539 10251
rect 3433 10149 3467 10183
rect 7297 10149 7331 10183
rect 8493 10149 8527 10183
rect 1685 10081 1719 10115
rect 4537 10081 4571 10115
rect 1409 10013 1443 10047
rect 3617 10013 3651 10047
rect 4905 10013 4939 10047
rect 6377 10013 6411 10047
rect 6929 10013 6963 10047
rect 7389 10013 7423 10047
rect 8033 10013 8067 10047
rect 8309 10013 8343 10047
rect 8861 10013 8895 10047
rect 1961 9945 1995 9979
rect 7113 9945 7147 9979
rect 7573 9945 7607 9979
rect 1593 9877 1627 9911
rect 4261 9877 4295 9911
rect 7757 9877 7791 9911
rect 8125 9877 8159 9911
rect 9505 9673 9539 9707
rect 8033 9605 8067 9639
rect 1225 9537 1259 9571
rect 4905 9537 4939 9571
rect 5549 9537 5583 9571
rect 6193 9537 6227 9571
rect 7113 9537 7147 9571
rect 7757 9537 7791 9571
rect 3065 9469 3099 9503
rect 3433 9469 3467 9503
rect 6469 9469 6503 9503
rect 7573 9469 7607 9503
rect 2973 9401 3007 9435
rect 6009 9401 6043 9435
rect 1488 9333 1522 9367
rect 5365 9333 5399 9367
rect 5825 9333 5859 9367
rect 7389 9333 7423 9367
rect 3065 9129 3099 9163
rect 4261 9129 4295 9163
rect 4629 9129 4663 9163
rect 8217 9129 8251 9163
rect 1501 9061 1535 9095
rect 2789 9061 2823 9095
rect 3341 9061 3375 9095
rect 5917 8993 5951 9027
rect 9137 8993 9171 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 1961 8925 1995 8959
rect 2237 8925 2271 8959
rect 2513 8925 2547 8959
rect 2605 8925 2639 8959
rect 2881 8925 2915 8959
rect 3249 8925 3283 8959
rect 3617 8925 3651 8959
rect 4353 8925 4387 8959
rect 4997 8925 5031 8959
rect 5273 8925 5307 8959
rect 6285 8925 6319 8959
rect 7757 8925 7791 8959
rect 8309 8925 8343 8959
rect 8861 8925 8895 8959
rect 1225 8789 1259 8823
rect 1777 8789 1811 8823
rect 2053 8789 2087 8823
rect 2329 8789 2363 8823
rect 4813 8789 4847 8823
rect 8493 8789 8527 8823
rect 2145 8585 2179 8619
rect 2421 8585 2455 8619
rect 2881 8585 2915 8619
rect 9137 8585 9171 8619
rect 2513 8517 2547 8551
rect 1409 8449 1443 8483
rect 1685 8449 1719 8483
rect 1961 8449 1995 8483
rect 2237 8449 2271 8483
rect 2697 8449 2731 8483
rect 2973 8449 3007 8483
rect 3525 8449 3559 8483
rect 4445 8449 4479 8483
rect 5181 8449 5215 8483
rect 6193 8449 6227 8483
rect 6377 8449 6411 8483
rect 6837 8449 6871 8483
rect 7205 8449 7239 8483
rect 8677 8449 8711 8483
rect 9229 8449 9263 8483
rect 3433 8381 3467 8415
rect 5457 8381 5491 8415
rect 4169 8313 4203 8347
rect 9413 8313 9447 8347
rect 1593 8245 1627 8279
rect 1869 8245 1903 8279
rect 3157 8245 3191 8279
rect 5089 8245 5123 8279
rect 6561 8245 6595 8279
rect 1501 8041 1535 8075
rect 1961 8041 1995 8075
rect 2881 8041 2915 8075
rect 3249 8041 3283 8075
rect 5549 8041 5583 8075
rect 7849 8041 7883 8075
rect 8585 8041 8619 8075
rect 8769 8041 8803 8075
rect 1685 7973 1719 8007
rect 3433 7973 3467 8007
rect 6929 7973 6963 8007
rect 9321 7905 9355 7939
rect 1317 7837 1351 7871
rect 1593 7837 1627 7871
rect 1869 7837 1903 7871
rect 2237 7837 2271 7871
rect 2513 7837 2547 7871
rect 2973 7837 3007 7871
rect 3801 7837 3835 7871
rect 5641 7837 5675 7871
rect 7665 7837 7699 7871
rect 7941 7837 7975 7871
rect 2697 7769 2731 7803
rect 4077 7769 4111 7803
rect 7481 7769 7515 7803
rect 9137 7769 9171 7803
rect 2329 7701 2363 7735
rect 9229 7701 9263 7735
rect 1225 7497 1259 7531
rect 1685 7497 1719 7531
rect 6009 7497 6043 7531
rect 8585 7497 8619 7531
rect 2145 7429 2179 7463
rect 6561 7429 6595 7463
rect 1409 7361 1443 7395
rect 1501 7361 1535 7395
rect 1777 7361 1811 7395
rect 2053 7361 2087 7395
rect 2513 7361 2547 7395
rect 4445 7361 4479 7395
rect 4997 7361 5031 7395
rect 5365 7361 5399 7395
rect 6285 7361 6319 7395
rect 8125 7361 8159 7395
rect 9045 7361 9079 7395
rect 2593 7293 2627 7327
rect 2973 7293 3007 7327
rect 8033 7293 8067 7327
rect 9137 7293 9171 7327
rect 9229 7293 9263 7327
rect 4905 7225 4939 7259
rect 1961 7157 1995 7191
rect 2329 7157 2363 7191
rect 5181 7157 5215 7191
rect 8401 7157 8435 7191
rect 8677 7157 8711 7191
rect 1942 6953 1976 6987
rect 8769 6953 8803 6987
rect 8585 6817 8619 6851
rect 9321 6817 9355 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 3617 6749 3651 6783
rect 4537 6749 4571 6783
rect 4905 6749 4939 6783
rect 6377 6749 6411 6783
rect 6929 6749 6963 6783
rect 7573 6749 7607 6783
rect 7849 6749 7883 6783
rect 7941 6749 7975 6783
rect 9229 6681 9263 6715
rect 1501 6613 1535 6647
rect 3433 6613 3467 6647
rect 4261 6613 4295 6647
rect 6837 6613 6871 6647
rect 7665 6613 7699 6647
rect 9137 6613 9171 6647
rect 1501 6409 1535 6443
rect 1961 6409 1995 6443
rect 1409 6273 1443 6307
rect 1685 6273 1719 6307
rect 1777 6273 1811 6307
rect 2053 6273 2087 6307
rect 2329 6273 2363 6307
rect 4537 6273 4571 6307
rect 6193 6273 6227 6307
rect 6745 6273 6779 6307
rect 8585 6273 8619 6307
rect 9321 6273 9355 6307
rect 2697 6205 2731 6239
rect 3065 6205 3099 6239
rect 4997 6205 5031 6239
rect 5181 6205 5215 6239
rect 5457 6205 5491 6239
rect 6653 6205 6687 6239
rect 7113 6205 7147 6239
rect 9137 6205 9171 6239
rect 1225 6137 1259 6171
rect 2513 6137 2547 6171
rect 2237 6069 2271 6103
rect 6285 6069 6319 6103
rect 8769 6069 8803 6103
rect 9045 6069 9079 6103
rect 9505 6069 9539 6103
rect 5549 5865 5583 5899
rect 5917 5797 5951 5831
rect 8769 5797 8803 5831
rect 1685 5729 1719 5763
rect 3617 5729 3651 5763
rect 5365 5729 5399 5763
rect 6653 5729 6687 5763
rect 6929 5729 6963 5763
rect 9321 5729 9355 5763
rect 1593 5661 1627 5695
rect 5457 5661 5491 5695
rect 6561 5661 6595 5695
rect 9137 5661 9171 5695
rect 1961 5593 1995 5627
rect 3893 5593 3927 5627
rect 6193 5593 6227 5627
rect 6377 5593 6411 5627
rect 1409 5525 1443 5559
rect 3433 5525 3467 5559
rect 8401 5525 8435 5559
rect 9229 5525 9263 5559
rect 8953 5321 8987 5355
rect 3433 5185 3467 5219
rect 5825 5185 5859 5219
rect 6377 5185 6411 5219
rect 8309 5185 8343 5219
rect 9229 5185 9263 5219
rect 3985 5117 4019 5151
rect 4353 5117 4387 5151
rect 6653 5117 6687 5151
rect 3525 4981 3559 5015
rect 3893 4981 3927 5015
rect 6285 4981 6319 5015
rect 8125 4981 8159 5015
rect 9413 4981 9447 5015
rect 5089 4777 5123 4811
rect 3341 4641 3375 4675
rect 3617 4641 3651 4675
rect 5825 4641 5859 4675
rect 7665 4641 7699 4675
rect 5181 4573 5215 4607
rect 5365 4573 5399 4607
rect 6101 4505 6135 4539
rect 7849 4505 7883 4539
rect 9505 4505 9539 4539
rect 5549 4437 5583 4471
rect 7573 4437 7607 4471
rect 4813 4233 4847 4267
rect 3525 4097 3559 4131
rect 4261 4097 4295 4131
rect 4997 4097 5031 4131
rect 5089 4097 5123 4131
rect 5733 4097 5767 4131
rect 7665 4097 7699 4131
rect 8309 4097 8343 4131
rect 9045 4097 9079 4131
rect 5825 4029 5859 4063
rect 6193 4029 6227 4063
rect 4721 3961 4755 3995
rect 8953 3961 8987 3995
rect 4169 3893 4203 3927
rect 4537 3893 4571 3927
rect 8125 3893 8159 3927
rect 9137 3893 9171 3927
rect 9505 3893 9539 3927
rect 3801 3689 3835 3723
rect 5365 3689 5399 3723
rect 8953 3689 8987 3723
rect 4077 3621 4111 3655
rect 6377 3621 6411 3655
rect 6837 3553 6871 3587
rect 3341 3485 3375 3519
rect 3617 3485 3651 3519
rect 3893 3485 3927 3519
rect 4169 3485 4203 3519
rect 4629 3485 4663 3519
rect 5549 3485 5583 3519
rect 5733 3485 5767 3519
rect 6469 3485 6503 3519
rect 8309 3485 8343 3519
rect 8861 3485 8895 3519
rect 4721 3417 4755 3451
rect 4905 3417 4939 3451
rect 3525 3349 3559 3383
rect 4353 3349 4387 3383
rect 4445 3349 4479 3383
rect 5089 3349 5123 3383
rect 8769 3349 8803 3383
rect 9321 3349 9355 3383
rect 5917 3145 5951 3179
rect 7297 3145 7331 3179
rect 9321 3145 9355 3179
rect 8769 3077 8803 3111
rect 3525 3009 3559 3043
rect 3617 3009 3651 3043
rect 3985 3009 4019 3043
rect 5457 3009 5491 3043
rect 6101 3009 6135 3043
rect 6653 3009 6687 3043
rect 7481 3009 7515 3043
rect 7849 3009 7883 3043
rect 8585 3009 8619 3043
rect 9505 3009 9539 3043
rect 8401 2941 8435 2975
rect 9045 2941 9079 2975
rect 3341 2873 3375 2907
rect 7665 2873 7699 2907
rect 6377 2805 6411 2839
rect 6561 2805 6595 2839
rect 8033 2805 8067 2839
rect 3341 2601 3375 2635
rect 4905 2601 4939 2635
rect 6285 2601 6319 2635
rect 7665 2601 7699 2635
rect 9413 2533 9447 2567
rect 7021 2465 7055 2499
rect 7941 2465 7975 2499
rect 3525 2397 3559 2431
rect 3801 2397 3835 2431
rect 4169 2397 4203 2431
rect 4629 2397 4663 2431
rect 5089 2397 5123 2431
rect 5273 2397 5307 2431
rect 5733 2397 5767 2431
rect 6101 2397 6135 2431
rect 6377 2397 6411 2431
rect 7297 2397 7331 2431
rect 7481 2397 7515 2431
rect 9321 2397 9355 2431
rect 3617 2261 3651 2295
rect 4445 2261 4479 2295
rect 5457 2261 5491 2295
rect 5917 2261 5951 2295
rect 7113 2261 7147 2295
rect 3893 2057 3927 2091
rect 4997 2057 5031 2091
rect 6193 2057 6227 2091
rect 6837 2057 6871 2091
rect 7113 2057 7147 2091
rect 7389 2057 7423 2091
rect 9229 2057 9263 2091
rect 6561 1989 6595 2023
rect 8861 1989 8895 2023
rect 9045 1989 9079 2023
rect 3617 1921 3651 1955
rect 4077 1921 4111 1955
rect 4905 1921 4939 1955
rect 5181 1921 5215 1955
rect 5457 1921 5491 1955
rect 5733 1921 5767 1955
rect 6009 1921 6043 1955
rect 7021 1921 7055 1955
rect 7297 1921 7331 1955
rect 7573 1921 7607 1955
rect 7849 1921 7883 1955
rect 8493 1921 8527 1955
rect 9505 1921 9539 1955
rect 4445 1853 4479 1887
rect 4721 1785 4755 1819
rect 5549 1785 5583 1819
rect 8033 1785 8067 1819
rect 8677 1785 8711 1819
rect 9321 1785 9355 1819
rect 5273 1717 5307 1751
rect 4445 1513 4479 1547
rect 4721 1513 4755 1547
rect 5273 1513 5307 1547
rect 4169 1445 4203 1479
rect 8953 1445 8987 1479
rect 9413 1445 9447 1479
rect 7573 1377 7607 1411
rect 3525 1309 3559 1343
rect 3801 1309 3835 1343
rect 4077 1309 4111 1343
rect 4353 1309 4387 1343
rect 4629 1309 4663 1343
rect 4905 1309 4939 1343
rect 5181 1309 5215 1343
rect 5457 1309 5491 1343
rect 5917 1309 5951 1343
rect 6193 1309 6227 1343
rect 6653 1309 6687 1343
rect 8585 1309 8619 1343
rect 8861 1309 8895 1343
rect 9137 1309 9171 1343
rect 3341 1173 3375 1207
rect 3617 1173 3651 1207
rect 3893 1173 3927 1207
rect 4997 1173 5031 1207
rect 5733 1173 5767 1207
rect 6009 1173 6043 1207
rect 6745 1173 6779 1207
rect 7205 1173 7239 1207
rect 7941 1173 7975 1207
rect 8401 1173 8435 1207
rect 8677 1173 8711 1207
rect 9229 1173 9263 1207
<< metal1 >>
rect 2130 11840 2136 11892
rect 2188 11880 2194 11892
rect 7006 11880 7012 11892
rect 2188 11852 7012 11880
rect 2188 11840 2194 11852
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 16666 11880 16672 11892
rect 13872 11852 16672 11880
rect 13872 11840 13878 11852
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 2774 11772 2780 11824
rect 2832 11812 2838 11824
rect 3786 11812 3792 11824
rect 2832 11784 3792 11812
rect 2832 11772 2838 11784
rect 3786 11772 3792 11784
rect 3844 11772 3850 11824
rect 3970 11772 3976 11824
rect 4028 11812 4034 11824
rect 5534 11812 5540 11824
rect 4028 11784 5540 11812
rect 4028 11772 4034 11784
rect 5534 11772 5540 11784
rect 5592 11772 5598 11824
rect 2958 11704 2964 11756
rect 3016 11744 3022 11756
rect 8662 11744 8668 11756
rect 3016 11716 8668 11744
rect 3016 11704 3022 11716
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 1486 11636 1492 11688
rect 1544 11676 1550 11688
rect 5442 11676 5448 11688
rect 1544 11648 5448 11676
rect 1544 11636 1550 11648
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 1302 11568 1308 11620
rect 1360 11608 1366 11620
rect 5534 11608 5540 11620
rect 1360 11580 5540 11608
rect 1360 11568 1366 11580
rect 5534 11568 5540 11580
rect 5592 11568 5598 11620
rect 5902 11568 5908 11620
rect 5960 11608 5966 11620
rect 6454 11608 6460 11620
rect 5960 11580 6460 11608
rect 5960 11568 5966 11580
rect 6454 11568 6460 11580
rect 6512 11568 6518 11620
rect 3142 11500 3148 11552
rect 3200 11540 3206 11552
rect 6362 11540 6368 11552
rect 3200 11512 6368 11540
rect 3200 11500 3206 11512
rect 6362 11500 6368 11512
rect 6420 11500 6426 11552
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 7566 11450
rect 7618 11398 7630 11450
rect 7682 11398 7694 11450
rect 7746 11398 7758 11450
rect 7810 11398 7822 11450
rect 7874 11398 9844 11450
rect 920 11376 9844 11398
rect 1302 11336 1308 11348
rect 1263 11308 1308 11336
rect 1302 11296 1308 11308
rect 1360 11296 1366 11348
rect 1765 11339 1823 11345
rect 1765 11305 1777 11339
rect 1811 11336 1823 11339
rect 4522 11336 4528 11348
rect 1811 11308 4528 11336
rect 1811 11305 1823 11308
rect 1765 11299 1823 11305
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 5813 11339 5871 11345
rect 5813 11305 5825 11339
rect 5859 11336 5871 11339
rect 8386 11336 8392 11348
rect 5859 11308 8392 11336
rect 5859 11305 5871 11308
rect 5813 11299 5871 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 8481 11339 8539 11345
rect 8481 11305 8493 11339
rect 8527 11336 8539 11339
rect 9306 11336 9312 11348
rect 8527 11308 9312 11336
rect 8527 11305 8539 11308
rect 8481 11299 8539 11305
rect 9306 11296 9312 11308
rect 9364 11296 9370 11348
rect 9401 11339 9459 11345
rect 9401 11305 9413 11339
rect 9447 11336 9459 11339
rect 10870 11336 10876 11348
rect 9447 11308 10876 11336
rect 9447 11305 9459 11308
rect 9401 11299 9459 11305
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 2041 11271 2099 11277
rect 2041 11237 2053 11271
rect 2087 11237 2099 11271
rect 2041 11231 2099 11237
rect 2056 11200 2084 11231
rect 2130 11228 2136 11280
rect 2188 11268 2194 11280
rect 2869 11271 2927 11277
rect 2188 11240 2233 11268
rect 2188 11228 2194 11240
rect 2869 11237 2881 11271
rect 2915 11237 2927 11271
rect 2869 11231 2927 11237
rect 2884 11200 2912 11231
rect 2958 11228 2964 11280
rect 3016 11268 3022 11280
rect 3016 11240 3061 11268
rect 3016 11228 3022 11240
rect 3142 11228 3148 11280
rect 3200 11268 3206 11280
rect 3237 11271 3295 11277
rect 3237 11268 3249 11271
rect 3200 11240 3249 11268
rect 3200 11228 3206 11240
rect 3237 11237 3249 11240
rect 3283 11237 3295 11271
rect 3237 11231 3295 11237
rect 3326 11228 3332 11280
rect 3384 11268 3390 11280
rect 6365 11271 6423 11277
rect 3384 11240 6316 11268
rect 3384 11228 3390 11240
rect 1596 11172 2084 11200
rect 2424 11172 2912 11200
rect 1486 11132 1492 11144
rect 1447 11104 1492 11132
rect 1486 11092 1492 11104
rect 1544 11092 1550 11144
rect 1596 11141 1624 11172
rect 1581 11135 1639 11141
rect 1581 11101 1593 11135
rect 1627 11101 1639 11135
rect 1854 11132 1860 11144
rect 1815 11104 1860 11132
rect 1581 11095 1639 11101
rect 1854 11092 1860 11104
rect 1912 11092 1918 11144
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2424 11141 2452 11172
rect 4338 11160 4344 11212
rect 4396 11160 4402 11212
rect 4433 11203 4491 11209
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 4890 11200 4896 11212
rect 4479 11172 4896 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 6288 11200 6316 11240
rect 6365 11237 6377 11271
rect 6411 11268 6423 11271
rect 7466 11268 7472 11280
rect 6411 11240 7472 11268
rect 6411 11237 6423 11240
rect 6365 11231 6423 11237
rect 7466 11228 7472 11240
rect 7524 11228 7530 11280
rect 7745 11271 7803 11277
rect 7745 11237 7757 11271
rect 7791 11268 7803 11271
rect 9582 11268 9588 11280
rect 7791 11240 9588 11268
rect 7791 11237 7803 11240
rect 7745 11231 7803 11237
rect 9582 11228 9588 11240
rect 9640 11228 9646 11280
rect 6730 11200 6736 11212
rect 6288 11172 6736 11200
rect 6730 11160 6736 11172
rect 6788 11160 6794 11212
rect 11146 11200 11152 11212
rect 8680 11172 11152 11200
rect 2317 11135 2375 11141
rect 2317 11132 2329 11135
rect 2280 11104 2329 11132
rect 2280 11092 2286 11104
rect 2317 11101 2329 11104
rect 2363 11101 2375 11135
rect 2317 11095 2375 11101
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11101 2743 11135
rect 2685 11095 2743 11101
rect 3145 11135 3203 11141
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 3326 11132 3332 11144
rect 3191 11104 3332 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 2700 11064 2728 11095
rect 3326 11092 3332 11104
rect 3384 11092 3390 11144
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 3602 11132 3608 11144
rect 3467 11104 3608 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 3789 11135 3847 11141
rect 3789 11101 3801 11135
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11132 4123 11135
rect 4356 11132 4384 11160
rect 4706 11132 4712 11144
rect 4111 11104 4384 11132
rect 4667 11104 4712 11132
rect 4111 11101 4123 11104
rect 4065 11095 4123 11101
rect 3804 11064 3832 11095
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11132 6055 11135
rect 6454 11132 6460 11144
rect 6043 11104 6460 11132
rect 6043 11101 6055 11104
rect 5997 11095 6055 11101
rect 2424 11036 3832 11064
rect 4249 11067 4307 11073
rect 2424 11008 2452 11036
rect 4249 11033 4261 11067
rect 4295 11064 4307 11067
rect 4338 11064 4344 11076
rect 4295 11036 4344 11064
rect 4295 11033 4307 11036
rect 4249 11027 4307 11033
rect 4338 11024 4344 11036
rect 4396 11024 4402 11076
rect 5736 11064 5764 11095
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 6546 11092 6552 11144
rect 6604 11132 6610 11144
rect 6604 11104 6649 11132
rect 6748 11104 7328 11132
rect 6604 11092 6610 11104
rect 6178 11064 6184 11076
rect 5736 11036 6184 11064
rect 6178 11024 6184 11036
rect 6236 11064 6242 11076
rect 6641 11067 6699 11073
rect 6641 11064 6653 11067
rect 6236 11036 6653 11064
rect 6236 11024 6242 11036
rect 6641 11033 6653 11036
rect 6687 11064 6699 11067
rect 6748 11064 6776 11104
rect 6687 11036 6776 11064
rect 6825 11067 6883 11073
rect 6687 11033 6699 11036
rect 6641 11027 6699 11033
rect 6825 11033 6837 11067
rect 6871 11033 6883 11067
rect 6825 11027 6883 11033
rect 7009 11067 7067 11073
rect 7009 11033 7021 11067
rect 7055 11064 7067 11067
rect 7098 11064 7104 11076
rect 7055 11036 7104 11064
rect 7055 11033 7067 11036
rect 7009 11027 7067 11033
rect 14 10956 20 11008
rect 72 10996 78 11008
rect 934 10996 940 11008
rect 72 10968 940 10996
rect 72 10956 78 10968
rect 934 10956 940 10968
rect 992 10956 998 11008
rect 2406 10956 2412 11008
rect 2464 10956 2470 11008
rect 2590 10996 2596 11008
rect 2551 10968 2596 10996
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 2682 10956 2688 11008
rect 2740 10996 2746 11008
rect 3973 10999 4031 11005
rect 3973 10996 3985 10999
rect 2740 10968 3985 10996
rect 2740 10956 2746 10968
rect 3973 10965 3985 10968
rect 4019 10965 4031 10999
rect 3973 10959 4031 10965
rect 4982 10956 4988 11008
rect 5040 10996 5046 11008
rect 5353 10999 5411 11005
rect 5353 10996 5365 10999
rect 5040 10968 5365 10996
rect 5040 10956 5046 10968
rect 5353 10965 5365 10968
rect 5399 10965 5411 10999
rect 5353 10959 5411 10965
rect 5537 10999 5595 11005
rect 5537 10965 5549 10999
rect 5583 10996 5595 10999
rect 5718 10996 5724 11008
rect 5583 10968 5724 10996
rect 5583 10965 5595 10968
rect 5537 10959 5595 10965
rect 5718 10956 5724 10968
rect 5776 10956 5782 11008
rect 6546 10956 6552 11008
rect 6604 10996 6610 11008
rect 6840 10996 6868 11027
rect 7098 11024 7104 11036
rect 7156 11024 7162 11076
rect 7300 11005 7328 11104
rect 7374 11092 7380 11144
rect 7432 11132 7438 11144
rect 7469 11135 7527 11141
rect 7469 11132 7481 11135
rect 7432 11104 7481 11132
rect 7432 11092 7438 11104
rect 7469 11101 7481 11104
rect 7515 11101 7527 11135
rect 7469 11095 7527 11101
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11132 7619 11135
rect 7834 11132 7840 11144
rect 7607 11104 7840 11132
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 7484 11064 7512 11095
rect 7834 11092 7840 11104
rect 7892 11092 7898 11144
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11132 7987 11135
rect 8018 11132 8024 11144
rect 7975 11104 8024 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 8018 11092 8024 11104
rect 8076 11092 8082 11144
rect 8294 11132 8300 11144
rect 8255 11104 8300 11132
rect 8294 11092 8300 11104
rect 8352 11092 8358 11144
rect 8478 11064 8484 11076
rect 7484 11036 8484 11064
rect 8478 11024 8484 11036
rect 8536 11024 8542 11076
rect 6604 10968 6868 10996
rect 7285 10999 7343 11005
rect 6604 10956 6610 10968
rect 7285 10965 7297 10999
rect 7331 10965 7343 10999
rect 7285 10959 7343 10965
rect 8113 10999 8171 11005
rect 8113 10965 8125 10999
rect 8159 10996 8171 10999
rect 8680 10996 8708 11172
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 8849 11135 8907 11141
rect 8849 11101 8861 11135
rect 8895 11132 8907 11135
rect 9122 11132 9128 11144
rect 8895 11104 9128 11132
rect 8895 11101 8907 11104
rect 8849 11095 8907 11101
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 8754 11024 8760 11076
rect 8812 11064 8818 11076
rect 9232 11064 9260 11095
rect 9306 11092 9312 11144
rect 9364 11132 9370 11144
rect 10410 11132 10416 11144
rect 9364 11104 10416 11132
rect 9364 11092 9370 11104
rect 10410 11092 10416 11104
rect 10468 11092 10474 11144
rect 10686 11064 10692 11076
rect 8812 11036 9260 11064
rect 9324 11036 10692 11064
rect 8812 11024 8818 11036
rect 8159 10968 8708 10996
rect 9033 10999 9091 11005
rect 8159 10965 8171 10968
rect 8113 10959 8171 10965
rect 9033 10965 9045 10999
rect 9079 10996 9091 10999
rect 9324 10996 9352 11036
rect 10686 11024 10692 11036
rect 10744 11024 10750 11076
rect 9079 10968 9352 10996
rect 9079 10965 9091 10968
rect 9033 10959 9091 10965
rect 920 10906 9844 10928
rect 920 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 5194 10906
rect 5246 10854 5258 10906
rect 5310 10854 5322 10906
rect 5374 10854 9844 10906
rect 920 10832 9844 10854
rect 2501 10795 2559 10801
rect 2501 10761 2513 10795
rect 2547 10792 2559 10795
rect 6086 10792 6092 10804
rect 2547 10764 6092 10792
rect 2547 10761 2559 10764
rect 2501 10755 2559 10761
rect 6086 10752 6092 10764
rect 6144 10752 6150 10804
rect 6196 10764 7604 10792
rect 2774 10680 2780 10692
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1213 10659 1271 10665
rect 1213 10656 1225 10659
rect 992 10628 1225 10656
rect 992 10616 998 10628
rect 1213 10625 1225 10628
rect 1259 10625 1271 10659
rect 1213 10619 1271 10625
rect 1946 10616 1952 10668
rect 2004 10656 2010 10668
rect 2225 10659 2283 10665
rect 2225 10656 2237 10659
rect 2004 10628 2237 10656
rect 2004 10616 2010 10628
rect 2225 10625 2237 10628
rect 2271 10625 2283 10659
rect 2225 10619 2283 10625
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10625 2375 10659
rect 2735 10652 2780 10680
rect 2774 10640 2780 10652
rect 2832 10640 2838 10692
rect 3878 10684 3884 10736
rect 3936 10684 3942 10736
rect 5074 10684 5080 10736
rect 5132 10724 5138 10736
rect 6196 10724 6224 10764
rect 5132 10696 6224 10724
rect 7576 10710 7604 10764
rect 5132 10684 5138 10696
rect 2317 10619 2375 10625
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 2332 10588 2360 10619
rect 4706 10616 4712 10668
rect 4764 10616 4770 10668
rect 4890 10656 4896 10668
rect 4851 10628 4896 10656
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10656 5043 10659
rect 5166 10656 5172 10668
rect 5031 10628 5172 10656
rect 5031 10625 5043 10628
rect 4985 10619 5043 10625
rect 5166 10616 5172 10628
rect 5224 10656 5230 10668
rect 5537 10659 5595 10665
rect 5537 10656 5549 10659
rect 5224 10628 5549 10656
rect 5224 10616 5230 10628
rect 5537 10625 5549 10628
rect 5583 10625 5595 10659
rect 5718 10656 5724 10668
rect 5679 10628 5724 10656
rect 5537 10619 5595 10625
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 6273 10659 6331 10665
rect 6273 10625 6285 10659
rect 6319 10656 6331 10659
rect 6546 10656 6552 10668
rect 6319 10628 6552 10656
rect 6319 10625 6331 10628
rect 6273 10619 6331 10625
rect 6546 10616 6552 10628
rect 6604 10656 6610 10668
rect 7282 10656 7288 10668
rect 6604 10628 7288 10656
rect 6604 10616 6610 10628
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 9030 10656 9036 10668
rect 8711 10628 9036 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 9217 10659 9275 10665
rect 9217 10625 9229 10659
rect 9263 10656 9275 10659
rect 16574 10656 16580 10668
rect 9263 10628 16580 10656
rect 9263 10625 9275 10628
rect 9217 10619 9275 10625
rect 2682 10588 2688 10600
rect 1728 10560 1992 10588
rect 2332 10560 2688 10588
rect 1728 10548 1734 10560
rect 1578 10480 1584 10532
rect 1636 10520 1642 10532
rect 1857 10523 1915 10529
rect 1857 10520 1869 10523
rect 1636 10492 1869 10520
rect 1636 10480 1642 10492
rect 1857 10489 1869 10492
rect 1903 10489 1915 10523
rect 1964 10520 1992 10560
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 2858 10591 2916 10597
rect 2858 10588 2870 10591
rect 2792 10560 2870 10588
rect 2792 10520 2820 10560
rect 2858 10557 2870 10560
rect 2904 10557 2916 10591
rect 2858 10551 2916 10557
rect 3510 10548 3516 10600
rect 3568 10588 3574 10600
rect 4617 10591 4675 10597
rect 4617 10588 4629 10591
rect 3568 10560 4629 10588
rect 3568 10548 3574 10560
rect 4617 10557 4629 10560
rect 4663 10588 4675 10591
rect 4724 10588 4752 10616
rect 5442 10588 5448 10600
rect 4663 10560 4752 10588
rect 5403 10560 5448 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 5868 10560 6837 10588
rect 5868 10548 5874 10560
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 7190 10588 7196 10600
rect 7151 10560 7196 10588
rect 6825 10551 6883 10557
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 1964 10492 2820 10520
rect 1857 10483 1915 10489
rect 4338 10480 4344 10532
rect 4396 10520 4402 10532
rect 5905 10523 5963 10529
rect 5905 10520 5917 10523
rect 4396 10492 5917 10520
rect 4396 10480 4402 10492
rect 5905 10489 5917 10492
rect 5951 10489 5963 10523
rect 5905 10483 5963 10489
rect 6270 10480 6276 10532
rect 6328 10520 6334 10532
rect 6733 10523 6791 10529
rect 6733 10520 6745 10523
rect 6328 10492 6745 10520
rect 6328 10480 6334 10492
rect 6733 10489 6745 10492
rect 6779 10489 6791 10523
rect 6733 10483 6791 10489
rect 8110 10480 8116 10532
rect 8168 10520 8174 10532
rect 9232 10520 9260 10619
rect 16574 10616 16580 10628
rect 16632 10616 16638 10668
rect 8168 10492 9260 10520
rect 8168 10480 8174 10492
rect 2038 10452 2044 10464
rect 1999 10424 2044 10452
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 2593 10455 2651 10461
rect 2593 10421 2605 10455
rect 2639 10452 2651 10455
rect 2958 10452 2964 10464
rect 2639 10424 2964 10452
rect 2639 10421 2651 10424
rect 2593 10415 2651 10421
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 3142 10461 3148 10464
rect 3132 10455 3148 10461
rect 3132 10421 3144 10455
rect 3132 10415 3148 10421
rect 3142 10412 3148 10415
rect 3200 10412 3206 10464
rect 4709 10455 4767 10461
rect 4709 10421 4721 10455
rect 4755 10452 4767 10455
rect 4890 10452 4896 10464
rect 4755 10424 4896 10452
rect 4755 10421 4767 10424
rect 4709 10415 4767 10421
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 5261 10455 5319 10461
rect 5261 10421 5273 10455
rect 5307 10452 5319 10455
rect 5994 10452 6000 10464
rect 5307 10424 6000 10452
rect 5307 10421 5319 10424
rect 5261 10415 5319 10421
rect 5994 10412 6000 10424
rect 6052 10452 6058 10464
rect 6365 10455 6423 10461
rect 6365 10452 6377 10455
rect 6052 10424 6377 10452
rect 6052 10412 6058 10424
rect 6365 10421 6377 10424
rect 6411 10421 6423 10455
rect 6365 10415 6423 10421
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 8938 10452 8944 10464
rect 6604 10424 8944 10452
rect 6604 10412 6610 10424
rect 8938 10412 8944 10424
rect 8996 10412 9002 10464
rect 9125 10455 9183 10461
rect 9125 10421 9137 10455
rect 9171 10452 9183 10455
rect 9214 10452 9220 10464
rect 9171 10424 9220 10452
rect 9171 10421 9183 10424
rect 9125 10415 9183 10421
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 9306 10412 9312 10464
rect 9364 10452 9370 10464
rect 9401 10455 9459 10461
rect 9401 10452 9413 10455
rect 9364 10424 9413 10452
rect 9364 10412 9370 10424
rect 9401 10421 9413 10424
rect 9447 10421 9459 10455
rect 9401 10415 9459 10421
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 7566 10362
rect 7618 10310 7630 10362
rect 7682 10310 7694 10362
rect 7746 10310 7758 10362
rect 7810 10310 7822 10362
rect 7874 10310 9844 10362
rect 920 10288 9844 10310
rect 2038 10208 2044 10260
rect 2096 10248 2102 10260
rect 2096 10220 6408 10248
rect 2096 10208 2102 10220
rect 3142 10140 3148 10192
rect 3200 10180 3206 10192
rect 3418 10180 3424 10192
rect 3200 10152 3424 10180
rect 3200 10140 3206 10152
rect 3418 10140 3424 10152
rect 3476 10140 3482 10192
rect 1670 10112 1676 10124
rect 1631 10084 1676 10112
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 1946 10072 1952 10124
rect 2004 10112 2010 10124
rect 4338 10112 4344 10124
rect 2004 10084 4344 10112
rect 2004 10072 2010 10084
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 4522 10112 4528 10124
rect 4483 10084 4528 10112
rect 4522 10072 4528 10084
rect 4580 10072 4586 10124
rect 5258 10112 5264 10124
rect 4908 10084 5264 10112
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 1578 10004 1584 10056
rect 1636 10004 1642 10056
rect 3602 10044 3608 10056
rect 3563 10016 3608 10044
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 4062 10044 4068 10056
rect 3804 10016 4068 10044
rect 1596 9976 1624 10004
rect 1949 9979 2007 9985
rect 1596 9948 1900 9976
rect 1486 9868 1492 9920
rect 1544 9908 1550 9920
rect 1581 9911 1639 9917
rect 1581 9908 1593 9911
rect 1544 9880 1593 9908
rect 1544 9868 1550 9880
rect 1581 9877 1593 9880
rect 1627 9877 1639 9911
rect 1872 9908 1900 9948
rect 1949 9945 1961 9979
rect 1995 9976 2007 9979
rect 2222 9976 2228 9988
rect 1995 9948 2228 9976
rect 1995 9945 2007 9948
rect 1949 9939 2007 9945
rect 2222 9936 2228 9948
rect 2280 9936 2286 9988
rect 3326 9976 3332 9988
rect 3174 9948 3332 9976
rect 3326 9936 3332 9948
rect 3384 9976 3390 9988
rect 3804 9976 3832 10016
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 4908 10053 4936 10084
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10013 4951 10047
rect 4893 10007 4951 10013
rect 5902 10004 5908 10056
rect 5960 10044 5966 10056
rect 6380 10053 6408 10220
rect 6546 10208 6552 10260
rect 6604 10248 6610 10260
rect 6825 10251 6883 10257
rect 6825 10248 6837 10251
rect 6604 10220 6837 10248
rect 6604 10208 6610 10220
rect 6825 10217 6837 10220
rect 6871 10217 6883 10251
rect 6825 10211 6883 10217
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 9493 10251 9551 10257
rect 9493 10248 9505 10251
rect 7248 10220 9505 10248
rect 7248 10208 7254 10220
rect 9493 10217 9505 10220
rect 9539 10217 9551 10251
rect 9493 10211 9551 10217
rect 6730 10140 6736 10192
rect 6788 10180 6794 10192
rect 7285 10183 7343 10189
rect 7285 10180 7297 10183
rect 6788 10152 7297 10180
rect 6788 10140 6794 10152
rect 7285 10149 7297 10152
rect 7331 10149 7343 10183
rect 7285 10143 7343 10149
rect 8481 10183 8539 10189
rect 8481 10149 8493 10183
rect 8527 10180 8539 10183
rect 11054 10180 11060 10192
rect 8527 10152 11060 10180
rect 8527 10149 8539 10152
rect 8481 10143 8539 10149
rect 11054 10140 11060 10152
rect 11112 10140 11118 10192
rect 6365 10047 6423 10053
rect 5960 10016 6132 10044
rect 5960 10004 5966 10016
rect 3384 9948 3832 9976
rect 3384 9936 3390 9948
rect 3878 9936 3884 9988
rect 3936 9976 3942 9988
rect 3936 9948 4568 9976
rect 3936 9936 3942 9948
rect 2958 9908 2964 9920
rect 1872 9880 2964 9908
rect 1581 9871 1639 9877
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 4249 9911 4307 9917
rect 4249 9908 4261 9911
rect 4212 9880 4261 9908
rect 4212 9868 4218 9880
rect 4249 9877 4261 9880
rect 4295 9877 4307 9911
rect 4540 9908 4568 9948
rect 5534 9936 5540 9988
rect 5592 9936 5598 9988
rect 6104 9976 6132 10016
rect 6365 10013 6377 10047
rect 6411 10013 6423 10047
rect 6914 10044 6920 10056
rect 6875 10016 6920 10044
rect 6365 10007 6423 10013
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 7024 10016 7389 10044
rect 7024 9976 7052 10016
rect 7377 10013 7389 10016
rect 7423 10013 7435 10047
rect 7377 10007 7435 10013
rect 7650 10004 7656 10056
rect 7708 10044 7714 10056
rect 8021 10047 8079 10053
rect 8021 10044 8033 10047
rect 7708 10016 8033 10044
rect 7708 10004 7714 10016
rect 8021 10013 8033 10016
rect 8067 10013 8079 10047
rect 8297 10047 8355 10053
rect 8297 10044 8309 10047
rect 8021 10007 8079 10013
rect 8128 10016 8309 10044
rect 6104 9948 7052 9976
rect 7101 9979 7159 9985
rect 7101 9945 7113 9979
rect 7147 9976 7159 9979
rect 7190 9976 7196 9988
rect 7147 9948 7196 9976
rect 7147 9945 7159 9948
rect 7101 9939 7159 9945
rect 7190 9936 7196 9948
rect 7248 9976 7254 9988
rect 7561 9979 7619 9985
rect 7561 9976 7573 9979
rect 7248 9948 7573 9976
rect 7248 9936 7254 9948
rect 7561 9945 7573 9948
rect 7607 9945 7619 9979
rect 7561 9939 7619 9945
rect 7745 9911 7803 9917
rect 7745 9908 7757 9911
rect 4540 9880 7757 9908
rect 4249 9871 4307 9877
rect 7745 9877 7757 9880
rect 7791 9877 7803 9911
rect 7745 9871 7803 9877
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 8128 9917 8156 10016
rect 8297 10013 8309 10016
rect 8343 10013 8355 10047
rect 8846 10044 8852 10056
rect 8807 10016 8852 10044
rect 8297 10007 8355 10013
rect 8846 10004 8852 10016
rect 8904 10004 8910 10056
rect 8113 9911 8171 9917
rect 8113 9908 8125 9911
rect 7892 9880 8125 9908
rect 7892 9868 7898 9880
rect 8113 9877 8125 9880
rect 8159 9877 8171 9911
rect 8113 9871 8171 9877
rect 920 9818 9844 9840
rect 920 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 5194 9818
rect 5246 9766 5258 9818
rect 5310 9766 5322 9818
rect 5374 9766 9844 9818
rect 920 9744 9844 9766
rect 1670 9664 1676 9716
rect 1728 9664 1734 9716
rect 2222 9664 2228 9716
rect 2280 9704 2286 9716
rect 8846 9704 8852 9716
rect 2280 9676 8852 9704
rect 2280 9664 2286 9676
rect 8846 9664 8852 9676
rect 8904 9704 8910 9716
rect 9493 9707 9551 9713
rect 9493 9704 9505 9707
rect 8904 9676 9505 9704
rect 8904 9664 8910 9676
rect 9493 9673 9505 9676
rect 9539 9673 9551 9707
rect 9493 9667 9551 9673
rect 1688 9636 1716 9664
rect 2774 9636 2780 9648
rect 1228 9608 1716 9636
rect 2714 9608 2780 9636
rect 1228 9577 1256 9608
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 3786 9596 3792 9648
rect 3844 9596 3850 9648
rect 5442 9596 5448 9648
rect 5500 9636 5506 9648
rect 5718 9636 5724 9648
rect 5500 9608 5724 9636
rect 5500 9596 5506 9608
rect 5718 9596 5724 9608
rect 5776 9596 5782 9648
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 8021 9639 8079 9645
rect 8021 9636 8033 9639
rect 6604 9608 8033 9636
rect 6604 9596 6610 9608
rect 8021 9605 8033 9608
rect 8067 9605 8079 9639
rect 8021 9599 8079 9605
rect 8478 9596 8484 9648
rect 8536 9596 8542 9648
rect 1213 9571 1271 9577
rect 1213 9537 1225 9571
rect 1259 9537 1271 9571
rect 3510 9568 3516 9580
rect 1213 9531 1271 9537
rect 2746 9540 3516 9568
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 2746 9500 2774 9540
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 4890 9568 4896 9580
rect 4851 9540 4896 9568
rect 4890 9528 4896 9540
rect 4948 9528 4954 9580
rect 5350 9528 5356 9580
rect 5408 9568 5414 9580
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 5408 9540 5549 9568
rect 5408 9528 5414 9540
rect 5537 9537 5549 9540
rect 5583 9537 5595 9571
rect 6178 9568 6184 9580
rect 5537 9531 5595 9537
rect 5644 9540 6184 9568
rect 5644 9512 5672 9540
rect 6178 9528 6184 9540
rect 6236 9528 6242 9580
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 6972 9540 7113 9568
rect 6972 9528 6978 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 7374 9528 7380 9580
rect 7432 9568 7438 9580
rect 7742 9568 7748 9580
rect 7432 9540 7604 9568
rect 7703 9540 7748 9568
rect 7432 9528 7438 9540
rect 3050 9500 3056 9512
rect 1636 9472 2774 9500
rect 3011 9472 3056 9500
rect 1636 9460 1642 9472
rect 3050 9460 3056 9472
rect 3108 9460 3114 9512
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9500 3479 9503
rect 4062 9500 4068 9512
rect 3467 9472 4068 9500
rect 3467 9469 3479 9472
rect 3421 9463 3479 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 5626 9460 5632 9512
rect 5684 9460 5690 9512
rect 5718 9460 5724 9512
rect 5776 9500 5782 9512
rect 7576 9509 7604 9540
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 5776 9472 6469 9500
rect 5776 9460 5782 9472
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 7561 9503 7619 9509
rect 6457 9463 6515 9469
rect 7116 9472 7328 9500
rect 2774 9392 2780 9444
rect 2832 9432 2838 9444
rect 2961 9435 3019 9441
rect 2961 9432 2973 9435
rect 2832 9404 2973 9432
rect 2832 9392 2838 9404
rect 2961 9401 2973 9404
rect 3007 9401 3019 9435
rect 5997 9435 6055 9441
rect 5997 9432 6009 9435
rect 2961 9395 3019 9401
rect 4356 9404 6009 9432
rect 1476 9367 1534 9373
rect 1476 9333 1488 9367
rect 1522 9364 1534 9367
rect 2038 9364 2044 9376
rect 1522 9336 2044 9364
rect 1522 9333 1534 9336
rect 1476 9327 1534 9333
rect 2038 9324 2044 9336
rect 2096 9324 2102 9376
rect 3142 9324 3148 9376
rect 3200 9364 3206 9376
rect 4356 9364 4384 9404
rect 5997 9401 6009 9404
rect 6043 9401 6055 9435
rect 5997 9395 6055 9401
rect 3200 9336 4384 9364
rect 5353 9367 5411 9373
rect 3200 9324 3206 9336
rect 5353 9333 5365 9367
rect 5399 9364 5411 9367
rect 5718 9364 5724 9376
rect 5399 9336 5724 9364
rect 5399 9333 5411 9336
rect 5353 9327 5411 9333
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9364 5871 9367
rect 5902 9364 5908 9376
rect 5859 9336 5908 9364
rect 5859 9333 5871 9336
rect 5813 9327 5871 9333
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 7116 9364 7144 9472
rect 7300 9432 7328 9472
rect 7561 9469 7573 9503
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 7760 9432 7788 9528
rect 7300 9404 7788 9432
rect 6236 9336 7144 9364
rect 6236 9324 6242 9336
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 7377 9367 7435 9373
rect 7377 9364 7389 9367
rect 7248 9336 7389 9364
rect 7248 9324 7254 9336
rect 7377 9333 7389 9336
rect 7423 9364 7435 9367
rect 8478 9364 8484 9376
rect 7423 9336 8484 9364
rect 7423 9333 7435 9336
rect 7377 9327 7435 9333
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 7566 9274
rect 7618 9222 7630 9274
rect 7682 9222 7694 9274
rect 7746 9222 7758 9274
rect 7810 9222 7822 9274
rect 7874 9222 9844 9274
rect 920 9200 9844 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 3050 9160 3056 9172
rect 1452 9132 2912 9160
rect 3011 9132 3056 9160
rect 1452 9120 1458 9132
rect 1489 9095 1547 9101
rect 1489 9061 1501 9095
rect 1535 9092 1547 9095
rect 1578 9092 1584 9104
rect 1535 9064 1584 9092
rect 1535 9061 1547 9064
rect 1489 9055 1547 9061
rect 1578 9052 1584 9064
rect 1636 9052 1642 9104
rect 2682 9092 2688 9104
rect 1688 9064 2688 9092
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 1578 8956 1584 8968
rect 1443 8928 1584 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 1578 8916 1584 8928
rect 1636 8916 1642 8968
rect 1688 8965 1716 9064
rect 2682 9052 2688 9064
rect 2740 9052 2746 9104
rect 2777 9095 2835 9101
rect 2777 9061 2789 9095
rect 2823 9061 2835 9095
rect 2884 9092 2912 9132
rect 3050 9120 3056 9132
rect 3108 9120 3114 9172
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 4249 9163 4307 9169
rect 4249 9160 4261 9163
rect 3660 9132 4261 9160
rect 3660 9120 3666 9132
rect 4249 9129 4261 9132
rect 4295 9129 4307 9163
rect 4249 9123 4307 9129
rect 4522 9120 4528 9172
rect 4580 9160 4586 9172
rect 4617 9163 4675 9169
rect 4617 9160 4629 9163
rect 4580 9132 4629 9160
rect 4580 9120 4586 9132
rect 4617 9129 4629 9132
rect 4663 9160 4675 9163
rect 5074 9160 5080 9172
rect 4663 9132 5080 9160
rect 4663 9129 4675 9132
rect 4617 9123 4675 9129
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5534 9120 5540 9172
rect 5592 9160 5598 9172
rect 8205 9163 8263 9169
rect 5592 9132 7788 9160
rect 5592 9120 5598 9132
rect 3329 9095 3387 9101
rect 3329 9092 3341 9095
rect 2884 9064 3341 9092
rect 2777 9055 2835 9061
rect 3329 9061 3341 9064
rect 3375 9061 3387 9095
rect 3329 9055 3387 9061
rect 2406 8984 2412 9036
rect 2464 9024 2470 9036
rect 2464 8996 2636 9024
rect 2464 8984 2470 8996
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8956 2007 8959
rect 2038 8956 2044 8968
rect 1995 8928 2044 8956
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 2222 8956 2228 8968
rect 2183 8928 2228 8956
rect 2222 8916 2228 8928
rect 2280 8916 2286 8968
rect 842 8848 848 8900
rect 900 8888 906 8900
rect 2424 8888 2452 8984
rect 2608 8965 2636 8996
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8925 2559 8959
rect 2501 8919 2559 8925
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8925 2651 8959
rect 2792 8956 2820 9055
rect 3878 9052 3884 9104
rect 3936 9092 3942 9104
rect 4798 9092 4804 9104
rect 3936 9064 4804 9092
rect 3936 9052 3942 9064
rect 4798 9052 4804 9064
rect 4856 9052 4862 9104
rect 4154 9024 4160 9036
rect 3252 8996 4160 9024
rect 3252 8968 3280 8996
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 4246 8984 4252 9036
rect 4304 9024 4310 9036
rect 5905 9027 5963 9033
rect 5905 9024 5917 9027
rect 4304 8996 5917 9024
rect 4304 8984 4310 8996
rect 5905 8993 5917 8996
rect 5951 8993 5963 9027
rect 5905 8987 5963 8993
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 2792 8928 2881 8956
rect 2593 8919 2651 8925
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 3234 8956 3240 8968
rect 3147 8928 3240 8956
rect 2869 8919 2927 8925
rect 900 8860 1808 8888
rect 900 8848 906 8860
rect 1210 8820 1216 8832
rect 1171 8792 1216 8820
rect 1210 8780 1216 8792
rect 1268 8780 1274 8832
rect 1780 8829 1808 8860
rect 1964 8860 2452 8888
rect 2516 8888 2544 8919
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3418 8916 3424 8968
rect 3476 8956 3482 8968
rect 3605 8959 3663 8965
rect 3605 8956 3617 8959
rect 3476 8928 3617 8956
rect 3476 8916 3482 8928
rect 3605 8925 3617 8928
rect 3651 8925 3663 8959
rect 3605 8919 3663 8925
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4341 8959 4399 8965
rect 4341 8956 4353 8959
rect 4120 8928 4353 8956
rect 4120 8916 4126 8928
rect 4341 8925 4353 8928
rect 4387 8956 4399 8959
rect 4430 8956 4436 8968
rect 4387 8928 4436 8956
rect 4387 8925 4399 8928
rect 4341 8919 4399 8925
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5000 8888 5028 8919
rect 5074 8916 5080 8968
rect 5132 8956 5138 8968
rect 5261 8959 5319 8965
rect 5261 8956 5273 8959
rect 5132 8928 5273 8956
rect 5132 8916 5138 8928
rect 5261 8925 5273 8928
rect 5307 8956 5319 8959
rect 6270 8956 6276 8968
rect 5307 8928 5764 8956
rect 6231 8928 6276 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 5626 8888 5632 8900
rect 2516 8860 4844 8888
rect 5000 8860 5632 8888
rect 1964 8832 1992 8860
rect 1765 8823 1823 8829
rect 1765 8789 1777 8823
rect 1811 8789 1823 8823
rect 1765 8783 1823 8789
rect 1946 8780 1952 8832
rect 2004 8780 2010 8832
rect 2041 8823 2099 8829
rect 2041 8789 2053 8823
rect 2087 8820 2099 8823
rect 2130 8820 2136 8832
rect 2087 8792 2136 8820
rect 2087 8789 2099 8792
rect 2041 8783 2099 8789
rect 2130 8780 2136 8792
rect 2188 8780 2194 8832
rect 2317 8823 2375 8829
rect 2317 8789 2329 8823
rect 2363 8820 2375 8823
rect 3786 8820 3792 8832
rect 2363 8792 3792 8820
rect 2363 8789 2375 8792
rect 2317 8783 2375 8789
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 4816 8829 4844 8860
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 4801 8823 4859 8829
rect 4801 8789 4813 8823
rect 4847 8789 4859 8823
rect 5736 8820 5764 8928
rect 6270 8916 6276 8928
rect 6328 8916 6334 8968
rect 7760 8965 7788 9132
rect 8205 9129 8217 9163
rect 8251 9160 8263 9163
rect 8294 9160 8300 9172
rect 8251 9132 8300 9160
rect 8251 9129 8263 9132
rect 8205 9123 8263 9129
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 8202 8984 8208 9036
rect 8260 9024 8266 9036
rect 8570 9024 8576 9036
rect 8260 8996 8576 9024
rect 8260 8984 8266 8996
rect 8570 8984 8576 8996
rect 8628 9024 8634 9036
rect 9125 9027 9183 9033
rect 9125 9024 9137 9027
rect 8628 8996 9137 9024
rect 8628 8984 8634 8996
rect 9125 8993 9137 8996
rect 9171 8993 9183 9027
rect 9125 8987 9183 8993
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8925 7803 8959
rect 7745 8919 7803 8925
rect 8018 8916 8024 8968
rect 8076 8956 8082 8968
rect 8297 8959 8355 8965
rect 8297 8956 8309 8959
rect 8076 8928 8309 8956
rect 8076 8916 8082 8928
rect 8297 8925 8309 8928
rect 8343 8925 8355 8959
rect 8846 8956 8852 8968
rect 8807 8928 8852 8956
rect 8297 8919 8355 8925
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 7006 8848 7012 8900
rect 7064 8848 7070 8900
rect 7190 8820 7196 8832
rect 5736 8792 7196 8820
rect 4801 8783 4859 8789
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 8481 8823 8539 8829
rect 8481 8789 8493 8823
rect 8527 8820 8539 8823
rect 9582 8820 9588 8832
rect 8527 8792 9588 8820
rect 8527 8789 8539 8792
rect 8481 8783 8539 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 920 8730 9844 8752
rect 920 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 5194 8730
rect 5246 8678 5258 8730
rect 5310 8678 5322 8730
rect 5374 8678 9844 8730
rect 920 8656 9844 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 1762 8616 1768 8628
rect 1452 8588 1768 8616
rect 1452 8576 1458 8588
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 2133 8619 2191 8625
rect 2133 8616 2145 8619
rect 1872 8588 2145 8616
rect 1394 8480 1400 8492
rect 1355 8452 1400 8480
rect 1394 8440 1400 8452
rect 1452 8440 1458 8492
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 1872 8480 1900 8588
rect 2133 8585 2145 8588
rect 2179 8585 2191 8619
rect 2133 8579 2191 8585
rect 2409 8619 2467 8625
rect 2409 8585 2421 8619
rect 2455 8585 2467 8619
rect 2409 8579 2467 8585
rect 1719 8452 1900 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 1946 8440 1952 8492
rect 2004 8480 2010 8492
rect 2225 8483 2283 8489
rect 2004 8452 2049 8480
rect 2004 8440 2010 8452
rect 2225 8449 2237 8483
rect 2271 8480 2283 8483
rect 2314 8480 2320 8492
rect 2271 8452 2320 8480
rect 2271 8449 2283 8452
rect 2225 8443 2283 8449
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 1762 8372 1768 8424
rect 1820 8412 1826 8424
rect 1964 8412 1992 8440
rect 2424 8412 2452 8579
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 2869 8619 2927 8625
rect 2869 8616 2881 8619
rect 2832 8588 2881 8616
rect 2832 8576 2838 8588
rect 2869 8585 2881 8588
rect 2915 8585 2927 8619
rect 5534 8616 5540 8628
rect 2869 8579 2927 8585
rect 3896 8588 5540 8616
rect 2501 8551 2559 8557
rect 2501 8517 2513 8551
rect 2547 8548 2559 8551
rect 3896 8548 3924 8588
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 7006 8616 7012 8628
rect 6788 8588 7012 8616
rect 6788 8576 6794 8588
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 7190 8576 7196 8628
rect 7248 8616 7254 8628
rect 8570 8616 8576 8628
rect 7248 8588 8576 8616
rect 7248 8576 7254 8588
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 9122 8616 9128 8628
rect 9083 8588 9128 8616
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 2547 8520 2636 8548
rect 2547 8517 2559 8520
rect 2501 8511 2559 8517
rect 2608 8424 2636 8520
rect 2700 8520 3924 8548
rect 2700 8489 2728 8520
rect 3970 8508 3976 8560
rect 4028 8548 4034 8560
rect 4706 8548 4712 8560
rect 4028 8520 4712 8548
rect 4028 8508 4034 8520
rect 4706 8508 4712 8520
rect 4764 8508 4770 8560
rect 4982 8508 4988 8560
rect 5040 8548 5046 8560
rect 5040 8520 5764 8548
rect 5040 8508 5046 8520
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 1820 8384 2452 8412
rect 1820 8372 1826 8384
rect 2590 8372 2596 8424
rect 2648 8372 2654 8424
rect 2406 8304 2412 8356
rect 2464 8344 2470 8356
rect 2698 8344 2726 8443
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 2961 8483 3019 8489
rect 2961 8480 2973 8483
rect 2832 8452 2973 8480
rect 2832 8440 2838 8452
rect 2961 8449 2973 8452
rect 3007 8449 3019 8483
rect 2961 8443 3019 8449
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8480 3571 8483
rect 3602 8480 3608 8492
rect 3559 8452 3608 8480
rect 3559 8449 3571 8452
rect 3513 8443 3571 8449
rect 3602 8440 3608 8452
rect 3660 8440 3666 8492
rect 4430 8480 4436 8492
rect 4391 8452 4436 8480
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5626 8480 5632 8492
rect 5215 8452 5632 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 5736 8480 5764 8520
rect 5902 8508 5908 8560
rect 5960 8548 5966 8560
rect 5960 8520 6408 8548
rect 5960 8508 5966 8520
rect 6380 8492 6408 8520
rect 7558 8508 7564 8560
rect 7616 8508 7622 8560
rect 6181 8483 6239 8489
rect 6181 8480 6193 8483
rect 5736 8452 6193 8480
rect 6181 8449 6193 8452
rect 6227 8449 6239 8483
rect 6362 8480 6368 8492
rect 6323 8452 6368 8480
rect 6181 8443 6239 8449
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 6822 8480 6828 8492
rect 6783 8452 6828 8480
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 7190 8480 7196 8492
rect 7151 8452 7196 8480
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 8662 8480 8668 8492
rect 8623 8452 8668 8480
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 9217 8483 9275 8489
rect 9217 8480 9229 8483
rect 8996 8452 9229 8480
rect 8996 8440 9002 8452
rect 9217 8449 9229 8452
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 2866 8372 2872 8424
rect 2924 8412 2930 8424
rect 3421 8415 3479 8421
rect 3421 8412 3433 8415
rect 2924 8384 3433 8412
rect 2924 8372 2930 8384
rect 3421 8381 3433 8384
rect 3467 8381 3479 8415
rect 3421 8375 3479 8381
rect 5445 8415 5503 8421
rect 5445 8381 5457 8415
rect 5491 8412 5503 8415
rect 5902 8412 5908 8424
rect 5491 8384 5908 8412
rect 5491 8381 5503 8384
rect 5445 8375 5503 8381
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 2464 8316 2726 8344
rect 2464 8304 2470 8316
rect 3326 8304 3332 8356
rect 3384 8344 3390 8356
rect 3786 8344 3792 8356
rect 3384 8316 3792 8344
rect 3384 8304 3390 8316
rect 3786 8304 3792 8316
rect 3844 8304 3850 8356
rect 4154 8344 4160 8356
rect 4115 8316 4160 8344
rect 4154 8304 4160 8316
rect 4212 8304 4218 8356
rect 4706 8304 4712 8356
rect 4764 8344 4770 8356
rect 6086 8344 6092 8356
rect 4764 8316 6092 8344
rect 4764 8304 4770 8316
rect 6086 8304 6092 8316
rect 6144 8304 6150 8356
rect 9401 8347 9459 8353
rect 9401 8313 9413 8347
rect 9447 8344 9459 8347
rect 10962 8344 10968 8356
rect 9447 8316 10968 8344
rect 9447 8313 9459 8316
rect 9401 8307 9459 8313
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 1578 8276 1584 8288
rect 1539 8248 1584 8276
rect 1578 8236 1584 8248
rect 1636 8236 1642 8288
rect 1857 8279 1915 8285
rect 1857 8245 1869 8279
rect 1903 8276 1915 8279
rect 1946 8276 1952 8288
rect 1903 8248 1952 8276
rect 1903 8245 1915 8248
rect 1857 8239 1915 8245
rect 1946 8236 1952 8248
rect 2004 8236 2010 8288
rect 3145 8279 3203 8285
rect 3145 8245 3157 8279
rect 3191 8276 3203 8279
rect 4246 8276 4252 8288
rect 3191 8248 4252 8276
rect 3191 8245 3203 8248
rect 3145 8239 3203 8245
rect 4246 8236 4252 8248
rect 4304 8276 4310 8288
rect 4522 8276 4528 8288
rect 4304 8248 4528 8276
rect 4304 8236 4310 8248
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 5077 8279 5135 8285
rect 5077 8245 5089 8279
rect 5123 8276 5135 8279
rect 5442 8276 5448 8288
rect 5123 8248 5448 8276
rect 5123 8245 5135 8248
rect 5077 8239 5135 8245
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 5534 8236 5540 8288
rect 5592 8276 5598 8288
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 5592 8248 6561 8276
rect 5592 8236 5598 8248
rect 6549 8245 6561 8248
rect 6595 8245 6607 8279
rect 6549 8239 6607 8245
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 7566 8186
rect 7618 8134 7630 8186
rect 7682 8134 7694 8186
rect 7746 8134 7758 8186
rect 7810 8134 7822 8186
rect 7874 8134 9844 8186
rect 920 8112 9844 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 1489 8075 1547 8081
rect 1489 8072 1501 8075
rect 1452 8044 1501 8072
rect 1452 8032 1458 8044
rect 1489 8041 1501 8044
rect 1535 8041 1547 8075
rect 1489 8035 1547 8041
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 1949 8075 2007 8081
rect 1949 8072 1961 8075
rect 1912 8044 1961 8072
rect 1912 8032 1918 8044
rect 1949 8041 1961 8044
rect 1995 8041 2007 8075
rect 1949 8035 2007 8041
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 2958 8072 2964 8084
rect 2915 8044 2964 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 2958 8032 2964 8044
rect 3016 8032 3022 8084
rect 3237 8075 3295 8081
rect 3237 8041 3249 8075
rect 3283 8072 3295 8075
rect 4246 8072 4252 8084
rect 3283 8044 4252 8072
rect 3283 8041 3295 8044
rect 3237 8035 3295 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4430 8032 4436 8084
rect 4488 8072 4494 8084
rect 4798 8072 4804 8084
rect 4488 8044 4804 8072
rect 4488 8032 4494 8044
rect 4798 8032 4804 8044
rect 4856 8072 4862 8084
rect 5537 8075 5595 8081
rect 5537 8072 5549 8075
rect 4856 8044 5549 8072
rect 4856 8032 4862 8044
rect 5537 8041 5549 8044
rect 5583 8041 5595 8075
rect 5537 8035 5595 8041
rect 6454 8032 6460 8084
rect 6512 8072 6518 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 6512 8044 7849 8072
rect 6512 8032 6518 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 8570 8072 8576 8084
rect 8531 8044 8576 8072
rect 7837 8035 7895 8041
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 8754 8072 8760 8084
rect 8715 8044 8760 8072
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 1673 8007 1731 8013
rect 1673 7973 1685 8007
rect 1719 8004 1731 8007
rect 2222 8004 2228 8016
rect 1719 7976 2228 8004
rect 1719 7973 1731 7976
rect 1673 7967 1731 7973
rect 2222 7964 2228 7976
rect 2280 7964 2286 8016
rect 3421 8007 3479 8013
rect 2700 7976 3372 8004
rect 1762 7936 1768 7948
rect 1320 7908 1768 7936
rect 1320 7877 1348 7908
rect 1762 7896 1768 7908
rect 1820 7896 1826 7948
rect 2700 7936 2728 7976
rect 2240 7908 2728 7936
rect 3344 7936 3372 7976
rect 3421 7973 3433 8007
rect 3467 8004 3479 8007
rect 3786 8004 3792 8016
rect 3467 7976 3792 8004
rect 3467 7973 3479 7976
rect 3421 7967 3479 7973
rect 3786 7964 3792 7976
rect 3844 7964 3850 8016
rect 6917 8007 6975 8013
rect 6917 8004 6929 8007
rect 5276 7976 6929 8004
rect 5276 7936 5304 7976
rect 6917 7973 6929 7976
rect 6963 8004 6975 8007
rect 7006 8004 7012 8016
rect 6963 7976 7012 8004
rect 6963 7973 6975 7976
rect 6917 7967 6975 7973
rect 7006 7964 7012 7976
rect 7064 7964 7070 8016
rect 7190 7964 7196 8016
rect 7248 8004 7254 8016
rect 7926 8004 7932 8016
rect 7248 7976 7932 8004
rect 7248 7964 7254 7976
rect 7926 7964 7932 7976
rect 7984 7964 7990 8016
rect 3344 7908 5304 7936
rect 1305 7871 1363 7877
rect 1305 7837 1317 7871
rect 1351 7837 1363 7871
rect 1305 7831 1363 7837
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 1854 7868 1860 7880
rect 1627 7840 1860 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 1854 7828 1860 7840
rect 1912 7828 1918 7880
rect 2240 7877 2268 7908
rect 9214 7896 9220 7948
rect 9272 7936 9278 7948
rect 9309 7939 9367 7945
rect 9309 7936 9321 7939
rect 9272 7908 9321 7936
rect 9272 7896 9278 7908
rect 9309 7905 9321 7908
rect 9355 7905 9367 7939
rect 9309 7899 9367 7905
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7837 2283 7871
rect 2225 7831 2283 7837
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7868 2559 7871
rect 2961 7871 3019 7877
rect 2961 7868 2973 7871
rect 2547 7840 2973 7868
rect 2547 7837 2559 7840
rect 2501 7831 2559 7837
rect 2961 7837 2973 7840
rect 3007 7868 3019 7871
rect 3050 7868 3056 7880
rect 3007 7840 3056 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 3050 7828 3056 7840
rect 3108 7828 3114 7880
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3344 7840 3801 7868
rect 2406 7760 2412 7812
rect 2464 7800 2470 7812
rect 2685 7803 2743 7809
rect 2685 7800 2697 7803
rect 2464 7772 2697 7800
rect 2464 7760 2470 7772
rect 2685 7769 2697 7772
rect 2731 7769 2743 7803
rect 2685 7763 2743 7769
rect 1670 7692 1676 7744
rect 1728 7732 1734 7744
rect 2317 7735 2375 7741
rect 2317 7732 2329 7735
rect 1728 7704 2329 7732
rect 1728 7692 1734 7704
rect 2317 7701 2329 7704
rect 2363 7732 2375 7735
rect 3344 7732 3372 7840
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 5626 7868 5632 7880
rect 5587 7840 5632 7868
rect 3789 7831 3847 7837
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 7282 7828 7288 7880
rect 7340 7868 7346 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7340 7840 7665 7868
rect 7340 7828 7346 7840
rect 7653 7837 7665 7840
rect 7699 7868 7711 7871
rect 7929 7871 7987 7877
rect 7699 7840 7880 7868
rect 7699 7837 7711 7840
rect 7653 7831 7711 7837
rect 4065 7803 4123 7809
rect 4065 7769 4077 7803
rect 4111 7769 4123 7803
rect 5994 7800 6000 7812
rect 5290 7772 6000 7800
rect 4065 7763 4123 7769
rect 2363 7704 3372 7732
rect 4080 7732 4108 7763
rect 5994 7760 6000 7772
rect 6052 7760 6058 7812
rect 7469 7803 7527 7809
rect 7469 7800 7481 7803
rect 6196 7772 7481 7800
rect 4246 7732 4252 7744
rect 4080 7704 4252 7732
rect 2363 7701 2375 7704
rect 2317 7695 2375 7701
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 4430 7692 4436 7744
rect 4488 7732 4494 7744
rect 6196 7732 6224 7772
rect 7469 7769 7481 7772
rect 7515 7800 7527 7803
rect 7742 7800 7748 7812
rect 7515 7772 7748 7800
rect 7515 7769 7527 7772
rect 7469 7763 7527 7769
rect 7742 7760 7748 7772
rect 7800 7760 7806 7812
rect 7852 7800 7880 7840
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8202 7868 8208 7880
rect 7975 7840 8208 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8202 7828 8208 7840
rect 8260 7828 8266 7880
rect 8478 7800 8484 7812
rect 7852 7772 8484 7800
rect 8478 7760 8484 7772
rect 8536 7760 8542 7812
rect 9125 7803 9183 7809
rect 9125 7769 9137 7803
rect 9171 7800 9183 7803
rect 9398 7800 9404 7812
rect 9171 7772 9404 7800
rect 9171 7769 9183 7772
rect 9125 7763 9183 7769
rect 9398 7760 9404 7772
rect 9456 7760 9462 7812
rect 4488 7704 6224 7732
rect 4488 7692 4494 7704
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 9217 7735 9275 7741
rect 9217 7732 9229 7735
rect 6604 7704 9229 7732
rect 6604 7692 6610 7704
rect 9217 7701 9229 7704
rect 9263 7701 9275 7735
rect 9217 7695 9275 7701
rect 920 7642 9844 7664
rect 920 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 5194 7642
rect 5246 7590 5258 7642
rect 5310 7590 5322 7642
rect 5374 7590 9844 7642
rect 920 7568 9844 7590
rect 1118 7488 1124 7540
rect 1176 7528 1182 7540
rect 1213 7531 1271 7537
rect 1213 7528 1225 7531
rect 1176 7500 1225 7528
rect 1176 7488 1182 7500
rect 1213 7497 1225 7500
rect 1259 7497 1271 7531
rect 1213 7491 1271 7497
rect 1673 7531 1731 7537
rect 1673 7497 1685 7531
rect 1719 7528 1731 7531
rect 5810 7528 5816 7540
rect 1719 7500 5816 7528
rect 1719 7497 1731 7500
rect 1673 7491 1731 7497
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 5997 7531 6055 7537
rect 5997 7497 6009 7531
rect 6043 7528 6055 7531
rect 6270 7528 6276 7540
rect 6043 7500 6276 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 8573 7531 8631 7537
rect 8573 7528 8585 7531
rect 6880 7500 8585 7528
rect 6880 7488 6886 7500
rect 8573 7497 8585 7500
rect 8619 7497 8631 7531
rect 8573 7491 8631 7497
rect 1026 7420 1032 7472
rect 1084 7460 1090 7472
rect 1854 7460 1860 7472
rect 1084 7432 1860 7460
rect 1084 7420 1090 7432
rect 1854 7420 1860 7432
rect 1912 7420 1918 7472
rect 2133 7463 2191 7469
rect 2133 7429 2145 7463
rect 2179 7460 2191 7463
rect 2179 7432 2636 7460
rect 2179 7429 2191 7432
rect 2133 7423 2191 7429
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7361 1455 7395
rect 1397 7355 1455 7361
rect 1412 7256 1440 7355
rect 1486 7352 1492 7404
rect 1544 7392 1550 7404
rect 1762 7392 1768 7404
rect 1544 7364 1589 7392
rect 1723 7364 1768 7392
rect 1544 7352 1550 7364
rect 1762 7352 1768 7364
rect 1820 7352 1826 7404
rect 1946 7352 1952 7404
rect 2004 7392 2010 7404
rect 2041 7395 2099 7401
rect 2041 7392 2053 7395
rect 2004 7364 2053 7392
rect 2004 7352 2010 7364
rect 2041 7361 2053 7364
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 2406 7352 2412 7404
rect 2464 7392 2470 7404
rect 2501 7395 2559 7401
rect 2501 7392 2513 7395
rect 2464 7364 2513 7392
rect 2464 7352 2470 7364
rect 2501 7361 2513 7364
rect 2547 7361 2559 7395
rect 2608 7392 2636 7432
rect 3510 7420 3516 7472
rect 3568 7420 3574 7472
rect 4798 7420 4804 7472
rect 4856 7460 4862 7472
rect 6549 7463 6607 7469
rect 6549 7460 6561 7463
rect 4856 7432 6561 7460
rect 4856 7420 4862 7432
rect 6549 7429 6561 7432
rect 6595 7429 6607 7463
rect 8294 7460 8300 7472
rect 7774 7432 8300 7460
rect 6549 7423 6607 7429
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 2608 7364 2728 7392
rect 2501 7355 2559 7361
rect 1578 7284 1584 7336
rect 1636 7324 1642 7336
rect 2581 7327 2639 7333
rect 2581 7324 2593 7327
rect 1636 7296 2593 7324
rect 1636 7284 1642 7296
rect 2581 7293 2593 7296
rect 2627 7293 2639 7327
rect 2581 7287 2639 7293
rect 2038 7256 2044 7268
rect 1412 7228 2044 7256
rect 2038 7216 2044 7228
rect 2096 7216 2102 7268
rect 1949 7191 2007 7197
rect 1949 7157 1961 7191
rect 1995 7188 2007 7191
rect 2222 7188 2228 7200
rect 1995 7160 2228 7188
rect 1995 7157 2007 7160
rect 1949 7151 2007 7157
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 2406 7188 2412 7200
rect 2363 7160 2412 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 2700 7188 2728 7364
rect 3878 7352 3884 7404
rect 3936 7392 3942 7404
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 3936 7364 4445 7392
rect 3936 7352 3942 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7392 5043 7395
rect 5353 7395 5411 7401
rect 5031 7364 5212 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 2958 7284 2964 7336
rect 3016 7324 3022 7336
rect 3016 7296 3061 7324
rect 3016 7284 3022 7296
rect 4522 7216 4528 7268
rect 4580 7256 4586 7268
rect 4798 7256 4804 7268
rect 4580 7228 4804 7256
rect 4580 7216 4586 7228
rect 4798 7216 4804 7228
rect 4856 7216 4862 7268
rect 4893 7259 4951 7265
rect 4893 7225 4905 7259
rect 4939 7256 4951 7259
rect 5000 7256 5028 7355
rect 4939 7228 5028 7256
rect 5184 7256 5212 7364
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 5442 7392 5448 7404
rect 5399 7364 5448 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 6178 7352 6184 7404
rect 6236 7392 6242 7404
rect 6273 7395 6331 7401
rect 6273 7392 6285 7395
rect 6236 7364 6285 7392
rect 6236 7352 6242 7364
rect 6273 7361 6285 7364
rect 6319 7361 6331 7395
rect 6273 7355 6331 7361
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 7892 7364 8125 7392
rect 7892 7352 7898 7364
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 9033 7395 9091 7401
rect 9033 7392 9045 7395
rect 8113 7355 8171 7361
rect 8220 7364 9045 7392
rect 6380 7296 7604 7324
rect 5534 7256 5540 7268
rect 5184 7228 5540 7256
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 5534 7216 5540 7228
rect 5592 7216 5598 7268
rect 5994 7216 6000 7268
rect 6052 7256 6058 7268
rect 6380 7256 6408 7296
rect 6052 7228 6408 7256
rect 7576 7256 7604 7296
rect 7926 7284 7932 7336
rect 7984 7324 7990 7336
rect 8021 7327 8079 7333
rect 8021 7324 8033 7327
rect 7984 7296 8033 7324
rect 7984 7284 7990 7296
rect 8021 7293 8033 7296
rect 8067 7293 8079 7327
rect 8021 7287 8079 7293
rect 8220 7256 8248 7364
rect 9033 7361 9045 7364
rect 9079 7361 9091 7395
rect 9033 7355 9091 7361
rect 9122 7324 9128 7336
rect 9083 7296 9128 7324
rect 9122 7284 9128 7296
rect 9180 7284 9186 7336
rect 9214 7284 9220 7336
rect 9272 7324 9278 7336
rect 9272 7296 9317 7324
rect 9272 7284 9278 7296
rect 7576 7228 8248 7256
rect 6052 7216 6058 7228
rect 2958 7188 2964 7200
rect 2700 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3602 7148 3608 7200
rect 3660 7188 3666 7200
rect 4430 7188 4436 7200
rect 3660 7160 4436 7188
rect 3660 7148 3666 7160
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 5169 7191 5227 7197
rect 5169 7157 5181 7191
rect 5215 7188 5227 7191
rect 6730 7188 6736 7200
rect 5215 7160 6736 7188
rect 5215 7157 5227 7160
rect 5169 7151 5227 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 8389 7191 8447 7197
rect 8389 7157 8401 7191
rect 8435 7188 8447 7191
rect 8570 7188 8576 7200
rect 8435 7160 8576 7188
rect 8435 7157 8447 7160
rect 8389 7151 8447 7157
rect 8570 7148 8576 7160
rect 8628 7148 8634 7200
rect 8662 7148 8668 7200
rect 8720 7188 8726 7200
rect 8720 7160 8765 7188
rect 8720 7148 8726 7160
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 7566 7098
rect 7618 7046 7630 7098
rect 7682 7046 7694 7098
rect 7746 7046 7758 7098
rect 7810 7046 7822 7098
rect 7874 7046 9844 7098
rect 920 7024 9844 7046
rect 934 6944 940 6996
rect 992 6984 998 6996
rect 1930 6987 1988 6993
rect 1930 6984 1942 6987
rect 992 6956 1942 6984
rect 992 6944 998 6956
rect 1930 6953 1942 6956
rect 1976 6953 1988 6987
rect 1930 6947 1988 6953
rect 2406 6944 2412 6996
rect 2464 6984 2470 6996
rect 2464 6956 6316 6984
rect 2464 6944 2470 6956
rect 6288 6916 6316 6956
rect 6822 6944 6828 6996
rect 6880 6984 6886 6996
rect 7374 6984 7380 6996
rect 6880 6956 7380 6984
rect 6880 6944 6886 6956
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 8757 6987 8815 6993
rect 8757 6953 8769 6987
rect 8803 6984 8815 6987
rect 9122 6984 9128 6996
rect 8803 6956 9128 6984
rect 8803 6953 8815 6956
rect 8757 6947 8815 6953
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 11146 6944 11152 6996
rect 11204 6984 11210 6996
rect 16666 6984 16672 6996
rect 11204 6956 16672 6984
rect 11204 6944 11210 6956
rect 16666 6944 16672 6956
rect 16724 6944 16730 6996
rect 6288 6888 6408 6916
rect 1946 6848 1952 6860
rect 1412 6820 1952 6848
rect 1412 6789 1440 6820
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 3694 6848 3700 6860
rect 3068 6820 3700 6848
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6749 1455 6783
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1397 6743 1455 6749
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 3068 6766 3096 6820
rect 3694 6808 3700 6820
rect 3752 6808 3758 6860
rect 4614 6808 4620 6860
rect 4672 6848 4678 6860
rect 4672 6820 5028 6848
rect 4672 6808 4678 6820
rect 5000 6792 5028 6820
rect 3510 6780 3516 6792
rect 3436 6752 3516 6780
rect 1578 6672 1584 6724
rect 1636 6712 1642 6724
rect 1636 6684 2176 6712
rect 1636 6672 1642 6684
rect 1489 6647 1547 6653
rect 1489 6613 1501 6647
rect 1535 6644 1547 6647
rect 2038 6644 2044 6656
rect 1535 6616 2044 6644
rect 1535 6613 1547 6616
rect 1489 6607 1547 6613
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 2148 6644 2176 6684
rect 2866 6644 2872 6656
rect 2148 6616 2872 6644
rect 2866 6604 2872 6616
rect 2924 6604 2930 6656
rect 3234 6604 3240 6656
rect 3292 6644 3298 6656
rect 3436 6653 3464 6752
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 4154 6780 4160 6792
rect 3651 6752 4160 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 4522 6780 4528 6792
rect 4483 6752 4528 6780
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 4890 6780 4896 6792
rect 4851 6752 4896 6780
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 4982 6740 4988 6792
rect 5040 6740 5046 6792
rect 6380 6789 6408 6888
rect 6454 6808 6460 6860
rect 6512 6848 6518 6860
rect 6512 6820 7880 6848
rect 6512 6808 6518 6820
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6780 6975 6783
rect 7006 6780 7012 6792
rect 6963 6752 7012 6780
rect 6963 6749 6975 6752
rect 6917 6743 6975 6749
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 7098 6740 7104 6792
rect 7156 6780 7162 6792
rect 7852 6789 7880 6820
rect 8202 6808 8208 6860
rect 8260 6848 8266 6860
rect 8573 6851 8631 6857
rect 8573 6848 8585 6851
rect 8260 6820 8585 6848
rect 8260 6808 8266 6820
rect 8573 6817 8585 6820
rect 8619 6817 8631 6851
rect 8573 6811 8631 6817
rect 9030 6808 9036 6860
rect 9088 6848 9094 6860
rect 9309 6851 9367 6857
rect 9309 6848 9321 6851
rect 9088 6820 9321 6848
rect 9088 6808 9094 6820
rect 9309 6817 9321 6820
rect 9355 6817 9367 6851
rect 9309 6811 9367 6817
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7156 6752 7573 6780
rect 7156 6740 7162 6752
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 7926 6740 7932 6792
rect 7984 6780 7990 6792
rect 7984 6752 8029 6780
rect 7984 6740 7990 6752
rect 6026 6684 7696 6712
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 3292 6616 3433 6644
rect 3292 6604 3298 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 3421 6607 3479 6613
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 4249 6647 4307 6653
rect 4249 6644 4261 6647
rect 3568 6616 4261 6644
rect 3568 6604 3574 6616
rect 4249 6613 4261 6616
rect 4295 6613 4307 6647
rect 4249 6607 4307 6613
rect 4982 6604 4988 6656
rect 5040 6644 5046 6656
rect 5626 6644 5632 6656
rect 5040 6616 5632 6644
rect 5040 6604 5046 6616
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 6546 6644 6552 6656
rect 5868 6616 6552 6644
rect 5868 6604 5874 6616
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 6825 6647 6883 6653
rect 6825 6613 6837 6647
rect 6871 6644 6883 6647
rect 7282 6644 7288 6656
rect 6871 6616 7288 6644
rect 6871 6613 6883 6616
rect 6825 6607 6883 6613
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 7668 6653 7696 6684
rect 8386 6672 8392 6724
rect 8444 6712 8450 6724
rect 8570 6712 8576 6724
rect 8444 6684 8576 6712
rect 8444 6672 8450 6684
rect 8570 6672 8576 6684
rect 8628 6672 8634 6724
rect 8846 6672 8852 6724
rect 8904 6712 8910 6724
rect 9217 6715 9275 6721
rect 9217 6712 9229 6715
rect 8904 6684 9229 6712
rect 8904 6672 8910 6684
rect 9217 6681 9229 6684
rect 9263 6681 9275 6715
rect 9217 6675 9275 6681
rect 7653 6647 7711 6653
rect 7653 6613 7665 6647
rect 7699 6613 7711 6647
rect 9122 6644 9128 6656
rect 9083 6616 9128 6644
rect 7653 6607 7711 6613
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 920 6554 9844 6576
rect 920 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 5194 6554
rect 5246 6502 5258 6554
rect 5310 6502 5322 6554
rect 5374 6502 9844 6554
rect 920 6480 9844 6502
rect 1489 6443 1547 6449
rect 1489 6409 1501 6443
rect 1535 6440 1547 6443
rect 1578 6440 1584 6452
rect 1535 6412 1584 6440
rect 1535 6409 1547 6412
rect 1489 6403 1547 6409
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 1762 6400 1768 6452
rect 1820 6440 1826 6452
rect 1949 6443 2007 6449
rect 1949 6440 1961 6443
rect 1820 6412 1961 6440
rect 1820 6400 1826 6412
rect 1949 6409 1961 6412
rect 1995 6409 2007 6443
rect 1949 6403 2007 6409
rect 2222 6400 2228 6452
rect 2280 6440 2286 6452
rect 6546 6440 6552 6452
rect 2280 6412 6552 6440
rect 2280 6400 2286 6412
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 8018 6440 8024 6452
rect 6656 6412 8024 6440
rect 3418 6332 3424 6384
rect 3476 6332 3482 6384
rect 6656 6372 6684 6412
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 5000 6344 6684 6372
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6304 1455 6307
rect 1486 6304 1492 6316
rect 1443 6276 1492 6304
rect 1443 6273 1455 6276
rect 1397 6267 1455 6273
rect 1486 6264 1492 6276
rect 1544 6264 1550 6316
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 1673 6307 1731 6313
rect 1673 6304 1685 6307
rect 1636 6276 1685 6304
rect 1636 6264 1642 6276
rect 1673 6273 1685 6276
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6273 1823 6307
rect 2038 6304 2044 6316
rect 1999 6276 2044 6304
rect 1765 6267 1823 6273
rect 1780 6236 1808 6267
rect 2038 6264 2044 6276
rect 2096 6264 2102 6316
rect 2317 6307 2375 6313
rect 2317 6273 2329 6307
rect 2363 6304 2375 6307
rect 2363 6276 2820 6304
rect 2363 6273 2375 6276
rect 2317 6267 2375 6273
rect 1780 6208 2268 6236
rect 1213 6171 1271 6177
rect 1213 6137 1225 6171
rect 1259 6168 1271 6171
rect 2130 6168 2136 6180
rect 1259 6140 2136 6168
rect 1259 6137 1271 6140
rect 1213 6131 1271 6137
rect 2130 6128 2136 6140
rect 2188 6128 2194 6180
rect 2240 6112 2268 6208
rect 2406 6196 2412 6248
rect 2464 6236 2470 6248
rect 2685 6239 2743 6245
rect 2685 6236 2697 6239
rect 2464 6208 2697 6236
rect 2464 6196 2470 6208
rect 2685 6205 2697 6208
rect 2731 6205 2743 6239
rect 2685 6199 2743 6205
rect 2498 6168 2504 6180
rect 2459 6140 2504 6168
rect 2498 6128 2504 6140
rect 2556 6128 2562 6180
rect 2590 6128 2596 6180
rect 2648 6128 2654 6180
rect 2222 6100 2228 6112
rect 2183 6072 2228 6100
rect 2222 6060 2228 6072
rect 2280 6060 2286 6112
rect 2406 6060 2412 6112
rect 2464 6100 2470 6112
rect 2608 6100 2636 6128
rect 2464 6072 2636 6100
rect 2792 6100 2820 6276
rect 3970 6264 3976 6316
rect 4028 6304 4034 6316
rect 4525 6307 4583 6313
rect 4525 6304 4537 6307
rect 4028 6276 4537 6304
rect 4028 6264 4034 6276
rect 4525 6273 4537 6276
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 3053 6239 3111 6245
rect 3053 6205 3065 6239
rect 3099 6236 3111 6239
rect 3510 6236 3516 6248
rect 3099 6208 3516 6236
rect 3099 6205 3111 6208
rect 3053 6199 3111 6205
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 5000 6245 5028 6344
rect 7466 6332 7472 6384
rect 7524 6332 7530 6384
rect 8404 6344 8708 6372
rect 5718 6264 5724 6316
rect 5776 6304 5782 6316
rect 6086 6304 6092 6316
rect 5776 6276 6092 6304
rect 5776 6264 5782 6276
rect 6086 6264 6092 6276
rect 6144 6304 6150 6316
rect 6181 6307 6239 6313
rect 6181 6304 6193 6307
rect 6144 6276 6193 6304
rect 6144 6264 6150 6276
rect 6181 6273 6193 6276
rect 6227 6273 6239 6307
rect 6181 6267 6239 6273
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 6604 6276 6745 6304
rect 6604 6264 6610 6276
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 8018 6264 8024 6316
rect 8076 6304 8082 6316
rect 8404 6304 8432 6344
rect 8570 6304 8576 6316
rect 8076 6276 8432 6304
rect 8531 6276 8576 6304
rect 8076 6264 8082 6276
rect 8570 6264 8576 6276
rect 8628 6264 8634 6316
rect 4985 6239 5043 6245
rect 4985 6205 4997 6239
rect 5031 6205 5043 6239
rect 5166 6236 5172 6248
rect 5127 6208 5172 6236
rect 4985 6199 5043 6205
rect 5166 6196 5172 6208
rect 5224 6196 5230 6248
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6236 5503 6239
rect 5626 6236 5632 6248
rect 5491 6208 5632 6236
rect 5491 6205 5503 6208
rect 5445 6199 5503 6205
rect 5626 6196 5632 6208
rect 5684 6196 5690 6248
rect 6270 6196 6276 6248
rect 6328 6236 6334 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 6328 6208 6653 6236
rect 6328 6196 6334 6208
rect 6641 6205 6653 6208
rect 6687 6205 6699 6239
rect 6641 6199 6699 6205
rect 7101 6239 7159 6245
rect 7101 6205 7113 6239
rect 7147 6236 7159 6239
rect 7466 6236 7472 6248
rect 7147 6208 7472 6236
rect 7147 6205 7159 6208
rect 7101 6199 7159 6205
rect 7466 6196 7472 6208
rect 7524 6196 7530 6248
rect 8680 6236 8708 6344
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 9309 6307 9367 6313
rect 9309 6304 9321 6307
rect 9088 6276 9321 6304
rect 9088 6264 9094 6276
rect 9309 6273 9321 6276
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8680 6208 9137 6236
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9125 6199 9183 6205
rect 8662 6168 8668 6180
rect 3988 6140 6408 6168
rect 3988 6100 4016 6140
rect 2792 6072 4016 6100
rect 2464 6060 2470 6072
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 6273 6103 6331 6109
rect 6273 6100 6285 6103
rect 5592 6072 6285 6100
rect 5592 6060 5598 6072
rect 6273 6069 6285 6072
rect 6319 6069 6331 6103
rect 6380 6100 6408 6140
rect 8036 6140 8668 6168
rect 8036 6100 8064 6140
rect 8662 6128 8668 6140
rect 8720 6128 8726 6180
rect 8754 6100 8760 6112
rect 6380 6072 8064 6100
rect 8715 6072 8760 6100
rect 6273 6063 6331 6069
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 9033 6103 9091 6109
rect 9033 6069 9045 6103
rect 9079 6100 9091 6103
rect 9214 6100 9220 6112
rect 9079 6072 9220 6100
rect 9079 6069 9091 6072
rect 9033 6063 9091 6069
rect 9214 6060 9220 6072
rect 9272 6060 9278 6112
rect 9490 6100 9496 6112
rect 9451 6072 9496 6100
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 7566 6010
rect 7618 5958 7630 6010
rect 7682 5958 7694 6010
rect 7746 5958 7758 6010
rect 7810 5958 7822 6010
rect 7874 5958 9844 6010
rect 920 5936 9844 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 1544 5868 5488 5896
rect 1544 5856 1550 5868
rect 1670 5760 1676 5772
rect 1631 5732 1676 5760
rect 1670 5720 1676 5732
rect 1728 5760 1734 5772
rect 3326 5760 3332 5772
rect 1728 5732 3332 5760
rect 1728 5720 1734 5732
rect 3326 5720 3332 5732
rect 3384 5760 3390 5772
rect 3605 5763 3663 5769
rect 3605 5760 3617 5763
rect 3384 5732 3617 5760
rect 3384 5720 3390 5732
rect 3605 5729 3617 5732
rect 3651 5729 3663 5763
rect 3605 5723 3663 5729
rect 4246 5720 4252 5772
rect 4304 5760 4310 5772
rect 5353 5763 5411 5769
rect 5353 5760 5365 5763
rect 4304 5732 5365 5760
rect 4304 5720 4310 5732
rect 5353 5729 5365 5732
rect 5399 5729 5411 5763
rect 5460 5760 5488 5868
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5592 5868 5637 5896
rect 5592 5856 5598 5868
rect 6086 5856 6092 5908
rect 6144 5896 6150 5908
rect 9490 5896 9496 5908
rect 6144 5868 9496 5896
rect 6144 5856 6150 5868
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 5905 5831 5963 5837
rect 5905 5797 5917 5831
rect 5951 5828 5963 5831
rect 6454 5828 6460 5840
rect 5951 5800 6460 5828
rect 5951 5797 5963 5800
rect 5905 5791 5963 5797
rect 6454 5788 6460 5800
rect 6512 5788 6518 5840
rect 8757 5831 8815 5837
rect 8757 5797 8769 5831
rect 8803 5828 8815 5831
rect 8846 5828 8852 5840
rect 8803 5800 8852 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 8846 5788 8852 5800
rect 8904 5788 8910 5840
rect 6086 5760 6092 5772
rect 5460 5732 6092 5760
rect 5353 5723 5411 5729
rect 6086 5720 6092 5732
rect 6144 5720 6150 5772
rect 6178 5720 6184 5772
rect 6236 5760 6242 5772
rect 6641 5763 6699 5769
rect 6641 5760 6653 5763
rect 6236 5732 6653 5760
rect 6236 5720 6242 5732
rect 6641 5729 6653 5732
rect 6687 5729 6699 5763
rect 6641 5723 6699 5729
rect 6917 5763 6975 5769
rect 6917 5729 6929 5763
rect 6963 5760 6975 5763
rect 7926 5760 7932 5772
rect 6963 5732 7932 5760
rect 6963 5729 6975 5732
rect 6917 5723 6975 5729
rect 7926 5720 7932 5732
rect 7984 5720 7990 5772
rect 8938 5720 8944 5772
rect 8996 5760 9002 5772
rect 9309 5763 9367 5769
rect 9309 5760 9321 5763
rect 8996 5732 9321 5760
rect 8996 5720 9002 5732
rect 9309 5729 9321 5732
rect 9355 5729 9367 5763
rect 9309 5723 9367 5729
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 5368 5664 5457 5692
rect 1949 5627 2007 5633
rect 1949 5593 1961 5627
rect 1995 5593 2007 5627
rect 3881 5627 3939 5633
rect 3174 5596 3832 5624
rect 1949 5587 2007 5593
rect 1397 5559 1455 5565
rect 1397 5525 1409 5559
rect 1443 5556 1455 5559
rect 1762 5556 1768 5568
rect 1443 5528 1768 5556
rect 1443 5525 1455 5528
rect 1397 5519 1455 5525
rect 1762 5516 1768 5528
rect 1820 5516 1826 5568
rect 1964 5556 1992 5587
rect 3234 5556 3240 5568
rect 1964 5528 3240 5556
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 3421 5559 3479 5565
rect 3421 5525 3433 5559
rect 3467 5556 3479 5559
rect 3602 5556 3608 5568
rect 3467 5528 3608 5556
rect 3467 5525 3479 5528
rect 3421 5519 3479 5525
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 3804 5556 3832 5596
rect 3881 5593 3893 5627
rect 3927 5624 3939 5627
rect 4154 5624 4160 5636
rect 3927 5596 4160 5624
rect 3927 5593 3939 5596
rect 3881 5587 3939 5593
rect 4154 5584 4160 5596
rect 4212 5584 4218 5636
rect 5166 5624 5172 5636
rect 5106 5596 5172 5624
rect 5166 5584 5172 5596
rect 5224 5584 5230 5636
rect 3970 5556 3976 5568
rect 3752 5528 3976 5556
rect 3752 5516 3758 5528
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 5368 5556 5396 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 5592 5664 6561 5692
rect 5592 5652 5598 5664
rect 6549 5661 6561 5664
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 8812 5664 9137 5692
rect 8812 5652 8818 5664
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 6086 5584 6092 5636
rect 6144 5624 6150 5636
rect 6181 5627 6239 5633
rect 6181 5624 6193 5627
rect 6144 5596 6193 5624
rect 6144 5584 6150 5596
rect 6181 5593 6193 5596
rect 6227 5593 6239 5627
rect 6181 5587 6239 5593
rect 6362 5584 6368 5636
rect 6420 5624 6426 5636
rect 8202 5624 8208 5636
rect 6420 5596 6513 5624
rect 8142 5596 8208 5624
rect 6420 5584 6426 5596
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 8662 5584 8668 5636
rect 8720 5624 8726 5636
rect 9030 5624 9036 5636
rect 8720 5596 9036 5624
rect 8720 5584 8726 5596
rect 9030 5584 9036 5596
rect 9088 5584 9094 5636
rect 4672 5528 5396 5556
rect 4672 5516 4678 5528
rect 5626 5516 5632 5568
rect 5684 5556 5690 5568
rect 6380 5556 6408 5584
rect 5684 5528 6408 5556
rect 8389 5559 8447 5565
rect 5684 5516 5690 5528
rect 8389 5525 8401 5559
rect 8435 5556 8447 5559
rect 8478 5556 8484 5568
rect 8435 5528 8484 5556
rect 8435 5525 8447 5528
rect 8389 5519 8447 5525
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 9122 5556 9128 5568
rect 8628 5528 9128 5556
rect 8628 5516 8634 5528
rect 9122 5516 9128 5528
rect 9180 5556 9186 5568
rect 9217 5559 9275 5565
rect 9217 5556 9229 5559
rect 9180 5528 9229 5556
rect 9180 5516 9186 5528
rect 9217 5525 9229 5528
rect 9263 5525 9275 5559
rect 9217 5519 9275 5525
rect 920 5466 9844 5488
rect 920 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 5194 5466
rect 5246 5414 5258 5466
rect 5310 5414 5322 5466
rect 5374 5414 9844 5466
rect 920 5392 9844 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 2406 5352 2412 5364
rect 1452 5324 2412 5352
rect 1452 5312 1458 5324
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 3694 5312 3700 5364
rect 3752 5352 3758 5364
rect 3878 5352 3884 5364
rect 3752 5324 3884 5352
rect 3752 5312 3758 5324
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 6086 5352 6092 5364
rect 3988 5324 6092 5352
rect 1946 5176 1952 5228
rect 2004 5216 2010 5228
rect 2590 5216 2596 5228
rect 2004 5188 2596 5216
rect 2004 5176 2010 5188
rect 2590 5176 2596 5188
rect 2648 5176 2654 5228
rect 2866 5176 2872 5228
rect 2924 5216 2930 5228
rect 3421 5219 3479 5225
rect 3421 5216 3433 5219
rect 2924 5188 3433 5216
rect 2924 5176 2930 5188
rect 3421 5185 3433 5188
rect 3467 5216 3479 5219
rect 3988 5216 4016 5324
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 7466 5312 7472 5364
rect 7524 5352 7530 5364
rect 8941 5355 8999 5361
rect 8941 5352 8953 5355
rect 7524 5324 8953 5352
rect 7524 5312 7530 5324
rect 8941 5321 8953 5324
rect 8987 5321 8999 5355
rect 8941 5315 8999 5321
rect 4798 5244 4804 5296
rect 4856 5244 4862 5296
rect 7926 5284 7932 5296
rect 7866 5256 7932 5284
rect 7926 5244 7932 5256
rect 7984 5284 7990 5296
rect 8202 5284 8208 5296
rect 7984 5256 8208 5284
rect 7984 5244 7990 5256
rect 8202 5244 8208 5256
rect 8260 5244 8266 5296
rect 5810 5216 5816 5228
rect 3467 5188 4016 5216
rect 5771 5188 5816 5216
rect 3467 5185 3479 5188
rect 3421 5179 3479 5185
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6236 5188 6377 5216
rect 6236 5176 6242 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5216 8355 5219
rect 8386 5216 8392 5228
rect 8343 5188 8392 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 8386 5176 8392 5188
rect 8444 5176 8450 5228
rect 9214 5216 9220 5228
rect 9175 5188 9220 5216
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 2222 5108 2228 5160
rect 2280 5148 2286 5160
rect 3970 5148 3976 5160
rect 2280 5120 3976 5148
rect 2280 5108 2286 5120
rect 3970 5108 3976 5120
rect 4028 5108 4034 5160
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 4080 5120 4353 5148
rect 3510 5012 3516 5024
rect 3471 4984 3516 5012
rect 3510 4972 3516 4984
rect 3568 4972 3574 5024
rect 3878 5012 3884 5024
rect 3839 4984 3884 5012
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 4080 5012 4108 5120
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5148 6699 5151
rect 6730 5148 6736 5160
rect 6687 5120 6736 5148
rect 6687 5117 6699 5120
rect 6641 5111 6699 5117
rect 6730 5108 6736 5120
rect 6788 5148 6794 5160
rect 8478 5148 8484 5160
rect 6788 5120 8484 5148
rect 6788 5108 6794 5120
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 6086 5040 6092 5092
rect 6144 5080 6150 5092
rect 6144 5052 6500 5080
rect 6144 5040 6150 5052
rect 5718 5012 5724 5024
rect 4080 4984 5724 5012
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 6273 5015 6331 5021
rect 6273 4981 6285 5015
rect 6319 5012 6331 5015
rect 6362 5012 6368 5024
rect 6319 4984 6368 5012
rect 6319 4981 6331 4984
rect 6273 4975 6331 4981
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 6472 5012 6500 5052
rect 8113 5015 8171 5021
rect 8113 5012 8125 5015
rect 6472 4984 8125 5012
rect 8113 4981 8125 4984
rect 8159 4981 8171 5015
rect 8113 4975 8171 4981
rect 9401 5015 9459 5021
rect 9401 4981 9413 5015
rect 9447 5012 9459 5015
rect 16666 5012 16672 5024
rect 9447 4984 16672 5012
rect 9447 4981 9459 4984
rect 9401 4975 9459 4981
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 3036 4922 9844 4944
rect 3036 4870 7566 4922
rect 7618 4870 7630 4922
rect 7682 4870 7694 4922
rect 7746 4870 7758 4922
rect 7810 4870 7822 4922
rect 7874 4870 9844 4922
rect 3036 4848 9844 4870
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4982 4808 4988 4820
rect 4212 4780 4988 4808
rect 4212 4768 4218 4780
rect 4982 4768 4988 4780
rect 5040 4808 5046 4820
rect 5077 4811 5135 4817
rect 5077 4808 5089 4811
rect 5040 4780 5089 4808
rect 5040 4768 5046 4780
rect 5077 4777 5089 4780
rect 5123 4777 5135 4811
rect 5077 4771 5135 4777
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 8294 4808 8300 4820
rect 5408 4780 8300 4808
rect 5408 4768 5414 4780
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 15194 4768 15200 4820
rect 15252 4808 15258 4820
rect 20622 4808 20628 4820
rect 15252 4780 20628 4808
rect 15252 4768 15258 4780
rect 20622 4768 20628 4780
rect 20680 4768 20686 4820
rect 3326 4672 3332 4684
rect 3287 4644 3332 4672
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 3602 4672 3608 4684
rect 3563 4644 3608 4672
rect 3602 4632 3608 4644
rect 3660 4632 3666 4684
rect 4154 4632 4160 4684
rect 4212 4672 4218 4684
rect 4798 4672 4804 4684
rect 4212 4644 4804 4672
rect 4212 4632 4218 4644
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 5626 4672 5632 4684
rect 5184 4644 5632 4672
rect 5184 4613 5212 4644
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 5813 4675 5871 4681
rect 5813 4641 5825 4675
rect 5859 4672 5871 4675
rect 6178 4672 6184 4684
rect 5859 4644 6184 4672
rect 5859 4641 5871 4644
rect 5813 4635 5871 4641
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6638 4632 6644 4684
rect 6696 4672 6702 4684
rect 7653 4675 7711 4681
rect 7653 4672 7665 4675
rect 6696 4644 7665 4672
rect 6696 4632 6702 4644
rect 7653 4641 7665 4644
rect 7699 4641 7711 4675
rect 7653 4635 7711 4641
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4573 5227 4607
rect 5350 4604 5356 4616
rect 5311 4576 5356 4604
rect 5169 4567 5227 4573
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 6089 4539 6147 4545
rect 3418 4428 3424 4480
rect 3476 4468 3482 4480
rect 4816 4468 4844 4522
rect 5460 4508 6040 4536
rect 5460 4468 5488 4508
rect 3476 4440 5488 4468
rect 5537 4471 5595 4477
rect 3476 4428 3482 4440
rect 5537 4437 5549 4471
rect 5583 4468 5595 4471
rect 5902 4468 5908 4480
rect 5583 4440 5908 4468
rect 5583 4437 5595 4440
rect 5537 4431 5595 4437
rect 5902 4428 5908 4440
rect 5960 4428 5966 4480
rect 6012 4468 6040 4508
rect 6089 4505 6101 4539
rect 6135 4536 6147 4539
rect 6178 4536 6184 4548
rect 6135 4508 6184 4536
rect 6135 4505 6147 4508
rect 6089 4499 6147 4505
rect 6178 4496 6184 4508
rect 6236 4496 6242 4548
rect 7650 4536 7656 4548
rect 7314 4522 7656 4536
rect 7300 4508 7656 4522
rect 7300 4468 7328 4508
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 7837 4539 7895 4545
rect 7837 4505 7849 4539
rect 7883 4536 7895 4539
rect 8570 4536 8576 4548
rect 7883 4508 8576 4536
rect 7883 4505 7895 4508
rect 7837 4499 7895 4505
rect 8570 4496 8576 4508
rect 8628 4496 8634 4548
rect 9493 4539 9551 4545
rect 9493 4505 9505 4539
rect 9539 4536 9551 4539
rect 9582 4536 9588 4548
rect 9539 4508 9588 4536
rect 9539 4505 9551 4508
rect 9493 4499 9551 4505
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 6012 4440 7328 4468
rect 7561 4471 7619 4477
rect 7561 4437 7573 4471
rect 7607 4468 7619 4471
rect 8202 4468 8208 4480
rect 7607 4440 8208 4468
rect 7607 4437 7619 4440
rect 7561 4431 7619 4437
rect 8202 4428 8208 4440
rect 8260 4428 8266 4480
rect 3036 4378 9844 4400
rect 3036 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 5194 4378
rect 5246 4326 5258 4378
rect 5310 4326 5322 4378
rect 5374 4326 9844 4378
rect 3036 4304 9844 4326
rect 4154 4224 4160 4276
rect 4212 4264 4218 4276
rect 4801 4267 4859 4273
rect 4801 4264 4813 4267
rect 4212 4236 4813 4264
rect 4212 4224 4218 4236
rect 4801 4233 4813 4236
rect 4847 4233 4859 4267
rect 4801 4227 4859 4233
rect 4982 4224 4988 4276
rect 5040 4264 5046 4276
rect 5040 4236 5396 4264
rect 5040 4224 5046 4236
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 3602 4128 3608 4140
rect 3559 4100 3608 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4706 4128 4712 4140
rect 4295 4100 4712 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4706 4088 4712 4100
rect 4764 4088 4770 4140
rect 4985 4131 5043 4137
rect 4985 4097 4997 4131
rect 5031 4097 5043 4131
rect 4985 4091 5043 4097
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5368 4128 5396 4236
rect 5626 4224 5632 4276
rect 5684 4264 5690 4276
rect 6178 4264 6184 4276
rect 5684 4236 6184 4264
rect 5684 4224 5690 4236
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 6822 4224 6828 4276
rect 6880 4264 6886 4276
rect 7098 4264 7104 4276
rect 6880 4236 7104 4264
rect 6880 4224 6886 4236
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 7466 4196 7472 4208
rect 7314 4168 7472 4196
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 5718 4128 5724 4140
rect 5123 4100 5396 4128
rect 5679 4100 5724 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 3878 4020 3884 4072
rect 3936 4060 3942 4072
rect 5000 4060 5028 4091
rect 5718 4088 5724 4100
rect 5776 4088 5782 4140
rect 7190 4088 7196 4140
rect 7248 4128 7254 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7248 4100 7665 4128
rect 7248 4088 7254 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 8297 4131 8355 4137
rect 8297 4128 8309 4131
rect 8260 4100 8309 4128
rect 8260 4088 8266 4100
rect 8297 4097 8309 4100
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8754 4088 8760 4140
rect 8812 4128 8818 4140
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8812 4100 9045 4128
rect 8812 4088 8818 4100
rect 9033 4097 9045 4100
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 3936 4032 5028 4060
rect 5813 4063 5871 4069
rect 3936 4020 3942 4032
rect 5813 4029 5825 4063
rect 5859 4060 5871 4063
rect 6086 4060 6092 4072
rect 5859 4032 6092 4060
rect 5859 4029 5871 4032
rect 5813 4023 5871 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6181 4063 6239 4069
rect 6181 4029 6193 4063
rect 6227 4060 6239 4063
rect 6822 4060 6828 4072
rect 6227 4032 6828 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 7984 4032 9168 4060
rect 7984 4020 7990 4032
rect 3510 3952 3516 4004
rect 3568 3992 3574 4004
rect 3568 3964 4568 3992
rect 3568 3952 3574 3964
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4540 3933 4568 3964
rect 4614 3952 4620 4004
rect 4672 3992 4678 4004
rect 4709 3995 4767 4001
rect 4709 3992 4721 3995
rect 4672 3964 4721 3992
rect 4672 3952 4678 3964
rect 4709 3961 4721 3964
rect 4755 3961 4767 3995
rect 4709 3955 4767 3961
rect 5166 3952 5172 4004
rect 5224 3992 5230 4004
rect 5534 3992 5540 4004
rect 5224 3964 5540 3992
rect 5224 3952 5230 3964
rect 5534 3952 5540 3964
rect 5592 3952 5598 4004
rect 7098 3952 7104 4004
rect 7156 3992 7162 4004
rect 8941 3995 8999 4001
rect 8941 3992 8953 3995
rect 7156 3964 8953 3992
rect 7156 3952 7162 3964
rect 8941 3961 8953 3964
rect 8987 3961 8999 3995
rect 8941 3955 8999 3961
rect 4157 3927 4215 3933
rect 4157 3924 4169 3927
rect 4120 3896 4169 3924
rect 4120 3884 4126 3896
rect 4157 3893 4169 3896
rect 4203 3893 4215 3927
rect 4157 3887 4215 3893
rect 4525 3927 4583 3933
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 5718 3924 5724 3936
rect 4571 3896 5724 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 6822 3924 6828 3936
rect 6512 3896 6828 3924
rect 6512 3884 6518 3896
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8846 3924 8852 3936
rect 8159 3896 8852 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8846 3884 8852 3896
rect 8904 3884 8910 3936
rect 9140 3933 9168 4032
rect 16574 3992 16580 4004
rect 16546 3952 16580 3992
rect 16632 3952 16638 4004
rect 9125 3927 9183 3933
rect 9125 3893 9137 3927
rect 9171 3893 9183 3927
rect 9125 3887 9183 3893
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 9272 3896 9505 3924
rect 9272 3884 9278 3896
rect 9493 3893 9505 3896
rect 9539 3893 9551 3927
rect 9493 3887 9551 3893
rect 3036 3834 9844 3856
rect 3036 3782 7566 3834
rect 7618 3782 7630 3834
rect 7682 3782 7694 3834
rect 7746 3782 7758 3834
rect 7810 3782 7822 3834
rect 7874 3782 9844 3834
rect 3036 3760 9844 3782
rect 3789 3723 3847 3729
rect 3789 3689 3801 3723
rect 3835 3720 3847 3723
rect 4522 3720 4528 3732
rect 3835 3692 4528 3720
rect 3835 3689 3847 3692
rect 3789 3683 3847 3689
rect 4522 3680 4528 3692
rect 4580 3680 4586 3732
rect 5353 3723 5411 3729
rect 5353 3689 5365 3723
rect 5399 3720 5411 3723
rect 5810 3720 5816 3732
rect 5399 3692 5816 3720
rect 5399 3689 5411 3692
rect 5353 3683 5411 3689
rect 5810 3680 5816 3692
rect 5868 3680 5874 3732
rect 6178 3680 6184 3732
rect 6236 3720 6242 3732
rect 8754 3720 8760 3732
rect 6236 3692 8760 3720
rect 6236 3680 6242 3692
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 8941 3723 8999 3729
rect 8941 3689 8953 3723
rect 8987 3689 8999 3723
rect 8941 3683 8999 3689
rect 4065 3655 4123 3661
rect 4065 3621 4077 3655
rect 4111 3621 4123 3655
rect 4065 3615 4123 3621
rect 2958 3476 2964 3528
rect 3016 3516 3022 3528
rect 3329 3519 3387 3525
rect 3329 3516 3341 3519
rect 3016 3488 3341 3516
rect 3016 3476 3022 3488
rect 3329 3485 3341 3488
rect 3375 3485 3387 3519
rect 3605 3519 3663 3525
rect 3605 3516 3617 3519
rect 3329 3479 3387 3485
rect 3528 3488 3617 3516
rect 3528 3389 3556 3488
rect 3605 3485 3617 3488
rect 3651 3485 3663 3519
rect 3605 3479 3663 3485
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3516 3939 3519
rect 3970 3516 3976 3528
rect 3927 3488 3976 3516
rect 3927 3485 3939 3488
rect 3881 3479 3939 3485
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 4080 3516 4108 3615
rect 4890 3612 4896 3664
rect 4948 3652 4954 3664
rect 6365 3655 6423 3661
rect 6365 3652 6377 3655
rect 4948 3624 6377 3652
rect 4948 3612 4954 3624
rect 6365 3621 6377 3624
rect 6411 3621 6423 3655
rect 6365 3615 6423 3621
rect 4246 3544 4252 3596
rect 4304 3584 4310 3596
rect 6825 3587 6883 3593
rect 4304 3556 5672 3584
rect 4304 3544 4310 3556
rect 4157 3519 4215 3525
rect 4157 3516 4169 3519
rect 4080 3488 4169 3516
rect 4157 3485 4169 3488
rect 4203 3485 4215 3519
rect 4614 3516 4620 3528
rect 4575 3488 4620 3516
rect 4157 3479 4215 3485
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 5166 3476 5172 3528
rect 5224 3516 5230 3528
rect 5537 3519 5595 3525
rect 5537 3516 5549 3519
rect 5224 3488 5549 3516
rect 5224 3476 5230 3488
rect 5537 3485 5549 3488
rect 5583 3485 5595 3519
rect 5644 3516 5672 3556
rect 6825 3553 6837 3587
rect 6871 3584 6883 3587
rect 7098 3584 7104 3596
rect 6871 3556 7104 3584
rect 6871 3553 6883 3556
rect 6825 3547 6883 3553
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5644 3488 5733 3516
rect 5537 3479 5595 3485
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 6454 3516 6460 3528
rect 6415 3488 6460 3516
rect 5721 3479 5779 3485
rect 6454 3476 6460 3488
rect 6512 3476 6518 3528
rect 8294 3516 8300 3528
rect 8255 3488 8300 3516
rect 8294 3476 8300 3488
rect 8352 3476 8358 3528
rect 8846 3516 8852 3528
rect 8807 3488 8852 3516
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 4706 3448 4712 3460
rect 4667 3420 4712 3448
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 4893 3451 4951 3457
rect 4893 3417 4905 3451
rect 4939 3448 4951 3451
rect 5350 3448 5356 3460
rect 4939 3420 5356 3448
rect 4939 3417 4951 3420
rect 4893 3411 4951 3417
rect 5350 3408 5356 3420
rect 5408 3448 5414 3460
rect 5408 3420 5580 3448
rect 5408 3408 5414 3420
rect 5552 3392 5580 3420
rect 7098 3408 7104 3460
rect 7156 3448 7162 3460
rect 7156 3420 7222 3448
rect 7156 3408 7162 3420
rect 3513 3383 3571 3389
rect 3513 3349 3525 3383
rect 3559 3349 3571 3383
rect 3513 3343 3571 3349
rect 3878 3340 3884 3392
rect 3936 3380 3942 3392
rect 4341 3383 4399 3389
rect 4341 3380 4353 3383
rect 3936 3352 4353 3380
rect 3936 3340 3942 3352
rect 4341 3349 4353 3352
rect 4387 3349 4399 3383
rect 4341 3343 4399 3349
rect 4430 3340 4436 3392
rect 4488 3380 4494 3392
rect 4488 3352 4533 3380
rect 4488 3340 4494 3352
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 5077 3383 5135 3389
rect 5077 3380 5089 3383
rect 5040 3352 5089 3380
rect 5040 3340 5046 3352
rect 5077 3349 5089 3352
rect 5123 3349 5135 3383
rect 5077 3343 5135 3349
rect 5534 3340 5540 3392
rect 5592 3340 5598 3392
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 8757 3383 8815 3389
rect 8757 3380 8769 3383
rect 8168 3352 8769 3380
rect 8168 3340 8174 3352
rect 8757 3349 8769 3352
rect 8803 3380 8815 3383
rect 8956 3380 8984 3683
rect 8803 3352 8984 3380
rect 8803 3349 8815 3352
rect 8757 3343 8815 3349
rect 9122 3340 9128 3392
rect 9180 3380 9186 3392
rect 9309 3383 9367 3389
rect 9309 3380 9321 3383
rect 9180 3352 9321 3380
rect 9180 3340 9186 3352
rect 9309 3349 9321 3352
rect 9355 3349 9367 3383
rect 9309 3343 9367 3349
rect 3036 3290 9844 3312
rect 3036 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 5194 3290
rect 5246 3238 5258 3290
rect 5310 3238 5322 3290
rect 5374 3238 9844 3290
rect 3036 3216 9844 3238
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 5905 3179 5963 3185
rect 4856 3148 5580 3176
rect 4856 3136 4862 3148
rect 4430 3068 4436 3120
rect 4488 3068 4494 3120
rect 3418 3000 3424 3052
rect 3476 3040 3482 3052
rect 3513 3043 3571 3049
rect 3513 3040 3525 3043
rect 3476 3012 3525 3040
rect 3476 3000 3482 3012
rect 3513 3009 3525 3012
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3040 3663 3043
rect 3878 3040 3884 3052
rect 3651 3012 3884 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3040 4031 3043
rect 4062 3040 4068 3052
rect 4019 3012 4068 3040
rect 4019 3009 4031 3012
rect 3973 3003 4031 3009
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 5442 3040 5448 3052
rect 5403 3012 5448 3040
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 3329 2907 3387 2913
rect 3329 2873 3341 2907
rect 3375 2904 3387 2907
rect 3510 2904 3516 2916
rect 3375 2876 3516 2904
rect 3375 2873 3387 2876
rect 3329 2867 3387 2873
rect 3510 2864 3516 2876
rect 3568 2864 3574 2916
rect 5552 2904 5580 3148
rect 5905 3145 5917 3179
rect 5951 3145 5963 3179
rect 5905 3139 5963 3145
rect 7285 3179 7343 3185
rect 7285 3145 7297 3179
rect 7331 3176 7343 3179
rect 7331 3148 7972 3176
rect 7331 3145 7343 3148
rect 7285 3139 7343 3145
rect 5920 3108 5948 3139
rect 7944 3108 7972 3148
rect 8294 3136 8300 3188
rect 8352 3176 8358 3188
rect 9309 3179 9367 3185
rect 9309 3176 9321 3179
rect 8352 3148 9321 3176
rect 8352 3136 8358 3148
rect 9309 3145 9321 3148
rect 9355 3145 9367 3179
rect 9309 3139 9367 3145
rect 8386 3108 8392 3120
rect 5920 3080 7880 3108
rect 7944 3080 8392 3108
rect 5810 3000 5816 3052
rect 5868 3040 5874 3052
rect 6089 3043 6147 3049
rect 6089 3040 6101 3043
rect 5868 3012 6101 3040
rect 5868 3000 5874 3012
rect 6089 3009 6101 3012
rect 6135 3009 6147 3043
rect 6089 3003 6147 3009
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3040 6699 3043
rect 6730 3040 6736 3052
rect 6687 3012 6736 3040
rect 6687 3009 6699 3012
rect 6641 3003 6699 3009
rect 6730 3000 6736 3012
rect 6788 3000 6794 3052
rect 7282 3000 7288 3052
rect 7340 3040 7346 3052
rect 7852 3049 7880 3080
rect 8386 3068 8392 3080
rect 8444 3068 8450 3120
rect 8754 3108 8760 3120
rect 8715 3080 8760 3108
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 9030 3068 9036 3120
rect 9088 3108 9094 3120
rect 11146 3108 11152 3120
rect 9088 3080 11152 3108
rect 9088 3068 9094 3080
rect 11146 3068 11152 3080
rect 11204 3068 11210 3120
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 7340 3012 7481 3040
rect 7340 3000 7346 3012
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 8573 3043 8631 3049
rect 8573 3040 8585 3043
rect 8260 3012 8585 3040
rect 8260 3000 8266 3012
rect 8573 3009 8585 3012
rect 8619 3009 8631 3043
rect 9490 3040 9496 3052
rect 9451 3012 9496 3040
rect 8573 3003 8631 3009
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 8389 2975 8447 2981
rect 7668 2944 8340 2972
rect 5368 2876 5580 2904
rect 5368 2848 5396 2876
rect 5718 2864 5724 2916
rect 5776 2904 5782 2916
rect 5776 2876 6684 2904
rect 5776 2864 5782 2876
rect 5350 2796 5356 2848
rect 5408 2796 5414 2848
rect 6380 2845 6408 2876
rect 6365 2839 6423 2845
rect 6365 2805 6377 2839
rect 6411 2805 6423 2839
rect 6546 2836 6552 2848
rect 6507 2808 6552 2836
rect 6365 2799 6423 2805
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 6656 2836 6684 2876
rect 6730 2864 6736 2916
rect 6788 2904 6794 2916
rect 7006 2904 7012 2916
rect 6788 2876 7012 2904
rect 6788 2864 6794 2876
rect 7006 2864 7012 2876
rect 7064 2864 7070 2916
rect 7558 2904 7564 2916
rect 7105 2876 7564 2904
rect 7105 2836 7133 2876
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 7668 2913 7696 2944
rect 7653 2907 7711 2913
rect 7653 2873 7665 2907
rect 7699 2873 7711 2907
rect 8312 2904 8340 2944
rect 8389 2941 8401 2975
rect 8435 2972 8447 2975
rect 9030 2972 9036 2984
rect 8435 2944 9036 2972
rect 8435 2941 8447 2944
rect 8389 2935 8447 2941
rect 9030 2932 9036 2944
rect 9088 2932 9094 2984
rect 16546 2904 16574 3952
rect 8312 2876 16574 2904
rect 7653 2867 7711 2873
rect 6656 2808 7133 2836
rect 8021 2839 8079 2845
rect 8021 2805 8033 2839
rect 8067 2836 8079 2839
rect 8202 2836 8208 2848
rect 8067 2808 8208 2836
rect 8067 2805 8079 2808
rect 8021 2799 8079 2805
rect 8202 2796 8208 2808
rect 8260 2796 8266 2848
rect 8478 2796 8484 2848
rect 8536 2836 8542 2848
rect 8662 2836 8668 2848
rect 8536 2808 8668 2836
rect 8536 2796 8542 2808
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 13906 2836 13912 2848
rect 13740 2808 13912 2836
rect 3036 2746 9844 2768
rect 3036 2694 7566 2746
rect 7618 2694 7630 2746
rect 7682 2694 7694 2746
rect 7746 2694 7758 2746
rect 7810 2694 7822 2746
rect 7874 2694 9844 2746
rect 10042 2728 10048 2780
rect 10100 2768 10106 2780
rect 13630 2768 13636 2780
rect 10100 2740 13636 2768
rect 10100 2728 10106 2740
rect 13630 2728 13636 2740
rect 13688 2728 13694 2780
rect 3036 2672 9844 2694
rect 9950 2660 9956 2712
rect 10008 2700 10014 2712
rect 13740 2700 13768 2808
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 10008 2672 13768 2700
rect 10008 2660 10014 2672
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 3602 2632 3608 2644
rect 3375 2604 3608 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 3602 2592 3608 2604
rect 3660 2592 3666 2644
rect 4893 2635 4951 2641
rect 4893 2601 4905 2635
rect 4939 2632 4951 2635
rect 5442 2632 5448 2644
rect 4939 2604 5448 2632
rect 4939 2601 4951 2604
rect 4893 2595 4951 2601
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 6273 2635 6331 2641
rect 6273 2601 6285 2635
rect 6319 2632 6331 2635
rect 6454 2632 6460 2644
rect 6319 2604 6460 2632
rect 6319 2601 6331 2604
rect 6273 2595 6331 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 7653 2635 7711 2641
rect 6656 2604 7052 2632
rect 3878 2524 3884 2576
rect 3936 2564 3942 2576
rect 5718 2564 5724 2576
rect 3936 2536 5724 2564
rect 3936 2524 3942 2536
rect 5718 2524 5724 2536
rect 5776 2524 5782 2576
rect 6362 2524 6368 2576
rect 6420 2564 6426 2576
rect 6656 2564 6684 2604
rect 6420 2536 6684 2564
rect 6420 2524 6426 2536
rect 6730 2524 6736 2576
rect 6788 2564 6794 2576
rect 7024 2564 7052 2604
rect 7653 2601 7665 2635
rect 7699 2632 7711 2635
rect 13538 2632 13544 2644
rect 7699 2604 13544 2632
rect 7699 2601 7711 2604
rect 7653 2595 7711 2601
rect 13538 2592 13544 2604
rect 13596 2592 13602 2644
rect 6788 2536 6960 2564
rect 7024 2536 7512 2564
rect 6788 2524 6794 2536
rect 3970 2456 3976 2508
rect 4028 2496 4034 2508
rect 4028 2468 5304 2496
rect 4028 2456 4034 2468
rect 3513 2431 3571 2437
rect 3513 2428 3525 2431
rect 2608 2400 3525 2428
rect 14 1504 20 1556
rect 72 1544 78 1556
rect 2608 1544 2636 2400
rect 3513 2397 3525 2400
rect 3559 2397 3571 2431
rect 3786 2428 3792 2440
rect 3747 2400 3792 2428
rect 3513 2391 3571 2397
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 4157 2431 4215 2437
rect 4157 2397 4169 2431
rect 4203 2428 4215 2431
rect 4614 2428 4620 2440
rect 4203 2400 4620 2428
rect 4203 2397 4215 2400
rect 4157 2391 4215 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4982 2388 4988 2440
rect 5040 2428 5046 2440
rect 5276 2437 5304 2468
rect 5994 2456 6000 2508
rect 6052 2496 6058 2508
rect 6932 2496 6960 2536
rect 7009 2499 7067 2505
rect 7009 2496 7021 2499
rect 6052 2468 6408 2496
rect 6932 2468 7021 2496
rect 6052 2456 6058 2468
rect 6380 2437 6408 2468
rect 7009 2465 7021 2468
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 7484 2437 7512 2536
rect 8294 2524 8300 2576
rect 8352 2564 8358 2576
rect 9214 2564 9220 2576
rect 8352 2536 9220 2564
rect 8352 2524 8358 2536
rect 9214 2524 9220 2536
rect 9272 2524 9278 2576
rect 9401 2567 9459 2573
rect 9401 2533 9413 2567
rect 9447 2564 9459 2567
rect 15194 2564 15200 2576
rect 9447 2536 15200 2564
rect 9447 2533 9459 2536
rect 9401 2527 9459 2533
rect 15194 2524 15200 2536
rect 15252 2524 15258 2576
rect 7926 2496 7932 2508
rect 7887 2468 7932 2496
rect 7926 2456 7932 2468
rect 7984 2456 7990 2508
rect 5077 2431 5135 2437
rect 5077 2428 5089 2431
rect 5040 2400 5089 2428
rect 5040 2388 5046 2400
rect 5077 2397 5089 2400
rect 5123 2397 5135 2431
rect 5077 2391 5135 2397
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2428 5319 2431
rect 5721 2431 5779 2437
rect 5721 2428 5733 2431
rect 5307 2400 5733 2428
rect 5307 2397 5319 2400
rect 5261 2391 5319 2397
rect 5721 2397 5733 2400
rect 5767 2397 5779 2431
rect 6089 2431 6147 2437
rect 6089 2428 6101 2431
rect 5721 2391 5779 2397
rect 5920 2400 6101 2428
rect 3234 2320 3240 2372
rect 3292 2360 3298 2372
rect 5626 2360 5632 2372
rect 3292 2332 5632 2360
rect 3292 2320 3298 2332
rect 5626 2320 5632 2332
rect 5684 2320 5690 2372
rect 2958 2252 2964 2304
rect 3016 2292 3022 2304
rect 3605 2295 3663 2301
rect 3605 2292 3617 2295
rect 3016 2264 3617 2292
rect 3016 2252 3022 2264
rect 3605 2261 3617 2264
rect 3651 2261 3663 2295
rect 4430 2292 4436 2304
rect 4391 2264 4436 2292
rect 3605 2255 3663 2261
rect 4430 2252 4436 2264
rect 4488 2252 4494 2304
rect 5445 2295 5503 2301
rect 5445 2261 5457 2295
rect 5491 2292 5503 2295
rect 5810 2292 5816 2304
rect 5491 2264 5816 2292
rect 5491 2261 5503 2264
rect 5445 2255 5503 2261
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 5920 2301 5948 2400
rect 6089 2397 6101 2400
rect 6135 2397 6147 2431
rect 6089 2391 6147 2397
rect 6365 2431 6423 2437
rect 6365 2397 6377 2431
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 6546 2320 6552 2372
rect 6604 2360 6610 2372
rect 7300 2360 7328 2391
rect 8570 2388 8576 2440
rect 8628 2428 8634 2440
rect 9214 2428 9220 2440
rect 8628 2400 9220 2428
rect 8628 2388 8634 2400
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 6604 2332 7328 2360
rect 6604 2320 6610 2332
rect 7558 2320 7564 2372
rect 7616 2360 7622 2372
rect 9324 2360 9352 2391
rect 22094 2360 22100 2372
rect 7616 2332 9352 2360
rect 16546 2332 22100 2360
rect 7616 2320 7622 2332
rect 5905 2295 5963 2301
rect 5905 2261 5917 2295
rect 5951 2261 5963 2295
rect 5905 2255 5963 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7156 2264 7201 2292
rect 7156 2252 7162 2264
rect 3036 2202 9844 2224
rect 3036 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 5194 2202
rect 5246 2150 5258 2202
rect 5310 2150 5322 2202
rect 5374 2150 9844 2202
rect 3036 2128 9844 2150
rect 3878 2088 3884 2100
rect 3839 2060 3884 2088
rect 3878 2048 3884 2060
rect 3936 2048 3942 2100
rect 4246 2048 4252 2100
rect 4304 2088 4310 2100
rect 4985 2091 5043 2097
rect 4985 2088 4997 2091
rect 4304 2060 4997 2088
rect 4304 2048 4310 2060
rect 4985 2057 4997 2060
rect 5031 2057 5043 2091
rect 4985 2051 5043 2057
rect 6086 2048 6092 2100
rect 6144 2088 6150 2100
rect 6181 2091 6239 2097
rect 6181 2088 6193 2091
rect 6144 2060 6193 2088
rect 6144 2048 6150 2060
rect 6181 2057 6193 2060
rect 6227 2057 6239 2091
rect 6181 2051 6239 2057
rect 6638 2048 6644 2100
rect 6696 2088 6702 2100
rect 6825 2091 6883 2097
rect 6825 2088 6837 2091
rect 6696 2060 6837 2088
rect 6696 2048 6702 2060
rect 6825 2057 6837 2060
rect 6871 2057 6883 2091
rect 6825 2051 6883 2057
rect 7101 2091 7159 2097
rect 7101 2057 7113 2091
rect 7147 2088 7159 2091
rect 7190 2088 7196 2100
rect 7147 2060 7196 2088
rect 7147 2057 7159 2060
rect 7101 2051 7159 2057
rect 7190 2048 7196 2060
rect 7248 2048 7254 2100
rect 7282 2048 7288 2100
rect 7340 2088 7346 2100
rect 7377 2091 7435 2097
rect 7377 2088 7389 2091
rect 7340 2060 7389 2088
rect 7340 2048 7346 2060
rect 7377 2057 7389 2060
rect 7423 2057 7435 2091
rect 8018 2088 8024 2100
rect 7377 2051 7435 2057
rect 7484 2060 8024 2088
rect 4522 1980 4528 2032
rect 4580 2020 4586 2032
rect 6549 2023 6607 2029
rect 4580 1992 5488 2020
rect 4580 1980 4586 1992
rect 3605 1955 3663 1961
rect 3605 1921 3617 1955
rect 3651 1952 3663 1955
rect 4065 1955 4123 1961
rect 4065 1952 4077 1955
rect 3651 1924 4077 1952
rect 3651 1921 3663 1924
rect 3605 1915 3663 1921
rect 4065 1921 4077 1924
rect 4111 1952 4123 1955
rect 4798 1952 4804 1964
rect 4111 1924 4804 1952
rect 4111 1921 4123 1924
rect 4065 1915 4123 1921
rect 4798 1912 4804 1924
rect 4856 1912 4862 1964
rect 4893 1955 4951 1961
rect 4893 1921 4905 1955
rect 4939 1921 4951 1955
rect 4893 1915 4951 1921
rect 4433 1887 4491 1893
rect 4433 1853 4445 1887
rect 4479 1884 4491 1887
rect 4908 1884 4936 1915
rect 4982 1912 4988 1964
rect 5040 1952 5046 1964
rect 5460 1961 5488 1992
rect 6549 1989 6561 2023
rect 6595 2020 6607 2023
rect 7484 2020 7512 2060
rect 8018 2048 8024 2060
rect 8076 2048 8082 2100
rect 9217 2091 9275 2097
rect 9217 2057 9229 2091
rect 9263 2088 9275 2091
rect 9490 2088 9496 2100
rect 9263 2060 9496 2088
rect 9263 2057 9275 2060
rect 9217 2051 9275 2057
rect 9490 2048 9496 2060
rect 9548 2048 9554 2100
rect 8294 2020 8300 2032
rect 6595 1992 7512 2020
rect 7576 1992 8300 2020
rect 6595 1989 6607 1992
rect 6549 1983 6607 1989
rect 5169 1955 5227 1961
rect 5169 1952 5181 1955
rect 5040 1924 5181 1952
rect 5040 1912 5046 1924
rect 5169 1921 5181 1924
rect 5215 1921 5227 1955
rect 5169 1915 5227 1921
rect 5445 1955 5503 1961
rect 5445 1921 5457 1955
rect 5491 1921 5503 1955
rect 5445 1915 5503 1921
rect 5534 1912 5540 1964
rect 5592 1952 5598 1964
rect 5721 1955 5779 1961
rect 5721 1952 5733 1955
rect 5592 1924 5733 1952
rect 5592 1912 5598 1924
rect 5721 1921 5733 1924
rect 5767 1921 5779 1955
rect 5721 1915 5779 1921
rect 5810 1912 5816 1964
rect 5868 1952 5874 1964
rect 7024 1961 7052 1992
rect 7576 1961 7604 1992
rect 8294 1980 8300 1992
rect 8352 1980 8358 2032
rect 8846 1980 8852 2032
rect 8904 2020 8910 2032
rect 9033 2023 9091 2029
rect 8904 1992 8949 2020
rect 8904 1980 8910 1992
rect 9033 1989 9045 2023
rect 9079 1989 9091 2023
rect 9033 1983 9091 1989
rect 5997 1955 6055 1961
rect 5997 1952 6009 1955
rect 5868 1924 6009 1952
rect 5868 1912 5874 1924
rect 5997 1921 6009 1924
rect 6043 1921 6055 1955
rect 5997 1915 6055 1921
rect 7009 1955 7067 1961
rect 7009 1921 7021 1955
rect 7055 1921 7067 1955
rect 7009 1915 7067 1921
rect 7285 1955 7343 1961
rect 7285 1921 7297 1955
rect 7331 1921 7343 1955
rect 7285 1915 7343 1921
rect 7561 1955 7619 1961
rect 7561 1921 7573 1955
rect 7607 1921 7619 1955
rect 7561 1915 7619 1921
rect 7837 1955 7895 1961
rect 7837 1921 7849 1955
rect 7883 1952 7895 1955
rect 8110 1952 8116 1964
rect 7883 1924 8116 1952
rect 7883 1921 7895 1924
rect 7837 1915 7895 1921
rect 4479 1856 5396 1884
rect 4479 1853 4491 1856
rect 4433 1847 4491 1853
rect 4709 1819 4767 1825
rect 4709 1785 4721 1819
rect 4755 1816 4767 1819
rect 5166 1816 5172 1828
rect 4755 1788 5172 1816
rect 4755 1785 4767 1788
rect 4709 1779 4767 1785
rect 5166 1776 5172 1788
rect 5224 1776 5230 1828
rect 4890 1708 4896 1760
rect 4948 1748 4954 1760
rect 5261 1751 5319 1757
rect 5261 1748 5273 1751
rect 4948 1720 5273 1748
rect 4948 1708 4954 1720
rect 5261 1717 5273 1720
rect 5307 1717 5319 1751
rect 5368 1748 5396 1856
rect 5902 1844 5908 1896
rect 5960 1884 5966 1896
rect 7300 1884 7328 1915
rect 8110 1912 8116 1924
rect 8168 1912 8174 1964
rect 8481 1955 8539 1961
rect 8481 1921 8493 1955
rect 8527 1952 8539 1955
rect 8588 1952 8708 1956
rect 8754 1952 8760 1964
rect 8527 1928 8760 1952
rect 8527 1924 8616 1928
rect 8680 1924 8760 1928
rect 8527 1921 8539 1924
rect 8481 1915 8539 1921
rect 8754 1912 8760 1924
rect 8812 1912 8818 1964
rect 5960 1856 7328 1884
rect 5960 1844 5966 1856
rect 7374 1844 7380 1896
rect 7432 1884 7438 1896
rect 9048 1884 9076 1983
rect 9398 1912 9404 1964
rect 9456 1952 9462 1964
rect 9493 1955 9551 1961
rect 9493 1952 9505 1955
rect 9456 1924 9505 1952
rect 9456 1912 9462 1924
rect 9493 1921 9505 1924
rect 9539 1921 9551 1955
rect 9493 1915 9551 1921
rect 16546 1884 16574 2332
rect 22094 2320 22100 2332
rect 22152 2320 22158 2372
rect 7432 1856 9076 1884
rect 12406 1856 16574 1884
rect 7432 1844 7438 1856
rect 5537 1819 5595 1825
rect 5537 1785 5549 1819
rect 5583 1816 5595 1819
rect 6178 1816 6184 1828
rect 5583 1788 6184 1816
rect 5583 1785 5595 1788
rect 5537 1779 5595 1785
rect 6178 1776 6184 1788
rect 6236 1776 6242 1828
rect 6730 1776 6736 1828
rect 6788 1816 6794 1828
rect 7558 1816 7564 1828
rect 6788 1788 7564 1816
rect 6788 1776 6794 1788
rect 7558 1776 7564 1788
rect 7616 1776 7622 1828
rect 8018 1816 8024 1828
rect 7979 1788 8024 1816
rect 8018 1776 8024 1788
rect 8076 1776 8082 1828
rect 8662 1816 8668 1828
rect 8623 1788 8668 1816
rect 8662 1776 8668 1788
rect 8720 1776 8726 1828
rect 9214 1776 9220 1828
rect 9272 1816 9278 1828
rect 9309 1819 9367 1825
rect 9309 1816 9321 1819
rect 9272 1788 9321 1816
rect 9272 1776 9278 1788
rect 9309 1785 9321 1788
rect 9355 1785 9367 1819
rect 9309 1779 9367 1785
rect 12406 1748 12434 1856
rect 13814 1776 13820 1828
rect 13872 1816 13878 1828
rect 16850 1816 16856 1828
rect 13872 1788 16856 1816
rect 13872 1776 13878 1788
rect 16850 1776 16856 1788
rect 16908 1776 16914 1828
rect 5368 1720 12434 1748
rect 5261 1711 5319 1717
rect 3036 1658 9844 1680
rect 3036 1606 7566 1658
rect 7618 1606 7630 1658
rect 7682 1606 7694 1658
rect 7746 1606 7758 1658
rect 7810 1606 7822 1658
rect 7874 1606 9844 1658
rect 3036 1584 9844 1606
rect 72 1516 2636 1544
rect 72 1504 78 1516
rect 3050 1504 3056 1556
rect 3108 1544 3114 1556
rect 4433 1547 4491 1553
rect 4433 1544 4445 1547
rect 3108 1516 4445 1544
rect 3108 1504 3114 1516
rect 4433 1513 4445 1516
rect 4479 1513 4491 1547
rect 4706 1544 4712 1556
rect 4667 1516 4712 1544
rect 4433 1507 4491 1513
rect 4706 1504 4712 1516
rect 4764 1504 4770 1556
rect 5261 1547 5319 1553
rect 5261 1513 5273 1547
rect 5307 1544 5319 1547
rect 5442 1544 5448 1556
rect 5307 1516 5448 1544
rect 5307 1513 5319 1516
rect 5261 1507 5319 1513
rect 5442 1504 5448 1516
rect 5500 1504 5506 1556
rect 10502 1544 10508 1556
rect 5552 1516 10508 1544
rect 3142 1436 3148 1488
rect 3200 1476 3206 1488
rect 4154 1476 4160 1488
rect 3200 1448 4016 1476
rect 4115 1448 4160 1476
rect 3200 1436 3206 1448
rect 750 1368 756 1420
rect 808 1408 814 1420
rect 3988 1408 4016 1448
rect 4154 1436 4160 1448
rect 4212 1436 4218 1488
rect 4798 1436 4804 1488
rect 4856 1476 4862 1488
rect 5552 1476 5580 1516
rect 10502 1504 10508 1516
rect 10560 1504 10566 1556
rect 4856 1448 5580 1476
rect 4856 1436 4862 1448
rect 5718 1436 5724 1488
rect 5776 1476 5782 1488
rect 8754 1476 8760 1488
rect 5776 1448 8760 1476
rect 5776 1436 5782 1448
rect 8754 1436 8760 1448
rect 8812 1436 8818 1488
rect 8938 1476 8944 1488
rect 8899 1448 8944 1476
rect 8938 1436 8944 1448
rect 8996 1436 9002 1488
rect 9401 1479 9459 1485
rect 9048 1448 9260 1476
rect 7561 1411 7619 1417
rect 808 1380 3924 1408
rect 3988 1380 4936 1408
rect 808 1368 814 1380
rect 3326 1300 3332 1352
rect 3384 1340 3390 1352
rect 3513 1343 3571 1349
rect 3513 1340 3525 1343
rect 3384 1312 3525 1340
rect 3384 1300 3390 1312
rect 3513 1309 3525 1312
rect 3559 1309 3571 1343
rect 3513 1303 3571 1309
rect 3694 1300 3700 1352
rect 3752 1340 3758 1352
rect 3789 1343 3847 1349
rect 3789 1340 3801 1343
rect 3752 1312 3801 1340
rect 3752 1300 3758 1312
rect 3789 1309 3801 1312
rect 3835 1309 3847 1343
rect 3896 1340 3924 1380
rect 4065 1343 4123 1349
rect 4065 1340 4077 1343
rect 3896 1312 4077 1340
rect 3789 1303 3847 1309
rect 4065 1309 4077 1312
rect 4111 1309 4123 1343
rect 4065 1303 4123 1309
rect 4341 1343 4399 1349
rect 4341 1309 4353 1343
rect 4387 1309 4399 1343
rect 4614 1340 4620 1352
rect 4575 1312 4620 1340
rect 4341 1303 4399 1309
rect 4356 1272 4384 1303
rect 4614 1300 4620 1312
rect 4672 1300 4678 1352
rect 4908 1349 4936 1380
rect 6564 1380 6868 1408
rect 4893 1343 4951 1349
rect 4893 1309 4905 1343
rect 4939 1309 4951 1343
rect 4893 1303 4951 1309
rect 5169 1343 5227 1349
rect 5169 1309 5181 1343
rect 5215 1340 5227 1343
rect 5350 1340 5356 1352
rect 5215 1312 5356 1340
rect 5215 1309 5227 1312
rect 5169 1303 5227 1309
rect 5350 1300 5356 1312
rect 5408 1300 5414 1352
rect 5445 1343 5503 1349
rect 5445 1309 5457 1343
rect 5491 1309 5503 1343
rect 5445 1303 5503 1309
rect 2746 1244 4384 1272
rect 2590 892 2596 944
rect 2648 932 2654 944
rect 2746 932 2774 1244
rect 4522 1232 4528 1284
rect 4580 1272 4586 1284
rect 5460 1272 5488 1303
rect 5626 1300 5632 1352
rect 5684 1340 5690 1352
rect 5905 1343 5963 1349
rect 5905 1340 5917 1343
rect 5684 1312 5917 1340
rect 5684 1300 5690 1312
rect 5905 1309 5917 1312
rect 5951 1309 5963 1343
rect 5905 1303 5963 1309
rect 6181 1343 6239 1349
rect 6181 1309 6193 1343
rect 6227 1340 6239 1343
rect 6564 1340 6592 1380
rect 6227 1312 6592 1340
rect 6227 1309 6239 1312
rect 6181 1303 6239 1309
rect 6638 1300 6644 1352
rect 6696 1340 6702 1352
rect 6840 1340 6868 1380
rect 7561 1377 7573 1411
rect 7607 1408 7619 1411
rect 7607 1380 8616 1408
rect 7607 1377 7619 1380
rect 7561 1371 7619 1377
rect 8294 1340 8300 1352
rect 6696 1312 6741 1340
rect 6840 1312 8300 1340
rect 6696 1300 6702 1312
rect 8294 1300 8300 1312
rect 8352 1300 8358 1352
rect 8588 1349 8616 1380
rect 8662 1368 8668 1420
rect 8720 1408 8726 1420
rect 9048 1408 9076 1448
rect 8720 1380 8900 1408
rect 8720 1368 8726 1380
rect 8573 1343 8631 1349
rect 8573 1309 8585 1343
rect 8619 1340 8631 1343
rect 8754 1340 8760 1352
rect 8619 1312 8760 1340
rect 8619 1309 8631 1312
rect 8573 1303 8631 1309
rect 8754 1300 8760 1312
rect 8812 1300 8818 1352
rect 8872 1349 8900 1380
rect 8956 1380 9076 1408
rect 8956 1352 8984 1380
rect 8849 1343 8907 1349
rect 8849 1309 8861 1343
rect 8895 1309 8907 1343
rect 8849 1303 8907 1309
rect 8938 1300 8944 1352
rect 8996 1300 9002 1352
rect 9122 1340 9128 1352
rect 9083 1312 9128 1340
rect 9122 1300 9128 1312
rect 9180 1300 9186 1352
rect 9232 1340 9260 1448
rect 9401 1445 9413 1479
rect 9447 1476 9459 1479
rect 9447 1448 16574 1476
rect 9447 1445 9459 1448
rect 9401 1439 9459 1445
rect 16546 1408 16574 1448
rect 16666 1408 16672 1420
rect 16546 1380 16672 1408
rect 16666 1368 16672 1380
rect 16724 1368 16730 1420
rect 9232 1312 16574 1340
rect 9950 1272 9956 1284
rect 4580 1244 5488 1272
rect 6012 1244 8800 1272
rect 4580 1232 4586 1244
rect 2866 1164 2872 1216
rect 2924 1204 2930 1216
rect 3329 1207 3387 1213
rect 3329 1204 3341 1207
rect 2924 1176 3341 1204
rect 2924 1164 2930 1176
rect 3329 1173 3341 1176
rect 3375 1173 3387 1207
rect 3602 1204 3608 1216
rect 3563 1176 3608 1204
rect 3329 1167 3387 1173
rect 3602 1164 3608 1176
rect 3660 1164 3666 1216
rect 3878 1204 3884 1216
rect 3839 1176 3884 1204
rect 3878 1164 3884 1176
rect 3936 1164 3942 1216
rect 4982 1204 4988 1216
rect 4943 1176 4988 1204
rect 4982 1164 4988 1176
rect 5040 1164 5046 1216
rect 5534 1164 5540 1216
rect 5592 1204 5598 1216
rect 6012 1213 6040 1244
rect 5721 1207 5779 1213
rect 5721 1204 5733 1207
rect 5592 1176 5733 1204
rect 5592 1164 5598 1176
rect 5721 1173 5733 1176
rect 5767 1173 5779 1207
rect 5721 1167 5779 1173
rect 5997 1207 6055 1213
rect 5997 1173 6009 1207
rect 6043 1173 6055 1207
rect 6730 1204 6736 1216
rect 6691 1176 6736 1204
rect 5997 1167 6055 1173
rect 6730 1164 6736 1176
rect 6788 1164 6794 1216
rect 7190 1204 7196 1216
rect 7151 1176 7196 1204
rect 7190 1164 7196 1176
rect 7248 1164 7254 1216
rect 7926 1204 7932 1216
rect 7887 1176 7932 1204
rect 7926 1164 7932 1176
rect 7984 1164 7990 1216
rect 8386 1204 8392 1216
rect 8347 1176 8392 1204
rect 8386 1164 8392 1176
rect 8444 1164 8450 1216
rect 8478 1164 8484 1216
rect 8536 1204 8542 1216
rect 8665 1207 8723 1213
rect 8665 1204 8677 1207
rect 8536 1176 8677 1204
rect 8536 1164 8542 1176
rect 8665 1173 8677 1176
rect 8711 1173 8723 1207
rect 8772 1204 8800 1244
rect 8956 1244 9956 1272
rect 8956 1204 8984 1244
rect 9950 1232 9956 1244
rect 10008 1232 10014 1284
rect 16546 1272 16574 1312
rect 16758 1272 16764 1284
rect 16546 1244 16764 1272
rect 16758 1232 16764 1244
rect 16816 1232 16822 1284
rect 8772 1176 8984 1204
rect 8665 1167 8723 1173
rect 9030 1164 9036 1216
rect 9088 1204 9094 1216
rect 9214 1204 9220 1216
rect 9088 1176 9220 1204
rect 9088 1164 9094 1176
rect 9214 1164 9220 1176
rect 9272 1164 9278 1216
rect 3036 1114 9844 1136
rect 3036 1062 5066 1114
rect 5118 1062 5130 1114
rect 5182 1062 5194 1114
rect 5246 1062 5258 1114
rect 5310 1062 5322 1114
rect 5374 1062 9844 1114
rect 3036 1040 9844 1062
rect 7190 960 7196 1012
rect 7248 1000 7254 1012
rect 9030 1000 9036 1012
rect 7248 972 9036 1000
rect 7248 960 7254 972
rect 9030 960 9036 972
rect 9088 960 9094 1012
rect 2648 904 2774 932
rect 2648 892 2654 904
rect 7926 892 7932 944
rect 7984 932 7990 944
rect 8662 932 8668 944
rect 7984 904 8668 932
rect 7984 892 7990 904
rect 8662 892 8668 904
rect 8720 932 8726 944
rect 16574 932 16580 944
rect 8720 904 16580 932
rect 8720 892 8726 904
rect 16574 892 16580 904
rect 16632 892 16638 944
rect 2314 824 2320 876
rect 2372 864 2378 876
rect 4614 864 4620 876
rect 2372 836 4620 864
rect 2372 824 2378 836
rect 4614 824 4620 836
rect 4672 824 4678 876
rect 8294 824 8300 876
rect 8352 864 8358 876
rect 9306 864 9312 876
rect 8352 836 9312 864
rect 8352 824 8358 836
rect 9306 824 9312 836
rect 9364 824 9370 876
rect 2406 756 2412 808
rect 2464 796 2470 808
rect 4522 796 4528 808
rect 2464 768 4528 796
rect 2464 756 2470 768
rect 4522 756 4528 768
rect 4580 756 4586 808
rect 3878 688 3884 740
rect 3936 728 3942 740
rect 5718 728 5724 740
rect 3936 700 5724 728
rect 3936 688 3942 700
rect 5718 688 5724 700
rect 5776 688 5782 740
<< via1 >>
rect 2136 11840 2188 11892
rect 7012 11840 7064 11892
rect 13820 11840 13872 11892
rect 16672 11840 16724 11892
rect 2780 11772 2832 11824
rect 3792 11772 3844 11824
rect 3976 11772 4028 11824
rect 5540 11772 5592 11824
rect 2964 11704 3016 11756
rect 8668 11704 8720 11756
rect 1492 11636 1544 11688
rect 5448 11636 5500 11688
rect 1308 11568 1360 11620
rect 5540 11568 5592 11620
rect 5908 11568 5960 11620
rect 6460 11568 6512 11620
rect 3148 11500 3200 11552
rect 6368 11500 6420 11552
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 7566 11398 7618 11450
rect 7630 11398 7682 11450
rect 7694 11398 7746 11450
rect 7758 11398 7810 11450
rect 7822 11398 7874 11450
rect 1308 11339 1360 11348
rect 1308 11305 1317 11339
rect 1317 11305 1351 11339
rect 1351 11305 1360 11339
rect 1308 11296 1360 11305
rect 4528 11296 4580 11348
rect 8392 11296 8444 11348
rect 9312 11296 9364 11348
rect 10876 11296 10928 11348
rect 2136 11271 2188 11280
rect 2136 11237 2145 11271
rect 2145 11237 2179 11271
rect 2179 11237 2188 11271
rect 2136 11228 2188 11237
rect 2964 11271 3016 11280
rect 2964 11237 2973 11271
rect 2973 11237 3007 11271
rect 3007 11237 3016 11271
rect 2964 11228 3016 11237
rect 3148 11228 3200 11280
rect 3332 11228 3384 11280
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 1860 11135 1912 11144
rect 1860 11101 1869 11135
rect 1869 11101 1903 11135
rect 1903 11101 1912 11135
rect 1860 11092 1912 11101
rect 2228 11092 2280 11144
rect 4344 11160 4396 11212
rect 4896 11160 4948 11212
rect 7472 11228 7524 11280
rect 9588 11228 9640 11280
rect 6736 11160 6788 11212
rect 3332 11092 3384 11144
rect 3608 11092 3660 11144
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 4344 11024 4396 11076
rect 6460 11092 6512 11144
rect 6552 11135 6604 11144
rect 6552 11101 6561 11135
rect 6561 11101 6595 11135
rect 6595 11101 6604 11135
rect 6552 11092 6604 11101
rect 6184 11024 6236 11076
rect 20 10956 72 11008
rect 940 10956 992 11008
rect 2412 10956 2464 11008
rect 2596 10999 2648 11008
rect 2596 10965 2605 10999
rect 2605 10965 2639 10999
rect 2639 10965 2648 10999
rect 2596 10956 2648 10965
rect 2688 10956 2740 11008
rect 4988 10956 5040 11008
rect 5724 10956 5776 11008
rect 6552 10956 6604 11008
rect 7104 11024 7156 11076
rect 7380 11092 7432 11144
rect 7840 11092 7892 11144
rect 8024 11092 8076 11144
rect 8300 11135 8352 11144
rect 8300 11101 8309 11135
rect 8309 11101 8343 11135
rect 8343 11101 8352 11135
rect 8300 11092 8352 11101
rect 8484 11024 8536 11076
rect 11152 11160 11204 11212
rect 9128 11092 9180 11144
rect 8760 11024 8812 11076
rect 9312 11092 9364 11144
rect 10416 11092 10468 11144
rect 10692 11024 10744 11076
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 5194 10854 5246 10906
rect 5258 10854 5310 10906
rect 5322 10854 5374 10906
rect 6092 10752 6144 10804
rect 2780 10683 2832 10692
rect 940 10616 992 10668
rect 1952 10616 2004 10668
rect 2780 10649 2789 10683
rect 2789 10649 2823 10683
rect 2823 10649 2832 10683
rect 2780 10640 2832 10649
rect 3884 10684 3936 10736
rect 5080 10684 5132 10736
rect 1676 10548 1728 10600
rect 4712 10616 4764 10668
rect 4896 10659 4948 10668
rect 4896 10625 4905 10659
rect 4905 10625 4939 10659
rect 4939 10625 4948 10659
rect 4896 10616 4948 10625
rect 5172 10616 5224 10668
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 6552 10616 6604 10668
rect 7288 10616 7340 10668
rect 9036 10616 9088 10668
rect 1584 10480 1636 10532
rect 2688 10548 2740 10600
rect 3516 10548 3568 10600
rect 5448 10591 5500 10600
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 5816 10548 5868 10600
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 4344 10480 4396 10532
rect 6276 10480 6328 10532
rect 8116 10480 8168 10532
rect 16580 10616 16632 10668
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 2964 10412 3016 10464
rect 3148 10455 3200 10464
rect 3148 10421 3178 10455
rect 3178 10421 3200 10455
rect 3148 10412 3200 10421
rect 4896 10412 4948 10464
rect 6000 10412 6052 10464
rect 6552 10412 6604 10464
rect 8944 10412 8996 10464
rect 9220 10412 9272 10464
rect 9312 10412 9364 10464
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 7566 10310 7618 10362
rect 7630 10310 7682 10362
rect 7694 10310 7746 10362
rect 7758 10310 7810 10362
rect 7822 10310 7874 10362
rect 2044 10208 2096 10260
rect 3148 10140 3200 10192
rect 3424 10183 3476 10192
rect 3424 10149 3433 10183
rect 3433 10149 3467 10183
rect 3467 10149 3476 10183
rect 3424 10140 3476 10149
rect 1676 10115 1728 10124
rect 1676 10081 1685 10115
rect 1685 10081 1719 10115
rect 1719 10081 1728 10115
rect 1676 10072 1728 10081
rect 1952 10072 2004 10124
rect 4344 10072 4396 10124
rect 4528 10115 4580 10124
rect 4528 10081 4537 10115
rect 4537 10081 4571 10115
rect 4571 10081 4580 10115
rect 4528 10072 4580 10081
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 1584 10004 1636 10056
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 3608 10004 3660 10013
rect 1492 9868 1544 9920
rect 2228 9936 2280 9988
rect 3332 9936 3384 9988
rect 4068 10004 4120 10056
rect 5264 10072 5316 10124
rect 5908 10004 5960 10056
rect 6552 10208 6604 10260
rect 7196 10208 7248 10260
rect 6736 10140 6788 10192
rect 11060 10140 11112 10192
rect 3884 9936 3936 9988
rect 2964 9868 3016 9920
rect 4160 9868 4212 9920
rect 5540 9936 5592 9988
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 7656 10004 7708 10056
rect 7196 9936 7248 9988
rect 7840 9868 7892 9920
rect 8852 10047 8904 10056
rect 8852 10013 8861 10047
rect 8861 10013 8895 10047
rect 8895 10013 8904 10047
rect 8852 10004 8904 10013
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 5194 9766 5246 9818
rect 5258 9766 5310 9818
rect 5322 9766 5374 9818
rect 1676 9664 1728 9716
rect 2228 9664 2280 9716
rect 8852 9664 8904 9716
rect 2780 9596 2832 9648
rect 3792 9596 3844 9648
rect 5448 9596 5500 9648
rect 5724 9596 5776 9648
rect 6552 9596 6604 9648
rect 8484 9596 8536 9648
rect 1584 9460 1636 9512
rect 3516 9528 3568 9580
rect 4896 9571 4948 9580
rect 4896 9537 4905 9571
rect 4905 9537 4939 9571
rect 4939 9537 4948 9571
rect 4896 9528 4948 9537
rect 5356 9528 5408 9580
rect 6184 9571 6236 9580
rect 6184 9537 6193 9571
rect 6193 9537 6227 9571
rect 6227 9537 6236 9571
rect 6184 9528 6236 9537
rect 6920 9528 6972 9580
rect 7380 9528 7432 9580
rect 7748 9571 7800 9580
rect 3056 9503 3108 9512
rect 3056 9469 3065 9503
rect 3065 9469 3099 9503
rect 3099 9469 3108 9503
rect 3056 9460 3108 9469
rect 4068 9460 4120 9512
rect 5632 9460 5684 9512
rect 5724 9460 5776 9512
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 2780 9392 2832 9444
rect 2044 9324 2096 9376
rect 3148 9324 3200 9376
rect 5724 9324 5776 9376
rect 5908 9324 5960 9376
rect 6184 9324 6236 9376
rect 7196 9324 7248 9376
rect 8484 9324 8536 9376
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 7566 9222 7618 9274
rect 7630 9222 7682 9274
rect 7694 9222 7746 9274
rect 7758 9222 7810 9274
rect 7822 9222 7874 9274
rect 1400 9120 1452 9172
rect 3056 9163 3108 9172
rect 1584 9052 1636 9104
rect 1584 8916 1636 8968
rect 2688 9052 2740 9104
rect 3056 9129 3065 9163
rect 3065 9129 3099 9163
rect 3099 9129 3108 9163
rect 3056 9120 3108 9129
rect 3608 9120 3660 9172
rect 4528 9120 4580 9172
rect 5080 9120 5132 9172
rect 5540 9120 5592 9172
rect 2412 8984 2464 9036
rect 2044 8916 2096 8968
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 848 8848 900 8900
rect 3884 9052 3936 9104
rect 4804 9052 4856 9104
rect 4160 8984 4212 9036
rect 4252 8984 4304 9036
rect 3240 8959 3292 8968
rect 1216 8823 1268 8832
rect 1216 8789 1225 8823
rect 1225 8789 1259 8823
rect 1259 8789 1268 8823
rect 1216 8780 1268 8789
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 3424 8916 3476 8968
rect 4068 8916 4120 8968
rect 4436 8916 4488 8968
rect 5080 8916 5132 8968
rect 6276 8959 6328 8968
rect 1952 8780 2004 8832
rect 2136 8780 2188 8832
rect 3792 8780 3844 8832
rect 5632 8848 5684 8900
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 8300 9120 8352 9172
rect 8208 8984 8260 9036
rect 8576 8984 8628 9036
rect 8024 8916 8076 8968
rect 8852 8959 8904 8968
rect 8852 8925 8861 8959
rect 8861 8925 8895 8959
rect 8895 8925 8904 8959
rect 8852 8916 8904 8925
rect 7012 8848 7064 8900
rect 7196 8780 7248 8832
rect 9588 8780 9640 8832
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 5194 8678 5246 8730
rect 5258 8678 5310 8730
rect 5322 8678 5374 8730
rect 1400 8576 1452 8628
rect 1768 8576 1820 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2320 8440 2372 8492
rect 1768 8372 1820 8424
rect 2780 8576 2832 8628
rect 5540 8576 5592 8628
rect 6736 8576 6788 8628
rect 7012 8576 7064 8628
rect 7196 8576 7248 8628
rect 8576 8576 8628 8628
rect 9128 8619 9180 8628
rect 9128 8585 9137 8619
rect 9137 8585 9171 8619
rect 9171 8585 9180 8619
rect 9128 8576 9180 8585
rect 3976 8508 4028 8560
rect 4712 8508 4764 8560
rect 4988 8508 5040 8560
rect 2596 8372 2648 8424
rect 2412 8304 2464 8356
rect 2780 8440 2832 8492
rect 3608 8440 3660 8492
rect 4436 8483 4488 8492
rect 4436 8449 4445 8483
rect 4445 8449 4479 8483
rect 4479 8449 4488 8483
rect 4436 8440 4488 8449
rect 5632 8440 5684 8492
rect 5908 8508 5960 8560
rect 7564 8508 7616 8560
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 8944 8440 8996 8492
rect 2872 8372 2924 8424
rect 5908 8372 5960 8424
rect 3332 8304 3384 8356
rect 3792 8304 3844 8356
rect 4160 8347 4212 8356
rect 4160 8313 4169 8347
rect 4169 8313 4203 8347
rect 4203 8313 4212 8347
rect 4160 8304 4212 8313
rect 4712 8304 4764 8356
rect 6092 8304 6144 8356
rect 10968 8304 11020 8356
rect 1584 8279 1636 8288
rect 1584 8245 1593 8279
rect 1593 8245 1627 8279
rect 1627 8245 1636 8279
rect 1584 8236 1636 8245
rect 1952 8236 2004 8288
rect 4252 8236 4304 8288
rect 4528 8236 4580 8288
rect 5448 8236 5500 8288
rect 5540 8236 5592 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 7566 8134 7618 8186
rect 7630 8134 7682 8186
rect 7694 8134 7746 8186
rect 7758 8134 7810 8186
rect 7822 8134 7874 8186
rect 1400 8032 1452 8084
rect 1860 8032 1912 8084
rect 2964 8032 3016 8084
rect 4252 8032 4304 8084
rect 4436 8032 4488 8084
rect 4804 8032 4856 8084
rect 6460 8032 6512 8084
rect 8576 8075 8628 8084
rect 8576 8041 8585 8075
rect 8585 8041 8619 8075
rect 8619 8041 8628 8075
rect 8576 8032 8628 8041
rect 8760 8075 8812 8084
rect 8760 8041 8769 8075
rect 8769 8041 8803 8075
rect 8803 8041 8812 8075
rect 8760 8032 8812 8041
rect 2228 7964 2280 8016
rect 1768 7896 1820 7948
rect 3792 7964 3844 8016
rect 7012 7964 7064 8016
rect 7196 7964 7248 8016
rect 7932 7964 7984 8016
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 9220 7896 9272 7948
rect 3056 7828 3108 7880
rect 2412 7760 2464 7812
rect 1676 7692 1728 7744
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 7288 7828 7340 7880
rect 6000 7760 6052 7812
rect 4252 7692 4304 7744
rect 4436 7692 4488 7744
rect 7748 7760 7800 7812
rect 8208 7828 8260 7880
rect 8484 7760 8536 7812
rect 9404 7760 9456 7812
rect 6552 7692 6604 7744
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 5194 7590 5246 7642
rect 5258 7590 5310 7642
rect 5322 7590 5374 7642
rect 1124 7488 1176 7540
rect 5816 7488 5868 7540
rect 6276 7488 6328 7540
rect 6828 7488 6880 7540
rect 1032 7420 1084 7472
rect 1860 7420 1912 7472
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1768 7395 1820 7404
rect 1492 7352 1544 7361
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 1952 7352 2004 7404
rect 2412 7352 2464 7404
rect 3516 7420 3568 7472
rect 4804 7420 4856 7472
rect 8300 7420 8352 7472
rect 1584 7284 1636 7336
rect 2044 7216 2096 7268
rect 2228 7148 2280 7200
rect 2412 7148 2464 7200
rect 3884 7352 3936 7404
rect 2964 7327 3016 7336
rect 2964 7293 2973 7327
rect 2973 7293 3007 7327
rect 3007 7293 3016 7327
rect 2964 7284 3016 7293
rect 4528 7216 4580 7268
rect 4804 7216 4856 7268
rect 5448 7352 5500 7404
rect 6184 7352 6236 7404
rect 7840 7352 7892 7404
rect 5540 7216 5592 7268
rect 6000 7216 6052 7268
rect 7932 7284 7984 7336
rect 9128 7327 9180 7336
rect 9128 7293 9137 7327
rect 9137 7293 9171 7327
rect 9171 7293 9180 7327
rect 9128 7284 9180 7293
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 2964 7148 3016 7200
rect 3608 7148 3660 7200
rect 4436 7148 4488 7200
rect 6736 7148 6788 7200
rect 8576 7148 8628 7200
rect 8668 7191 8720 7200
rect 8668 7157 8677 7191
rect 8677 7157 8711 7191
rect 8711 7157 8720 7191
rect 8668 7148 8720 7157
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 7566 7046 7618 7098
rect 7630 7046 7682 7098
rect 7694 7046 7746 7098
rect 7758 7046 7810 7098
rect 7822 7046 7874 7098
rect 940 6944 992 6996
rect 2412 6944 2464 6996
rect 6828 6944 6880 6996
rect 7380 6944 7432 6996
rect 9128 6944 9180 6996
rect 11152 6944 11204 6996
rect 16672 6944 16724 6996
rect 1952 6808 2004 6860
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 3700 6808 3752 6860
rect 4620 6808 4672 6860
rect 1584 6672 1636 6724
rect 2044 6604 2096 6656
rect 2872 6604 2924 6656
rect 3240 6604 3292 6656
rect 3516 6740 3568 6792
rect 4160 6740 4212 6792
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 4988 6740 5040 6792
rect 6460 6808 6512 6860
rect 7012 6740 7064 6792
rect 7104 6740 7156 6792
rect 8208 6808 8260 6860
rect 9036 6808 9088 6860
rect 7932 6783 7984 6792
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 3516 6604 3568 6656
rect 4988 6604 5040 6656
rect 5632 6604 5684 6656
rect 5816 6604 5868 6656
rect 6552 6604 6604 6656
rect 7288 6604 7340 6656
rect 8392 6672 8444 6724
rect 8576 6672 8628 6724
rect 8852 6672 8904 6724
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 5194 6502 5246 6554
rect 5258 6502 5310 6554
rect 5322 6502 5374 6554
rect 1584 6400 1636 6452
rect 1768 6400 1820 6452
rect 2228 6400 2280 6452
rect 6552 6400 6604 6452
rect 3424 6332 3476 6384
rect 8024 6400 8076 6452
rect 1492 6264 1544 6316
rect 1584 6264 1636 6316
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 2136 6128 2188 6180
rect 2412 6196 2464 6248
rect 2504 6171 2556 6180
rect 2504 6137 2513 6171
rect 2513 6137 2547 6171
rect 2547 6137 2556 6171
rect 2504 6128 2556 6137
rect 2596 6128 2648 6180
rect 2228 6103 2280 6112
rect 2228 6069 2237 6103
rect 2237 6069 2271 6103
rect 2271 6069 2280 6103
rect 2228 6060 2280 6069
rect 2412 6060 2464 6112
rect 3976 6264 4028 6316
rect 3516 6196 3568 6248
rect 7472 6332 7524 6384
rect 5724 6264 5776 6316
rect 6092 6264 6144 6316
rect 6552 6264 6604 6316
rect 8024 6264 8076 6316
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 5172 6239 5224 6248
rect 5172 6205 5181 6239
rect 5181 6205 5215 6239
rect 5215 6205 5224 6239
rect 5172 6196 5224 6205
rect 5632 6196 5684 6248
rect 6276 6196 6328 6248
rect 7472 6196 7524 6248
rect 9036 6264 9088 6316
rect 5540 6060 5592 6112
rect 8668 6128 8720 6180
rect 8760 6103 8812 6112
rect 8760 6069 8769 6103
rect 8769 6069 8803 6103
rect 8803 6069 8812 6103
rect 8760 6060 8812 6069
rect 9220 6060 9272 6112
rect 9496 6103 9548 6112
rect 9496 6069 9505 6103
rect 9505 6069 9539 6103
rect 9539 6069 9548 6103
rect 9496 6060 9548 6069
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 7566 5958 7618 6010
rect 7630 5958 7682 6010
rect 7694 5958 7746 6010
rect 7758 5958 7810 6010
rect 7822 5958 7874 6010
rect 1492 5856 1544 5908
rect 1676 5763 1728 5772
rect 1676 5729 1685 5763
rect 1685 5729 1719 5763
rect 1719 5729 1728 5763
rect 1676 5720 1728 5729
rect 3332 5720 3384 5772
rect 4252 5720 4304 5772
rect 5540 5899 5592 5908
rect 5540 5865 5549 5899
rect 5549 5865 5583 5899
rect 5583 5865 5592 5899
rect 5540 5856 5592 5865
rect 6092 5856 6144 5908
rect 9496 5856 9548 5908
rect 6460 5788 6512 5840
rect 8852 5788 8904 5840
rect 6092 5720 6144 5772
rect 6184 5720 6236 5772
rect 7932 5720 7984 5772
rect 8944 5720 8996 5772
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 1768 5516 1820 5568
rect 3240 5516 3292 5568
rect 3608 5516 3660 5568
rect 3700 5516 3752 5568
rect 4160 5584 4212 5636
rect 5172 5584 5224 5636
rect 3976 5516 4028 5568
rect 4620 5516 4672 5568
rect 5540 5652 5592 5704
rect 8760 5652 8812 5704
rect 6092 5584 6144 5636
rect 6368 5627 6420 5636
rect 6368 5593 6377 5627
rect 6377 5593 6411 5627
rect 6411 5593 6420 5627
rect 6368 5584 6420 5593
rect 8208 5584 8260 5636
rect 8668 5584 8720 5636
rect 9036 5584 9088 5636
rect 5632 5516 5684 5568
rect 8484 5516 8536 5568
rect 8576 5516 8628 5568
rect 9128 5516 9180 5568
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 5194 5414 5246 5466
rect 5258 5414 5310 5466
rect 5322 5414 5374 5466
rect 1400 5312 1452 5364
rect 2412 5312 2464 5364
rect 3700 5312 3752 5364
rect 3884 5312 3936 5364
rect 1952 5176 2004 5228
rect 2596 5176 2648 5228
rect 2872 5176 2924 5228
rect 6092 5312 6144 5364
rect 7472 5312 7524 5364
rect 4804 5244 4856 5296
rect 7932 5244 7984 5296
rect 8208 5244 8260 5296
rect 5816 5219 5868 5228
rect 5816 5185 5825 5219
rect 5825 5185 5859 5219
rect 5859 5185 5868 5219
rect 5816 5176 5868 5185
rect 6184 5176 6236 5228
rect 8392 5176 8444 5228
rect 9220 5219 9272 5228
rect 9220 5185 9229 5219
rect 9229 5185 9263 5219
rect 9263 5185 9272 5219
rect 9220 5176 9272 5185
rect 2228 5108 2280 5160
rect 3976 5151 4028 5160
rect 3976 5117 3985 5151
rect 3985 5117 4019 5151
rect 4019 5117 4028 5151
rect 3976 5108 4028 5117
rect 3516 5015 3568 5024
rect 3516 4981 3525 5015
rect 3525 4981 3559 5015
rect 3559 4981 3568 5015
rect 3516 4972 3568 4981
rect 3884 5015 3936 5024
rect 3884 4981 3893 5015
rect 3893 4981 3927 5015
rect 3927 4981 3936 5015
rect 3884 4972 3936 4981
rect 6736 5108 6788 5160
rect 8484 5108 8536 5160
rect 6092 5040 6144 5092
rect 5724 4972 5776 5024
rect 6368 4972 6420 5024
rect 16672 4972 16724 5024
rect 7566 4870 7618 4922
rect 7630 4870 7682 4922
rect 7694 4870 7746 4922
rect 7758 4870 7810 4922
rect 7822 4870 7874 4922
rect 4160 4768 4212 4820
rect 4988 4768 5040 4820
rect 5356 4768 5408 4820
rect 8300 4768 8352 4820
rect 15200 4768 15252 4820
rect 20628 4768 20680 4820
rect 3332 4675 3384 4684
rect 3332 4641 3341 4675
rect 3341 4641 3375 4675
rect 3375 4641 3384 4675
rect 3332 4632 3384 4641
rect 3608 4675 3660 4684
rect 3608 4641 3617 4675
rect 3617 4641 3651 4675
rect 3651 4641 3660 4675
rect 3608 4632 3660 4641
rect 4160 4632 4212 4684
rect 4804 4632 4856 4684
rect 5632 4632 5684 4684
rect 6184 4632 6236 4684
rect 6644 4632 6696 4684
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 3424 4428 3476 4480
rect 5908 4428 5960 4480
rect 6184 4496 6236 4548
rect 7656 4496 7708 4548
rect 8576 4496 8628 4548
rect 9588 4496 9640 4548
rect 8208 4428 8260 4480
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 5194 4326 5246 4378
rect 5258 4326 5310 4378
rect 5322 4326 5374 4378
rect 4160 4224 4212 4276
rect 4988 4224 5040 4276
rect 3608 4088 3660 4140
rect 4712 4088 4764 4140
rect 5632 4224 5684 4276
rect 6184 4224 6236 4276
rect 6828 4224 6880 4276
rect 7104 4224 7156 4276
rect 7472 4156 7524 4208
rect 5724 4131 5776 4140
rect 3884 4020 3936 4072
rect 5724 4097 5733 4131
rect 5733 4097 5767 4131
rect 5767 4097 5776 4131
rect 5724 4088 5776 4097
rect 7196 4088 7248 4140
rect 8208 4088 8260 4140
rect 8760 4088 8812 4140
rect 6092 4020 6144 4072
rect 6828 4020 6880 4072
rect 7932 4020 7984 4072
rect 3516 3952 3568 4004
rect 4068 3884 4120 3936
rect 4620 3952 4672 4004
rect 5172 3952 5224 4004
rect 5540 3952 5592 4004
rect 7104 3952 7156 4004
rect 5724 3884 5776 3936
rect 6460 3884 6512 3936
rect 6828 3884 6880 3936
rect 8852 3884 8904 3936
rect 16580 3952 16632 4004
rect 9220 3884 9272 3936
rect 7566 3782 7618 3834
rect 7630 3782 7682 3834
rect 7694 3782 7746 3834
rect 7758 3782 7810 3834
rect 7822 3782 7874 3834
rect 4528 3680 4580 3732
rect 5816 3680 5868 3732
rect 6184 3680 6236 3732
rect 8760 3680 8812 3732
rect 2964 3476 3016 3528
rect 3976 3476 4028 3528
rect 4896 3612 4948 3664
rect 4252 3544 4304 3596
rect 4620 3519 4672 3528
rect 4620 3485 4629 3519
rect 4629 3485 4663 3519
rect 4663 3485 4672 3519
rect 4620 3476 4672 3485
rect 5172 3476 5224 3528
rect 7104 3544 7156 3596
rect 6460 3519 6512 3528
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 8300 3519 8352 3528
rect 8300 3485 8309 3519
rect 8309 3485 8343 3519
rect 8343 3485 8352 3519
rect 8300 3476 8352 3485
rect 8852 3519 8904 3528
rect 8852 3485 8861 3519
rect 8861 3485 8895 3519
rect 8895 3485 8904 3519
rect 8852 3476 8904 3485
rect 4712 3451 4764 3460
rect 4712 3417 4721 3451
rect 4721 3417 4755 3451
rect 4755 3417 4764 3451
rect 4712 3408 4764 3417
rect 5356 3408 5408 3460
rect 7104 3408 7156 3460
rect 3884 3340 3936 3392
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 4988 3340 5040 3392
rect 5540 3340 5592 3392
rect 8116 3340 8168 3392
rect 9128 3340 9180 3392
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 5194 3238 5246 3290
rect 5258 3238 5310 3290
rect 5322 3238 5374 3290
rect 4804 3136 4856 3188
rect 4436 3068 4488 3120
rect 3424 3000 3476 3052
rect 3884 3000 3936 3052
rect 4068 3000 4120 3052
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 3516 2864 3568 2916
rect 8300 3136 8352 3188
rect 5816 3000 5868 3052
rect 6736 3000 6788 3052
rect 7288 3000 7340 3052
rect 8392 3068 8444 3120
rect 8760 3111 8812 3120
rect 8760 3077 8769 3111
rect 8769 3077 8803 3111
rect 8803 3077 8812 3111
rect 8760 3068 8812 3077
rect 9036 3068 9088 3120
rect 11152 3068 11204 3120
rect 8208 3000 8260 3052
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9496 3000 9548 3009
rect 5724 2864 5776 2916
rect 5356 2796 5408 2848
rect 6552 2839 6604 2848
rect 6552 2805 6561 2839
rect 6561 2805 6595 2839
rect 6595 2805 6604 2839
rect 6552 2796 6604 2805
rect 6736 2864 6788 2916
rect 7012 2864 7064 2916
rect 7564 2864 7616 2916
rect 9036 2975 9088 2984
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 8208 2796 8260 2848
rect 8484 2796 8536 2848
rect 8668 2796 8720 2848
rect 7566 2694 7618 2746
rect 7630 2694 7682 2746
rect 7694 2694 7746 2746
rect 7758 2694 7810 2746
rect 7822 2694 7874 2746
rect 10048 2728 10100 2780
rect 13636 2728 13688 2780
rect 9956 2660 10008 2712
rect 13912 2796 13964 2848
rect 3608 2592 3660 2644
rect 5448 2592 5500 2644
rect 6460 2592 6512 2644
rect 3884 2524 3936 2576
rect 5724 2524 5776 2576
rect 6368 2524 6420 2576
rect 6736 2524 6788 2576
rect 13544 2592 13596 2644
rect 3976 2456 4028 2508
rect 20 1504 72 1556
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 4988 2388 5040 2440
rect 6000 2456 6052 2508
rect 8300 2524 8352 2576
rect 9220 2524 9272 2576
rect 15200 2524 15252 2576
rect 7932 2499 7984 2508
rect 7932 2465 7941 2499
rect 7941 2465 7975 2499
rect 7975 2465 7984 2499
rect 7932 2456 7984 2465
rect 3240 2320 3292 2372
rect 5632 2320 5684 2372
rect 2964 2252 3016 2304
rect 4436 2295 4488 2304
rect 4436 2261 4445 2295
rect 4445 2261 4479 2295
rect 4479 2261 4488 2295
rect 4436 2252 4488 2261
rect 5816 2252 5868 2304
rect 6552 2320 6604 2372
rect 8576 2388 8628 2440
rect 9220 2388 9272 2440
rect 7564 2320 7616 2372
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 5194 2150 5246 2202
rect 5258 2150 5310 2202
rect 5322 2150 5374 2202
rect 3884 2091 3936 2100
rect 3884 2057 3893 2091
rect 3893 2057 3927 2091
rect 3927 2057 3936 2091
rect 3884 2048 3936 2057
rect 4252 2048 4304 2100
rect 6092 2048 6144 2100
rect 6644 2048 6696 2100
rect 7196 2048 7248 2100
rect 7288 2048 7340 2100
rect 4528 1980 4580 2032
rect 4804 1912 4856 1964
rect 4988 1912 5040 1964
rect 8024 2048 8076 2100
rect 9496 2048 9548 2100
rect 5540 1912 5592 1964
rect 5816 1912 5868 1964
rect 8300 1980 8352 2032
rect 8852 2023 8904 2032
rect 8852 1989 8861 2023
rect 8861 1989 8895 2023
rect 8895 1989 8904 2023
rect 8852 1980 8904 1989
rect 5172 1776 5224 1828
rect 4896 1708 4948 1760
rect 5908 1844 5960 1896
rect 8116 1912 8168 1964
rect 8760 1912 8812 1964
rect 7380 1844 7432 1896
rect 9404 1912 9456 1964
rect 22100 2320 22152 2372
rect 6184 1776 6236 1828
rect 6736 1776 6788 1828
rect 7564 1776 7616 1828
rect 8024 1819 8076 1828
rect 8024 1785 8033 1819
rect 8033 1785 8067 1819
rect 8067 1785 8076 1819
rect 8024 1776 8076 1785
rect 8668 1819 8720 1828
rect 8668 1785 8677 1819
rect 8677 1785 8711 1819
rect 8711 1785 8720 1819
rect 8668 1776 8720 1785
rect 9220 1776 9272 1828
rect 13820 1776 13872 1828
rect 16856 1776 16908 1828
rect 7566 1606 7618 1658
rect 7630 1606 7682 1658
rect 7694 1606 7746 1658
rect 7758 1606 7810 1658
rect 7822 1606 7874 1658
rect 3056 1504 3108 1556
rect 4712 1547 4764 1556
rect 4712 1513 4721 1547
rect 4721 1513 4755 1547
rect 4755 1513 4764 1547
rect 4712 1504 4764 1513
rect 5448 1504 5500 1556
rect 3148 1436 3200 1488
rect 4160 1479 4212 1488
rect 756 1368 808 1420
rect 4160 1445 4169 1479
rect 4169 1445 4203 1479
rect 4203 1445 4212 1479
rect 4160 1436 4212 1445
rect 4804 1436 4856 1488
rect 10508 1504 10560 1556
rect 5724 1436 5776 1488
rect 8760 1436 8812 1488
rect 8944 1479 8996 1488
rect 8944 1445 8953 1479
rect 8953 1445 8987 1479
rect 8987 1445 8996 1479
rect 8944 1436 8996 1445
rect 3332 1300 3384 1352
rect 3700 1300 3752 1352
rect 4620 1343 4672 1352
rect 4620 1309 4629 1343
rect 4629 1309 4663 1343
rect 4663 1309 4672 1343
rect 4620 1300 4672 1309
rect 5356 1300 5408 1352
rect 2596 892 2648 944
rect 4528 1232 4580 1284
rect 5632 1300 5684 1352
rect 6644 1343 6696 1352
rect 6644 1309 6653 1343
rect 6653 1309 6687 1343
rect 6687 1309 6696 1343
rect 6644 1300 6696 1309
rect 8300 1300 8352 1352
rect 8668 1368 8720 1420
rect 8760 1300 8812 1352
rect 8944 1300 8996 1352
rect 9128 1343 9180 1352
rect 9128 1309 9137 1343
rect 9137 1309 9171 1343
rect 9171 1309 9180 1343
rect 9128 1300 9180 1309
rect 16672 1368 16724 1420
rect 2872 1164 2924 1216
rect 3608 1207 3660 1216
rect 3608 1173 3617 1207
rect 3617 1173 3651 1207
rect 3651 1173 3660 1207
rect 3608 1164 3660 1173
rect 3884 1207 3936 1216
rect 3884 1173 3893 1207
rect 3893 1173 3927 1207
rect 3927 1173 3936 1207
rect 3884 1164 3936 1173
rect 4988 1207 5040 1216
rect 4988 1173 4997 1207
rect 4997 1173 5031 1207
rect 5031 1173 5040 1207
rect 4988 1164 5040 1173
rect 5540 1164 5592 1216
rect 6736 1207 6788 1216
rect 6736 1173 6745 1207
rect 6745 1173 6779 1207
rect 6779 1173 6788 1207
rect 6736 1164 6788 1173
rect 7196 1207 7248 1216
rect 7196 1173 7205 1207
rect 7205 1173 7239 1207
rect 7239 1173 7248 1207
rect 7196 1164 7248 1173
rect 7932 1207 7984 1216
rect 7932 1173 7941 1207
rect 7941 1173 7975 1207
rect 7975 1173 7984 1207
rect 7932 1164 7984 1173
rect 8392 1207 8444 1216
rect 8392 1173 8401 1207
rect 8401 1173 8435 1207
rect 8435 1173 8444 1207
rect 8392 1164 8444 1173
rect 8484 1164 8536 1216
rect 9956 1232 10008 1284
rect 16764 1232 16816 1284
rect 9036 1164 9088 1216
rect 9220 1207 9272 1216
rect 9220 1173 9229 1207
rect 9229 1173 9263 1207
rect 9263 1173 9272 1207
rect 9220 1164 9272 1173
rect 5066 1062 5118 1114
rect 5130 1062 5182 1114
rect 5194 1062 5246 1114
rect 5258 1062 5310 1114
rect 5322 1062 5374 1114
rect 7196 960 7248 1012
rect 9036 960 9088 1012
rect 7932 892 7984 944
rect 8668 892 8720 944
rect 16580 892 16632 944
rect 2320 824 2372 876
rect 4620 824 4672 876
rect 8300 824 8352 876
rect 9312 824 9364 876
rect 2412 756 2464 808
rect 4528 756 4580 808
rect 3884 688 3936 740
rect 5724 688 5776 740
<< metal2 >>
rect 1789 13984 2149 13994
rect 1789 13966 4333 13984
rect 1789 13450 1817 13966
rect 2119 13956 4333 13966
rect 4305 13712 4333 13956
rect 1688 13422 1817 13450
rect 4249 13684 4333 13712
rect 5356 13932 9630 13960
rect 4249 13456 4277 13684
rect 4249 13428 4418 13456
rect 938 12200 994 13000
rect 1398 12200 1454 13000
rect 952 11014 980 12200
rect 1308 11620 1360 11626
rect 1308 11562 1360 11568
rect 1320 11354 1348 11562
rect 1308 11348 1360 11354
rect 1308 11290 1360 11296
rect 20 11008 72 11014
rect 20 10950 72 10956
rect 940 11008 992 11014
rect 940 10950 992 10956
rect 32 1562 60 10950
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 754 9616 810 9625
rect 754 9551 810 9560
rect 20 1556 72 1562
rect 20 1498 72 1504
rect 768 1426 796 9551
rect 952 9489 980 10610
rect 1412 10146 1440 12200
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1504 11150 1532 11630
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1688 10606 1716 13422
rect 1858 12200 1914 13000
rect 2318 12200 2374 13000
rect 2778 12200 2834 13000
rect 3238 12200 3294 13000
rect 3698 12200 3754 13000
rect 4158 12200 4214 13000
rect 1872 11234 1900 12200
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2148 11286 2176 11834
rect 1780 11206 1900 11234
rect 2136 11280 2188 11286
rect 2136 11222 2188 11228
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1584 10532 1636 10538
rect 1584 10474 1636 10480
rect 1044 10118 1440 10146
rect 938 9480 994 9489
rect 938 9415 994 9424
rect 848 8900 900 8906
rect 848 8842 900 8848
rect 860 6497 888 8842
rect 952 7002 980 9415
rect 1044 7478 1072 10118
rect 1596 10062 1624 10474
rect 1688 10130 1716 10542
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1412 9178 1440 9998
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1398 9072 1454 9081
rect 1398 9007 1454 9016
rect 1412 8922 1440 9007
rect 1136 8894 1440 8922
rect 1136 7546 1164 8894
rect 1216 8832 1268 8838
rect 1216 8774 1268 8780
rect 1228 7585 1256 8774
rect 1400 8628 1452 8634
rect 1320 8588 1400 8616
rect 1320 7970 1348 8588
rect 1400 8570 1452 8576
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8090 1440 8434
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1320 7942 1440 7970
rect 1214 7576 1270 7585
rect 1124 7540 1176 7546
rect 1214 7511 1270 7520
rect 1124 7482 1176 7488
rect 1032 7472 1084 7478
rect 1032 7414 1084 7420
rect 940 6996 992 7002
rect 940 6938 992 6944
rect 846 6488 902 6497
rect 846 6423 902 6432
rect 1412 5370 1440 7942
rect 1504 7410 1532 9862
rect 1688 9722 1716 10066
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 9110 1624 9454
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1596 8537 1624 8910
rect 1582 8528 1638 8537
rect 1582 8463 1638 8472
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1596 7342 1624 8230
rect 1688 7750 1716 9658
rect 1780 8634 1808 11206
rect 1860 11144 1912 11150
rect 1860 11086 1912 11092
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1780 7954 1808 8366
rect 1872 8090 1900 11086
rect 2134 10704 2190 10713
rect 1952 10668 2004 10674
rect 2134 10639 2190 10648
rect 1952 10610 2004 10616
rect 1964 10130 1992 10610
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2056 10266 2084 10406
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 2148 9674 2176 10639
rect 2240 10169 2268 11086
rect 2226 10160 2282 10169
rect 2226 10095 2282 10104
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 2240 9722 2268 9930
rect 2056 9646 2176 9674
rect 2228 9716 2280 9722
rect 2228 9658 2280 9664
rect 2056 9382 2084 9646
rect 2044 9376 2096 9382
rect 2044 9318 2096 9324
rect 2044 8968 2096 8974
rect 2228 8968 2280 8974
rect 2044 8910 2096 8916
rect 2226 8936 2228 8945
rect 2280 8936 2282 8945
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1964 8498 1992 8774
rect 2056 8673 2084 8910
rect 2226 8871 2282 8880
rect 2136 8832 2188 8838
rect 2134 8800 2136 8809
rect 2188 8800 2190 8809
rect 2134 8735 2190 8744
rect 2042 8664 2098 8673
rect 2332 8616 2360 12200
rect 2792 11830 2820 12200
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2566 11452 2874 11472
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11376 2874 11396
rect 2976 11286 3004 11698
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3160 11286 3188 11494
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2424 9042 2452 10950
rect 2608 10849 2636 10950
rect 2594 10840 2650 10849
rect 2594 10775 2650 10784
rect 2700 10606 2728 10950
rect 2780 10692 2832 10698
rect 2780 10634 2832 10640
rect 2688 10600 2740 10606
rect 2792 10577 2820 10634
rect 2688 10542 2740 10548
rect 2778 10568 2834 10577
rect 2778 10503 2834 10512
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 2566 10364 2874 10384
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10288 2874 10308
rect 2976 10305 3004 10406
rect 2962 10296 3018 10305
rect 2962 10231 3018 10240
rect 3160 10198 3188 10406
rect 3148 10192 3200 10198
rect 3054 10160 3110 10169
rect 3148 10134 3200 10140
rect 3054 10095 3110 10104
rect 2964 9920 3016 9926
rect 2870 9888 2926 9897
rect 2964 9862 3016 9868
rect 2870 9823 2926 9832
rect 2778 9752 2834 9761
rect 2778 9687 2834 9696
rect 2792 9654 2820 9687
rect 2780 9648 2832 9654
rect 2884 9625 2912 9823
rect 2780 9590 2832 9596
rect 2870 9616 2926 9625
rect 2870 9551 2926 9560
rect 2778 9480 2834 9489
rect 2778 9415 2780 9424
rect 2832 9415 2834 9424
rect 2780 9386 2832 9392
rect 2566 9276 2874 9296
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9200 2874 9220
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2412 9036 2464 9042
rect 2412 8978 2464 8984
rect 2700 8945 2728 9046
rect 2502 8936 2558 8945
rect 2686 8936 2742 8945
rect 2558 8894 2636 8922
rect 2502 8871 2558 8880
rect 2608 8786 2636 8894
rect 2686 8871 2742 8880
rect 2608 8758 2912 8786
rect 2042 8599 2098 8608
rect 2148 8588 2360 8616
rect 2778 8664 2834 8673
rect 2778 8599 2780 8608
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 2042 8392 2098 8401
rect 2042 8327 2098 8336
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1964 8129 1992 8230
rect 1950 8120 2006 8129
rect 1860 8084 1912 8090
rect 1950 8055 2006 8064
rect 1860 8026 1912 8032
rect 1858 7984 1914 7993
rect 1768 7948 1820 7954
rect 1858 7919 1914 7928
rect 1768 7890 1820 7896
rect 1872 7886 1900 7919
rect 1860 7880 1912 7886
rect 1912 7840 1992 7868
rect 1860 7822 1912 7828
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1688 6798 1716 7686
rect 1860 7472 1912 7478
rect 1860 7414 1912 7420
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 1596 6458 1624 6666
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1582 6352 1638 6361
rect 1492 6316 1544 6322
rect 1582 6287 1584 6296
rect 1492 6258 1544 6264
rect 1636 6287 1638 6296
rect 1584 6258 1636 6264
rect 1504 5914 1532 6258
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1688 5778 1716 6734
rect 1780 6458 1808 7346
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1766 5808 1822 5817
rect 1676 5772 1728 5778
rect 1872 5794 1900 7414
rect 1964 7410 1992 7840
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1964 6866 1992 7346
rect 2056 7274 2084 8327
rect 2044 7268 2096 7274
rect 2044 7210 2096 7216
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 2044 6656 2096 6662
rect 2044 6598 2096 6604
rect 2056 6322 2084 6598
rect 2044 6316 2096 6322
rect 2148 6304 2176 8588
rect 2832 8599 2834 8608
rect 2780 8570 2832 8576
rect 2320 8492 2372 8498
rect 2240 8452 2320 8480
rect 2240 8022 2268 8452
rect 2320 8434 2372 8440
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2412 8356 2464 8362
rect 2412 8298 2464 8304
rect 2318 8120 2374 8129
rect 2318 8055 2374 8064
rect 2228 8016 2280 8022
rect 2228 7958 2280 7964
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2240 6458 2268 7142
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2332 6338 2360 8055
rect 2424 7818 2452 8298
rect 2608 8276 2636 8366
rect 2792 8276 2820 8434
rect 2884 8430 2912 8758
rect 2976 8616 3004 9862
rect 3068 9602 3096 10095
rect 3068 9574 3188 9602
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3068 9178 3096 9454
rect 3160 9382 3188 9574
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 3252 9058 3280 12200
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 3344 11150 3372 11222
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3514 10704 3570 10713
rect 3514 10639 3570 10648
rect 3528 10606 3556 10639
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3620 10441 3648 11086
rect 3606 10432 3662 10441
rect 3606 10367 3662 10376
rect 3424 10192 3476 10198
rect 3424 10134 3476 10140
rect 3332 9988 3384 9994
rect 3332 9930 3384 9936
rect 3344 9761 3372 9930
rect 3330 9752 3386 9761
rect 3330 9687 3386 9696
rect 3160 9030 3280 9058
rect 2976 8588 3096 8616
rect 2962 8528 3018 8537
rect 2962 8463 3018 8472
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2492 8248 2820 8276
rect 2492 8072 2520 8248
rect 2566 8188 2874 8208
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8112 2874 8132
rect 2976 8090 3004 8463
rect 2964 8084 3016 8090
rect 2492 8044 2544 8072
rect 2412 7812 2464 7818
rect 2412 7754 2464 7760
rect 2410 7440 2466 7449
rect 2410 7375 2412 7384
rect 2464 7375 2466 7384
rect 2412 7346 2464 7352
rect 2412 7200 2464 7206
rect 2516 7188 2544 8044
rect 2964 8026 3016 8032
rect 3068 7970 3096 8588
rect 2976 7942 3096 7970
rect 2976 7342 3004 7942
rect 3056 7880 3108 7886
rect 3056 7822 3108 7828
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2412 7142 2464 7148
rect 2492 7160 2544 7188
rect 2964 7200 3016 7206
rect 2424 7002 2452 7142
rect 2412 6996 2464 7002
rect 2492 6984 2520 7160
rect 2964 7142 3016 7148
rect 2566 7100 2874 7120
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7024 2874 7044
rect 2492 6956 2636 6984
rect 2412 6938 2464 6944
rect 2502 6624 2558 6633
rect 2502 6559 2558 6568
rect 2332 6310 2452 6338
rect 2148 6276 2268 6304
rect 2044 6258 2096 6264
rect 2134 6216 2190 6225
rect 2240 6202 2268 6276
rect 2424 6254 2452 6310
rect 2412 6248 2464 6254
rect 2240 6174 2360 6202
rect 2412 6190 2464 6196
rect 2516 6186 2544 6559
rect 2608 6186 2636 6956
rect 2870 6896 2926 6905
rect 2870 6831 2926 6840
rect 2884 6662 2912 6831
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2134 6151 2136 6160
rect 2188 6151 2190 6160
rect 2136 6122 2188 6128
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 1872 5766 1992 5794
rect 1766 5743 1822 5752
rect 1676 5714 1728 5720
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 1596 4729 1624 5646
rect 1780 5574 1808 5743
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1964 5234 1992 5766
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 2240 5166 2268 6054
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 1582 4720 1638 4729
rect 1582 4655 1638 4664
rect 756 1420 808 1426
rect 756 1362 808 1368
rect 2332 882 2360 6174
rect 2504 6180 2556 6186
rect 2504 6122 2556 6128
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5896 2452 6054
rect 2566 6012 2874 6032
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5936 2874 5956
rect 2424 5868 2544 5896
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2320 876 2372 882
rect 2320 818 2372 824
rect 2424 814 2452 5306
rect 2516 1873 2544 5868
rect 2778 5672 2834 5681
rect 2778 5607 2834 5616
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2502 1864 2558 1873
rect 2502 1799 2558 1808
rect 2608 950 2636 5170
rect 2792 2774 2820 5607
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2884 3346 2912 5170
rect 2976 3534 3004 7142
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2884 3318 3004 3346
rect 2792 2746 2912 2774
rect 2884 1222 2912 2746
rect 2976 2310 3004 3318
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 3068 1562 3096 7822
rect 3056 1556 3108 1562
rect 3056 1498 3108 1504
rect 3160 1494 3188 9030
rect 3436 8974 3464 10134
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3240 8968 3292 8974
rect 3424 8968 3476 8974
rect 3240 8910 3292 8916
rect 3330 8936 3386 8945
rect 3252 8242 3280 8910
rect 3424 8910 3476 8916
rect 3330 8871 3386 8880
rect 3344 8362 3372 8871
rect 3422 8800 3478 8809
rect 3422 8735 3478 8744
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3252 8214 3372 8242
rect 3344 7993 3372 8214
rect 3330 7984 3386 7993
rect 3330 7919 3386 7928
rect 3330 7712 3386 7721
rect 3330 7647 3386 7656
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3252 5574 3280 6598
rect 3344 6236 3372 7647
rect 3436 6390 3464 8735
rect 3528 7478 3556 9522
rect 3620 9178 3648 9998
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3516 7472 3568 7478
rect 3516 7414 3568 7420
rect 3620 7324 3648 8434
rect 3712 7562 3740 12200
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 3804 9738 3832 11766
rect 3882 11112 3938 11121
rect 3882 11047 3938 11056
rect 3896 10742 3924 11047
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 3882 10568 3938 10577
rect 3882 10503 3938 10512
rect 3896 9994 3924 10503
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 3804 9710 3924 9738
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3804 8838 3832 9590
rect 3896 9110 3924 9710
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3988 8650 4016 11766
rect 4066 11112 4122 11121
rect 4066 11047 4122 11056
rect 4080 10062 4108 11047
rect 4068 10056 4120 10062
rect 4172 10033 4200 12200
rect 4390 11384 4418 13428
rect 4618 12200 4674 13000
rect 5078 12200 5134 13000
rect 4390 11356 4478 11384
rect 4450 11234 4478 11356
rect 4540 11354 4568 11506
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4344 11212 4396 11218
rect 4450 11206 4568 11234
rect 4344 11154 4396 11160
rect 4368 11140 4396 11154
rect 4368 11112 4476 11140
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4250 10840 4306 10849
rect 4250 10775 4306 10784
rect 4068 9998 4120 10004
rect 4158 10024 4214 10033
rect 4158 9959 4214 9968
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4068 9512 4120 9518
rect 4172 9466 4200 9862
rect 4120 9460 4200 9466
rect 4068 9454 4200 9460
rect 4080 9438 4200 9454
rect 4264 9042 4292 10775
rect 4356 10713 4384 11018
rect 4342 10704 4398 10713
rect 4342 10639 4398 10648
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 4356 10130 4384 10474
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4342 10024 4398 10033
rect 4342 9959 4398 9968
rect 4160 9036 4212 9042
rect 4160 8978 4212 8984
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4068 8968 4120 8974
rect 4172 8945 4200 8978
rect 4068 8910 4120 8916
rect 4158 8936 4214 8945
rect 3896 8622 4016 8650
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3804 8022 3832 8298
rect 3792 8016 3844 8022
rect 3792 7958 3844 7964
rect 3896 7721 3924 8622
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3882 7712 3938 7721
rect 3882 7647 3938 7656
rect 3882 7576 3938 7585
rect 3712 7534 3832 7562
rect 3528 7296 3648 7324
rect 3528 6798 3556 7296
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3424 6384 3476 6390
rect 3424 6326 3476 6332
rect 3528 6254 3556 6598
rect 3516 6248 3568 6254
rect 3344 6208 3464 6236
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3238 5400 3294 5409
rect 3238 5335 3294 5344
rect 3252 2378 3280 5335
rect 3344 4690 3372 5714
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3436 4570 3464 6208
rect 3516 6190 3568 6196
rect 3514 5944 3570 5953
rect 3514 5879 3570 5888
rect 3528 5030 3556 5879
rect 3620 5681 3648 7142
rect 3700 6860 3752 6866
rect 3700 6802 3752 6808
rect 3606 5672 3662 5681
rect 3606 5607 3662 5616
rect 3712 5574 3740 6802
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3344 4542 3464 4570
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 3148 1488 3200 1494
rect 3148 1430 3200 1436
rect 3344 1358 3372 4542
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3436 3058 3464 4422
rect 3528 4010 3556 4966
rect 3620 4690 3648 5510
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 3620 4146 3648 4626
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 3514 3360 3570 3369
rect 3514 3295 3570 3304
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3528 2922 3556 3295
rect 3606 2952 3662 2961
rect 3516 2916 3568 2922
rect 3606 2887 3662 2896
rect 3516 2858 3568 2864
rect 3620 2650 3648 2887
rect 3608 2644 3660 2650
rect 3608 2586 3660 2592
rect 3606 1728 3662 1737
rect 3606 1663 3662 1672
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 3620 1222 3648 1663
rect 3712 1358 3740 5306
rect 3804 2446 3832 7534
rect 3882 7511 3938 7520
rect 3896 7410 3924 7511
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3988 6848 4016 8502
rect 3896 6820 4016 6848
rect 3896 5370 3924 6820
rect 3974 6488 4030 6497
rect 3974 6423 4030 6432
rect 3988 6322 4016 6423
rect 3976 6316 4028 6322
rect 3976 6258 4028 6264
rect 3974 5672 4030 5681
rect 3974 5607 4030 5616
rect 3988 5574 4016 5607
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 4078 3924 4966
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3988 3534 4016 5102
rect 4080 4162 4108 8910
rect 4158 8871 4214 8880
rect 4160 8356 4212 8362
rect 4160 8298 4212 8304
rect 4172 6798 4200 8298
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4264 8090 4292 8230
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4264 5778 4292 7686
rect 4252 5772 4304 5778
rect 4252 5714 4304 5720
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4172 4826 4200 5578
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4172 4282 4200 4626
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4080 4134 4200 4162
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 3058 3924 3334
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3896 2106 3924 2518
rect 3988 2514 4016 3470
rect 4080 3058 4108 3878
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 3884 2100 3936 2106
rect 3884 2042 3936 2048
rect 4172 1494 4200 4134
rect 4264 3602 4292 5714
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4250 3496 4306 3505
rect 4250 3431 4306 3440
rect 4264 2106 4292 3431
rect 4356 2938 4384 9959
rect 4448 8974 4476 11112
rect 4540 10130 4568 11206
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4448 8090 4476 8434
rect 4540 8294 4568 9114
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4526 8120 4582 8129
rect 4436 8084 4488 8090
rect 4526 8055 4582 8064
rect 4436 8026 4488 8032
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 7206 4476 7686
rect 4540 7274 4568 8055
rect 4528 7268 4580 7274
rect 4528 7210 4580 7216
rect 4436 7200 4488 7206
rect 4632 7154 4660 12200
rect 5092 11336 5120 12200
rect 4816 11308 5120 11336
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4724 10674 4752 11086
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4710 10568 4766 10577
rect 4710 10503 4766 10512
rect 4724 9489 4752 10503
rect 4710 9480 4766 9489
rect 4710 9415 4766 9424
rect 4816 9194 4844 11308
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4908 10674 4936 11154
rect 5000 11014 5028 11119
rect 5356 11056 5384 13932
rect 5538 12200 5594 13000
rect 5998 12200 6054 13000
rect 6458 12200 6514 13000
rect 5552 11830 5580 12200
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5460 11150 5488 11630
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5908 11620 5960 11626
rect 5908 11562 5960 11568
rect 5552 11270 5580 11562
rect 5552 11242 5620 11270
rect 5460 11122 5528 11150
rect 5356 11028 5454 11056
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 5066 10908 5374 10928
rect 5066 10906 5072 10908
rect 5128 10906 5152 10908
rect 5208 10906 5232 10908
rect 5288 10906 5312 10908
rect 5368 10906 5374 10908
rect 5128 10854 5130 10906
rect 5310 10854 5312 10906
rect 5066 10852 5072 10854
rect 5128 10852 5152 10854
rect 5208 10852 5232 10854
rect 5288 10852 5312 10854
rect 5368 10852 5374 10854
rect 5066 10832 5374 10852
rect 5426 10798 5454 11028
rect 5000 10770 5454 10798
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 5000 10577 5028 10770
rect 5080 10736 5132 10742
rect 5500 10694 5528 11122
rect 5080 10678 5132 10684
rect 4986 10568 5042 10577
rect 4986 10503 5042 10512
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 9586 4936 10406
rect 5092 10010 5120 10678
rect 5172 10668 5224 10674
rect 5172 10610 5224 10616
rect 5460 10666 5528 10694
rect 5184 10033 5212 10610
rect 5460 10606 5488 10666
rect 5448 10600 5500 10606
rect 5262 10568 5318 10577
rect 5592 10572 5620 11242
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5736 10674 5764 10950
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5448 10542 5500 10548
rect 5552 10544 5620 10572
rect 5262 10503 5318 10512
rect 5276 10130 5304 10503
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5000 9982 5120 10010
rect 5170 10024 5226 10033
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 5000 9217 5028 9982
rect 5552 9994 5580 10544
rect 5630 10296 5686 10305
rect 5630 10231 5686 10240
rect 5170 9959 5226 9968
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5066 9820 5374 9840
rect 5066 9818 5072 9820
rect 5128 9818 5152 9820
rect 5208 9818 5232 9820
rect 5288 9818 5312 9820
rect 5368 9818 5374 9820
rect 5128 9766 5130 9818
rect 5310 9766 5312 9818
rect 5066 9764 5072 9766
rect 5128 9764 5152 9766
rect 5208 9764 5232 9766
rect 5288 9764 5312 9766
rect 5368 9764 5374 9766
rect 5066 9744 5374 9764
rect 5078 9688 5134 9697
rect 5644 9674 5672 10231
rect 5736 9897 5764 10610
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5722 9888 5778 9897
rect 5722 9823 5778 9832
rect 5134 9646 5304 9674
rect 5078 9623 5134 9632
rect 4724 9166 4844 9194
rect 4986 9208 5042 9217
rect 4724 8566 4752 9166
rect 4986 9143 5042 9152
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4436 7142 4488 7148
rect 4540 7126 4660 7154
rect 4540 6882 4568 7126
rect 4448 6854 4568 6882
rect 4620 6860 4672 6866
rect 4448 3618 4476 6854
rect 4620 6802 4672 6808
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 3738 4568 6734
rect 4632 5574 4660 6802
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4632 4185 4660 5510
rect 4724 4264 4752 8298
rect 4816 8265 4844 9046
rect 5092 8974 5120 9114
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5276 8820 5304 9646
rect 5448 9648 5500 9654
rect 5354 9616 5410 9625
rect 5448 9590 5500 9596
rect 5552 9646 5672 9674
rect 5736 9654 5764 9823
rect 5724 9648 5776 9654
rect 5354 9551 5356 9560
rect 5408 9551 5410 9560
rect 5356 9522 5408 9528
rect 5368 8956 5396 9522
rect 5460 9058 5488 9590
rect 5552 9178 5580 9646
rect 5724 9590 5776 9596
rect 5632 9512 5684 9518
rect 5724 9512 5776 9518
rect 5632 9454 5684 9460
rect 5722 9480 5724 9489
rect 5776 9480 5778 9489
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5460 9030 5580 9058
rect 5368 8928 5488 8956
rect 4908 8792 5304 8820
rect 4802 8256 4858 8265
rect 4802 8191 4858 8200
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4816 7478 4844 8026
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4816 5409 4844 7210
rect 4908 7041 4936 8792
rect 5066 8732 5374 8752
rect 5066 8730 5072 8732
rect 5128 8730 5152 8732
rect 5208 8730 5232 8732
rect 5288 8730 5312 8732
rect 5368 8730 5374 8732
rect 5128 8678 5130 8730
rect 5310 8678 5312 8730
rect 5066 8676 5072 8678
rect 5128 8676 5152 8678
rect 5208 8676 5232 8678
rect 5288 8676 5312 8678
rect 5368 8676 5374 8678
rect 5066 8656 5374 8676
rect 5460 8616 5488 8928
rect 5552 8634 5580 9030
rect 5644 8906 5672 9454
rect 5722 9415 5778 9424
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5368 8588 5488 8616
rect 5540 8628 5592 8634
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 4894 7032 4950 7041
rect 4894 6967 4950 6976
rect 5000 6798 5028 8502
rect 5368 7857 5396 8588
rect 5540 8570 5592 8576
rect 5644 8498 5672 8842
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5354 7848 5410 7857
rect 5354 7783 5410 7792
rect 5066 7644 5374 7664
rect 5066 7642 5072 7644
rect 5128 7642 5152 7644
rect 5208 7642 5232 7644
rect 5288 7642 5312 7644
rect 5368 7642 5374 7644
rect 5128 7590 5130 7642
rect 5310 7590 5312 7642
rect 5066 7588 5072 7590
rect 5128 7588 5152 7590
rect 5208 7588 5232 7590
rect 5288 7588 5312 7590
rect 5368 7588 5374 7590
rect 5066 7568 5374 7588
rect 5460 7410 5488 8230
rect 5552 7449 5580 8230
rect 5630 7984 5686 7993
rect 5630 7919 5686 7928
rect 5644 7886 5672 7919
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5630 7712 5686 7721
rect 5630 7647 5686 7656
rect 5538 7440 5594 7449
rect 5448 7404 5500 7410
rect 5538 7375 5594 7384
rect 5448 7346 5500 7352
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5446 7032 5502 7041
rect 5446 6967 5502 6976
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4988 6792 5040 6798
rect 4988 6734 5040 6740
rect 4802 5400 4858 5409
rect 4802 5335 4858 5344
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4816 4690 4844 5238
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4724 4236 4844 4264
rect 4618 4176 4674 4185
rect 4618 4111 4674 4120
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4448 3590 4568 3618
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4448 3126 4476 3334
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4356 2910 4476 2938
rect 4448 2825 4476 2910
rect 4434 2816 4490 2825
rect 4434 2751 4490 2760
rect 4434 2408 4490 2417
rect 4434 2343 4490 2352
rect 4448 2310 4476 2343
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 4252 2100 4304 2106
rect 4252 2042 4304 2048
rect 4540 2038 4568 3590
rect 4632 3534 4660 3946
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 4724 3466 4752 4082
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4618 3088 4674 3097
rect 4618 3023 4674 3032
rect 4632 2446 4660 3023
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4528 2032 4580 2038
rect 4528 1974 4580 1980
rect 4724 1562 4752 3402
rect 4816 3194 4844 4236
rect 4908 3670 4936 6734
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5000 5352 5028 6598
rect 5066 6556 5374 6576
rect 5066 6554 5072 6556
rect 5128 6554 5152 6556
rect 5208 6554 5232 6556
rect 5288 6554 5312 6556
rect 5368 6554 5374 6556
rect 5128 6502 5130 6554
rect 5310 6502 5312 6554
rect 5066 6500 5072 6502
rect 5128 6500 5152 6502
rect 5208 6500 5232 6502
rect 5288 6500 5312 6502
rect 5368 6500 5374 6502
rect 5066 6480 5374 6500
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 5184 5681 5212 6190
rect 5170 5672 5226 5681
rect 5170 5607 5172 5616
rect 5224 5607 5226 5616
rect 5172 5578 5224 5584
rect 5184 5547 5212 5578
rect 5066 5468 5374 5488
rect 5066 5466 5072 5468
rect 5128 5466 5152 5468
rect 5208 5466 5232 5468
rect 5288 5466 5312 5468
rect 5368 5466 5374 5468
rect 5128 5414 5130 5466
rect 5310 5414 5312 5466
rect 5066 5412 5072 5414
rect 5128 5412 5152 5414
rect 5208 5412 5232 5414
rect 5288 5412 5312 5414
rect 5368 5412 5374 5414
rect 5066 5392 5374 5412
rect 5000 5324 5212 5352
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 5000 4282 5028 4762
rect 5184 4593 5212 5324
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5368 4622 5396 4762
rect 5356 4616 5408 4622
rect 5170 4584 5226 4593
rect 5460 4593 5488 6967
rect 5552 6118 5580 7210
rect 5644 6662 5672 7647
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5736 6322 5764 9318
rect 5828 7546 5856 10542
rect 5920 10169 5948 11562
rect 6012 10554 6040 12200
rect 6472 11626 6500 12200
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 6090 10840 6146 10849
rect 6090 10775 6092 10784
rect 6144 10775 6146 10784
rect 6092 10746 6144 10752
rect 6012 10526 6132 10554
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5906 10160 5962 10169
rect 5906 10095 5962 10104
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5920 9761 5948 9998
rect 5906 9752 5962 9761
rect 5906 9687 5962 9696
rect 6012 9602 6040 10406
rect 5920 9574 6040 9602
rect 5920 9382 5948 9574
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 8566 5948 9318
rect 5998 9208 6054 9217
rect 5998 9143 6054 9152
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 5908 8424 5960 8430
rect 6012 8401 6040 9143
rect 5908 8366 5960 8372
rect 5998 8392 6054 8401
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5632 6248 5684 6254
rect 5828 6225 5856 6598
rect 5632 6190 5684 6196
rect 5814 6216 5870 6225
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5538 5944 5594 5953
rect 5538 5879 5540 5888
rect 5592 5879 5594 5888
rect 5540 5850 5592 5856
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5356 4558 5408 4564
rect 5446 4584 5502 4593
rect 5170 4519 5226 4528
rect 5368 4468 5396 4558
rect 5446 4519 5502 4528
rect 5368 4440 5488 4468
rect 5066 4380 5374 4400
rect 5066 4378 5072 4380
rect 5128 4378 5152 4380
rect 5208 4378 5232 4380
rect 5288 4378 5312 4380
rect 5368 4378 5374 4380
rect 5128 4326 5130 4378
rect 5310 4326 5312 4378
rect 5066 4324 5072 4326
rect 5128 4324 5152 4326
rect 5208 4324 5232 4326
rect 5288 4324 5312 4326
rect 5368 4324 5374 4326
rect 5066 4304 5374 4324
rect 4988 4276 5040 4282
rect 5460 4264 5488 4440
rect 4988 4218 5040 4224
rect 5368 4236 5488 4264
rect 4986 4176 5042 4185
rect 4986 4111 5042 4120
rect 4896 3664 4948 3670
rect 4896 3606 4948 3612
rect 5000 3516 5028 4111
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5184 3534 5212 3946
rect 4908 3488 5028 3516
rect 5172 3528 5224 3534
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4908 3074 4936 3488
rect 5172 3470 5224 3476
rect 5368 3466 5396 4236
rect 5446 4176 5502 4185
rect 5446 4111 5502 4120
rect 5356 3460 5408 3466
rect 5356 3402 5408 3408
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4816 3046 4936 3074
rect 4816 2122 4844 3046
rect 4894 2816 4950 2825
rect 4894 2751 4950 2760
rect 4908 2258 4936 2751
rect 5000 2446 5028 3334
rect 5066 3292 5374 3312
rect 5066 3290 5072 3292
rect 5128 3290 5152 3292
rect 5208 3290 5232 3292
rect 5288 3290 5312 3292
rect 5368 3290 5374 3292
rect 5128 3238 5130 3290
rect 5310 3238 5312 3290
rect 5066 3236 5072 3238
rect 5128 3236 5152 3238
rect 5208 3236 5232 3238
rect 5288 3236 5312 3238
rect 5368 3236 5374 3238
rect 5066 3216 5374 3236
rect 5460 3176 5488 4111
rect 5552 4010 5580 5646
rect 5644 5574 5672 6190
rect 5814 6151 5870 6160
rect 5920 5953 5948 8366
rect 6104 8362 6132 10526
rect 6196 9586 6224 11018
rect 6276 10532 6328 10538
rect 6276 10474 6328 10480
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 5998 8327 6054 8336
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 5998 7848 6054 7857
rect 5998 7783 6000 7792
rect 6052 7783 6054 7792
rect 6000 7754 6052 7760
rect 6196 7410 6224 9318
rect 6288 9217 6316 10474
rect 6274 9208 6330 9217
rect 6274 9143 6330 9152
rect 6380 9081 6408 11494
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6552 11144 6604 11150
rect 6604 11104 6684 11132
rect 6552 11086 6604 11092
rect 6366 9072 6422 9081
rect 6366 9007 6422 9016
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6288 7546 6316 8910
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 5906 5944 5962 5953
rect 5906 5879 5962 5888
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5644 4282 5672 4626
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5630 4176 5686 4185
rect 5736 4146 5764 4966
rect 5630 4111 5686 4120
rect 5724 4140 5776 4146
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5276 3148 5488 3176
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5276 2292 5304 3148
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5368 2530 5396 2790
rect 5460 2650 5488 2994
rect 5552 2825 5580 3334
rect 5538 2816 5594 2825
rect 5538 2751 5594 2760
rect 5644 2768 5672 4111
rect 5724 4082 5776 4088
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5736 2922 5764 3878
rect 5828 3738 5856 5170
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5644 2740 5764 2768
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5736 2582 5764 2740
rect 5724 2576 5776 2582
rect 5368 2502 5580 2530
rect 5724 2518 5776 2524
rect 5276 2264 5488 2292
rect 4908 2230 5028 2258
rect 4816 2094 4936 2122
rect 4804 1964 4856 1970
rect 4804 1906 4856 1912
rect 4712 1556 4764 1562
rect 4712 1498 4764 1504
rect 4816 1494 4844 1906
rect 4908 1766 4936 2094
rect 5000 1970 5028 2230
rect 5066 2204 5374 2224
rect 5066 2202 5072 2204
rect 5128 2202 5152 2204
rect 5208 2202 5232 2204
rect 5288 2202 5312 2204
rect 5368 2202 5374 2204
rect 5128 2150 5130 2202
rect 5310 2150 5312 2202
rect 5066 2148 5072 2150
rect 5128 2148 5152 2150
rect 5208 2148 5232 2150
rect 5288 2148 5312 2150
rect 5368 2148 5374 2150
rect 5066 2128 5374 2148
rect 5170 2000 5226 2009
rect 4988 1964 5040 1970
rect 5170 1935 5226 1944
rect 4988 1906 5040 1912
rect 5184 1834 5212 1935
rect 5172 1828 5224 1834
rect 5172 1770 5224 1776
rect 4896 1760 4948 1766
rect 4896 1702 4948 1708
rect 5460 1562 5488 2264
rect 5552 1970 5580 2502
rect 5828 2394 5856 2994
rect 5632 2372 5684 2378
rect 5632 2314 5684 2320
rect 5736 2366 5856 2394
rect 5540 1964 5592 1970
rect 5540 1906 5592 1912
rect 5538 1864 5594 1873
rect 5538 1799 5594 1808
rect 5448 1556 5500 1562
rect 5448 1498 5500 1504
rect 4160 1488 4212 1494
rect 4160 1430 4212 1436
rect 4804 1488 4856 1494
rect 4804 1430 4856 1436
rect 3700 1352 3752 1358
rect 3700 1294 3752 1300
rect 4620 1352 4672 1358
rect 5356 1352 5408 1358
rect 4620 1294 4672 1300
rect 4986 1320 5042 1329
rect 4528 1284 4580 1290
rect 4528 1226 4580 1232
rect 2872 1216 2924 1222
rect 2872 1158 2924 1164
rect 3608 1216 3660 1222
rect 3608 1158 3660 1164
rect 3884 1216 3936 1222
rect 3884 1158 3936 1164
rect 2596 944 2648 950
rect 2596 886 2648 892
rect 2412 808 2464 814
rect 2412 750 2464 756
rect 3896 746 3924 1158
rect 4540 814 4568 1226
rect 4632 882 4660 1294
rect 5408 1300 5488 1306
rect 5356 1294 5488 1300
rect 5368 1278 5488 1294
rect 4986 1255 5042 1264
rect 5000 1222 5028 1255
rect 4988 1216 5040 1222
rect 5460 1193 5488 1278
rect 5552 1222 5580 1799
rect 5644 1358 5672 2314
rect 5736 1494 5764 2366
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5828 1970 5856 2246
rect 5816 1964 5868 1970
rect 5816 1906 5868 1912
rect 5920 1902 5948 4422
rect 6012 4321 6040 7210
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6104 6225 6132 6258
rect 6090 6216 6146 6225
rect 6090 6151 6146 6160
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 6104 5778 6132 5850
rect 6196 5778 6224 7346
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 6104 5370 6132 5578
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6196 5234 6224 5714
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 6104 4570 6132 5034
rect 6196 4690 6224 5170
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6104 4554 6224 4570
rect 6104 4548 6236 4554
rect 6104 4542 6184 4548
rect 5998 4312 6054 4321
rect 5998 4247 6054 4256
rect 6104 4162 6132 4542
rect 6184 4490 6236 4496
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6012 4134 6132 4162
rect 6012 2514 6040 4134
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6104 2106 6132 4014
rect 6196 3738 6224 4218
rect 6184 3732 6236 3738
rect 6184 3674 6236 3680
rect 6092 2100 6144 2106
rect 6092 2042 6144 2048
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 6196 1834 6224 3674
rect 6288 2145 6316 6190
rect 6380 5642 6408 8434
rect 6472 8090 6500 11086
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6564 10674 6592 10950
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6564 10266 6592 10406
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6564 7834 6592 9590
rect 6656 8480 6684 11104
rect 6748 10198 6776 11154
rect 6826 10840 6882 10849
rect 6826 10775 6882 10784
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6734 10024 6790 10033
rect 6734 9959 6790 9968
rect 6748 8634 6776 9959
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6840 8498 6868 10775
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6932 9586 6960 9998
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6828 8492 6880 8498
rect 6656 8452 6776 8480
rect 6748 8378 6776 8452
rect 6828 8434 6880 8440
rect 6748 8350 6868 8378
rect 6564 7806 6684 7834
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6472 5846 6500 6802
rect 6564 6662 6592 7686
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6564 6322 6592 6394
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6380 2582 6408 4966
rect 6656 4808 6684 7806
rect 6840 7546 6868 8350
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6748 6497 6776 7142
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6734 6488 6790 6497
rect 6734 6423 6790 6432
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6472 4780 6684 4808
rect 6472 3942 6500 4780
rect 6644 4684 6696 4690
rect 6644 4626 6696 4632
rect 6550 4448 6606 4457
rect 6550 4383 6606 4392
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6472 2650 6500 3470
rect 6564 2961 6592 4383
rect 6550 2952 6606 2961
rect 6550 2887 6606 2896
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6368 2576 6420 2582
rect 6368 2518 6420 2524
rect 6564 2378 6592 2790
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 6274 2136 6330 2145
rect 6656 2106 6684 4626
rect 6748 3058 6776 5102
rect 6840 4457 6868 6938
rect 6826 4448 6882 4457
rect 6826 4383 6882 4392
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 6840 4078 6868 4218
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6748 2582 6776 2858
rect 6736 2576 6788 2582
rect 6736 2518 6788 2524
rect 6274 2071 6330 2080
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6184 1828 6236 1834
rect 6184 1770 6236 1776
rect 5724 1488 5776 1494
rect 5724 1430 5776 1436
rect 5632 1352 5684 1358
rect 5632 1294 5684 1300
rect 5540 1216 5592 1222
rect 4988 1158 5040 1164
rect 5446 1184 5502 1193
rect 5066 1116 5374 1136
rect 5540 1158 5592 1164
rect 5446 1119 5502 1128
rect 5066 1114 5072 1116
rect 5128 1114 5152 1116
rect 5208 1114 5232 1116
rect 5288 1114 5312 1116
rect 5368 1114 5374 1116
rect 5128 1062 5130 1114
rect 5310 1062 5312 1114
rect 5066 1060 5072 1062
rect 5128 1060 5152 1062
rect 5208 1060 5232 1062
rect 5288 1060 5312 1062
rect 5368 1060 5374 1062
rect 5066 1040 5374 1060
rect 4620 876 4672 882
rect 4620 818 4672 824
rect 4528 808 4580 814
rect 4528 750 4580 756
rect 5736 746 5764 1430
rect 6656 1358 6684 2042
rect 6840 2009 6868 3878
rect 6826 2000 6882 2009
rect 6826 1935 6882 1944
rect 6736 1828 6788 1834
rect 6736 1770 6788 1776
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 6748 1222 6776 1770
rect 6932 1737 6960 9522
rect 7024 8906 7052 11834
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 7566 11452 7874 11472
rect 7566 11450 7572 11452
rect 7628 11450 7652 11452
rect 7708 11450 7732 11452
rect 7788 11450 7812 11452
rect 7868 11450 7874 11452
rect 7628 11398 7630 11450
rect 7810 11398 7812 11450
rect 7566 11396 7572 11398
rect 7628 11396 7652 11398
rect 7708 11396 7732 11398
rect 7788 11396 7812 11398
rect 7868 11396 7874 11398
rect 7566 11376 7874 11396
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7380 11144 7432 11150
rect 7378 11112 7380 11121
rect 7432 11112 7434 11121
rect 7104 11076 7156 11082
rect 7378 11047 7434 11056
rect 7104 11018 7156 11024
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7024 8022 7052 8570
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 7116 6916 7144 11018
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7208 10266 7236 10542
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7208 9897 7236 9930
rect 7194 9888 7250 9897
rect 7194 9823 7250 9832
rect 7300 9466 7328 10610
rect 7378 10432 7434 10441
rect 7378 10367 7434 10376
rect 7392 9586 7420 10367
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7300 9438 7420 9466
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7286 9344 7342 9353
rect 7208 8838 7236 9318
rect 7286 9279 7342 9288
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7208 8498 7236 8570
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 7208 6984 7236 7958
rect 7300 7886 7328 9279
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7392 7002 7420 9438
rect 7380 6996 7432 7002
rect 7208 6956 7328 6984
rect 7116 6888 7236 6916
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7024 2922 7052 6734
rect 7116 4282 7144 6734
rect 7208 6361 7236 6888
rect 7300 6746 7328 6956
rect 7380 6938 7432 6944
rect 7300 6718 7420 6746
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7194 6352 7250 6361
rect 7194 6287 7250 6296
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7104 4004 7156 4010
rect 7104 3946 7156 3952
rect 7116 3602 7144 3946
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 7116 2310 7144 3402
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7208 2106 7236 4082
rect 7300 3058 7328 6598
rect 7392 5817 7420 6718
rect 7484 6390 7512 11222
rect 7840 11144 7892 11150
rect 8024 11144 8076 11150
rect 7892 11104 7972 11132
rect 7840 11086 7892 11092
rect 7566 10364 7874 10384
rect 7566 10362 7572 10364
rect 7628 10362 7652 10364
rect 7708 10362 7732 10364
rect 7788 10362 7812 10364
rect 7868 10362 7874 10364
rect 7628 10310 7630 10362
rect 7810 10310 7812 10362
rect 7566 10308 7572 10310
rect 7628 10308 7652 10310
rect 7708 10308 7732 10310
rect 7788 10308 7812 10310
rect 7868 10308 7874 10310
rect 7566 10288 7874 10308
rect 7656 10056 7708 10062
rect 7654 10024 7656 10033
rect 7708 10024 7710 10033
rect 7654 9959 7710 9968
rect 7840 9920 7892 9926
rect 7760 9868 7840 9874
rect 7760 9862 7892 9868
rect 7760 9846 7880 9862
rect 7760 9586 7788 9846
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7566 9276 7874 9296
rect 7566 9274 7572 9276
rect 7628 9274 7652 9276
rect 7708 9274 7732 9276
rect 7788 9274 7812 9276
rect 7868 9274 7874 9276
rect 7628 9222 7630 9274
rect 7810 9222 7812 9274
rect 7566 9220 7572 9222
rect 7628 9220 7652 9222
rect 7708 9220 7732 9222
rect 7788 9220 7812 9222
rect 7868 9220 7874 9222
rect 7566 9200 7874 9220
rect 7562 9072 7618 9081
rect 7562 9007 7618 9016
rect 7576 8566 7604 9007
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7566 8188 7874 8208
rect 7566 8186 7572 8188
rect 7628 8186 7652 8188
rect 7708 8186 7732 8188
rect 7788 8186 7812 8188
rect 7868 8186 7874 8188
rect 7628 8134 7630 8186
rect 7810 8134 7812 8186
rect 7566 8132 7572 8134
rect 7628 8132 7652 8134
rect 7708 8132 7732 8134
rect 7788 8132 7812 8134
rect 7868 8132 7874 8134
rect 7566 8112 7874 8132
rect 7944 8022 7972 11104
rect 8024 11086 8076 11092
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8036 9058 8064 11086
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 8128 9217 8156 10474
rect 8114 9208 8170 9217
rect 8312 9178 8340 11086
rect 8114 9143 8170 9152
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8036 9030 8156 9058
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7760 7392 7788 7754
rect 7840 7404 7892 7410
rect 7760 7364 7840 7392
rect 7840 7346 7892 7352
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7566 7100 7874 7120
rect 7566 7098 7572 7100
rect 7628 7098 7652 7100
rect 7708 7098 7732 7100
rect 7788 7098 7812 7100
rect 7868 7098 7874 7100
rect 7628 7046 7630 7098
rect 7810 7046 7812 7098
rect 7566 7044 7572 7046
rect 7628 7044 7652 7046
rect 7708 7044 7732 7046
rect 7788 7044 7812 7046
rect 7868 7044 7874 7046
rect 7566 7024 7874 7044
rect 7944 6798 7972 7278
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7378 5808 7434 5817
rect 7378 5743 7434 5752
rect 7484 5370 7512 6190
rect 7566 6012 7874 6032
rect 7566 6010 7572 6012
rect 7628 6010 7652 6012
rect 7708 6010 7732 6012
rect 7788 6010 7812 6012
rect 7868 6010 7874 6012
rect 7628 5958 7630 6010
rect 7810 5958 7812 6010
rect 7566 5956 7572 5958
rect 7628 5956 7652 5958
rect 7708 5956 7732 5958
rect 7788 5956 7812 5958
rect 7868 5956 7874 5958
rect 7566 5936 7874 5956
rect 7944 5778 7972 6734
rect 8036 6458 8064 8910
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8036 6225 8064 6258
rect 8022 6216 8078 6225
rect 8022 6151 8078 6160
rect 8022 5808 8078 5817
rect 7932 5772 7984 5778
rect 8022 5743 8078 5752
rect 7932 5714 7984 5720
rect 7472 5364 7524 5370
rect 7472 5306 7524 5312
rect 7932 5296 7984 5302
rect 7932 5238 7984 5244
rect 7566 4924 7874 4944
rect 7566 4922 7572 4924
rect 7628 4922 7652 4924
rect 7708 4922 7732 4924
rect 7788 4922 7812 4924
rect 7868 4922 7874 4924
rect 7628 4870 7630 4922
rect 7810 4870 7812 4922
rect 7566 4868 7572 4870
rect 7628 4868 7652 4870
rect 7708 4868 7732 4870
rect 7788 4868 7812 4870
rect 7868 4868 7874 4870
rect 7566 4848 7874 4868
rect 7378 4720 7434 4729
rect 7378 4655 7434 4664
rect 7392 3233 7420 4655
rect 7656 4548 7708 4554
rect 7944 4536 7972 5238
rect 7708 4508 7972 4536
rect 7656 4490 7708 4496
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7378 3224 7434 3233
rect 7378 3159 7434 3168
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7484 2938 7512 4150
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7566 3836 7874 3856
rect 7566 3834 7572 3836
rect 7628 3834 7652 3836
rect 7708 3834 7732 3836
rect 7788 3834 7812 3836
rect 7868 3834 7874 3836
rect 7628 3782 7630 3834
rect 7810 3782 7812 3834
rect 7566 3780 7572 3782
rect 7628 3780 7652 3782
rect 7708 3780 7732 3782
rect 7788 3780 7812 3782
rect 7868 3780 7874 3782
rect 7566 3760 7874 3780
rect 7300 2910 7512 2938
rect 7564 2916 7616 2922
rect 7300 2106 7328 2910
rect 7944 2904 7972 4014
rect 7616 2876 7972 2904
rect 7564 2858 7616 2864
rect 7378 2816 7434 2825
rect 7378 2751 7434 2760
rect 7196 2100 7248 2106
rect 7196 2042 7248 2048
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 7392 1902 7420 2751
rect 7566 2748 7874 2768
rect 7566 2746 7572 2748
rect 7628 2746 7652 2748
rect 7708 2746 7732 2748
rect 7788 2746 7812 2748
rect 7868 2746 7874 2748
rect 7628 2694 7630 2746
rect 7810 2694 7812 2746
rect 7566 2692 7572 2694
rect 7628 2692 7652 2694
rect 7708 2692 7732 2694
rect 7788 2692 7812 2694
rect 7868 2692 7874 2694
rect 7566 2672 7874 2692
rect 7930 2544 7986 2553
rect 7930 2479 7932 2488
rect 7984 2479 7986 2488
rect 7932 2450 7984 2456
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 7380 1896 7432 1902
rect 7380 1838 7432 1844
rect 7576 1834 7604 2314
rect 8036 2106 8064 5743
rect 8128 3505 8156 9030
rect 8208 9036 8260 9042
rect 8260 8996 8340 9024
rect 8208 8978 8260 8984
rect 8208 7880 8260 7886
rect 8312 7857 8340 8996
rect 8208 7822 8260 7828
rect 8298 7848 8354 7857
rect 8220 6866 8248 7822
rect 8298 7783 8354 7792
rect 8312 7478 8340 7783
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8312 6610 8340 7414
rect 8404 6730 8432 11290
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8496 9654 8524 11018
rect 8484 9648 8536 9654
rect 8536 9608 8616 9636
rect 8484 9590 8536 9596
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8496 7970 8524 9318
rect 8588 9042 8616 9608
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8588 8090 8616 8570
rect 8680 8498 8708 11698
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9324 11150 9352 11290
rect 9602 11286 9630 13932
rect 10170 12452 11008 12480
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8772 8090 8800 11018
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8864 9722 8892 9998
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8864 8401 8892 8910
rect 8956 8498 8984 10406
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8850 8392 8906 8401
rect 8850 8327 8906 8336
rect 9048 8242 9076 10610
rect 9140 8634 9168 11086
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9312 10464 9364 10470
rect 10170 10424 10198 12452
rect 10506 12336 10562 12345
rect 10506 12271 10562 12280
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 9312 10406 9364 10412
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 8956 8214 9076 8242
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8496 7942 8616 7970
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 8220 6582 8340 6610
rect 8220 5681 8248 6582
rect 8496 6474 8524 7754
rect 8588 7206 8616 7942
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8312 6446 8524 6474
rect 8206 5672 8262 5681
rect 8206 5607 8208 5616
rect 8260 5607 8262 5616
rect 8208 5578 8260 5584
rect 8220 5302 8248 5578
rect 8208 5296 8260 5302
rect 8208 5238 8260 5244
rect 8312 4826 8340 6446
rect 8588 6322 8616 6666
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8680 6186 8708 7142
rect 8956 6905 8984 8214
rect 9232 7954 9260 10406
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9232 7342 9260 7890
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9140 7002 9168 7278
rect 9128 6996 9180 7002
rect 9128 6938 9180 6944
rect 8942 6896 8998 6905
rect 8942 6831 8998 6840
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8772 5710 8800 6054
rect 8864 5846 8892 6666
rect 9048 6322 9076 6802
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8852 5840 8904 5846
rect 8852 5782 8904 5788
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8220 4146 8248 4422
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8114 3496 8170 3505
rect 8114 3431 8170 3440
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8024 2100 8076 2106
rect 8024 2042 8076 2048
rect 8128 1970 8156 3334
rect 8220 3058 8248 4082
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8312 3194 8340 3470
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8404 3126 8432 5170
rect 8496 5166 8524 5510
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8588 4978 8616 5510
rect 8496 4950 8616 4978
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8496 2938 8524 4950
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8404 2910 8524 2938
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8220 2553 8248 2790
rect 8300 2576 8352 2582
rect 8206 2544 8262 2553
rect 8300 2518 8352 2524
rect 8206 2479 8262 2488
rect 8312 2038 8340 2518
rect 8300 2032 8352 2038
rect 8300 1974 8352 1980
rect 8116 1964 8168 1970
rect 8116 1906 8168 1912
rect 8022 1864 8078 1873
rect 7564 1828 7616 1834
rect 8022 1799 8024 1808
rect 7564 1770 7616 1776
rect 8076 1799 8078 1808
rect 8024 1770 8076 1776
rect 6918 1728 6974 1737
rect 6918 1663 6974 1672
rect 7566 1660 7874 1680
rect 7566 1658 7572 1660
rect 7628 1658 7652 1660
rect 7708 1658 7732 1660
rect 7788 1658 7812 1660
rect 7868 1658 7874 1660
rect 7628 1606 7630 1658
rect 7810 1606 7812 1658
rect 7566 1604 7572 1606
rect 7628 1604 7652 1606
rect 7708 1604 7732 1606
rect 7788 1604 7812 1606
rect 7868 1604 7874 1606
rect 7566 1584 7874 1604
rect 8300 1352 8352 1358
rect 8300 1294 8352 1300
rect 6736 1216 6788 1222
rect 6736 1158 6788 1164
rect 7196 1216 7248 1222
rect 7196 1158 7248 1164
rect 7932 1216 7984 1222
rect 7932 1158 7984 1164
rect 7208 1018 7236 1158
rect 7196 1012 7248 1018
rect 7196 954 7248 960
rect 7944 950 7972 1158
rect 7932 944 7984 950
rect 7932 886 7984 892
rect 8312 882 8340 1294
rect 8404 1222 8432 2910
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8496 1222 8524 2790
rect 8588 2446 8616 4490
rect 8680 2854 8708 5578
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8772 3738 8800 4082
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8864 3534 8892 3878
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 8758 3224 8814 3233
rect 8758 3159 8814 3168
rect 8772 3126 8800 3159
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8864 2774 8892 3470
rect 8772 2746 8892 2774
rect 8666 2680 8722 2689
rect 8666 2615 8722 2624
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8680 1834 8708 2615
rect 8772 1970 8800 2746
rect 8852 2032 8904 2038
rect 8852 1974 8904 1980
rect 8760 1964 8812 1970
rect 8760 1906 8812 1912
rect 8864 1850 8892 1974
rect 8668 1828 8720 1834
rect 8668 1770 8720 1776
rect 8772 1822 8892 1850
rect 8772 1494 8800 1822
rect 8956 1494 8984 5714
rect 9048 5642 9076 6258
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 9140 5574 9168 6598
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9232 5234 9260 6054
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9036 3120 9088 3126
rect 9034 3088 9036 3097
rect 9088 3088 9090 3097
rect 9034 3023 9090 3032
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 8760 1488 8812 1494
rect 8760 1430 8812 1436
rect 8944 1488 8996 1494
rect 8944 1430 8996 1436
rect 8668 1420 8720 1426
rect 8668 1362 8720 1368
rect 8392 1216 8444 1222
rect 8392 1158 8444 1164
rect 8484 1216 8536 1222
rect 8484 1158 8536 1164
rect 8680 950 8708 1362
rect 8760 1352 8812 1358
rect 8944 1352 8996 1358
rect 8812 1312 8944 1340
rect 8760 1294 8812 1300
rect 8944 1294 8996 1300
rect 9048 1222 9076 2926
rect 9140 1358 9168 3334
rect 9232 2582 9260 3878
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9232 1834 9260 2382
rect 9220 1828 9272 1834
rect 9220 1770 9272 1776
rect 9128 1352 9180 1358
rect 9128 1294 9180 1300
rect 9036 1216 9088 1222
rect 9036 1158 9088 1164
rect 9220 1216 9272 1222
rect 9220 1158 9272 1164
rect 9048 1018 9076 1158
rect 9232 1057 9260 1158
rect 9218 1048 9274 1057
rect 9036 1012 9088 1018
rect 9218 983 9274 992
rect 9036 954 9088 960
rect 8668 944 8720 950
rect 8668 886 8720 892
rect 9324 882 9352 10406
rect 9600 10396 10198 10424
rect 9600 10305 9628 10396
rect 9586 10296 9642 10305
rect 9586 10231 9642 10240
rect 9678 9072 9734 9081
rect 9678 9007 9734 9016
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9416 3482 9444 7754
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5914 9536 6054
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9600 5409 9628 8774
rect 9692 7993 9720 9007
rect 9678 7984 9734 7993
rect 9678 7919 9734 7928
rect 10428 7449 10456 11086
rect 10414 7440 10470 7449
rect 10414 7375 10470 7384
rect 9586 5400 9642 5409
rect 9586 5335 9642 5344
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9600 3618 9628 4490
rect 9600 3590 9720 3618
rect 9416 3454 9628 3482
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9402 2136 9458 2145
rect 9508 2106 9536 2994
rect 9600 2417 9628 3454
rect 9586 2408 9642 2417
rect 9586 2343 9642 2352
rect 9402 2071 9458 2080
rect 9496 2100 9548 2106
rect 9416 1970 9444 2071
rect 9496 2042 9548 2048
rect 9404 1964 9456 1970
rect 9404 1906 9456 1912
rect 9692 921 9720 3590
rect 10048 2780 10100 2786
rect 10048 2722 10100 2728
rect 9956 2712 10008 2718
rect 9956 2654 10008 2660
rect 9968 1290 9996 2654
rect 10060 1329 10088 2722
rect 10520 1562 10548 12271
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10704 7857 10732 11018
rect 10690 7848 10746 7857
rect 10690 7783 10746 7792
rect 10888 7041 10916 11290
rect 10980 8362 11008 12452
rect 13818 11928 13874 11937
rect 13818 11863 13820 11872
rect 13872 11863 13874 11872
rect 16672 11892 16724 11898
rect 13820 11834 13872 11840
rect 16672 11834 16724 11840
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11060 10192 11112 10198
rect 11060 10134 11112 10140
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10874 7032 10930 7041
rect 10874 6967 10930 6976
rect 10966 4992 11022 5001
rect 10966 4927 11022 4936
rect 10508 1556 10560 1562
rect 10508 1498 10560 1504
rect 10046 1320 10102 1329
rect 9956 1284 10008 1290
rect 10046 1255 10102 1264
rect 9956 1226 10008 1232
rect 9678 912 9734 921
rect 8300 876 8352 882
rect 8300 818 8352 824
rect 9312 876 9364 882
rect 9678 847 9734 856
rect 9312 818 9364 824
rect 10976 760 11004 4927
rect 11072 1193 11100 10134
rect 11164 8673 11192 11154
rect 13818 11112 13874 11121
rect 13874 11070 13952 11098
rect 13818 11047 13874 11056
rect 13818 9480 13874 9489
rect 13818 9415 13874 9424
rect 11150 8664 11206 8673
rect 11150 8599 11206 8608
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11164 3126 11192 6938
rect 13450 4176 13506 4185
rect 13450 4111 13506 4120
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 13464 2689 13492 4111
rect 13542 3360 13598 3369
rect 13542 3295 13598 3304
rect 13450 2680 13506 2689
rect 13556 2650 13584 3295
rect 13832 3074 13860 9415
rect 13648 3046 13860 3074
rect 13648 2786 13676 3046
rect 13924 2854 13952 11070
rect 16578 10704 16634 10713
rect 16578 10639 16580 10648
rect 16632 10639 16634 10648
rect 16580 10610 16632 10616
rect 16684 7002 16712 11834
rect 20718 11520 20774 11529
rect 20718 11455 20774 11464
rect 20732 9194 20760 11455
rect 22098 9888 22154 9897
rect 22098 9823 22154 9832
rect 20640 9166 20760 9194
rect 16672 6996 16724 7002
rect 16672 6938 16724 6944
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 13636 2780 13688 2786
rect 13636 2722 13688 2728
rect 13450 2615 13506 2624
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 15212 2582 15240 4762
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16592 2961 16620 3946
rect 16684 3777 16712 4966
rect 20640 4826 20668 9166
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 16854 4584 16910 4593
rect 16854 4519 16910 4528
rect 16670 3768 16726 3777
rect 16670 3703 16726 3712
rect 16578 2952 16634 2961
rect 16578 2887 16634 2896
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 16762 2136 16818 2145
rect 16762 2071 16818 2080
rect 13818 1864 13874 1873
rect 13818 1799 13820 1808
rect 13872 1799 13874 1808
rect 13820 1770 13872 1776
rect 16578 1728 16634 1737
rect 16578 1663 16634 1672
rect 11058 1184 11114 1193
rect 11058 1119 11114 1128
rect 16592 950 16620 1663
rect 16672 1420 16724 1426
rect 16672 1362 16724 1368
rect 16580 944 16632 950
rect 16580 886 16632 892
rect 16684 760 16712 1362
rect 16776 1290 16804 2071
rect 16868 1834 16896 4519
rect 22112 2378 22140 9823
rect 22100 2372 22152 2378
rect 22100 2314 22152 2320
rect 16856 1828 16908 1834
rect 16856 1770 16908 1776
rect 16764 1284 16816 1290
rect 16764 1226 16816 1232
rect 3884 740 3936 746
rect 3884 682 3936 688
rect 5724 740 5776 746
rect 10976 732 16712 760
rect 5724 682 5776 688
rect 16684 513 16712 732
rect 16670 504 16726 513
rect 16670 439 16726 448
<< via2 >>
rect 754 9560 810 9616
rect 938 9424 994 9480
rect 1398 9016 1454 9072
rect 1214 7520 1270 7576
rect 846 6432 902 6488
rect 1582 8472 1638 8528
rect 2134 10648 2190 10704
rect 2226 10104 2282 10160
rect 2226 8916 2228 8936
rect 2228 8916 2280 8936
rect 2280 8916 2282 8936
rect 2226 8880 2282 8916
rect 2134 8780 2136 8800
rect 2136 8780 2188 8800
rect 2188 8780 2190 8800
rect 2134 8744 2190 8780
rect 2042 8608 2098 8664
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2594 10784 2650 10840
rect 2778 10512 2834 10568
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2962 10240 3018 10296
rect 3054 10104 3110 10160
rect 2870 9832 2926 9888
rect 2778 9696 2834 9752
rect 2870 9560 2926 9616
rect 2778 9444 2834 9480
rect 2778 9424 2780 9444
rect 2780 9424 2832 9444
rect 2832 9424 2834 9444
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2502 8880 2558 8936
rect 2686 8880 2742 8936
rect 2778 8628 2834 8664
rect 2778 8608 2780 8628
rect 2780 8608 2832 8628
rect 2832 8608 2834 8628
rect 2042 8336 2098 8392
rect 1950 8064 2006 8120
rect 1858 7928 1914 7984
rect 1582 6316 1638 6352
rect 1582 6296 1584 6316
rect 1584 6296 1636 6316
rect 1636 6296 1638 6316
rect 1766 5752 1822 5808
rect 2318 8064 2374 8120
rect 3514 10648 3570 10704
rect 3606 10376 3662 10432
rect 3330 9696 3386 9752
rect 2962 8472 3018 8528
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2410 7404 2466 7440
rect 2410 7384 2412 7404
rect 2412 7384 2464 7404
rect 2464 7384 2466 7404
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 2502 6568 2558 6624
rect 2134 6180 2190 6216
rect 2134 6160 2136 6180
rect 2136 6160 2188 6180
rect 2188 6160 2190 6180
rect 2870 6840 2926 6896
rect 1582 4664 1638 4720
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 2778 5616 2834 5672
rect 2502 1808 2558 1864
rect 3330 8880 3386 8936
rect 3422 8744 3478 8800
rect 3330 7928 3386 7984
rect 3330 7656 3386 7712
rect 3882 11056 3938 11112
rect 3882 10512 3938 10568
rect 4066 11056 4122 11112
rect 4250 10784 4306 10840
rect 4158 9968 4214 10024
rect 4342 10648 4398 10704
rect 4342 9968 4398 10024
rect 3882 7656 3938 7712
rect 3238 5344 3294 5400
rect 3514 5888 3570 5944
rect 3606 5616 3662 5672
rect 3514 3304 3570 3360
rect 3606 2896 3662 2952
rect 3606 1672 3662 1728
rect 3882 7520 3938 7576
rect 3974 6432 4030 6488
rect 3974 5616 4030 5672
rect 4158 8880 4214 8936
rect 4250 3440 4306 3496
rect 4526 8064 4582 8120
rect 4710 10512 4766 10568
rect 4710 9424 4766 9480
rect 5072 10906 5128 10908
rect 5152 10906 5208 10908
rect 5232 10906 5288 10908
rect 5312 10906 5368 10908
rect 5072 10854 5118 10906
rect 5118 10854 5128 10906
rect 5152 10854 5182 10906
rect 5182 10854 5194 10906
rect 5194 10854 5208 10906
rect 5232 10854 5246 10906
rect 5246 10854 5258 10906
rect 5258 10854 5288 10906
rect 5312 10854 5322 10906
rect 5322 10854 5368 10906
rect 5072 10852 5128 10854
rect 5152 10852 5208 10854
rect 5232 10852 5288 10854
rect 5312 10852 5368 10854
rect 4986 10512 5042 10568
rect 5262 10512 5318 10568
rect 5170 9968 5226 10024
rect 5630 10240 5686 10296
rect 5072 9818 5128 9820
rect 5152 9818 5208 9820
rect 5232 9818 5288 9820
rect 5312 9818 5368 9820
rect 5072 9766 5118 9818
rect 5118 9766 5128 9818
rect 5152 9766 5182 9818
rect 5182 9766 5194 9818
rect 5194 9766 5208 9818
rect 5232 9766 5246 9818
rect 5246 9766 5258 9818
rect 5258 9766 5288 9818
rect 5312 9766 5322 9818
rect 5322 9766 5368 9818
rect 5072 9764 5128 9766
rect 5152 9764 5208 9766
rect 5232 9764 5288 9766
rect 5312 9764 5368 9766
rect 5078 9632 5134 9688
rect 5722 9832 5778 9888
rect 4986 9152 5042 9208
rect 5354 9580 5410 9616
rect 5354 9560 5356 9580
rect 5356 9560 5408 9580
rect 5408 9560 5410 9580
rect 5722 9460 5724 9480
rect 5724 9460 5776 9480
rect 5776 9460 5778 9480
rect 4802 8200 4858 8256
rect 5072 8730 5128 8732
rect 5152 8730 5208 8732
rect 5232 8730 5288 8732
rect 5312 8730 5368 8732
rect 5072 8678 5118 8730
rect 5118 8678 5128 8730
rect 5152 8678 5182 8730
rect 5182 8678 5194 8730
rect 5194 8678 5208 8730
rect 5232 8678 5246 8730
rect 5246 8678 5258 8730
rect 5258 8678 5288 8730
rect 5312 8678 5322 8730
rect 5322 8678 5368 8730
rect 5072 8676 5128 8678
rect 5152 8676 5208 8678
rect 5232 8676 5288 8678
rect 5312 8676 5368 8678
rect 5722 9424 5778 9460
rect 4894 6976 4950 7032
rect 5354 7792 5410 7848
rect 5072 7642 5128 7644
rect 5152 7642 5208 7644
rect 5232 7642 5288 7644
rect 5312 7642 5368 7644
rect 5072 7590 5118 7642
rect 5118 7590 5128 7642
rect 5152 7590 5182 7642
rect 5182 7590 5194 7642
rect 5194 7590 5208 7642
rect 5232 7590 5246 7642
rect 5246 7590 5258 7642
rect 5258 7590 5288 7642
rect 5312 7590 5322 7642
rect 5322 7590 5368 7642
rect 5072 7588 5128 7590
rect 5152 7588 5208 7590
rect 5232 7588 5288 7590
rect 5312 7588 5368 7590
rect 5630 7928 5686 7984
rect 5630 7656 5686 7712
rect 5538 7384 5594 7440
rect 5446 6976 5502 7032
rect 4802 5344 4858 5400
rect 4618 4120 4674 4176
rect 4434 2760 4490 2816
rect 4434 2352 4490 2408
rect 4618 3032 4674 3088
rect 5072 6554 5128 6556
rect 5152 6554 5208 6556
rect 5232 6554 5288 6556
rect 5312 6554 5368 6556
rect 5072 6502 5118 6554
rect 5118 6502 5128 6554
rect 5152 6502 5182 6554
rect 5182 6502 5194 6554
rect 5194 6502 5208 6554
rect 5232 6502 5246 6554
rect 5246 6502 5258 6554
rect 5258 6502 5288 6554
rect 5312 6502 5322 6554
rect 5322 6502 5368 6554
rect 5072 6500 5128 6502
rect 5152 6500 5208 6502
rect 5232 6500 5288 6502
rect 5312 6500 5368 6502
rect 5170 5636 5226 5672
rect 5170 5616 5172 5636
rect 5172 5616 5224 5636
rect 5224 5616 5226 5636
rect 5072 5466 5128 5468
rect 5152 5466 5208 5468
rect 5232 5466 5288 5468
rect 5312 5466 5368 5468
rect 5072 5414 5118 5466
rect 5118 5414 5128 5466
rect 5152 5414 5182 5466
rect 5182 5414 5194 5466
rect 5194 5414 5208 5466
rect 5232 5414 5246 5466
rect 5246 5414 5258 5466
rect 5258 5414 5288 5466
rect 5312 5414 5322 5466
rect 5322 5414 5368 5466
rect 5072 5412 5128 5414
rect 5152 5412 5208 5414
rect 5232 5412 5288 5414
rect 5312 5412 5368 5414
rect 5170 4528 5226 4584
rect 6090 10804 6146 10840
rect 6090 10784 6092 10804
rect 6092 10784 6144 10804
rect 6144 10784 6146 10804
rect 5906 10104 5962 10160
rect 5906 9696 5962 9752
rect 5998 9152 6054 9208
rect 5538 5908 5594 5944
rect 5538 5888 5540 5908
rect 5540 5888 5592 5908
rect 5592 5888 5594 5908
rect 5446 4528 5502 4584
rect 5072 4378 5128 4380
rect 5152 4378 5208 4380
rect 5232 4378 5288 4380
rect 5312 4378 5368 4380
rect 5072 4326 5118 4378
rect 5118 4326 5128 4378
rect 5152 4326 5182 4378
rect 5182 4326 5194 4378
rect 5194 4326 5208 4378
rect 5232 4326 5246 4378
rect 5246 4326 5258 4378
rect 5258 4326 5288 4378
rect 5312 4326 5322 4378
rect 5322 4326 5368 4378
rect 5072 4324 5128 4326
rect 5152 4324 5208 4326
rect 5232 4324 5288 4326
rect 5312 4324 5368 4326
rect 4986 4120 5042 4176
rect 5446 4120 5502 4176
rect 4894 2760 4950 2816
rect 5072 3290 5128 3292
rect 5152 3290 5208 3292
rect 5232 3290 5288 3292
rect 5312 3290 5368 3292
rect 5072 3238 5118 3290
rect 5118 3238 5128 3290
rect 5152 3238 5182 3290
rect 5182 3238 5194 3290
rect 5194 3238 5208 3290
rect 5232 3238 5246 3290
rect 5246 3238 5258 3290
rect 5258 3238 5288 3290
rect 5312 3238 5322 3290
rect 5322 3238 5368 3290
rect 5072 3236 5128 3238
rect 5152 3236 5208 3238
rect 5232 3236 5288 3238
rect 5312 3236 5368 3238
rect 5814 6160 5870 6216
rect 5998 8336 6054 8392
rect 5998 7812 6054 7848
rect 5998 7792 6000 7812
rect 6000 7792 6052 7812
rect 6052 7792 6054 7812
rect 6274 9152 6330 9208
rect 6366 9016 6422 9072
rect 5906 5888 5962 5944
rect 5630 4120 5686 4176
rect 5538 2760 5594 2816
rect 5072 2202 5128 2204
rect 5152 2202 5208 2204
rect 5232 2202 5288 2204
rect 5312 2202 5368 2204
rect 5072 2150 5118 2202
rect 5118 2150 5128 2202
rect 5152 2150 5182 2202
rect 5182 2150 5194 2202
rect 5194 2150 5208 2202
rect 5232 2150 5246 2202
rect 5246 2150 5258 2202
rect 5258 2150 5288 2202
rect 5312 2150 5322 2202
rect 5322 2150 5368 2202
rect 5072 2148 5128 2150
rect 5152 2148 5208 2150
rect 5232 2148 5288 2150
rect 5312 2148 5368 2150
rect 5170 1944 5226 2000
rect 5538 1808 5594 1864
rect 4986 1264 5042 1320
rect 6090 6160 6146 6216
rect 5998 4256 6054 4312
rect 6826 10784 6882 10840
rect 6734 9968 6790 10024
rect 6734 6432 6790 6488
rect 6550 4392 6606 4448
rect 6550 2896 6606 2952
rect 6274 2080 6330 2136
rect 6826 4392 6882 4448
rect 5446 1128 5502 1184
rect 5072 1114 5128 1116
rect 5152 1114 5208 1116
rect 5232 1114 5288 1116
rect 5312 1114 5368 1116
rect 5072 1062 5118 1114
rect 5118 1062 5128 1114
rect 5152 1062 5182 1114
rect 5182 1062 5194 1114
rect 5194 1062 5208 1114
rect 5232 1062 5246 1114
rect 5246 1062 5258 1114
rect 5258 1062 5288 1114
rect 5312 1062 5322 1114
rect 5322 1062 5368 1114
rect 5072 1060 5128 1062
rect 5152 1060 5208 1062
rect 5232 1060 5288 1062
rect 5312 1060 5368 1062
rect 6826 1944 6882 2000
rect 7572 11450 7628 11452
rect 7652 11450 7708 11452
rect 7732 11450 7788 11452
rect 7812 11450 7868 11452
rect 7572 11398 7618 11450
rect 7618 11398 7628 11450
rect 7652 11398 7682 11450
rect 7682 11398 7694 11450
rect 7694 11398 7708 11450
rect 7732 11398 7746 11450
rect 7746 11398 7758 11450
rect 7758 11398 7788 11450
rect 7812 11398 7822 11450
rect 7822 11398 7868 11450
rect 7572 11396 7628 11398
rect 7652 11396 7708 11398
rect 7732 11396 7788 11398
rect 7812 11396 7868 11398
rect 7378 11092 7380 11112
rect 7380 11092 7432 11112
rect 7432 11092 7434 11112
rect 7378 11056 7434 11092
rect 7194 9832 7250 9888
rect 7378 10376 7434 10432
rect 7286 9288 7342 9344
rect 7194 6296 7250 6352
rect 7572 10362 7628 10364
rect 7652 10362 7708 10364
rect 7732 10362 7788 10364
rect 7812 10362 7868 10364
rect 7572 10310 7618 10362
rect 7618 10310 7628 10362
rect 7652 10310 7682 10362
rect 7682 10310 7694 10362
rect 7694 10310 7708 10362
rect 7732 10310 7746 10362
rect 7746 10310 7758 10362
rect 7758 10310 7788 10362
rect 7812 10310 7822 10362
rect 7822 10310 7868 10362
rect 7572 10308 7628 10310
rect 7652 10308 7708 10310
rect 7732 10308 7788 10310
rect 7812 10308 7868 10310
rect 7654 10004 7656 10024
rect 7656 10004 7708 10024
rect 7708 10004 7710 10024
rect 7654 9968 7710 10004
rect 7572 9274 7628 9276
rect 7652 9274 7708 9276
rect 7732 9274 7788 9276
rect 7812 9274 7868 9276
rect 7572 9222 7618 9274
rect 7618 9222 7628 9274
rect 7652 9222 7682 9274
rect 7682 9222 7694 9274
rect 7694 9222 7708 9274
rect 7732 9222 7746 9274
rect 7746 9222 7758 9274
rect 7758 9222 7788 9274
rect 7812 9222 7822 9274
rect 7822 9222 7868 9274
rect 7572 9220 7628 9222
rect 7652 9220 7708 9222
rect 7732 9220 7788 9222
rect 7812 9220 7868 9222
rect 7562 9016 7618 9072
rect 7572 8186 7628 8188
rect 7652 8186 7708 8188
rect 7732 8186 7788 8188
rect 7812 8186 7868 8188
rect 7572 8134 7618 8186
rect 7618 8134 7628 8186
rect 7652 8134 7682 8186
rect 7682 8134 7694 8186
rect 7694 8134 7708 8186
rect 7732 8134 7746 8186
rect 7746 8134 7758 8186
rect 7758 8134 7788 8186
rect 7812 8134 7822 8186
rect 7822 8134 7868 8186
rect 7572 8132 7628 8134
rect 7652 8132 7708 8134
rect 7732 8132 7788 8134
rect 7812 8132 7868 8134
rect 8114 9152 8170 9208
rect 7572 7098 7628 7100
rect 7652 7098 7708 7100
rect 7732 7098 7788 7100
rect 7812 7098 7868 7100
rect 7572 7046 7618 7098
rect 7618 7046 7628 7098
rect 7652 7046 7682 7098
rect 7682 7046 7694 7098
rect 7694 7046 7708 7098
rect 7732 7046 7746 7098
rect 7746 7046 7758 7098
rect 7758 7046 7788 7098
rect 7812 7046 7822 7098
rect 7822 7046 7868 7098
rect 7572 7044 7628 7046
rect 7652 7044 7708 7046
rect 7732 7044 7788 7046
rect 7812 7044 7868 7046
rect 7378 5752 7434 5808
rect 7572 6010 7628 6012
rect 7652 6010 7708 6012
rect 7732 6010 7788 6012
rect 7812 6010 7868 6012
rect 7572 5958 7618 6010
rect 7618 5958 7628 6010
rect 7652 5958 7682 6010
rect 7682 5958 7694 6010
rect 7694 5958 7708 6010
rect 7732 5958 7746 6010
rect 7746 5958 7758 6010
rect 7758 5958 7788 6010
rect 7812 5958 7822 6010
rect 7822 5958 7868 6010
rect 7572 5956 7628 5958
rect 7652 5956 7708 5958
rect 7732 5956 7788 5958
rect 7812 5956 7868 5958
rect 8022 6160 8078 6216
rect 8022 5752 8078 5808
rect 7572 4922 7628 4924
rect 7652 4922 7708 4924
rect 7732 4922 7788 4924
rect 7812 4922 7868 4924
rect 7572 4870 7618 4922
rect 7618 4870 7628 4922
rect 7652 4870 7682 4922
rect 7682 4870 7694 4922
rect 7694 4870 7708 4922
rect 7732 4870 7746 4922
rect 7746 4870 7758 4922
rect 7758 4870 7788 4922
rect 7812 4870 7822 4922
rect 7822 4870 7868 4922
rect 7572 4868 7628 4870
rect 7652 4868 7708 4870
rect 7732 4868 7788 4870
rect 7812 4868 7868 4870
rect 7378 4664 7434 4720
rect 7378 3168 7434 3224
rect 7572 3834 7628 3836
rect 7652 3834 7708 3836
rect 7732 3834 7788 3836
rect 7812 3834 7868 3836
rect 7572 3782 7618 3834
rect 7618 3782 7628 3834
rect 7652 3782 7682 3834
rect 7682 3782 7694 3834
rect 7694 3782 7708 3834
rect 7732 3782 7746 3834
rect 7746 3782 7758 3834
rect 7758 3782 7788 3834
rect 7812 3782 7822 3834
rect 7822 3782 7868 3834
rect 7572 3780 7628 3782
rect 7652 3780 7708 3782
rect 7732 3780 7788 3782
rect 7812 3780 7868 3782
rect 7378 2760 7434 2816
rect 7572 2746 7628 2748
rect 7652 2746 7708 2748
rect 7732 2746 7788 2748
rect 7812 2746 7868 2748
rect 7572 2694 7618 2746
rect 7618 2694 7628 2746
rect 7652 2694 7682 2746
rect 7682 2694 7694 2746
rect 7694 2694 7708 2746
rect 7732 2694 7746 2746
rect 7746 2694 7758 2746
rect 7758 2694 7788 2746
rect 7812 2694 7822 2746
rect 7822 2694 7868 2746
rect 7572 2692 7628 2694
rect 7652 2692 7708 2694
rect 7732 2692 7788 2694
rect 7812 2692 7868 2694
rect 7930 2508 7986 2544
rect 7930 2488 7932 2508
rect 7932 2488 7984 2508
rect 7984 2488 7986 2508
rect 8298 7792 8354 7848
rect 8850 8336 8906 8392
rect 10506 12280 10562 12336
rect 8206 5636 8262 5672
rect 8206 5616 8208 5636
rect 8208 5616 8260 5636
rect 8260 5616 8262 5636
rect 8942 6840 8998 6896
rect 8114 3440 8170 3496
rect 8206 2488 8262 2544
rect 8022 1828 8078 1864
rect 8022 1808 8024 1828
rect 8024 1808 8076 1828
rect 8076 1808 8078 1828
rect 6918 1672 6974 1728
rect 7572 1658 7628 1660
rect 7652 1658 7708 1660
rect 7732 1658 7788 1660
rect 7812 1658 7868 1660
rect 7572 1606 7618 1658
rect 7618 1606 7628 1658
rect 7652 1606 7682 1658
rect 7682 1606 7694 1658
rect 7694 1606 7708 1658
rect 7732 1606 7746 1658
rect 7746 1606 7758 1658
rect 7758 1606 7788 1658
rect 7812 1606 7822 1658
rect 7822 1606 7868 1658
rect 7572 1604 7628 1606
rect 7652 1604 7708 1606
rect 7732 1604 7788 1606
rect 7812 1604 7868 1606
rect 8758 3168 8814 3224
rect 8666 2624 8722 2680
rect 9034 3068 9036 3088
rect 9036 3068 9088 3088
rect 9088 3068 9090 3088
rect 9034 3032 9090 3068
rect 9218 992 9274 1048
rect 9586 10240 9642 10296
rect 9678 9016 9734 9072
rect 9678 7928 9734 7984
rect 10414 7384 10470 7440
rect 9586 5344 9642 5400
rect 9402 2080 9458 2136
rect 9586 2352 9642 2408
rect 10690 7792 10746 7848
rect 13818 11892 13874 11928
rect 13818 11872 13820 11892
rect 13820 11872 13872 11892
rect 13872 11872 13874 11892
rect 10874 6976 10930 7032
rect 10966 4936 11022 4992
rect 10046 1264 10102 1320
rect 9678 856 9734 912
rect 13818 11056 13874 11112
rect 13818 9424 13874 9480
rect 11150 8608 11206 8664
rect 13450 4120 13506 4176
rect 13542 3304 13598 3360
rect 13450 2624 13506 2680
rect 16578 10668 16634 10704
rect 16578 10648 16580 10668
rect 16580 10648 16632 10668
rect 16632 10648 16634 10668
rect 20718 11464 20774 11520
rect 22098 9832 22154 9888
rect 16854 4528 16910 4584
rect 16670 3712 16726 3768
rect 16578 2896 16634 2952
rect 16762 2080 16818 2136
rect 13818 1828 13874 1864
rect 13818 1808 13820 1828
rect 13820 1808 13872 1828
rect 13872 1808 13874 1828
rect 16578 1672 16634 1728
rect 11058 1128 11114 1184
rect 16670 448 16726 504
<< metal3 >>
rect 10501 12338 10567 12341
rect 14000 12338 34000 12368
rect 10501 12336 34000 12338
rect 10501 12280 10506 12336
rect 10562 12280 34000 12336
rect 10501 12278 34000 12280
rect 10501 12275 10567 12278
rect 14000 12248 34000 12278
rect 13813 11930 13879 11933
rect 14000 11930 34000 11960
rect 13813 11928 34000 11930
rect 13813 11872 13818 11928
rect 13874 11872 34000 11928
rect 13813 11870 34000 11872
rect 13813 11867 13879 11870
rect 14000 11840 34000 11870
rect 14000 11520 34000 11552
rect 14000 11464 20718 11520
rect 20774 11464 34000 11520
rect 2560 11456 2880 11457
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 11391 2880 11392
rect 7560 11456 7880 11457
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 14000 11432 34000 11464
rect 7560 11391 7880 11392
rect 3877 11114 3943 11117
rect 4061 11114 4127 11117
rect 7373 11114 7439 11117
rect 3877 11112 7439 11114
rect 3877 11056 3882 11112
rect 3938 11056 4066 11112
rect 4122 11056 7378 11112
rect 7434 11056 7439 11112
rect 3877 11054 7439 11056
rect 3877 11051 3943 11054
rect 4061 11051 4127 11054
rect 7373 11051 7439 11054
rect 13813 11114 13879 11117
rect 14000 11114 34000 11144
rect 13813 11112 34000 11114
rect 13813 11056 13818 11112
rect 13874 11056 34000 11112
rect 13813 11054 34000 11056
rect 13813 11051 13879 11054
rect 14000 11024 34000 11054
rect 5060 10912 5380 10913
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 10847 5380 10848
rect 2589 10842 2655 10845
rect 4245 10842 4311 10845
rect 2589 10840 4311 10842
rect 2589 10784 2594 10840
rect 2650 10784 4250 10840
rect 4306 10784 4311 10840
rect 2589 10782 4311 10784
rect 2589 10779 2655 10782
rect 4245 10779 4311 10782
rect 6085 10842 6151 10845
rect 6821 10842 6887 10845
rect 6085 10840 6887 10842
rect 6085 10784 6090 10840
rect 6146 10784 6826 10840
rect 6882 10784 6887 10840
rect 6085 10782 6887 10784
rect 6085 10779 6151 10782
rect 6821 10779 6887 10782
rect 2129 10706 2195 10709
rect 3509 10706 3575 10709
rect 2129 10704 3575 10706
rect 2129 10648 2134 10704
rect 2190 10648 3514 10704
rect 3570 10648 3575 10704
rect 2129 10646 3575 10648
rect 2129 10643 2195 10646
rect 3509 10643 3575 10646
rect 4337 10706 4403 10709
rect 4337 10704 4722 10706
rect 4337 10648 4342 10704
rect 4398 10648 4722 10704
rect 4337 10646 4722 10648
rect 4337 10643 4403 10646
rect 4662 10573 4722 10646
rect 14000 10704 34000 10736
rect 14000 10648 16578 10704
rect 16634 10648 34000 10704
rect 14000 10616 34000 10648
rect 2773 10570 2839 10573
rect 3877 10570 3943 10573
rect 2773 10568 3943 10570
rect 2773 10512 2778 10568
rect 2834 10512 3882 10568
rect 3938 10512 3943 10568
rect 2773 10510 3943 10512
rect 4662 10568 4771 10573
rect 4662 10512 4710 10568
rect 4766 10512 4771 10568
rect 4662 10510 4771 10512
rect 2773 10507 2839 10510
rect 3877 10507 3943 10510
rect 4705 10507 4771 10510
rect 4981 10570 5047 10573
rect 5257 10570 5323 10573
rect 4981 10568 5323 10570
rect 4981 10512 4986 10568
rect 5042 10512 5262 10568
rect 5318 10512 5323 10568
rect 4981 10510 5323 10512
rect 4981 10507 5047 10510
rect 5257 10507 5323 10510
rect 3601 10434 3667 10437
rect 7373 10434 7439 10437
rect 3601 10432 7439 10434
rect 3601 10376 3606 10432
rect 3662 10376 7378 10432
rect 7434 10376 7439 10432
rect 3601 10374 7439 10376
rect 3601 10371 3667 10374
rect 7373 10371 7439 10374
rect 2560 10368 2880 10369
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 10303 2880 10304
rect 7560 10368 7880 10369
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 10303 7880 10304
rect 2957 10298 3023 10301
rect 5625 10298 5691 10301
rect 2957 10296 5691 10298
rect 2957 10240 2962 10296
rect 3018 10240 5630 10296
rect 5686 10240 5691 10296
rect 2957 10238 5691 10240
rect 2957 10235 3023 10238
rect 5625 10235 5691 10238
rect 9581 10298 9647 10301
rect 14000 10298 34000 10328
rect 9581 10296 34000 10298
rect 9581 10240 9586 10296
rect 9642 10240 34000 10296
rect 9581 10238 34000 10240
rect 9581 10235 9647 10238
rect 14000 10208 34000 10238
rect 2221 10162 2287 10165
rect 3049 10162 3115 10165
rect 5901 10162 5967 10165
rect 2221 10160 3115 10162
rect 2221 10104 2226 10160
rect 2282 10104 3054 10160
rect 3110 10104 3115 10160
rect 2221 10102 3115 10104
rect 2221 10099 2287 10102
rect 3049 10099 3115 10102
rect 3190 10160 5967 10162
rect 3190 10104 5906 10160
rect 5962 10104 5967 10160
rect 3190 10102 5967 10104
rect 2865 9890 2931 9893
rect 3190 9890 3250 10102
rect 5901 10099 5967 10102
rect 4153 10026 4219 10029
rect 4337 10026 4403 10029
rect 5165 10026 5231 10029
rect 4153 10024 4403 10026
rect 4153 9968 4158 10024
rect 4214 9968 4342 10024
rect 4398 9968 4403 10024
rect 4153 9966 4403 9968
rect 4153 9963 4219 9966
rect 4337 9963 4403 9966
rect 4846 10024 5231 10026
rect 4846 9968 5170 10024
rect 5226 9968 5231 10024
rect 4846 9966 5231 9968
rect 2865 9888 3250 9890
rect 2865 9832 2870 9888
rect 2926 9832 3250 9888
rect 2865 9830 3250 9832
rect 2865 9827 2931 9830
rect 2773 9754 2839 9757
rect 3325 9754 3391 9757
rect 2773 9752 3391 9754
rect 2773 9696 2778 9752
rect 2834 9696 3330 9752
rect 3386 9696 3391 9752
rect 2773 9694 3391 9696
rect 2773 9691 2839 9694
rect 3325 9691 3391 9694
rect 4846 9690 4906 9966
rect 5165 9963 5231 9966
rect 6729 10026 6795 10029
rect 7649 10026 7715 10029
rect 6729 10024 7715 10026
rect 6729 9968 6734 10024
rect 6790 9968 7654 10024
rect 7710 9968 7715 10024
rect 6729 9966 7715 9968
rect 6729 9963 6795 9966
rect 7649 9963 7715 9966
rect 5717 9890 5783 9893
rect 7189 9890 7255 9893
rect 5717 9888 7255 9890
rect 5717 9832 5722 9888
rect 5778 9832 7194 9888
rect 7250 9832 7255 9888
rect 5717 9830 7255 9832
rect 5717 9827 5783 9830
rect 7189 9827 7255 9830
rect 14000 9888 34000 9920
rect 14000 9832 22098 9888
rect 22154 9832 34000 9888
rect 5060 9824 5380 9825
rect 5060 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5228 9824
rect 5292 9760 5308 9824
rect 5372 9760 5380 9824
rect 14000 9800 34000 9832
rect 5060 9759 5380 9760
rect 5901 9754 5967 9757
rect 5766 9752 5967 9754
rect 5766 9696 5906 9752
rect 5962 9696 5967 9752
rect 5766 9694 5967 9696
rect 5073 9690 5139 9693
rect 4846 9688 5139 9690
rect 4846 9632 5078 9688
rect 5134 9632 5139 9688
rect 4846 9630 5139 9632
rect 5073 9627 5139 9630
rect 749 9618 815 9621
rect 2865 9618 2931 9621
rect 749 9616 2931 9618
rect 749 9560 754 9616
rect 810 9560 2870 9616
rect 2926 9560 2931 9616
rect 749 9558 2931 9560
rect 749 9555 815 9558
rect 2865 9555 2931 9558
rect 5349 9618 5415 9621
rect 5766 9618 5826 9694
rect 5901 9691 5967 9694
rect 5349 9616 5826 9618
rect 5349 9560 5354 9616
rect 5410 9560 5826 9616
rect 5349 9558 5826 9560
rect 5349 9555 5415 9558
rect 933 9482 999 9485
rect 2773 9482 2839 9485
rect 933 9480 2839 9482
rect 933 9424 938 9480
rect 994 9424 2778 9480
rect 2834 9424 2839 9480
rect 933 9422 2839 9424
rect 933 9419 999 9422
rect 2773 9419 2839 9422
rect 4705 9482 4771 9485
rect 5717 9482 5783 9485
rect 4705 9480 5783 9482
rect 4705 9424 4710 9480
rect 4766 9424 5722 9480
rect 5778 9424 5783 9480
rect 4705 9422 5783 9424
rect 4705 9419 4771 9422
rect 5717 9419 5783 9422
rect 13813 9482 13879 9485
rect 14000 9482 34000 9512
rect 13813 9480 34000 9482
rect 13813 9424 13818 9480
rect 13874 9424 34000 9480
rect 13813 9422 34000 9424
rect 13813 9419 13879 9422
rect 5720 9346 5780 9419
rect 14000 9392 34000 9422
rect 7281 9346 7347 9349
rect 5720 9344 7347 9346
rect 5720 9288 7286 9344
rect 7342 9288 7347 9344
rect 5720 9286 7347 9288
rect 7281 9283 7347 9286
rect 2560 9280 2880 9281
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9215 2880 9216
rect 7560 9280 7880 9281
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 9215 7880 9216
rect 4981 9210 5047 9213
rect 3006 9208 5047 9210
rect 3006 9152 4986 9208
rect 5042 9152 5047 9208
rect 3006 9150 5047 9152
rect 1393 9074 1459 9077
rect 3006 9074 3066 9150
rect 4981 9147 5047 9150
rect 5993 9210 6059 9213
rect 6269 9210 6335 9213
rect 5993 9208 6335 9210
rect 5993 9152 5998 9208
rect 6054 9152 6274 9208
rect 6330 9152 6335 9208
rect 5993 9150 6335 9152
rect 5993 9147 6059 9150
rect 6269 9147 6335 9150
rect 8109 9208 8175 9213
rect 8109 9152 8114 9208
rect 8170 9152 8175 9208
rect 8109 9147 8175 9152
rect 1393 9072 3066 9074
rect 1393 9016 1398 9072
rect 1454 9016 3066 9072
rect 1393 9014 3066 9016
rect 6361 9074 6427 9077
rect 7557 9074 7623 9077
rect 6361 9072 7623 9074
rect 6361 9016 6366 9072
rect 6422 9016 7562 9072
rect 7618 9016 7623 9072
rect 6361 9014 7623 9016
rect 1393 9011 1459 9014
rect 6361 9011 6427 9014
rect 7557 9011 7623 9014
rect 2221 8938 2287 8941
rect 2497 8938 2563 8941
rect 2221 8936 2563 8938
rect 2221 8880 2226 8936
rect 2282 8880 2502 8936
rect 2558 8880 2563 8936
rect 2221 8878 2563 8880
rect 2221 8875 2287 8878
rect 2497 8875 2563 8878
rect 2681 8938 2747 8941
rect 3325 8938 3391 8941
rect 2681 8936 3391 8938
rect 2681 8880 2686 8936
rect 2742 8880 3330 8936
rect 3386 8880 3391 8936
rect 2681 8878 3391 8880
rect 2681 8875 2747 8878
rect 3325 8875 3391 8878
rect 4153 8938 4219 8941
rect 8112 8938 8172 9147
rect 9673 9074 9739 9077
rect 14000 9074 34000 9104
rect 9673 9072 34000 9074
rect 9673 9016 9678 9072
rect 9734 9016 34000 9072
rect 9673 9014 34000 9016
rect 9673 9011 9739 9014
rect 14000 8984 34000 9014
rect 4153 8936 8172 8938
rect 4153 8880 4158 8936
rect 4214 8880 8172 8936
rect 4153 8878 8172 8880
rect 4153 8875 4219 8878
rect 2129 8802 2195 8805
rect 3417 8802 3483 8805
rect 2129 8800 3483 8802
rect 2129 8744 2134 8800
rect 2190 8744 3422 8800
rect 3478 8744 3483 8800
rect 2129 8742 3483 8744
rect 2129 8739 2195 8742
rect 3417 8739 3483 8742
rect 5060 8736 5380 8737
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 8671 5380 8672
rect 2037 8666 2103 8669
rect 2773 8666 2839 8669
rect 2037 8664 2839 8666
rect 2037 8608 2042 8664
rect 2098 8608 2778 8664
rect 2834 8608 2839 8664
rect 2037 8606 2839 8608
rect 2037 8603 2103 8606
rect 2773 8603 2839 8606
rect 11145 8666 11211 8669
rect 14000 8666 34000 8696
rect 11145 8664 34000 8666
rect 11145 8608 11150 8664
rect 11206 8608 34000 8664
rect 11145 8606 34000 8608
rect 11145 8603 11211 8606
rect 14000 8576 34000 8606
rect 1577 8530 1643 8533
rect 2957 8530 3023 8533
rect 1577 8528 3023 8530
rect 1577 8472 1582 8528
rect 1638 8472 2962 8528
rect 3018 8472 3023 8528
rect 1577 8470 3023 8472
rect 1577 8467 1643 8470
rect 2957 8467 3023 8470
rect 2037 8394 2103 8397
rect 5993 8394 6059 8397
rect 2037 8392 6059 8394
rect 2037 8336 2042 8392
rect 2098 8336 5998 8392
rect 6054 8336 6059 8392
rect 2037 8334 6059 8336
rect 2037 8331 2103 8334
rect 5993 8331 6059 8334
rect 8845 8394 8911 8397
rect 8845 8392 13922 8394
rect 8845 8336 8850 8392
rect 8906 8336 13922 8392
rect 8845 8334 13922 8336
rect 8845 8331 8911 8334
rect 4797 8258 4863 8261
rect 4524 8256 4863 8258
rect 4524 8200 4802 8256
rect 4858 8200 4863 8256
rect 4524 8198 4863 8200
rect 13862 8258 13922 8334
rect 14000 8258 34000 8288
rect 13862 8198 34000 8258
rect 2560 8192 2880 8193
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 8127 2880 8128
rect 4524 8125 4584 8198
rect 4797 8195 4863 8198
rect 7560 8192 7880 8193
rect 7560 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7880 8192
rect 14000 8168 34000 8198
rect 7560 8127 7880 8128
rect 1945 8122 2011 8125
rect 2313 8122 2379 8125
rect 1945 8120 2379 8122
rect 1945 8064 1950 8120
rect 2006 8064 2318 8120
rect 2374 8064 2379 8120
rect 1945 8062 2379 8064
rect 1945 8059 2011 8062
rect 2313 8059 2379 8062
rect 4521 8120 4587 8125
rect 4521 8064 4526 8120
rect 4582 8064 4587 8120
rect 4521 8059 4587 8064
rect 1853 7986 1919 7989
rect 3325 7986 3391 7989
rect 1853 7984 3391 7986
rect 1853 7928 1858 7984
rect 1914 7928 3330 7984
rect 3386 7928 3391 7984
rect 1853 7926 3391 7928
rect 1853 7923 1919 7926
rect 3325 7923 3391 7926
rect 5625 7986 5691 7989
rect 9673 7986 9739 7989
rect 5625 7984 9739 7986
rect 5625 7928 5630 7984
rect 5686 7928 9678 7984
rect 9734 7928 9739 7984
rect 5625 7926 9739 7928
rect 5625 7923 5691 7926
rect 9673 7923 9739 7926
rect 5349 7850 5415 7853
rect 5993 7850 6059 7853
rect 8293 7850 8359 7853
rect 5349 7848 5688 7850
rect 5349 7792 5354 7848
rect 5410 7792 5688 7848
rect 5349 7790 5688 7792
rect 5349 7787 5415 7790
rect 5628 7717 5688 7790
rect 5993 7848 8359 7850
rect 5993 7792 5998 7848
rect 6054 7792 8298 7848
rect 8354 7792 8359 7848
rect 5993 7790 8359 7792
rect 5993 7787 6059 7790
rect 8293 7787 8359 7790
rect 10685 7850 10751 7853
rect 14000 7850 34000 7880
rect 10685 7848 34000 7850
rect 10685 7792 10690 7848
rect 10746 7792 34000 7848
rect 10685 7790 34000 7792
rect 10685 7787 10751 7790
rect 14000 7760 34000 7790
rect 3325 7714 3391 7717
rect 3877 7714 3943 7717
rect 3325 7712 3943 7714
rect 3325 7656 3330 7712
rect 3386 7656 3882 7712
rect 3938 7656 3943 7712
rect 3325 7654 3943 7656
rect 3325 7651 3391 7654
rect 3877 7651 3943 7654
rect 5625 7712 5691 7717
rect 5625 7656 5630 7712
rect 5686 7656 5691 7712
rect 5625 7651 5691 7656
rect 5060 7648 5380 7649
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 7583 5380 7584
rect 1209 7578 1275 7581
rect 3877 7578 3943 7581
rect 1209 7576 3943 7578
rect 1209 7520 1214 7576
rect 1270 7520 3882 7576
rect 3938 7520 3943 7576
rect 1209 7518 3943 7520
rect 1209 7515 1275 7518
rect 3877 7515 3943 7518
rect 2405 7442 2471 7445
rect 5533 7442 5599 7445
rect 2405 7440 5599 7442
rect 2405 7384 2410 7440
rect 2466 7384 5538 7440
rect 5594 7384 5599 7440
rect 2405 7382 5599 7384
rect 2405 7379 2471 7382
rect 5533 7379 5599 7382
rect 10409 7442 10475 7445
rect 14000 7442 34000 7472
rect 10409 7440 34000 7442
rect 10409 7384 10414 7440
rect 10470 7384 34000 7440
rect 10409 7382 34000 7384
rect 10409 7379 10475 7382
rect 14000 7352 34000 7382
rect 2560 7104 2880 7105
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 7039 2880 7040
rect 7560 7104 7880 7105
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 7039 7880 7040
rect 4889 7034 4955 7037
rect 5441 7034 5507 7037
rect 4889 7032 5507 7034
rect 4889 6976 4894 7032
rect 4950 6976 5446 7032
rect 5502 6976 5507 7032
rect 4889 6974 5507 6976
rect 4889 6971 4955 6974
rect 5441 6971 5507 6974
rect 10869 7034 10935 7037
rect 14000 7034 34000 7064
rect 10869 7032 34000 7034
rect 10869 6976 10874 7032
rect 10930 6976 34000 7032
rect 10869 6974 34000 6976
rect 10869 6971 10935 6974
rect 14000 6944 34000 6974
rect 2865 6898 2931 6901
rect 8937 6898 9003 6901
rect 2865 6896 9003 6898
rect 2865 6840 2870 6896
rect 2926 6840 8942 6896
rect 8998 6840 9003 6896
rect 2865 6838 9003 6840
rect 2865 6835 2931 6838
rect 8937 6835 9003 6838
rect 2730 6702 12450 6762
rect 2497 6626 2563 6629
rect 2730 6626 2790 6702
rect 2497 6624 2790 6626
rect 2497 6568 2502 6624
rect 2558 6568 2790 6624
rect 2497 6566 2790 6568
rect 12390 6626 12450 6702
rect 14000 6626 34000 6656
rect 12390 6566 34000 6626
rect 2497 6563 2563 6566
rect 5060 6560 5380 6561
rect 5060 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5228 6560
rect 5292 6496 5308 6560
rect 5372 6496 5380 6560
rect 14000 6536 34000 6566
rect 5060 6495 5380 6496
rect 841 6490 907 6493
rect 3969 6490 4035 6493
rect 841 6488 4035 6490
rect 841 6432 846 6488
rect 902 6432 3974 6488
rect 4030 6432 4035 6488
rect 841 6430 4035 6432
rect 841 6427 907 6430
rect 3969 6427 4035 6430
rect 6729 6490 6795 6493
rect 6729 6488 9690 6490
rect 6729 6432 6734 6488
rect 6790 6432 9690 6488
rect 6729 6430 9690 6432
rect 6729 6427 6795 6430
rect 1577 6354 1643 6357
rect 7189 6354 7255 6357
rect 1577 6352 7255 6354
rect 1577 6296 1582 6352
rect 1638 6296 7194 6352
rect 7250 6296 7255 6352
rect 1577 6294 7255 6296
rect 1577 6291 1643 6294
rect 7189 6291 7255 6294
rect 2129 6218 2195 6221
rect 5809 6218 5875 6221
rect 2129 6216 5875 6218
rect 2129 6160 2134 6216
rect 2190 6160 5814 6216
rect 5870 6160 5875 6216
rect 2129 6158 5875 6160
rect 2129 6155 2195 6158
rect 5809 6155 5875 6158
rect 6085 6218 6151 6221
rect 8017 6218 8083 6221
rect 6085 6216 8083 6218
rect 6085 6160 6090 6216
rect 6146 6160 8022 6216
rect 8078 6160 8083 6216
rect 6085 6158 8083 6160
rect 9630 6218 9690 6430
rect 14000 6218 34000 6248
rect 9630 6158 34000 6218
rect 6085 6155 6151 6158
rect 8017 6155 8083 6158
rect 14000 6128 34000 6158
rect 2560 6016 2880 6017
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 5951 2880 5952
rect 7560 6016 7880 6017
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 5951 7880 5952
rect 3509 5946 3575 5949
rect 5533 5946 5599 5949
rect 5901 5946 5967 5949
rect 3509 5944 5967 5946
rect 3509 5888 3514 5944
rect 3570 5888 5538 5944
rect 5594 5888 5906 5944
rect 5962 5888 5967 5944
rect 3509 5886 5967 5888
rect 3509 5883 3575 5886
rect 5533 5883 5599 5886
rect 5901 5883 5967 5886
rect 1761 5810 1827 5813
rect 7373 5810 7439 5813
rect 1761 5808 7439 5810
rect 1761 5752 1766 5808
rect 1822 5752 7378 5808
rect 7434 5752 7439 5808
rect 1761 5750 7439 5752
rect 1761 5747 1827 5750
rect 7373 5747 7439 5750
rect 8017 5810 8083 5813
rect 14000 5810 34000 5840
rect 8017 5808 34000 5810
rect 8017 5752 8022 5808
rect 8078 5752 34000 5808
rect 8017 5750 34000 5752
rect 8017 5747 8083 5750
rect 14000 5720 34000 5750
rect 2773 5674 2839 5677
rect 3601 5674 3667 5677
rect 2773 5672 3667 5674
rect 2773 5616 2778 5672
rect 2834 5616 3606 5672
rect 3662 5616 3667 5672
rect 2773 5614 3667 5616
rect 2773 5611 2839 5614
rect 3601 5611 3667 5614
rect 3969 5674 4035 5677
rect 5165 5674 5231 5677
rect 8201 5674 8267 5677
rect 3969 5672 8267 5674
rect 3969 5616 3974 5672
rect 4030 5616 5170 5672
rect 5226 5616 8206 5672
rect 8262 5616 8267 5672
rect 3969 5614 8267 5616
rect 3969 5611 4035 5614
rect 5165 5611 5231 5614
rect 8201 5611 8267 5614
rect 5060 5472 5380 5473
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 5407 5380 5408
rect 3233 5402 3299 5405
rect 4797 5402 4863 5405
rect 3233 5400 4863 5402
rect 3233 5344 3238 5400
rect 3294 5344 4802 5400
rect 4858 5344 4863 5400
rect 3233 5342 4863 5344
rect 3233 5339 3299 5342
rect 4797 5339 4863 5342
rect 9581 5402 9647 5405
rect 14000 5402 34000 5432
rect 9581 5400 34000 5402
rect 9581 5344 9586 5400
rect 9642 5344 34000 5400
rect 9581 5342 34000 5344
rect 9581 5339 9647 5342
rect 14000 5312 34000 5342
rect 10961 4994 11027 4997
rect 14000 4994 34000 5024
rect 10961 4992 34000 4994
rect 10961 4936 10966 4992
rect 11022 4936 34000 4992
rect 10961 4934 34000 4936
rect 10961 4931 11027 4934
rect 7560 4928 7880 4929
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 14000 4904 34000 4934
rect 7560 4863 7880 4864
rect 1577 4722 1643 4725
rect 7373 4722 7439 4725
rect 1577 4720 7439 4722
rect 1577 4664 1582 4720
rect 1638 4664 7378 4720
rect 7434 4664 7439 4720
rect 1577 4662 7439 4664
rect 1577 4659 1643 4662
rect 7373 4659 7439 4662
rect 5165 4586 5231 4589
rect 4846 4584 5231 4586
rect 4846 4528 5170 4584
rect 5226 4528 5231 4584
rect 4846 4526 5231 4528
rect 4613 4178 4679 4181
rect 4248 4176 4679 4178
rect 4248 4120 4618 4176
rect 4674 4120 4679 4176
rect 4248 4118 4679 4120
rect 4846 4178 4906 4526
rect 5165 4523 5231 4526
rect 5441 4584 5507 4589
rect 5441 4528 5446 4584
rect 5502 4528 5507 4584
rect 5441 4523 5507 4528
rect 14000 4584 34000 4616
rect 14000 4528 16854 4584
rect 16910 4528 34000 4584
rect 5060 4384 5380 4385
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 4319 5380 4320
rect 5444 4181 5504 4523
rect 14000 4496 34000 4528
rect 6545 4450 6611 4453
rect 6821 4450 6887 4453
rect 6545 4448 6887 4450
rect 6545 4392 6550 4448
rect 6606 4392 6826 4448
rect 6882 4392 6887 4448
rect 6545 4390 6887 4392
rect 6545 4387 6611 4390
rect 6821 4387 6887 4390
rect 5993 4312 6059 4317
rect 5993 4256 5998 4312
rect 6054 4256 6059 4312
rect 5993 4251 6059 4256
rect 4981 4178 5047 4181
rect 4846 4176 5047 4178
rect 4846 4120 4986 4176
rect 5042 4120 5047 4176
rect 4846 4118 5047 4120
rect 4248 3501 4308 4118
rect 4613 4115 4679 4118
rect 4981 4115 5047 4118
rect 5441 4176 5507 4181
rect 5441 4120 5446 4176
rect 5502 4120 5507 4176
rect 5441 4115 5507 4120
rect 5625 4178 5691 4181
rect 5996 4178 6056 4251
rect 5625 4176 6056 4178
rect 5625 4120 5630 4176
rect 5686 4120 6056 4176
rect 5625 4118 6056 4120
rect 13445 4178 13511 4181
rect 14000 4178 34000 4208
rect 13445 4176 34000 4178
rect 13445 4120 13450 4176
rect 13506 4120 34000 4176
rect 13445 4118 34000 4120
rect 5625 4115 5691 4118
rect 13445 4115 13511 4118
rect 14000 4088 34000 4118
rect 7560 3840 7880 3841
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 3775 7880 3776
rect 14000 3768 34000 3800
rect 14000 3712 16670 3768
rect 16726 3712 34000 3768
rect 14000 3680 34000 3712
rect 4245 3496 4311 3501
rect 8109 3498 8175 3501
rect 4245 3440 4250 3496
rect 4306 3440 4311 3496
rect 4245 3435 4311 3440
rect 4846 3496 8175 3498
rect 4846 3440 8114 3496
rect 8170 3440 8175 3496
rect 4846 3438 8175 3440
rect 3509 3362 3575 3365
rect 4846 3362 4906 3438
rect 8109 3435 8175 3438
rect 3509 3360 4906 3362
rect 2454 2546 2514 3332
rect 3509 3304 3514 3360
rect 3570 3304 4906 3360
rect 3509 3302 4906 3304
rect 13537 3362 13603 3365
rect 14000 3362 34000 3392
rect 13537 3360 34000 3362
rect 13537 3304 13542 3360
rect 13598 3304 34000 3360
rect 13537 3302 34000 3304
rect 3509 3299 3575 3302
rect 13537 3299 13603 3302
rect 5060 3296 5380 3297
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 14000 3272 34000 3302
rect 5060 3231 5380 3232
rect 7373 3226 7439 3229
rect 8753 3226 8819 3229
rect 7373 3224 8819 3226
rect 7373 3168 7378 3224
rect 7434 3168 8758 3224
rect 8814 3168 8819 3224
rect 7373 3166 8819 3168
rect 7373 3163 7439 3166
rect 8753 3163 8819 3166
rect 4613 3090 4679 3093
rect 9029 3090 9095 3093
rect 4613 3088 9095 3090
rect 4613 3032 4618 3088
rect 4674 3032 9034 3088
rect 9090 3032 9095 3088
rect 4613 3030 9095 3032
rect 4613 3027 4679 3030
rect 9029 3027 9095 3030
rect 3601 2954 3667 2957
rect 6545 2954 6611 2957
rect 3601 2952 6611 2954
rect 3601 2896 3606 2952
rect 3662 2896 6550 2952
rect 6606 2896 6611 2952
rect 3601 2894 6611 2896
rect 3601 2891 3667 2894
rect 6545 2891 6611 2894
rect 14000 2952 34000 2984
rect 14000 2896 16578 2952
rect 16634 2896 34000 2952
rect 14000 2864 34000 2896
rect 4429 2818 4495 2821
rect 4889 2818 4955 2821
rect 4429 2816 4955 2818
rect 4429 2760 4434 2816
rect 4490 2760 4894 2816
rect 4950 2760 4955 2816
rect 4429 2758 4955 2760
rect 4429 2755 4495 2758
rect 4889 2755 4955 2758
rect 5533 2818 5599 2821
rect 7373 2818 7439 2821
rect 5533 2816 7439 2818
rect 5533 2760 5538 2816
rect 5594 2760 7378 2816
rect 7434 2760 7439 2816
rect 5533 2758 7439 2760
rect 5533 2755 5599 2758
rect 7373 2755 7439 2758
rect 7560 2752 7880 2753
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 2687 7880 2688
rect 8661 2682 8727 2685
rect 13445 2682 13511 2685
rect 8661 2680 13511 2682
rect 8661 2624 8666 2680
rect 8722 2624 13450 2680
rect 13506 2624 13511 2680
rect 8661 2622 13511 2624
rect 8661 2619 8727 2622
rect 13445 2619 13511 2622
rect 7925 2546 7991 2549
rect 2454 2544 7991 2546
rect 2454 2488 7930 2544
rect 7986 2488 7991 2544
rect 2454 2486 7991 2488
rect 7925 2483 7991 2486
rect 8201 2546 8267 2549
rect 14000 2546 34000 2576
rect 8201 2544 34000 2546
rect 8201 2488 8206 2544
rect 8262 2488 34000 2544
rect 8201 2486 34000 2488
rect 8201 2483 8267 2486
rect 14000 2456 34000 2486
rect 4429 2410 4495 2413
rect 9581 2410 9647 2413
rect 4429 2408 9647 2410
rect 4429 2352 4434 2408
rect 4490 2352 9586 2408
rect 9642 2352 9647 2408
rect 4429 2350 9647 2352
rect 4429 2347 4495 2350
rect 9581 2347 9647 2350
rect 5060 2208 5380 2209
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 2143 5380 2144
rect 6269 2138 6335 2141
rect 9397 2138 9463 2141
rect 6269 2136 9463 2138
rect 6269 2080 6274 2136
rect 6330 2080 9402 2136
rect 9458 2080 9463 2136
rect 6269 2078 9463 2080
rect 6269 2075 6335 2078
rect 9397 2075 9463 2078
rect 14000 2136 34000 2168
rect 14000 2080 16762 2136
rect 16818 2080 34000 2136
rect 14000 2048 34000 2080
rect 5165 2002 5231 2005
rect 6821 2002 6887 2005
rect 5165 2000 6887 2002
rect 5165 1944 5170 2000
rect 5226 1944 6826 2000
rect 6882 1944 6887 2000
rect 5165 1942 6887 1944
rect 5165 1939 5231 1942
rect 6821 1939 6887 1942
rect 2497 1866 2563 1869
rect 5533 1866 5599 1869
rect 2497 1864 5599 1866
rect 2497 1808 2502 1864
rect 2558 1808 5538 1864
rect 5594 1808 5599 1864
rect 2497 1806 5599 1808
rect 2497 1803 2563 1806
rect 5533 1803 5599 1806
rect 8017 1866 8083 1869
rect 13813 1866 13879 1869
rect 8017 1864 13879 1866
rect 8017 1808 8022 1864
rect 8078 1808 13818 1864
rect 13874 1808 13879 1864
rect 8017 1806 13879 1808
rect 8017 1803 8083 1806
rect 13813 1803 13879 1806
rect 3601 1730 3667 1733
rect 6913 1730 6979 1733
rect 3601 1728 6979 1730
rect 3601 1672 3606 1728
rect 3662 1672 6918 1728
rect 6974 1672 6979 1728
rect 3601 1670 6979 1672
rect 3601 1667 3667 1670
rect 6913 1667 6979 1670
rect 14000 1728 34000 1760
rect 14000 1672 16578 1728
rect 16634 1672 34000 1728
rect 7560 1664 7880 1665
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 14000 1640 34000 1672
rect 7560 1599 7880 1600
rect 4981 1322 5047 1325
rect 10041 1322 10107 1325
rect 14000 1322 34000 1352
rect 4981 1320 10107 1322
rect 4981 1264 4986 1320
rect 5042 1264 10046 1320
rect 10102 1264 10107 1320
rect 4981 1262 10107 1264
rect 4981 1259 5047 1262
rect 10041 1259 10107 1262
rect 12390 1262 34000 1322
rect 5441 1186 5507 1189
rect 11053 1186 11119 1189
rect 5441 1184 11119 1186
rect 5441 1128 5446 1184
rect 5502 1128 11058 1184
rect 11114 1128 11119 1184
rect 5441 1126 11119 1128
rect 5441 1123 5507 1126
rect 11053 1123 11119 1126
rect 5060 1120 5380 1121
rect 5060 1056 5068 1120
rect 5132 1056 5148 1120
rect 5212 1056 5228 1120
rect 5292 1056 5308 1120
rect 5372 1056 5380 1120
rect 5060 1055 5380 1056
rect 9213 1050 9279 1053
rect 12390 1050 12450 1262
rect 14000 1232 34000 1262
rect 9213 1048 12450 1050
rect 9213 992 9218 1048
rect 9274 992 12450 1048
rect 9213 990 12450 992
rect 9213 987 9279 990
rect 9673 914 9739 917
rect 14000 914 34000 944
rect 9673 912 34000 914
rect 9673 856 9678 912
rect 9734 856 34000 912
rect 9673 854 34000 856
rect 9673 851 9739 854
rect 14000 824 34000 854
rect 14000 504 34000 536
rect 14000 448 16670 504
rect 16726 448 34000 504
rect 14000 416 34000 448
<< via3 >>
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 7568 11452 7632 11456
rect 7568 11396 7572 11452
rect 7572 11396 7628 11452
rect 7628 11396 7632 11452
rect 7568 11392 7632 11396
rect 7648 11452 7712 11456
rect 7648 11396 7652 11452
rect 7652 11396 7708 11452
rect 7708 11396 7712 11452
rect 7648 11392 7712 11396
rect 7728 11452 7792 11456
rect 7728 11396 7732 11452
rect 7732 11396 7788 11452
rect 7788 11396 7792 11452
rect 7728 11392 7792 11396
rect 7808 11452 7872 11456
rect 7808 11396 7812 11452
rect 7812 11396 7868 11452
rect 7868 11396 7872 11452
rect 7808 11392 7872 11396
rect 5068 10908 5132 10912
rect 5068 10852 5072 10908
rect 5072 10852 5128 10908
rect 5128 10852 5132 10908
rect 5068 10848 5132 10852
rect 5148 10908 5212 10912
rect 5148 10852 5152 10908
rect 5152 10852 5208 10908
rect 5208 10852 5212 10908
rect 5148 10848 5212 10852
rect 5228 10908 5292 10912
rect 5228 10852 5232 10908
rect 5232 10852 5288 10908
rect 5288 10852 5292 10908
rect 5228 10848 5292 10852
rect 5308 10908 5372 10912
rect 5308 10852 5312 10908
rect 5312 10852 5368 10908
rect 5368 10852 5372 10908
rect 5308 10848 5372 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 7568 10364 7632 10368
rect 7568 10308 7572 10364
rect 7572 10308 7628 10364
rect 7628 10308 7632 10364
rect 7568 10304 7632 10308
rect 7648 10364 7712 10368
rect 7648 10308 7652 10364
rect 7652 10308 7708 10364
rect 7708 10308 7712 10364
rect 7648 10304 7712 10308
rect 7728 10364 7792 10368
rect 7728 10308 7732 10364
rect 7732 10308 7788 10364
rect 7788 10308 7792 10364
rect 7728 10304 7792 10308
rect 7808 10364 7872 10368
rect 7808 10308 7812 10364
rect 7812 10308 7868 10364
rect 7868 10308 7872 10364
rect 7808 10304 7872 10308
rect 5068 9820 5132 9824
rect 5068 9764 5072 9820
rect 5072 9764 5128 9820
rect 5128 9764 5132 9820
rect 5068 9760 5132 9764
rect 5148 9820 5212 9824
rect 5148 9764 5152 9820
rect 5152 9764 5208 9820
rect 5208 9764 5212 9820
rect 5148 9760 5212 9764
rect 5228 9820 5292 9824
rect 5228 9764 5232 9820
rect 5232 9764 5288 9820
rect 5288 9764 5292 9820
rect 5228 9760 5292 9764
rect 5308 9820 5372 9824
rect 5308 9764 5312 9820
rect 5312 9764 5368 9820
rect 5368 9764 5372 9820
rect 5308 9760 5372 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 7568 9276 7632 9280
rect 7568 9220 7572 9276
rect 7572 9220 7628 9276
rect 7628 9220 7632 9276
rect 7568 9216 7632 9220
rect 7648 9276 7712 9280
rect 7648 9220 7652 9276
rect 7652 9220 7708 9276
rect 7708 9220 7712 9276
rect 7648 9216 7712 9220
rect 7728 9276 7792 9280
rect 7728 9220 7732 9276
rect 7732 9220 7788 9276
rect 7788 9220 7792 9276
rect 7728 9216 7792 9220
rect 7808 9276 7872 9280
rect 7808 9220 7812 9276
rect 7812 9220 7868 9276
rect 7868 9220 7872 9276
rect 7808 9216 7872 9220
rect 5068 8732 5132 8736
rect 5068 8676 5072 8732
rect 5072 8676 5128 8732
rect 5128 8676 5132 8732
rect 5068 8672 5132 8676
rect 5148 8732 5212 8736
rect 5148 8676 5152 8732
rect 5152 8676 5208 8732
rect 5208 8676 5212 8732
rect 5148 8672 5212 8676
rect 5228 8732 5292 8736
rect 5228 8676 5232 8732
rect 5232 8676 5288 8732
rect 5288 8676 5292 8732
rect 5228 8672 5292 8676
rect 5308 8732 5372 8736
rect 5308 8676 5312 8732
rect 5312 8676 5368 8732
rect 5368 8676 5372 8732
rect 5308 8672 5372 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 7568 8188 7632 8192
rect 7568 8132 7572 8188
rect 7572 8132 7628 8188
rect 7628 8132 7632 8188
rect 7568 8128 7632 8132
rect 7648 8188 7712 8192
rect 7648 8132 7652 8188
rect 7652 8132 7708 8188
rect 7708 8132 7712 8188
rect 7648 8128 7712 8132
rect 7728 8188 7792 8192
rect 7728 8132 7732 8188
rect 7732 8132 7788 8188
rect 7788 8132 7792 8188
rect 7728 8128 7792 8132
rect 7808 8188 7872 8192
rect 7808 8132 7812 8188
rect 7812 8132 7868 8188
rect 7868 8132 7872 8188
rect 7808 8128 7872 8132
rect 5068 7644 5132 7648
rect 5068 7588 5072 7644
rect 5072 7588 5128 7644
rect 5128 7588 5132 7644
rect 5068 7584 5132 7588
rect 5148 7644 5212 7648
rect 5148 7588 5152 7644
rect 5152 7588 5208 7644
rect 5208 7588 5212 7644
rect 5148 7584 5212 7588
rect 5228 7644 5292 7648
rect 5228 7588 5232 7644
rect 5232 7588 5288 7644
rect 5288 7588 5292 7644
rect 5228 7584 5292 7588
rect 5308 7644 5372 7648
rect 5308 7588 5312 7644
rect 5312 7588 5368 7644
rect 5368 7588 5372 7644
rect 5308 7584 5372 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 7568 7100 7632 7104
rect 7568 7044 7572 7100
rect 7572 7044 7628 7100
rect 7628 7044 7632 7100
rect 7568 7040 7632 7044
rect 7648 7100 7712 7104
rect 7648 7044 7652 7100
rect 7652 7044 7708 7100
rect 7708 7044 7712 7100
rect 7648 7040 7712 7044
rect 7728 7100 7792 7104
rect 7728 7044 7732 7100
rect 7732 7044 7788 7100
rect 7788 7044 7792 7100
rect 7728 7040 7792 7044
rect 7808 7100 7872 7104
rect 7808 7044 7812 7100
rect 7812 7044 7868 7100
rect 7868 7044 7872 7100
rect 7808 7040 7872 7044
rect 5068 6556 5132 6560
rect 5068 6500 5072 6556
rect 5072 6500 5128 6556
rect 5128 6500 5132 6556
rect 5068 6496 5132 6500
rect 5148 6556 5212 6560
rect 5148 6500 5152 6556
rect 5152 6500 5208 6556
rect 5208 6500 5212 6556
rect 5148 6496 5212 6500
rect 5228 6556 5292 6560
rect 5228 6500 5232 6556
rect 5232 6500 5288 6556
rect 5288 6500 5292 6556
rect 5228 6496 5292 6500
rect 5308 6556 5372 6560
rect 5308 6500 5312 6556
rect 5312 6500 5368 6556
rect 5368 6500 5372 6556
rect 5308 6496 5372 6500
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 7568 6012 7632 6016
rect 7568 5956 7572 6012
rect 7572 5956 7628 6012
rect 7628 5956 7632 6012
rect 7568 5952 7632 5956
rect 7648 6012 7712 6016
rect 7648 5956 7652 6012
rect 7652 5956 7708 6012
rect 7708 5956 7712 6012
rect 7648 5952 7712 5956
rect 7728 6012 7792 6016
rect 7728 5956 7732 6012
rect 7732 5956 7788 6012
rect 7788 5956 7792 6012
rect 7728 5952 7792 5956
rect 7808 6012 7872 6016
rect 7808 5956 7812 6012
rect 7812 5956 7868 6012
rect 7868 5956 7872 6012
rect 7808 5952 7872 5956
rect 5068 5468 5132 5472
rect 5068 5412 5072 5468
rect 5072 5412 5128 5468
rect 5128 5412 5132 5468
rect 5068 5408 5132 5412
rect 5148 5468 5212 5472
rect 5148 5412 5152 5468
rect 5152 5412 5208 5468
rect 5208 5412 5212 5468
rect 5148 5408 5212 5412
rect 5228 5468 5292 5472
rect 5228 5412 5232 5468
rect 5232 5412 5288 5468
rect 5288 5412 5292 5468
rect 5228 5408 5292 5412
rect 5308 5468 5372 5472
rect 5308 5412 5312 5468
rect 5312 5412 5368 5468
rect 5368 5412 5372 5468
rect 5308 5408 5372 5412
rect 7568 4924 7632 4928
rect 7568 4868 7572 4924
rect 7572 4868 7628 4924
rect 7628 4868 7632 4924
rect 7568 4864 7632 4868
rect 7648 4924 7712 4928
rect 7648 4868 7652 4924
rect 7652 4868 7708 4924
rect 7708 4868 7712 4924
rect 7648 4864 7712 4868
rect 7728 4924 7792 4928
rect 7728 4868 7732 4924
rect 7732 4868 7788 4924
rect 7788 4868 7792 4924
rect 7728 4864 7792 4868
rect 7808 4924 7872 4928
rect 7808 4868 7812 4924
rect 7812 4868 7868 4924
rect 7868 4868 7872 4924
rect 7808 4864 7872 4868
rect 5068 4380 5132 4384
rect 5068 4324 5072 4380
rect 5072 4324 5128 4380
rect 5128 4324 5132 4380
rect 5068 4320 5132 4324
rect 5148 4380 5212 4384
rect 5148 4324 5152 4380
rect 5152 4324 5208 4380
rect 5208 4324 5212 4380
rect 5148 4320 5212 4324
rect 5228 4380 5292 4384
rect 5228 4324 5232 4380
rect 5232 4324 5288 4380
rect 5288 4324 5292 4380
rect 5228 4320 5292 4324
rect 5308 4380 5372 4384
rect 5308 4324 5312 4380
rect 5312 4324 5368 4380
rect 5368 4324 5372 4380
rect 5308 4320 5372 4324
rect 7568 3836 7632 3840
rect 7568 3780 7572 3836
rect 7572 3780 7628 3836
rect 7628 3780 7632 3836
rect 7568 3776 7632 3780
rect 7648 3836 7712 3840
rect 7648 3780 7652 3836
rect 7652 3780 7708 3836
rect 7708 3780 7712 3836
rect 7648 3776 7712 3780
rect 7728 3836 7792 3840
rect 7728 3780 7732 3836
rect 7732 3780 7788 3836
rect 7788 3780 7792 3836
rect 7728 3776 7792 3780
rect 7808 3836 7872 3840
rect 7808 3780 7812 3836
rect 7812 3780 7868 3836
rect 7868 3780 7872 3836
rect 7808 3776 7872 3780
rect 5068 3292 5132 3296
rect 5068 3236 5072 3292
rect 5072 3236 5128 3292
rect 5128 3236 5132 3292
rect 5068 3232 5132 3236
rect 5148 3292 5212 3296
rect 5148 3236 5152 3292
rect 5152 3236 5208 3292
rect 5208 3236 5212 3292
rect 5148 3232 5212 3236
rect 5228 3292 5292 3296
rect 5228 3236 5232 3292
rect 5232 3236 5288 3292
rect 5288 3236 5292 3292
rect 5228 3232 5292 3236
rect 5308 3292 5372 3296
rect 5308 3236 5312 3292
rect 5312 3236 5368 3292
rect 5368 3236 5372 3292
rect 5308 3232 5372 3236
rect 7568 2748 7632 2752
rect 7568 2692 7572 2748
rect 7572 2692 7628 2748
rect 7628 2692 7632 2748
rect 7568 2688 7632 2692
rect 7648 2748 7712 2752
rect 7648 2692 7652 2748
rect 7652 2692 7708 2748
rect 7708 2692 7712 2748
rect 7648 2688 7712 2692
rect 7728 2748 7792 2752
rect 7728 2692 7732 2748
rect 7732 2692 7788 2748
rect 7788 2692 7792 2748
rect 7728 2688 7792 2692
rect 7808 2748 7872 2752
rect 7808 2692 7812 2748
rect 7812 2692 7868 2748
rect 7868 2692 7872 2748
rect 7808 2688 7872 2692
rect 5068 2204 5132 2208
rect 5068 2148 5072 2204
rect 5072 2148 5128 2204
rect 5128 2148 5132 2204
rect 5068 2144 5132 2148
rect 5148 2204 5212 2208
rect 5148 2148 5152 2204
rect 5152 2148 5208 2204
rect 5208 2148 5212 2204
rect 5148 2144 5212 2148
rect 5228 2204 5292 2208
rect 5228 2148 5232 2204
rect 5232 2148 5288 2204
rect 5288 2148 5292 2204
rect 5228 2144 5292 2148
rect 5308 2204 5372 2208
rect 5308 2148 5312 2204
rect 5312 2148 5368 2204
rect 5368 2148 5372 2204
rect 5308 2144 5372 2148
rect 7568 1660 7632 1664
rect 7568 1604 7572 1660
rect 7572 1604 7628 1660
rect 7628 1604 7632 1660
rect 7568 1600 7632 1604
rect 7648 1660 7712 1664
rect 7648 1604 7652 1660
rect 7652 1604 7708 1660
rect 7708 1604 7712 1660
rect 7648 1600 7712 1604
rect 7728 1660 7792 1664
rect 7728 1604 7732 1660
rect 7732 1604 7788 1660
rect 7788 1604 7792 1660
rect 7728 1600 7792 1604
rect 7808 1660 7872 1664
rect 7808 1604 7812 1660
rect 7812 1604 7868 1660
rect 7868 1604 7872 1660
rect 7808 1600 7872 1604
rect 5068 1116 5132 1120
rect 5068 1060 5072 1116
rect 5072 1060 5128 1116
rect 5128 1060 5132 1116
rect 5068 1056 5132 1060
rect 5148 1116 5212 1120
rect 5148 1060 5152 1116
rect 5152 1060 5208 1116
rect 5208 1060 5212 1116
rect 5148 1056 5212 1060
rect 5228 1116 5292 1120
rect 5228 1060 5232 1116
rect 5232 1060 5288 1116
rect 5288 1060 5292 1116
rect 5228 1056 5292 1060
rect 5308 1116 5372 1120
rect 5308 1060 5312 1116
rect 5312 1060 5368 1116
rect 5368 1060 5372 1116
rect 5308 1056 5372 1060
<< metal4 >>
rect 2560 11456 2880 11472
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 8218 2880 9216
rect 2560 8192 2602 8218
rect 2838 8192 2880 8218
rect 2560 8128 2568 8192
rect 2872 8128 2880 8192
rect 2560 7982 2602 8128
rect 2838 7982 2880 8128
rect 2560 7104 2880 7982
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 4838 2880 5952
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1088 2880 1222
rect 3560 9266 3880 11424
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3560 5886 3880 9030
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 3560 2506 3880 5650
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 3560 1088 3880 2270
rect 5060 10912 5380 11472
rect 7560 11456 7880 11472
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 9908 5380 10848
rect 5060 9824 5102 9908
rect 5338 9824 5380 9908
rect 5060 9760 5068 9824
rect 5372 9760 5380 9824
rect 5060 9672 5102 9760
rect 5338 9672 5380 9760
rect 5060 8736 5380 9672
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 7648 5380 8672
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 6560 5380 7584
rect 5060 6496 5068 6560
rect 5132 6528 5148 6560
rect 5212 6528 5228 6560
rect 5292 6528 5308 6560
rect 5372 6496 5380 6560
rect 5060 6292 5102 6496
rect 5338 6292 5380 6496
rect 5060 5472 5380 6292
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 4384 5380 5408
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 3296 5380 4320
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 5060 3148 5380 3232
rect 5060 2912 5102 3148
rect 5338 2912 5380 3148
rect 5060 2208 5380 2912
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 1120 5380 2144
rect 5060 1056 5068 1120
rect 5132 1056 5148 1120
rect 5212 1056 5228 1120
rect 5292 1056 5308 1120
rect 5372 1056 5380 1120
rect 6060 10956 6380 11424
rect 6060 10720 6102 10956
rect 6338 10720 6380 10956
rect 6060 7576 6380 10720
rect 6060 7340 6102 7576
rect 6338 7340 6380 7576
rect 6060 4196 6380 7340
rect 6060 3960 6102 4196
rect 6338 3960 6380 4196
rect 6060 1088 6380 3960
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 7560 10368 7880 11392
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 9280 7880 10304
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 8218 7880 9216
rect 7560 8192 7602 8218
rect 7838 8192 7880 8218
rect 7560 8128 7568 8192
rect 7872 8128 7880 8192
rect 7560 7982 7602 8128
rect 7838 7982 7880 8128
rect 7560 7104 7880 7982
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 6016 7880 7040
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 4928 7880 5952
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 7560 4838 7880 4864
rect 7560 4602 7602 4838
rect 7838 4602 7880 4838
rect 7560 3840 7880 4602
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 2752 7880 3776
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 1664 7880 2688
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 7560 1458 7880 1600
rect 7560 1222 7602 1458
rect 7838 1222 7880 1458
rect 5060 1040 5380 1056
rect 7560 1040 7880 1222
rect 8560 9266 8880 11424
rect 8560 9030 8602 9266
rect 8838 9030 8880 9266
rect 8560 5886 8880 9030
rect 8560 5650 8602 5886
rect 8838 5650 8880 5886
rect 8560 2506 8880 5650
rect 8560 2270 8602 2506
rect 8838 2270 8880 2506
rect 8560 1088 8880 2270
<< via4 >>
rect 2602 8192 2838 8218
rect 2602 8128 2632 8192
rect 2632 8128 2648 8192
rect 2648 8128 2712 8192
rect 2712 8128 2728 8192
rect 2728 8128 2792 8192
rect 2792 8128 2808 8192
rect 2808 8128 2838 8192
rect 2602 7982 2838 8128
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 2602 1222 2838 1458
rect 3602 9030 3838 9266
rect 3602 5650 3838 5886
rect 3602 2270 3838 2506
rect 5102 9824 5338 9908
rect 5102 9760 5132 9824
rect 5132 9760 5148 9824
rect 5148 9760 5212 9824
rect 5212 9760 5228 9824
rect 5228 9760 5292 9824
rect 5292 9760 5308 9824
rect 5308 9760 5338 9824
rect 5102 9672 5338 9760
rect 5102 6496 5132 6528
rect 5132 6496 5148 6528
rect 5148 6496 5212 6528
rect 5212 6496 5228 6528
rect 5228 6496 5292 6528
rect 5292 6496 5308 6528
rect 5308 6496 5338 6528
rect 5102 6292 5338 6496
rect 5102 2912 5338 3148
rect 6102 10720 6338 10956
rect 6102 7340 6338 7576
rect 6102 3960 6338 4196
rect 7602 8192 7838 8218
rect 7602 8128 7632 8192
rect 7632 8128 7648 8192
rect 7648 8128 7712 8192
rect 7712 8128 7728 8192
rect 7728 8128 7792 8192
rect 7792 8128 7808 8192
rect 7808 8128 7838 8192
rect 7602 7982 7838 8128
rect 7602 4602 7838 4838
rect 7602 1222 7838 1458
rect 8602 9030 8838 9266
rect 8602 5650 8838 5886
rect 8602 2270 8838 2506
<< metal5 >>
rect 920 10956 9844 10998
rect 920 10720 6102 10956
rect 6338 10720 9844 10956
rect 920 10678 9844 10720
rect 920 9908 9844 9950
rect 920 9672 5102 9908
rect 5338 9672 9844 9908
rect 920 9630 9844 9672
rect 920 9266 9844 9308
rect 920 9030 3602 9266
rect 3838 9030 8602 9266
rect 8838 9030 9844 9266
rect 920 8988 9844 9030
rect 920 8218 9844 8260
rect 920 7982 2602 8218
rect 2838 7982 7602 8218
rect 7838 7982 9844 8218
rect 920 7940 9844 7982
rect 920 7576 9844 7618
rect 920 7340 6102 7576
rect 6338 7340 9844 7576
rect 920 7298 9844 7340
rect 920 6528 9844 6570
rect 920 6292 5102 6528
rect 5338 6292 9844 6528
rect 920 6250 9844 6292
rect 920 5886 9844 5928
rect 920 5650 3602 5886
rect 3838 5650 8602 5886
rect 8838 5650 9844 5886
rect 920 5608 9844 5650
rect 920 4838 9844 4880
rect 920 4602 2602 4838
rect 2838 4602 7602 4838
rect 7838 4602 9844 4838
rect 920 4560 9844 4602
rect 920 4196 9844 4238
rect 920 3960 2018 4196
rect 2254 3960 6102 4196
rect 6338 3960 9844 4196
rect 920 3918 9844 3960
rect 920 3148 9844 3190
rect 920 2912 5102 3148
rect 5338 2912 9844 3148
rect 920 2870 9844 2912
rect 920 2506 9844 2548
rect 920 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 8602 2506
rect 8838 2270 9844 2506
rect 920 2228 9844 2270
rect 920 1458 9844 1500
rect 920 1222 2602 1458
rect 2838 1222 7602 1458
rect 7838 1222 9844 1458
rect 920 1180 9844 1222
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform -1 0 8004 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1659391890
transform -1 0 7636 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1659391890
transform -1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1659391890
transform 1 0 7084 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1659391890
transform -1 0 6624 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1659391890
transform -1 0 4232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1659391890
transform -1 0 3680 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1659391890
transform 1 0 4324 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 5520 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 6256 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 6900 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69
timestamp 1659391890
transform 1 0 7268 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73
timestamp 1659391890
transform 1 0 7636 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1659391890
transform 1 0 8004 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80
timestamp 1659391890
transform 1 0 8280 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1659391890
transform 1 0 9476 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1659391890
transform 1 0 3312 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_30
timestamp 1659391890
transform 1 0 3680 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1659391890
transform 1 0 4140 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp 1659391890
transform 1 0 4508 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1659391890
transform 1 0 5796 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_58
timestamp 1659391890
transform 1 0 6256 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1659391890
transform 1 0 6624 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_73
timestamp 1659391890
transform 1 0 7636 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_80
timestamp 1659391890
transform 1 0 8280 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1659391890
transform 1 0 3864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_36
timestamp 1659391890
transform 1 0 4232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1659391890
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_46
timestamp 1659391890
transform 1 0 5152 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_50
timestamp 1659391890
transform 1 0 5520 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_55
timestamp 1659391890
transform 1 0 5980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_70
timestamp 1659391890
transform 1 0 7360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_75
timestamp 1659391890
transform 1 0 7820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1659391890
transform 1 0 5980 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_70
timestamp 1659391890
transform 1 0 7360 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_80
timestamp 1659391890
transform 1 0 8280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_86
timestamp 1659391890
transform 1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_90
timestamp 1659391890
transform 1 0 9200 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_46
timestamp 1659391890
transform 1 0 5152 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_92
timestamp 1659391890
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_26
timestamp 1659391890
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_52
timestamp 1659391890
transform 1 0 5704 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_26
timestamp 1659391890
transform 1 0 3312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_88
timestamp 1659391890
transform 1 0 9016 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1659391890
transform 1 0 1196 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_55
timestamp 1659391890
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1659391890
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_45
timestamp 1659391890
transform 1 0 5060 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1659391890
transform 1 0 1196 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_37
timestamp 1659391890
transform 1 0 4324 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1659391890
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_93
timestamp 1659391890
transform 1 0 9476 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1659391890
transform 1 0 1196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1659391890
transform 1 0 3588 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1659391890
transform 1 0 1196 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_36
timestamp 1659391890
transform 1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1659391890
transform 1 0 6624 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_24
timestamp 1659391890
transform 1 0 3128 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_43
timestamp 1659391890
transform 1 0 4876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_49
timestamp 1659391890
transform 1 0 5428 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_73
timestamp 1659391890
transform 1 0 7636 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_3
timestamp 1659391890
transform 1 0 1196 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_37
timestamp 1659391890
transform 1 0 4324 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_75
timestamp 1659391890
transform 1 0 7820 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1659391890
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_11
timestamp 1659391890
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1659391890
transform 1 0 5980 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1659391890
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1659391890
transform 1 0 1196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1659391890
transform 1 0 3588 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_39
timestamp 1659391890
transform 1 0 4508 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_49
timestamp 1659391890
transform 1 0 5428 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_57
timestamp 1659391890
transform 1 0 6164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_67
timestamp 1659391890
transform 1 0 7084 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1659391890
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1659391890
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1659391890
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1659391890
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1659391890
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1659391890
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1659391890
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1659391890
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1659391890
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1659391890
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1659391890
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1659391890
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1659391890
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1659391890
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1659391890
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1659391890
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1659391890
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1659391890
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1659391890
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1659391890
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1659391890
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1659391890
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1659391890
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1659391890
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1659391890
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1659391890
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1659391890
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1659391890
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1659391890
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1659391890
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1659391890
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1659391890
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1659391890
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1659391890
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1659391890
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1659391890
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1659391890
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1659391890
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1659391890
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1659391890
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1659391890
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1659391890
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1659391890
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1659391890
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1659391890
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1659391890
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1659391890
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1659391890
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1659391890
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1659391890
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1659391890
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1659391890
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1659391890
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1659391890
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1659391890
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1659391890
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1659391890
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1659391890
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1659391890
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1659391890
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1659391890
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1659391890
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1659391890
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1659391890
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1659391890
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 7268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 5152 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 5428 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1659391890
transform 1 0 7636 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _112_
timestamp 1659391890
transform 1 0 5152 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 6164 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1659391890
transform 1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115__1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115__2
timestamp 1659391890
transform 1 0 3220 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115__3
timestamp 1659391890
transform 1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115__4
timestamp 1659391890
transform 1 0 1564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115__5
timestamp 1659391890
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _116_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _117_
timestamp 1659391890
transform 1 0 3404 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1659391890
transform 1 0 4784 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _119_
timestamp 1659391890
transform 1 0 6164 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1659391890
transform 1 0 5336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _121_
timestamp 1659391890
transform 1 0 3864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _122_
timestamp 1659391890
transform 1 0 4140 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _123_
timestamp 1659391890
transform 1 0 4232 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1659391890
transform 1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _125_
timestamp 1659391890
transform 1 0 6164 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _126_
timestamp 1659391890
transform 1 0 4692 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1659391890
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _128_
timestamp 1659391890
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _129_
timestamp 1659391890
transform 1 0 6072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _130_
timestamp 1659391890
transform 1 0 6072 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1659391890
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _132_
timestamp 1659391890
transform 1 0 8832 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1659391890
transform 1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _134_
timestamp 1659391890
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _135_
timestamp 1659391890
transform 1 0 5980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _136_
timestamp 1659391890
transform 1 0 9016 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1659391890
transform 1 0 7360 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _138_
timestamp 1659391890
transform 1 0 5152 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1659391890
transform 1 0 7084 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _140_
timestamp 1659391890
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _141_
timestamp 1659391890
transform 1 0 1748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _142_
timestamp 1659391890
transform 1 0 4968 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _143_
timestamp 1659391890
transform 1 0 8096 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1659391890
transform 1 0 6348 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _145_
timestamp 1659391890
transform 1 0 7452 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1659391890
transform 1 0 5796 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _147_
timestamp 1659391890
transform 1 0 2208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _148_
timestamp 1659391890
transform 1 0 2576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _149_
timestamp 1659391890
transform 1 0 2852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _150_
timestamp 1659391890
transform 1 0 4324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1659391890
transform 1 0 2300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _152_
timestamp 1659391890
transform 1 0 4048 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1659391890
transform 1 0 4692 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _154_
timestamp 1659391890
transform 1 0 1932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _155_
timestamp 1659391890
transform 1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _156_
timestamp 1659391890
transform 1 0 2944 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1659391890
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1659391890
transform 1 0 5520 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _159_
timestamp 1659391890
transform 1 0 2484 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1659391890
transform 1 0 1748 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _161_
timestamp 1659391890
transform 1 0 1288 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _162_
timestamp 1659391890
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _163_
timestamp 1659391890
transform 1 0 2944 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1659391890
transform 1 0 1472 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _165_
timestamp 1659391890
transform 1 0 2484 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1659391890
transform 1 0 1196 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _167_
timestamp 1659391890
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _168_
timestamp 1659391890
transform 1 0 2300 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _169_
timestamp 1659391890
transform 1 0 7084 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1659391890
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _171_
timestamp 1659391890
transform 1 0 6900 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _172_
timestamp 1659391890
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _173_
timestamp 1659391890
transform 1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _174_
timestamp 1659391890
transform 1 0 2392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _175_
timestamp 1659391890
transform 1 0 5520 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _176_
timestamp 1659391890
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _177_
timestamp 1659391890
transform 1 0 7360 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _178_
timestamp 1659391890
transform 1 0 2576 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _179_
timestamp 1659391890
transform 1 0 1840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _180_
timestamp 1659391890
transform 1 0 1564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _181_
timestamp 1659391890
transform 1 0 4968 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1659391890
transform 1 0 1288 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _183_
timestamp 1659391890
transform 1 0 5520 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 1659391890
transform 1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _185_
timestamp 1659391890
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _186_
timestamp 1659391890
transform 1 0 1472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _187_
timestamp 1659391890
transform 1 0 6256 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 1659391890
transform 1 0 1196 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _189_
timestamp 1659391890
transform 1 0 6624 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 1659391890
transform 1 0 1472 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _191_
timestamp 1659391890
transform 1 0 6164 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 1659391890
transform 1 0 9292 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 9108 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1659391890
transform 1 0 1196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _195_
timestamp 1659391890
transform 1 0 8832 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1659391890
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _197_
timestamp 1659391890
transform 1 0 6624 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _198_
timestamp 1659391890
transform 1 0 8372 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _199_
timestamp 1659391890
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _200_
timestamp 1659391890
transform 1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _201_
timestamp 1659391890
transform 1 0 3588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _202_
timestamp 1659391890
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _203_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 8280 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _204_
timestamp 1659391890
transform 1 0 9200 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 8740 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _206_
timestamp 1659391890
transform 1 0 8740 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _207_
timestamp 1659391890
transform 1 0 8740 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 1659391890
transform 1 0 8648 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 7636 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfbbn_1  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 6808 0 -1 10880
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _211_
timestamp 1659391890
transform 1 0 4508 0 1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _212_
timestamp 1659391890
transform 1 0 5888 0 1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _213_
timestamp 1659391890
transform 1 0 6808 0 -1 8704
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _214_
timestamp 1659391890
transform 1 0 2576 0 -1 7616
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _215_
timestamp 1659391890
transform 1 0 2668 0 -1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _216_
timestamp 1659391890
transform 1 0 3036 0 -1 9792
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _217_
timestamp 1659391890
transform 1 0 6716 0 -1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _218_
timestamp 1659391890
transform 1 0 5796 0 -1 4352
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _219_
timestamp 1659391890
transform 1 0 6440 0 1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _220_
timestamp 1659391890
transform 1 0 3588 0 -1 3264
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _221_
timestamp 1659391890
transform 1 0 3956 0 -1 5440
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbn_1  _222_
timestamp 1659391890
transform 1 0 4508 0 1 6528
box -38 -48 2430 592
use sky130_fd_sc_hd__dfrtp_1  _223_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 7728 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _224_
timestamp 1659391890
transform 1 0 1656 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _225_
timestamp 1659391890
transform 1 0 2852 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _226_
timestamp 1659391890
transform 1 0 1196 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _227_
timestamp 1659391890
transform 1 0 1656 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _228_
timestamp 1659391890
transform 1 0 1656 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _229_
timestamp 1659391890
transform 1 0 3312 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _230_
timestamp 1659391890
transform 1 0 3588 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _231_
timestamp 1659391890
transform 1 0 3772 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _232_
timestamp 1659391890
transform 1 0 6256 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _233_
timestamp 1659391890
transform 1 0 6624 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _234_
timestamp 1659391890
transform 1 0 6348 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _235_
timestamp 1659391890
transform 1 0 5796 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 5612 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_clock
timestamp 1659391890
transform 1 0 7912 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 9200 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 7912 0 1 2176
box -38 -48 1694 592
use gpio_logic_high  gpio_logic_high
timestamp 1638030917
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1659391890
transform 1 0 3588 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1659391890
transform 1 0 3588 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1659391890
transform 1 0 5336 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1659391890
transform 1 0 6900 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1659391890
transform 1 0 8280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1659391890
transform 1 0 1196 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1659391890
transform 1 0 8280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1659391890
transform 1 0 3496 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1659391890
transform 1 0 4692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1659391890
transform 1 0 8832 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1659391890
transform 1 0 5060 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1659391890
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1659391890
transform 1 0 5704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1659391890
transform 1 0 4416 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1659391890
transform 1 0 3496 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1659391890
transform 1 0 6624 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1659391890
transform 1 0 3588 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1659391890
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1659391890
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1659391890
transform 1 0 3312 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1659391890
transform 1 0 5520 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1659391890
transform 1 0 3864 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1659391890
transform 1 0 4140 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1659391890
transform 1 0 5244 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1659391890
transform 1 0 4416 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1659391890
transform 1 0 5704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1659391890
transform 1 0 4692 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1659391890
transform 1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1659391890
transform 1 0 4968 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1659391890
transform 1 0 5244 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1659391890
transform 1 0 3588 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1659391890
transform 1 0 8648 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1659391890
transform 1 0 8372 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1659391890
transform 1 0 6808 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1659391890
transform 1 0 8740 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1659391890
transform 1 0 4692 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1659391890
transform 1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1659391890
transform 1 0 3864 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1659391890
transform 1 0 7820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1659391890
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1659391890
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1659391890
transform 1 0 9200 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1659391890
transform 1 0 8464 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1659391890
transform 1 0 7820 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1659391890
transform 1 0 9200 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1659391890
transform 1 0 8280 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1659391890
transform 1 0 4968 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1659391890
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1659391890
transform 1 0 9200 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1659391890
transform 1 0 8280 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1659391890
transform 1 0 8832 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1659391890
transform 1 0 7912 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output35
timestamp 1659391890
transform 1 0 4968 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1659391890
transform 1 0 7544 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output37
timestamp 1659391890
transform 1 0 5980 0 1 1088
box -38 -48 314 592
<< labels >>
rlabel metal2 s 938 12200 994 13000 6 gpio_defaults[0]
port 0 nsew signal input
rlabel metal2 s 5538 12200 5594 13000 6 gpio_defaults[10]
port 1 nsew signal input
rlabel metal2 s 5998 12200 6054 13000 6 gpio_defaults[11]
port 2 nsew signal input
rlabel metal2 s 6458 12200 6514 13000 6 gpio_defaults[12]
port 3 nsew signal input
rlabel metal2 s 1398 12200 1454 13000 6 gpio_defaults[1]
port 4 nsew signal input
rlabel metal2 s 1858 12200 1914 13000 6 gpio_defaults[2]
port 5 nsew signal input
rlabel metal2 s 2318 12200 2374 13000 6 gpio_defaults[3]
port 6 nsew signal input
rlabel metal2 s 2778 12200 2834 13000 6 gpio_defaults[4]
port 7 nsew signal input
rlabel metal2 s 3238 12200 3294 13000 6 gpio_defaults[5]
port 8 nsew signal input
rlabel metal2 s 3698 12200 3754 13000 6 gpio_defaults[6]
port 9 nsew signal input
rlabel metal2 s 4158 12200 4214 13000 6 gpio_defaults[7]
port 10 nsew signal input
rlabel metal2 s 4618 12200 4674 13000 6 gpio_defaults[8]
port 11 nsew signal input
rlabel metal2 s 5078 12200 5134 13000 6 gpio_defaults[9]
port 12 nsew signal input
rlabel metal3 s 14000 824 34000 944 6 mgmt_gpio_in
port 13 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 14 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 15 nsew signal input
rlabel metal3 s 14000 1232 34000 1352 6 one
port 16 nsew signal tristate
rlabel metal3 s 14000 2456 34000 2576 6 pad_gpio_ana_en
port 17 nsew signal tristate
rlabel metal3 s 14000 2864 34000 2984 6 pad_gpio_ana_pol
port 18 nsew signal tristate
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_sel
port 19 nsew signal tristate
rlabel metal3 s 14000 3680 34000 3800 6 pad_gpio_dm[0]
port 20 nsew signal tristate
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[1]
port 21 nsew signal tristate
rlabel metal3 s 14000 4496 34000 4616 6 pad_gpio_dm[2]
port 22 nsew signal tristate
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_holdover
port 23 nsew signal tristate
rlabel metal3 s 14000 5312 34000 5432 6 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
rlabel metal3 s 14000 5720 34000 5840 6 pad_gpio_in
port 25 nsew signal input
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_inenb
port 26 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_out
port 27 nsew signal tristate
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_outenb
port 28 nsew signal tristate
rlabel metal3 s 14000 7352 34000 7472 6 pad_gpio_slow_sel
port 29 nsew signal tristate
rlabel metal3 s 14000 7760 34000 7880 6 pad_gpio_vtrip_sel
port 30 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 resetn
port 31 nsew signal input
rlabel metal3 s 14000 8576 34000 8696 6 resetn_out
port 32 nsew signal tristate
rlabel metal3 s 14000 8984 34000 9104 6 serial_clock
port 33 nsew signal input
rlabel metal3 s 14000 9392 34000 9512 6 serial_clock_out
port 34 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 serial_data_in
port 35 nsew signal input
rlabel metal3 s 14000 10616 34000 10736 6 serial_load
port 37 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_load_out
port 38 nsew signal tristate
rlabel metal3 s 14000 11432 34000 11552 6 user_gpio_in
port 39 nsew signal tristate
rlabel metal3 s 14000 11840 34000 11960 6 user_gpio_oeb
port 40 nsew signal input
rlabel metal3 s 14000 12248 34000 12368 6 user_gpio_out
port 41 nsew signal input
rlabel metal5 s 920 1180 9844 1500 6 vccd
port 42 nsew power input
rlabel metal5 s 920 4560 9844 4880 6 vccd
port 42 nsew power input
rlabel metal5 s 920 7940 9844 8260 6 vccd
port 42 nsew power input
rlabel metal4 s 2560 1088 2880 11472 6 vccd
port 42 nsew power input
rlabel metal4 s 7560 1040 7880 11472 6 vccd
port 42 nsew power input
rlabel metal5 s 920 2228 9844 2548 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 5608 9844 5928 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 8988 9844 9308 6 vccd1
port 43 nsew power input
rlabel metal4 s 3560 1088 3880 11424 6 vccd1
port 43 nsew power input
rlabel metal4 s 8560 1088 8880 11424 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 2870 9844 3190 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 6250 9844 6570 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 9630 9844 9950 6 vssd
port 44 nsew ground input
rlabel metal4 s 5060 1040 5380 11472 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 3918 9844 4238 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 7298 9844 7618 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 10678 9844 10998 6 vssd1
port 45 nsew ground input
rlabel metal4 s 6060 1088 6380 11424 6 vssd1
port 45 nsew ground input
rlabel metal3 s 14000 416 34000 536 6 zero
port 46 nsew signal tristate
rlabel metal3 s 14000 10208 34000 10328 6 serial_data_out
port 36 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
