magic
tech sky130A
magscale 1 2
timestamp 1637791793
<< isosubstrate >>
rect 707553 886338 709093 889314
rect 8741 806938 10281 809914
rect 8741 763738 10281 766714
rect 8741 720538 10281 723514
rect 707553 705738 709093 708714
rect 8741 677338 10281 680314
rect 707553 660538 709093 663514
rect 8741 634138 10281 637114
rect 707553 615538 709093 618514
rect 8741 590938 10281 593914
rect 707553 570338 709093 573314
rect 8741 547738 10281 550714
rect 707553 525338 709093 528314
rect 707553 481338 709093 484314
rect 8741 420138 10281 423114
rect 707553 393138 709093 396114
rect 8741 376938 10281 379914
rect 707553 347938 709093 350914
rect 8741 333738 10281 336714
rect 707553 302938 709093 305914
rect 8741 290538 10281 293514
rect 707553 257938 709093 260914
rect 8741 247338 10281 250314
rect 193956 239226 214438 241244
rect 263310 241106 334156 246966
rect 386584 241220 387574 242376
rect 394166 241200 394996 242362
rect 707553 212738 709093 215714
rect 8741 204138 10281 207114
rect 707553 167738 709093 170714
rect 707553 122538 709093 125514
rect 142084 47031 145468 49885
rect 650094 46832 661434 55344
<< metal1 >>
rect 483566 1004640 483572 1004692
rect 483624 1004680 483630 1004692
rect 483624 1004652 518496 1004680
rect 483624 1004640 483630 1004652
rect 655514 896996 655520 897048
rect 655572 897036 655578 897048
rect 676030 897036 676036 897048
rect 655572 897008 676036 897036
rect 655572 896996 655578 897008
rect 676030 896996 676036 897008
rect 676088 896996 676094 897048
rect 673362 894616 673368 894668
rect 673420 894656 673426 894668
rect 675846 894656 675852 894668
rect 673420 894628 675852 894656
rect 673420 894616 673426 894628
rect 675846 894616 675852 894628
rect 675904 894616 675910 894668
rect 655422 894480 655428 894532
rect 655480 894520 655486 894532
rect 676030 894520 676036 894532
rect 655480 894492 676036 894520
rect 655480 894480 655486 894492
rect 676030 894480 676036 894492
rect 676088 894480 676094 894532
rect 670510 894412 670516 894464
rect 670568 894452 670574 894464
rect 676122 894452 676128 894464
rect 670568 894424 676128 894452
rect 670568 894412 670574 894424
rect 676122 894412 676128 894424
rect 676180 894412 676186 894464
rect 655698 894344 655704 894396
rect 655756 894384 655762 894396
rect 675938 894384 675944 894396
rect 655756 894356 675944 894384
rect 655756 894344 655762 894356
rect 675938 894344 675944 894356
rect 675996 894344 676002 894396
rect 670602 893800 670608 893852
rect 670660 893840 670666 893852
rect 676030 893840 676036 893852
rect 670660 893812 676036 893840
rect 670660 893800 670666 893812
rect 676030 893800 676036 893812
rect 676088 893800 676094 893852
rect 670418 892984 670424 893036
rect 670476 893024 670482 893036
rect 676030 893024 676036 893036
rect 670476 892996 676036 893024
rect 670476 892984 670482 892996
rect 676030 892984 676036 892996
rect 676088 892984 676094 893036
rect 674282 891488 674288 891540
rect 674340 891528 674346 891540
rect 676030 891528 676036 891540
rect 674340 891500 676036 891528
rect 674340 891488 674346 891500
rect 676030 891488 676036 891500
rect 676088 891488 676094 891540
rect 674742 890672 674748 890724
rect 674800 890712 674806 890724
rect 676030 890712 676036 890724
rect 674800 890684 676036 890712
rect 674800 890672 674806 890684
rect 676030 890672 676036 890684
rect 676088 890672 676094 890724
rect 674558 888768 674564 888820
rect 674616 888808 674622 888820
rect 675938 888808 675944 888820
rect 674616 888780 675944 888808
rect 674616 888768 674622 888780
rect 675938 888768 675944 888780
rect 675996 888768 676002 888820
rect 675018 888700 675024 888752
rect 675076 888740 675082 888752
rect 676030 888740 676036 888752
rect 675076 888712 676036 888740
rect 675076 888700 675082 888712
rect 676030 888700 676036 888712
rect 676088 888700 676094 888752
rect 673822 887816 673828 887868
rect 673880 887856 673886 887868
rect 676030 887856 676036 887868
rect 673880 887828 676036 887856
rect 673880 887816 673886 887828
rect 676030 887816 676036 887828
rect 676088 887816 676094 887868
rect 673730 886048 673736 886100
rect 673788 886088 673794 886100
rect 675938 886088 675944 886100
rect 673788 886060 675944 886088
rect 673788 886048 673794 886060
rect 675938 886048 675944 886060
rect 675996 886048 676002 886100
rect 674466 885980 674472 886032
rect 674524 886020 674530 886032
rect 676030 886020 676036 886032
rect 674524 885992 676036 886020
rect 674524 885980 674530 885992
rect 676030 885980 676036 885992
rect 676088 885980 676094 886032
rect 655606 883260 655612 883312
rect 655664 883300 655670 883312
rect 675386 883300 675392 883312
rect 655664 883272 675392 883300
rect 655664 883260 655670 883272
rect 675386 883260 675392 883272
rect 675444 883260 675450 883312
rect 671982 883192 671988 883244
rect 672040 883232 672046 883244
rect 679526 883232 679532 883244
rect 672040 883204 679532 883232
rect 672040 883192 672046 883204
rect 679526 883192 679532 883204
rect 679584 883192 679590 883244
rect 675294 883124 675300 883176
rect 675352 883164 675358 883176
rect 678974 883164 678980 883176
rect 675352 883136 678980 883164
rect 675352 883124 675358 883136
rect 678974 883124 678980 883136
rect 679032 883124 679038 883176
rect 675754 883056 675760 883108
rect 675812 883096 675818 883108
rect 679342 883096 679348 883108
rect 675812 883068 679348 883096
rect 675812 883056 675818 883068
rect 679342 883056 679348 883068
rect 679400 883056 679406 883108
rect 674834 882988 674840 883040
rect 674892 883028 674898 883040
rect 679618 883028 679624 883040
rect 674892 883000 679624 883028
rect 674892 882988 674898 883000
rect 679618 882988 679624 883000
rect 679676 882988 679682 883040
rect 674926 880404 674932 880456
rect 674984 880444 674990 880456
rect 679066 880444 679072 880456
rect 674984 880416 679072 880444
rect 674984 880404 674990 880416
rect 679066 880404 679072 880416
rect 679124 880404 679130 880456
rect 675202 880336 675208 880388
rect 675260 880376 675266 880388
rect 679158 880376 679164 880388
rect 675260 880348 679164 880376
rect 675260 880336 675266 880348
rect 679158 880336 679164 880348
rect 679216 880336 679222 880388
rect 675110 880268 675116 880320
rect 675168 880308 675174 880320
rect 679250 880308 679256 880320
rect 675168 880280 679256 880308
rect 675168 880268 675174 880280
rect 679250 880268 679256 880280
rect 679308 880268 679314 880320
rect 674650 880200 674656 880252
rect 674708 880240 674714 880252
rect 679434 880240 679440 880252
rect 674708 880212 679440 880240
rect 674708 880200 674714 880212
rect 679434 880200 679440 880212
rect 679492 880200 679498 880252
rect 675754 878364 675760 878416
rect 675812 878364 675818 878416
rect 675772 877804 675800 878364
rect 675754 877752 675760 877804
rect 675812 877752 675818 877804
rect 674834 877276 674840 877328
rect 674892 877316 674898 877328
rect 675294 877316 675300 877328
rect 674892 877288 675300 877316
rect 674892 877276 674898 877288
rect 675294 877276 675300 877288
rect 675352 877276 675358 877328
rect 674650 873740 674656 873792
rect 674708 873780 674714 873792
rect 675110 873780 675116 873792
rect 674708 873752 675116 873780
rect 674708 873740 674714 873752
rect 675110 873740 675116 873752
rect 675168 873740 675174 873792
rect 673730 873604 673736 873656
rect 673788 873644 673794 873656
rect 674650 873644 674656 873656
rect 673788 873616 674656 873644
rect 673788 873604 673794 873616
rect 674650 873604 674656 873616
rect 674708 873604 674714 873656
rect 675018 872720 675024 872772
rect 675076 872720 675082 872772
rect 675036 872568 675064 872720
rect 675018 872516 675024 872568
rect 675076 872516 675082 872568
rect 674742 872448 674748 872500
rect 674800 872488 674806 872500
rect 675202 872488 675208 872500
rect 674800 872460 675208 872488
rect 674800 872448 674806 872460
rect 675202 872448 675208 872460
rect 675260 872448 675266 872500
rect 673822 872312 673828 872364
rect 673880 872352 673886 872364
rect 674742 872352 674748 872364
rect 673880 872324 674748 872352
rect 673880 872312 673886 872324
rect 674742 872312 674748 872324
rect 674800 872312 674806 872364
rect 655790 872176 655796 872228
rect 655848 872216 655854 872228
rect 675110 872216 675116 872228
rect 655848 872188 675116 872216
rect 655848 872176 655854 872188
rect 675110 872176 675116 872188
rect 675168 872176 675174 872228
rect 674466 869932 674472 869984
rect 674524 869972 674530 869984
rect 675202 869972 675208 869984
rect 674524 869944 675208 869972
rect 674524 869932 674530 869944
rect 675202 869932 675208 869944
rect 675260 869932 675266 869984
rect 674742 869388 674748 869440
rect 674800 869428 674806 869440
rect 675202 869428 675208 869440
rect 674800 869400 675208 869428
rect 674800 869388 674806 869400
rect 675202 869388 675208 869400
rect 675260 869388 675266 869440
rect 674650 868708 674656 868760
rect 674708 868748 674714 868760
rect 675202 868748 675208 868760
rect 674708 868720 675208 868748
rect 674708 868708 674714 868720
rect 675202 868708 675208 868720
rect 675260 868708 675266 868760
rect 674558 867552 674564 867604
rect 674616 867592 674622 867604
rect 675110 867592 675116 867604
rect 674616 867564 675116 867592
rect 674616 867552 674622 867564
rect 675110 867552 675116 867564
rect 675168 867552 675174 867604
rect 674282 865716 674288 865768
rect 674340 865756 674346 865768
rect 675202 865756 675208 865768
rect 674340 865728 675208 865756
rect 674340 865716 674346 865728
rect 675202 865716 675208 865728
rect 675260 865716 675266 865768
rect 656802 863812 656808 863864
rect 656860 863852 656866 863864
rect 675110 863852 675116 863864
rect 656860 863824 675116 863852
rect 656860 863812 656866 863824
rect 675110 863812 675116 863824
rect 675168 863812 675174 863864
rect 41782 817640 41788 817692
rect 41840 817680 41846 817692
rect 50982 817680 50988 817692
rect 41840 817652 50988 817680
rect 41840 817640 41846 817652
rect 50982 817640 50988 817652
rect 51040 817640 51046 817692
rect 41782 817232 41788 817284
rect 41840 817272 41846 817284
rect 48314 817272 48320 817284
rect 41840 817244 48320 817272
rect 41840 817232 41846 817244
rect 48314 817232 48320 817244
rect 48372 817232 48378 817284
rect 41782 808256 41788 808308
rect 41840 808296 41846 808308
rect 43530 808296 43536 808308
rect 41840 808268 43536 808296
rect 41840 808256 41846 808268
rect 43530 808256 43536 808268
rect 43588 808256 43594 808308
rect 42334 805944 42340 805996
rect 42392 805984 42398 805996
rect 62114 805984 62120 805996
rect 42392 805956 62120 805984
rect 42392 805944 42398 805956
rect 62114 805944 62120 805956
rect 62172 805944 62178 805996
rect 41874 805876 41880 805928
rect 41932 805916 41938 805928
rect 43346 805916 43352 805928
rect 41932 805888 43352 805916
rect 41932 805876 41938 805888
rect 43346 805876 43352 805888
rect 43404 805876 43410 805928
rect 41966 804244 41972 804296
rect 42024 804284 42030 804296
rect 43254 804284 43260 804296
rect 42024 804256 43260 804284
rect 42024 804244 42030 804256
rect 43254 804244 43260 804256
rect 43312 804244 43318 804296
rect 42334 800436 42340 800488
rect 42392 800476 42398 800488
rect 58250 800476 58256 800488
rect 42392 800448 58256 800476
rect 42392 800436 42398 800448
rect 58250 800436 58256 800448
rect 58308 800436 58314 800488
rect 42242 799280 42248 799332
rect 42300 799320 42306 799332
rect 42702 799320 42708 799332
rect 42300 799292 42708 799320
rect 42300 799280 42306 799292
rect 42702 799280 42708 799292
rect 42760 799280 42766 799332
rect 42334 796832 42340 796884
rect 42392 796872 42398 796884
rect 42610 796872 42616 796884
rect 42392 796844 42616 796872
rect 42392 796832 42398 796844
rect 42610 796832 42616 796844
rect 42668 796832 42674 796884
rect 42242 794996 42248 795048
rect 42300 795036 42306 795048
rect 42886 795036 42892 795048
rect 42300 795008 42892 795036
rect 42300 794996 42306 795008
rect 42886 794996 42892 795008
rect 42944 794996 42950 795048
rect 42702 794860 42708 794912
rect 42760 794900 42766 794912
rect 42886 794900 42892 794912
rect 42760 794872 42892 794900
rect 42760 794860 42766 794872
rect 42886 794860 42892 794872
rect 42944 794860 42950 794912
rect 42150 794248 42156 794300
rect 42208 794288 42214 794300
rect 43254 794288 43260 794300
rect 42208 794260 43260 794288
rect 42208 794248 42214 794260
rect 43254 794248 43260 794260
rect 43312 794248 43318 794300
rect 42150 793772 42156 793824
rect 42208 793812 42214 793824
rect 43530 793812 43536 793824
rect 42208 793784 43536 793812
rect 42208 793772 42214 793784
rect 43530 793772 43536 793784
rect 43588 793772 43594 793824
rect 42242 792616 42248 792668
rect 42300 792656 42306 792668
rect 43070 792656 43076 792668
rect 42300 792628 43076 792656
rect 42300 792616 42306 792628
rect 43070 792616 43076 792628
rect 43128 792616 43134 792668
rect 655514 792140 655520 792192
rect 655572 792180 655578 792192
rect 675386 792180 675392 792192
rect 655572 792152 675392 792180
rect 655572 792140 655578 792152
rect 675386 792140 675392 792152
rect 675444 792140 675450 792192
rect 42150 790644 42156 790696
rect 42208 790684 42214 790696
rect 43346 790684 43352 790696
rect 42208 790656 43352 790684
rect 42208 790644 42214 790656
rect 43346 790644 43352 790656
rect 43404 790644 43410 790696
rect 42150 790100 42156 790152
rect 42208 790140 42214 790152
rect 43898 790140 43904 790152
rect 42208 790112 43904 790140
rect 42208 790100 42214 790112
rect 43898 790100 43904 790112
rect 43956 790100 43962 790152
rect 42334 789352 42340 789404
rect 42392 789392 42398 789404
rect 58066 789392 58072 789404
rect 42392 789364 58072 789392
rect 42392 789352 42398 789364
rect 58066 789352 58072 789364
rect 58124 789352 58130 789404
rect 42426 789284 42432 789336
rect 42484 789324 42490 789336
rect 58526 789324 58532 789336
rect 42484 789296 58532 789324
rect 42484 789284 42490 789296
rect 58526 789284 58532 789296
rect 58584 789284 58590 789336
rect 42150 789216 42156 789268
rect 42208 789256 42214 789268
rect 43806 789256 43812 789268
rect 42208 789228 43812 789256
rect 42208 789216 42214 789228
rect 43806 789216 43812 789228
rect 43864 789216 43870 789268
rect 42150 788808 42156 788860
rect 42208 788848 42214 788860
rect 42886 788848 42892 788860
rect 42208 788820 42892 788848
rect 42208 788808 42214 788820
rect 42886 788808 42892 788820
rect 42944 788808 42950 788860
rect 42150 786972 42156 787024
rect 42208 787012 42214 787024
rect 43438 787012 43444 787024
rect 42208 786984 43444 787012
rect 42208 786972 42214 786984
rect 43438 786972 43444 786984
rect 43496 786972 43502 787024
rect 48314 786564 48320 786616
rect 48372 786604 48378 786616
rect 58434 786604 58440 786616
rect 48372 786576 58440 786604
rect 48372 786564 48378 786576
rect 58434 786564 58440 786576
rect 58492 786564 58498 786616
rect 50982 786496 50988 786548
rect 51040 786536 51046 786548
rect 58526 786536 58532 786548
rect 51040 786508 58532 786536
rect 51040 786496 51046 786508
rect 58526 786496 58532 786508
rect 58584 786496 58590 786548
rect 42058 786224 42064 786276
rect 42116 786264 42122 786276
rect 43714 786264 43720 786276
rect 42116 786236 43720 786264
rect 42116 786224 42122 786236
rect 43714 786224 43720 786236
rect 43772 786224 43778 786276
rect 673730 784728 673736 784780
rect 673788 784768 673794 784780
rect 675110 784768 675116 784780
rect 673788 784740 675116 784768
rect 673788 784728 673794 784740
rect 675110 784728 675116 784740
rect 675168 784728 675174 784780
rect 656526 783844 656532 783896
rect 656584 783884 656590 783896
rect 674650 783884 674656 783896
rect 656584 783856 674656 783884
rect 656584 783844 656590 783856
rect 674650 783844 674656 783856
rect 674708 783844 674714 783896
rect 673638 780920 673644 780972
rect 673696 780960 673702 780972
rect 675202 780960 675208 780972
rect 673696 780932 675208 780960
rect 673696 780920 673702 780932
rect 675202 780920 675208 780932
rect 675260 780920 675266 780972
rect 674558 780104 674564 780156
rect 674616 780144 674622 780156
rect 675478 780144 675484 780156
rect 674616 780116 675484 780144
rect 674616 780104 674622 780116
rect 675478 780104 675484 780116
rect 675536 780104 675542 780156
rect 675018 780036 675024 780088
rect 675076 780036 675082 780088
rect 675036 779748 675064 780036
rect 675018 779696 675024 779748
rect 675076 779696 675082 779748
rect 674650 779560 674656 779612
rect 674708 779600 674714 779612
rect 675110 779600 675116 779612
rect 674708 779572 675116 779600
rect 674708 779560 674714 779572
rect 675110 779560 675116 779572
rect 675168 779560 675174 779612
rect 674282 779084 674288 779136
rect 674340 779124 674346 779136
rect 675202 779124 675208 779136
rect 674340 779096 675208 779124
rect 674340 779084 674346 779096
rect 675202 779084 675208 779096
rect 675260 779084 675266 779136
rect 673822 778608 673828 778660
rect 673880 778648 673886 778660
rect 675202 778648 675208 778660
rect 673880 778620 675208 778648
rect 673880 778608 673886 778620
rect 675202 778608 675208 778620
rect 675260 778608 675266 778660
rect 674466 777316 674472 777368
rect 674524 777356 674530 777368
rect 675386 777356 675392 777368
rect 674524 777328 675392 777356
rect 674524 777316 674530 777328
rect 675386 777316 675392 777328
rect 675444 777316 675450 777368
rect 654962 775480 654968 775532
rect 655020 775520 655026 775532
rect 675110 775520 675116 775532
rect 655020 775492 675116 775520
rect 655020 775480 655026 775492
rect 675110 775480 675116 775492
rect 675168 775480 675174 775532
rect 41506 774732 41512 774784
rect 41564 774772 41570 774784
rect 53742 774772 53748 774784
rect 41564 774744 53748 774772
rect 41564 774732 41570 774744
rect 53742 774732 53748 774744
rect 53800 774732 53806 774784
rect 41506 773848 41512 773900
rect 41564 773888 41570 773900
rect 50982 773888 50988 773900
rect 41564 773860 50988 773888
rect 41564 773848 41570 773860
rect 50982 773848 50988 773860
rect 51040 773848 51046 773900
rect 41506 773440 41512 773492
rect 41564 773480 41570 773492
rect 45462 773480 45468 773492
rect 41564 773452 45468 773480
rect 41564 773440 41570 773452
rect 45462 773440 45468 773452
rect 45520 773440 45526 773492
rect 675018 773372 675024 773424
rect 675076 773412 675082 773424
rect 675662 773412 675668 773424
rect 675076 773384 675668 773412
rect 675076 773372 675082 773384
rect 675662 773372 675668 773384
rect 675720 773372 675726 773424
rect 674742 773304 674748 773356
rect 674800 773344 674806 773356
rect 675754 773344 675760 773356
rect 674800 773316 675760 773344
rect 674800 773304 674806 773316
rect 675754 773304 675760 773316
rect 675812 773304 675818 773356
rect 674834 769632 674840 769684
rect 674892 769672 674898 769684
rect 675294 769672 675300 769684
rect 674892 769644 675300 769672
rect 674892 769632 674898 769644
rect 675294 769632 675300 769644
rect 675352 769632 675358 769684
rect 42426 767388 42432 767440
rect 42484 767428 42490 767440
rect 48222 767428 48228 767440
rect 42484 767400 48228 767428
rect 42484 767388 42490 767400
rect 48222 767388 48228 767400
rect 48280 767388 48286 767440
rect 38286 764464 38292 764516
rect 38344 764504 38350 764516
rect 42242 764504 42248 764516
rect 38344 764476 42248 764504
rect 38344 764464 38350 764476
rect 42242 764464 42248 764476
rect 42300 764464 42306 764516
rect 41598 762832 41604 762884
rect 41656 762872 41662 762884
rect 48314 762872 48320 762884
rect 41656 762844 48320 762872
rect 41656 762832 41662 762844
rect 48314 762832 48320 762844
rect 48372 762832 48378 762884
rect 38194 761676 38200 761728
rect 38252 761716 38258 761728
rect 42150 761716 42156 761728
rect 38252 761688 42156 761716
rect 38252 761676 38258 761688
rect 42150 761676 42156 761688
rect 42208 761676 42214 761728
rect 41506 759296 41512 759348
rect 41564 759336 41570 759348
rect 43530 759336 43536 759348
rect 41564 759308 43536 759336
rect 41564 759296 41570 759308
rect 43530 759296 43536 759308
rect 43588 759296 43594 759348
rect 42702 759092 42708 759144
rect 42760 759132 42766 759144
rect 43346 759132 43352 759144
rect 42760 759104 43352 759132
rect 42760 759092 42766 759104
rect 43346 759092 43352 759104
rect 43404 759092 43410 759144
rect 38562 758956 38568 759008
rect 38620 758996 38626 759008
rect 42702 758996 42708 759008
rect 38620 758968 42708 758996
rect 38620 758956 38626 758968
rect 42702 758956 42708 758968
rect 42760 758956 42766 759008
rect 43898 757732 43904 757784
rect 43956 757772 43962 757784
rect 44174 757772 44180 757784
rect 43956 757744 44180 757772
rect 43956 757732 43962 757744
rect 44174 757732 44180 757744
rect 44232 757732 44238 757784
rect 43622 757596 43628 757648
rect 43680 757636 43686 757648
rect 43898 757636 43904 757648
rect 43680 757608 43904 757636
rect 43680 757596 43686 757608
rect 43898 757596 43904 757608
rect 43956 757596 43962 757648
rect 42426 757460 42432 757512
rect 42484 757500 42490 757512
rect 43622 757500 43628 757512
rect 42484 757472 43628 757500
rect 42484 757460 42490 757472
rect 43622 757460 43628 757472
rect 43680 757460 43686 757512
rect 42150 756984 42156 757036
rect 42208 757024 42214 757036
rect 44266 757024 44272 757036
rect 42208 756996 44272 757024
rect 42208 756984 42214 756996
rect 44266 756984 44272 756996
rect 44324 756984 44330 757036
rect 42242 756236 42248 756288
rect 42300 756276 42306 756288
rect 59262 756276 59268 756288
rect 42300 756248 59268 756276
rect 42300 756236 42306 756248
rect 59262 756236 59268 756248
rect 59320 756236 59326 756288
rect 42150 754876 42156 754928
rect 42208 754916 42214 754928
rect 42334 754916 42340 754928
rect 42208 754888 42340 754916
rect 42208 754876 42214 754888
rect 42334 754876 42340 754888
rect 42392 754876 42398 754928
rect 42334 754264 42340 754316
rect 42392 754304 42398 754316
rect 43070 754304 43076 754316
rect 42392 754276 43076 754304
rect 42392 754264 42398 754276
rect 43070 754264 43076 754276
rect 43128 754264 43134 754316
rect 43162 754196 43168 754248
rect 43220 754196 43226 754248
rect 43180 753976 43208 754196
rect 43162 753924 43168 753976
rect 43220 753924 43226 753976
rect 42150 753312 42156 753364
rect 42208 753352 42214 753364
rect 43254 753352 43260 753364
rect 42208 753324 43260 753352
rect 42208 753312 42214 753324
rect 43254 753312 43260 753324
rect 43312 753312 43318 753364
rect 42150 753040 42156 753092
rect 42208 753080 42214 753092
rect 43162 753080 43168 753092
rect 42208 753052 43168 753080
rect 42208 753040 42214 753052
rect 43162 753040 43168 753052
rect 43220 753040 43226 753092
rect 42242 751748 42248 751800
rect 42300 751788 42306 751800
rect 42702 751788 42708 751800
rect 42300 751760 42708 751788
rect 42300 751748 42306 751760
rect 42702 751748 42708 751760
rect 42760 751748 42766 751800
rect 42242 751204 42248 751256
rect 42300 751244 42306 751256
rect 43346 751244 43352 751256
rect 42300 751216 43352 751244
rect 42300 751204 42306 751216
rect 43346 751204 43352 751216
rect 43404 751204 43410 751256
rect 42150 751068 42156 751120
rect 42208 751108 42214 751120
rect 43070 751108 43076 751120
rect 42208 751080 43076 751108
rect 42208 751068 42214 751080
rect 43070 751068 43076 751080
rect 43128 751068 43134 751120
rect 43346 751068 43352 751120
rect 43404 751108 43410 751120
rect 44082 751108 44088 751120
rect 43404 751080 44088 751108
rect 43404 751068 43410 751080
rect 44082 751068 44088 751080
rect 44140 751068 44146 751120
rect 42058 750592 42064 750644
rect 42116 750632 42122 750644
rect 43530 750632 43536 750644
rect 42116 750604 43536 750632
rect 42116 750592 42122 750604
rect 43530 750592 43536 750604
rect 43588 750592 43594 750644
rect 42242 749368 42248 749420
rect 42300 749408 42306 749420
rect 43806 749408 43812 749420
rect 42300 749380 43812 749408
rect 42300 749368 42306 749380
rect 43806 749368 43812 749380
rect 43864 749368 43870 749420
rect 655974 747940 655980 747992
rect 656032 747980 656038 747992
rect 675386 747980 675392 747992
rect 656032 747952 675392 747980
rect 656032 747940 656038 747952
rect 675386 747940 675392 747952
rect 675444 747940 675450 747992
rect 43254 747872 43260 747924
rect 43312 747912 43318 747924
rect 58434 747912 58440 747924
rect 43312 747884 58440 747912
rect 43312 747872 43318 747884
rect 58434 747872 58440 747884
rect 58492 747872 58498 747924
rect 42150 747464 42156 747516
rect 42208 747504 42214 747516
rect 43530 747504 43536 747516
rect 42208 747476 43536 747504
rect 42208 747464 42214 747476
rect 43530 747464 43536 747476
rect 43588 747464 43594 747516
rect 42242 746240 42248 746292
rect 42300 746280 42306 746292
rect 43990 746280 43996 746292
rect 42300 746252 43996 746280
rect 42300 746240 42306 746252
rect 43990 746240 43996 746252
rect 44048 746240 44054 746292
rect 42426 745220 42432 745272
rect 42484 745260 42490 745272
rect 58434 745260 58440 745272
rect 42484 745232 58440 745260
rect 42484 745220 42490 745232
rect 58434 745220 58440 745232
rect 58492 745220 58498 745272
rect 45462 745152 45468 745204
rect 45520 745192 45526 745204
rect 58526 745192 58532 745204
rect 45520 745164 58532 745192
rect 45520 745152 45526 745164
rect 58526 745152 58532 745164
rect 58584 745152 58590 745204
rect 42334 745084 42340 745136
rect 42392 745124 42398 745136
rect 43346 745124 43352 745136
rect 42392 745096 43352 745124
rect 42392 745084 42398 745096
rect 43346 745084 43352 745096
rect 43404 745084 43410 745136
rect 673546 744132 673552 744184
rect 673604 744172 673610 744184
rect 675754 744172 675760 744184
rect 673604 744144 675760 744172
rect 673604 744132 673610 744144
rect 675754 744132 675760 744144
rect 675812 744132 675818 744184
rect 42334 743248 42340 743300
rect 42392 743288 42398 743300
rect 43898 743288 43904 743300
rect 42392 743260 43904 743288
rect 42392 743248 42398 743260
rect 43898 743248 43904 743260
rect 43956 743248 43962 743300
rect 42150 743044 42156 743096
rect 42208 743084 42214 743096
rect 44082 743084 44088 743096
rect 42208 743056 44088 743084
rect 42208 743044 42214 743056
rect 44082 743044 44088 743056
rect 44140 743044 44146 743096
rect 50982 742364 50988 742416
rect 51040 742404 51046 742416
rect 58434 742404 58440 742416
rect 51040 742376 58440 742404
rect 51040 742364 51046 742376
rect 58434 742364 58440 742376
rect 58492 742364 58498 742416
rect 53742 742296 53748 742348
rect 53800 742336 53806 742348
rect 57974 742336 57980 742348
rect 53800 742308 57980 742336
rect 53800 742296 53806 742308
rect 57974 742296 57980 742308
rect 58032 742296 58038 742348
rect 674558 737264 674564 737316
rect 674616 737304 674622 737316
rect 675202 737304 675208 737316
rect 674616 737276 675208 737304
rect 674616 737264 674622 737276
rect 675202 737264 675208 737276
rect 675260 737264 675266 737316
rect 655146 736992 655152 737044
rect 655204 737032 655210 737044
rect 675202 737032 675208 737044
rect 655204 737004 675208 737032
rect 655204 736992 655210 737004
rect 675202 736992 675208 737004
rect 675260 736992 675266 737044
rect 656066 736924 656072 736976
rect 656124 736964 656130 736976
rect 674834 736964 674840 736976
rect 656124 736936 674840 736964
rect 656124 736924 656130 736936
rect 674834 736924 674840 736936
rect 674892 736924 674898 736976
rect 674650 735632 674656 735684
rect 674708 735672 674714 735684
rect 675386 735672 675392 735684
rect 674708 735644 675392 735672
rect 674708 735632 674714 735644
rect 675386 735632 675392 735644
rect 675444 735632 675450 735684
rect 674742 734748 674748 734800
rect 674800 734788 674806 734800
rect 675386 734788 675392 734800
rect 674800 734760 675392 734788
rect 674800 734748 674806 734760
rect 675386 734748 675392 734760
rect 675444 734748 675450 734800
rect 673822 734136 673828 734188
rect 673880 734176 673886 734188
rect 675386 734176 675392 734188
rect 673880 734148 675392 734176
rect 673880 734136 673886 734148
rect 675386 734136 675392 734148
rect 675444 734136 675450 734188
rect 673546 733864 673552 733916
rect 673604 733904 673610 733916
rect 675386 733904 675392 733916
rect 673604 733876 675392 733904
rect 673604 733864 673610 733876
rect 675386 733864 675392 733876
rect 675444 733864 675450 733916
rect 675294 733796 675300 733848
rect 675352 733796 675358 733848
rect 675312 733508 675340 733796
rect 675294 733456 675300 733508
rect 675352 733456 675358 733508
rect 673454 732300 673460 732352
rect 673512 732340 673518 732352
rect 675386 732340 675392 732352
rect 673512 732312 675392 732340
rect 673512 732300 673518 732312
rect 675386 732300 675392 732312
rect 675444 732300 675450 732352
rect 674834 732028 674840 732080
rect 674892 732068 674898 732080
rect 675386 732068 675392 732080
rect 674892 732040 675392 732068
rect 674892 732028 674898 732040
rect 675386 732028 675392 732040
rect 675444 732028 675450 732080
rect 41506 731076 41512 731128
rect 41564 731116 41570 731128
rect 43622 731116 43628 731128
rect 41564 731088 43628 731116
rect 41564 731076 41570 731088
rect 43622 731076 43628 731088
rect 43680 731076 43686 731128
rect 674742 730464 674748 730516
rect 674800 730504 674806 730516
rect 675386 730504 675392 730516
rect 674800 730476 675392 730504
rect 674800 730464 674806 730476
rect 675386 730464 675392 730476
rect 675444 730464 675450 730516
rect 674650 728804 674656 728816
rect 674576 728776 674656 728804
rect 674576 728192 674604 728776
rect 674650 728764 674656 728776
rect 674708 728764 674714 728816
rect 674650 728628 674656 728680
rect 674708 728668 674714 728680
rect 675386 728668 675392 728680
rect 674708 728640 675392 728668
rect 674708 728628 674714 728640
rect 675386 728628 675392 728640
rect 675444 728628 675450 728680
rect 674484 728164 674604 728192
rect 674484 727988 674512 728164
rect 674558 728084 674564 728136
rect 674616 728124 674622 728136
rect 676122 728124 676128 728136
rect 674616 728096 676128 728124
rect 674616 728084 674622 728096
rect 676122 728084 676128 728096
rect 676180 728084 676186 728136
rect 675202 728016 675208 728068
rect 675260 728056 675266 728068
rect 678974 728056 678980 728068
rect 675260 728028 678980 728056
rect 675260 728016 675266 728028
rect 678974 728016 678980 728028
rect 679032 728016 679038 728068
rect 674558 727988 674564 728000
rect 674484 727960 674564 727988
rect 674558 727948 674564 727960
rect 674616 727948 674622 728000
rect 673270 727880 673276 727932
rect 673328 727920 673334 727932
rect 675202 727920 675208 727932
rect 673328 727892 675208 727920
rect 673328 727880 673334 727892
rect 675202 727880 675208 727892
rect 675260 727880 675266 727932
rect 674834 727812 674840 727864
rect 674892 727852 674898 727864
rect 675110 727852 675116 727864
rect 674892 727824 675116 727852
rect 674892 727812 674898 727824
rect 675110 727812 675116 727824
rect 675168 727812 675174 727864
rect 673546 718836 673552 718888
rect 673604 718876 673610 718888
rect 675570 718876 675576 718888
rect 673604 718848 675576 718876
rect 673604 718836 673610 718848
rect 675570 718836 675576 718848
rect 675628 718836 675634 718888
rect 673454 718700 673460 718752
rect 673512 718740 673518 718752
rect 674650 718740 674656 718752
rect 673512 718712 674656 718740
rect 673512 718700 673518 718712
rect 674650 718700 674656 718712
rect 674708 718700 674714 718752
rect 41506 717612 41512 717664
rect 41564 717652 41570 717664
rect 53742 717652 53748 717664
rect 41564 717624 53748 717652
rect 41564 717612 41570 717624
rect 53742 717612 53748 717624
rect 53800 717612 53806 717664
rect 41414 717476 41420 717528
rect 41472 717516 41478 717528
rect 43530 717516 43536 717528
rect 41472 717488 43536 717516
rect 41472 717476 41478 717488
rect 43530 717476 43536 717488
rect 43588 717476 43594 717528
rect 670510 715408 670516 715420
rect 670508 715380 670516 715408
rect 670510 715368 670516 715380
rect 670568 715408 670574 715420
rect 676030 715408 676036 715420
rect 670568 715380 676036 715408
rect 670568 715368 670574 715380
rect 676030 715368 676036 715380
rect 676088 715368 676094 715420
rect 655790 715232 655796 715284
rect 655848 715272 655854 715284
rect 675938 715272 675944 715284
rect 655848 715244 675944 715272
rect 655848 715232 655854 715244
rect 675938 715232 675944 715244
rect 675996 715232 676002 715284
rect 655606 715096 655612 715148
rect 655664 715136 655670 715148
rect 675754 715136 675760 715148
rect 655664 715108 675760 715136
rect 655664 715096 655670 715108
rect 675754 715096 675760 715108
rect 675812 715096 675818 715148
rect 655422 714960 655428 715012
rect 655480 715000 655486 715012
rect 675846 715000 675852 715012
rect 655480 714972 675852 715000
rect 655480 714960 655486 714972
rect 675846 714960 675852 714972
rect 675904 714960 675910 715012
rect 675202 714892 675208 714944
rect 675260 714932 675266 714944
rect 675754 714932 675760 714944
rect 675260 714904 675760 714932
rect 675260 714892 675266 714904
rect 675754 714892 675760 714904
rect 675812 714892 675818 714944
rect 42426 714824 42432 714876
rect 42484 714864 42490 714876
rect 59354 714864 59360 714876
rect 42484 714836 59360 714864
rect 42484 714824 42490 714836
rect 59354 714824 59360 714836
rect 59412 714824 59418 714876
rect 670510 714824 670516 714876
rect 670568 714864 670574 714876
rect 676030 714864 676036 714876
rect 670568 714836 676036 714864
rect 670568 714824 670574 714836
rect 676030 714824 676036 714836
rect 676088 714824 676094 714876
rect 673362 714484 673368 714536
rect 673420 714524 673426 714536
rect 676030 714524 676036 714536
rect 673420 714496 676036 714524
rect 673420 714484 673426 714496
rect 676030 714484 676036 714496
rect 676088 714484 676094 714536
rect 43162 714144 43168 714196
rect 43220 714184 43226 714196
rect 44358 714184 44364 714196
rect 43220 714156 44364 714184
rect 43220 714144 43226 714156
rect 44358 714144 44364 714156
rect 44416 714144 44422 714196
rect 673270 714008 673276 714060
rect 673328 714048 673334 714060
rect 676030 714048 676036 714060
rect 673328 714020 676036 714048
rect 673328 714008 673334 714020
rect 676030 714008 676036 714020
rect 676088 714008 676094 714060
rect 41782 713804 41788 713856
rect 41840 713804 41846 713856
rect 41800 713584 41828 713804
rect 41782 713532 41788 713584
rect 41840 713532 41846 713584
rect 669866 713436 669872 713448
rect 669862 713408 669872 713436
rect 669866 713396 669872 713408
rect 669924 713436 669930 713448
rect 670418 713436 670424 713448
rect 669924 713408 670424 713436
rect 669924 713396 669930 713408
rect 670418 713396 670424 713408
rect 670476 713396 670482 713448
rect 676030 712552 676036 712564
rect 670666 712524 676036 712552
rect 670666 712428 670694 712524
rect 676030 712512 676036 712524
rect 676088 712512 676094 712564
rect 670602 712416 670608 712428
rect 670598 712388 670608 712416
rect 670602 712376 670608 712388
rect 670660 712388 670694 712428
rect 670660 712376 670666 712388
rect 669866 712308 669872 712360
rect 669924 712348 669930 712360
rect 675938 712348 675944 712360
rect 669924 712320 675944 712348
rect 669924 712308 669930 712320
rect 675938 712308 675944 712320
rect 675996 712308 676002 712360
rect 43806 712240 43812 712292
rect 43864 712280 43870 712292
rect 44266 712280 44272 712292
rect 43864 712252 44272 712280
rect 43864 712240 43870 712252
rect 44266 712240 44272 712252
rect 44324 712240 44330 712292
rect 670326 712240 670332 712292
rect 670384 712280 670390 712292
rect 676030 712280 676036 712292
rect 670384 712252 676036 712280
rect 670384 712240 670390 712252
rect 676030 712240 676036 712252
rect 676088 712240 676094 712292
rect 670418 712172 670424 712224
rect 670476 712212 670482 712224
rect 675846 712212 675852 712224
rect 670476 712184 675852 712212
rect 670476 712172 670482 712184
rect 675846 712172 675852 712184
rect 675904 712172 675910 712224
rect 43806 712104 43812 712156
rect 43864 712144 43870 712156
rect 59262 712144 59268 712156
rect 43864 712116 59268 712144
rect 43864 712104 43870 712116
rect 59262 712104 59268 712116
rect 59320 712104 59326 712156
rect 675018 712104 675024 712156
rect 675076 712144 675082 712156
rect 675938 712144 675944 712156
rect 675076 712116 675944 712144
rect 675076 712104 675082 712116
rect 675938 712104 675944 712116
rect 675996 712104 676002 712156
rect 42150 711696 42156 711748
rect 42208 711736 42214 711748
rect 43346 711736 43352 711748
rect 42208 711708 43352 711736
rect 42208 711696 42214 711708
rect 43346 711696 43352 711708
rect 43404 711696 43410 711748
rect 673730 711492 673736 711544
rect 673788 711532 673794 711544
rect 676030 711532 676036 711544
rect 673788 711504 676036 711532
rect 673788 711492 673794 711504
rect 676030 711492 676036 711504
rect 676088 711492 676094 711544
rect 42150 710880 42156 710932
rect 42208 710920 42214 710932
rect 42426 710920 42432 710932
rect 42208 710892 42432 710920
rect 42208 710880 42214 710892
rect 42426 710880 42432 710892
rect 42484 710880 42490 710932
rect 42334 710268 42340 710320
rect 42392 710308 42398 710320
rect 42702 710308 42708 710320
rect 42392 710280 42708 710308
rect 42392 710268 42398 710280
rect 42702 710268 42708 710280
rect 42760 710268 42766 710320
rect 42702 710132 42708 710184
rect 42760 710172 42766 710184
rect 43254 710172 43260 710184
rect 42760 710144 43260 710172
rect 42760 710132 42766 710144
rect 43254 710132 43260 710144
rect 43312 710132 43318 710184
rect 43438 709860 43444 709912
rect 43496 709900 43502 709912
rect 43898 709900 43904 709912
rect 43496 709872 43904 709900
rect 43496 709860 43502 709872
rect 43898 709860 43904 709872
rect 43956 709860 43962 709912
rect 43346 709792 43352 709844
rect 43404 709832 43410 709844
rect 43990 709832 43996 709844
rect 43404 709804 43996 709832
rect 43404 709792 43410 709804
rect 43990 709792 43996 709804
rect 44048 709792 44054 709844
rect 43990 709588 43996 709640
rect 44048 709628 44054 709640
rect 44266 709628 44272 709640
rect 44048 709600 44272 709628
rect 44048 709588 44054 709600
rect 44266 709588 44272 709600
rect 44324 709588 44330 709640
rect 44082 709520 44088 709572
rect 44140 709560 44146 709572
rect 44358 709560 44364 709572
rect 44140 709532 44364 709560
rect 44140 709520 44146 709532
rect 44358 709520 44364 709532
rect 44416 709520 44422 709572
rect 43806 709424 43812 709436
rect 42260 709396 43812 709424
rect 42260 709368 42288 709396
rect 43806 709384 43812 709396
rect 43864 709384 43870 709436
rect 42242 709316 42248 709368
rect 42300 709316 42306 709368
rect 674466 708840 674472 708892
rect 674524 708880 674530 708892
rect 676030 708880 676036 708892
rect 674524 708852 676036 708880
rect 674524 708840 674530 708852
rect 676030 708840 676036 708852
rect 676088 708840 676094 708892
rect 42150 708568 42156 708620
rect 42208 708608 42214 708620
rect 43622 708608 43628 708620
rect 42208 708580 43628 708608
rect 42208 708568 42214 708580
rect 43622 708568 43628 708580
rect 43680 708568 43686 708620
rect 674282 708228 674288 708280
rect 674340 708268 674346 708280
rect 676030 708268 676036 708280
rect 674340 708240 676036 708268
rect 674340 708228 674346 708240
rect 676030 708228 676036 708240
rect 676088 708228 676094 708280
rect 673638 707820 673644 707872
rect 673696 707860 673702 707872
rect 676030 707860 676036 707872
rect 673696 707832 676036 707860
rect 673696 707820 673702 707832
rect 676030 707820 676036 707832
rect 676088 707820 676094 707872
rect 42426 706732 42432 706784
rect 42484 706772 42490 706784
rect 43438 706772 43444 706784
rect 42484 706744 43444 706772
rect 42484 706732 42490 706744
rect 43438 706732 43444 706744
rect 43496 706732 43502 706784
rect 42242 706188 42248 706240
rect 42300 706228 42306 706240
rect 43530 706228 43536 706240
rect 42300 706200 43536 706228
rect 42300 706188 42306 706200
rect 43530 706188 43536 706200
rect 43588 706188 43594 706240
rect 42334 705916 42340 705968
rect 42392 705956 42398 705968
rect 43254 705956 43260 705968
rect 42392 705928 43260 705956
rect 42392 705916 42398 705928
rect 43254 705916 43260 705928
rect 43312 705916 43318 705968
rect 672074 705100 672080 705152
rect 672132 705140 672138 705152
rect 676030 705140 676036 705152
rect 672132 705112 676036 705140
rect 672132 705100 672138 705112
rect 676030 705100 676036 705112
rect 676088 705100 676094 705152
rect 42058 704216 42064 704268
rect 42116 704256 42122 704268
rect 42702 704256 42708 704268
rect 42116 704228 42708 704256
rect 42116 704216 42122 704228
rect 42702 704216 42708 704228
rect 42760 704216 42766 704268
rect 42426 703808 42432 703860
rect 42484 703848 42490 703860
rect 58526 703848 58532 703860
rect 42484 703820 58532 703848
rect 42484 703808 42490 703820
rect 58526 703808 58532 703820
rect 58584 703808 58590 703860
rect 655974 703808 655980 703860
rect 656032 703848 656038 703860
rect 675386 703848 675392 703860
rect 656032 703820 675392 703848
rect 656032 703808 656038 703820
rect 675386 703808 675392 703820
rect 675444 703808 675450 703860
rect 42334 702448 42340 702500
rect 42392 702488 42398 702500
rect 43346 702488 43352 702500
rect 42392 702460 43352 702488
rect 42392 702448 42398 702460
rect 43346 702448 43352 702460
rect 43404 702448 43410 702500
rect 42334 701904 42340 701956
rect 42392 701944 42398 701956
rect 43806 701944 43812 701956
rect 42392 701916 43812 701944
rect 42392 701904 42398 701916
rect 43806 701904 43812 701916
rect 43864 701904 43870 701956
rect 42242 701768 42248 701820
rect 42300 701808 42306 701820
rect 44082 701808 44088 701820
rect 42300 701780 44088 701808
rect 42300 701768 42306 701780
rect 44082 701768 44088 701780
rect 44140 701768 44146 701820
rect 42334 699388 42340 699440
rect 42392 699428 42398 699440
rect 43990 699428 43996 699440
rect 42392 699400 43996 699428
rect 42392 699388 42398 699400
rect 43990 699388 43996 699400
rect 44048 699388 44054 699440
rect 654226 692860 654232 692912
rect 654284 692900 654290 692912
rect 675202 692900 675208 692912
rect 654284 692872 675208 692900
rect 654284 692860 654290 692872
rect 675202 692860 675208 692872
rect 675260 692860 675266 692912
rect 673730 690140 673736 690192
rect 673788 690180 673794 690192
rect 675294 690180 675300 690192
rect 673788 690152 675300 690180
rect 673788 690140 673794 690152
rect 675294 690140 675300 690152
rect 675352 690140 675358 690192
rect 654134 690004 654140 690056
rect 654192 690044 654198 690056
rect 675294 690044 675300 690056
rect 654192 690016 675300 690044
rect 654192 690004 654198 690016
rect 675294 690004 675300 690016
rect 675352 690004 675358 690056
rect 673638 689120 673644 689172
rect 673696 689160 673702 689172
rect 675478 689160 675484 689172
rect 673696 689132 675484 689160
rect 673696 689120 673702 689132
rect 675478 689120 675484 689132
rect 675536 689120 675542 689172
rect 675202 688712 675208 688764
rect 675260 688752 675266 688764
rect 675478 688752 675484 688764
rect 675260 688724 675484 688752
rect 675260 688712 675266 688724
rect 675478 688712 675484 688724
rect 675536 688712 675542 688764
rect 673362 688576 673368 688628
rect 673420 688616 673426 688628
rect 675386 688616 675392 688628
rect 673420 688588 675392 688616
rect 673420 688576 673426 688588
rect 675386 688576 675392 688588
rect 675444 688576 675450 688628
rect 41506 688304 41512 688356
rect 41564 688344 41570 688356
rect 53834 688344 53840 688356
rect 41564 688316 53840 688344
rect 41564 688304 41570 688316
rect 53834 688304 53840 688316
rect 53892 688304 53898 688356
rect 673546 687828 673552 687880
rect 673604 687868 673610 687880
rect 675110 687868 675116 687880
rect 673604 687840 675116 687868
rect 673604 687828 673610 687840
rect 675110 687828 675116 687840
rect 675168 687828 675174 687880
rect 41782 687624 41788 687676
rect 41840 687664 41846 687676
rect 50982 687664 50988 687676
rect 41840 687636 50988 687664
rect 41840 687624 41846 687636
rect 50982 687624 50988 687636
rect 51040 687624 51046 687676
rect 674466 687284 674472 687336
rect 674524 687324 674530 687336
rect 675386 687324 675392 687336
rect 674524 687296 675392 687324
rect 674524 687284 674530 687296
rect 675386 687284 675392 687296
rect 675444 687284 675450 687336
rect 41782 687216 41788 687268
rect 41840 687256 41846 687268
rect 45738 687256 45744 687268
rect 41840 687228 45744 687256
rect 41840 687216 41846 687228
rect 45738 687216 45744 687228
rect 45796 687216 45802 687268
rect 675110 684224 675116 684276
rect 675168 684224 675174 684276
rect 675202 684224 675208 684276
rect 675260 684224 675266 684276
rect 675018 684020 675024 684072
rect 675076 684060 675082 684072
rect 675128 684060 675156 684224
rect 675076 684032 675156 684060
rect 675076 684020 675082 684032
rect 675220 683936 675248 684224
rect 674282 683884 674288 683936
rect 674340 683924 674346 683936
rect 675018 683924 675024 683936
rect 674340 683896 675024 683924
rect 674340 683884 674346 683896
rect 675018 683884 675024 683896
rect 675076 683884 675082 683936
rect 675202 683884 675208 683936
rect 675260 683884 675266 683936
rect 675110 683612 675116 683664
rect 675168 683652 675174 683664
rect 675386 683652 675392 683664
rect 675168 683624 675392 683652
rect 675168 683612 675174 683624
rect 675386 683612 675392 683624
rect 675444 683612 675450 683664
rect 673730 680348 673736 680400
rect 673788 680388 673794 680400
rect 674282 680388 674288 680400
rect 673788 680360 674288 680388
rect 673788 680348 673794 680360
rect 674282 680348 674288 680360
rect 674340 680348 674346 680400
rect 675294 678920 675300 678972
rect 675352 678960 675358 678972
rect 679066 678960 679072 678972
rect 675352 678932 679072 678960
rect 675352 678920 675358 678932
rect 679066 678920 679072 678932
rect 679124 678920 679130 678972
rect 41782 678580 41788 678632
rect 41840 678620 41846 678632
rect 44082 678620 44088 678632
rect 41840 678592 44088 678620
rect 41840 678580 41846 678592
rect 44082 678580 44088 678592
rect 44140 678580 44146 678632
rect 41782 676608 41788 676660
rect 41840 676648 41846 676660
rect 43162 676648 43168 676660
rect 41840 676620 43168 676648
rect 41840 676608 41846 676620
rect 43162 676608 43168 676620
rect 43220 676608 43226 676660
rect 5534 675724 5540 675776
rect 5592 675764 5598 675776
rect 30558 675764 30564 675776
rect 5592 675736 30564 675764
rect 5592 675724 5598 675736
rect 30558 675724 30564 675736
rect 30616 675724 30622 675776
rect 5442 674772 5448 674824
rect 5500 674812 5506 674824
rect 43346 674812 43352 674824
rect 5500 674784 43352 674812
rect 5500 674772 5506 674784
rect 43346 674772 43352 674784
rect 43404 674772 43410 674824
rect 43070 672528 43076 672580
rect 43128 672568 43134 672580
rect 43530 672568 43536 672580
rect 43128 672540 43536 672568
rect 43128 672528 43134 672540
rect 43530 672528 43536 672540
rect 43588 672528 43594 672580
rect 41874 672392 41880 672444
rect 41932 672432 41938 672444
rect 43070 672432 43076 672444
rect 41932 672404 43076 672432
rect 41932 672392 41938 672404
rect 43070 672392 43076 672404
rect 43128 672392 43134 672444
rect 43438 672120 43444 672172
rect 43496 672160 43502 672172
rect 43990 672160 43996 672172
rect 43496 672132 43996 672160
rect 43496 672120 43502 672132
rect 43990 672120 43996 672132
rect 44048 672120 44054 672172
rect 43254 671984 43260 672036
rect 43312 672024 43318 672036
rect 43438 672024 43444 672036
rect 43312 671996 43444 672024
rect 43312 671984 43318 671996
rect 43438 671984 43444 671996
rect 43496 671984 43502 672036
rect 42334 671780 42340 671832
rect 42392 671820 42398 671832
rect 43162 671820 43168 671832
rect 42392 671792 43168 671820
rect 42392 671780 42398 671792
rect 43162 671780 43168 671792
rect 43220 671780 43226 671832
rect 655882 670896 655888 670948
rect 655940 670936 655946 670948
rect 676214 670936 676220 670948
rect 655940 670908 676220 670936
rect 655940 670896 655946 670908
rect 676214 670896 676220 670908
rect 676272 670896 676278 670948
rect 43530 670828 43536 670880
rect 43588 670868 43594 670880
rect 43990 670868 43996 670880
rect 43588 670840 43996 670868
rect 43588 670828 43594 670840
rect 43990 670828 43996 670840
rect 44048 670828 44054 670880
rect 42334 670760 42340 670812
rect 42392 670800 42398 670812
rect 60642 670800 60648 670812
rect 42392 670772 60648 670800
rect 42392 670760 42398 670772
rect 60642 670760 60648 670772
rect 60700 670760 60706 670812
rect 655698 670760 655704 670812
rect 655756 670800 655762 670812
rect 676030 670800 676036 670812
rect 655756 670772 676036 670800
rect 655756 670760 655762 670772
rect 676030 670760 676036 670772
rect 676088 670760 676094 670812
rect 42426 670692 42432 670744
rect 42484 670732 42490 670744
rect 43530 670732 43536 670744
rect 42484 670704 43536 670732
rect 42484 670692 42490 670704
rect 43530 670692 43536 670704
rect 43588 670692 43594 670744
rect 43714 670624 43720 670676
rect 43772 670664 43778 670676
rect 44266 670664 44272 670676
rect 43772 670636 44272 670664
rect 43772 670624 43778 670636
rect 44266 670624 44272 670636
rect 44324 670624 44330 670676
rect 41782 670556 41788 670608
rect 41840 670556 41846 670608
rect 41800 670404 41828 670556
rect 41782 670352 41788 670404
rect 41840 670352 41846 670404
rect 673270 669332 673276 669384
rect 673328 669372 673334 669384
rect 676030 669372 676036 669384
rect 673328 669344 676036 669372
rect 673328 669332 673334 669344
rect 676030 669332 676036 669344
rect 676088 669332 676094 669384
rect 669590 669304 669596 669316
rect 669588 669276 669596 669304
rect 669590 669264 669596 669276
rect 669648 669304 669654 669316
rect 670510 669304 670516 669316
rect 669648 669276 670516 669304
rect 669648 669264 669654 669276
rect 670510 669264 670516 669276
rect 670568 669264 670574 669316
rect 669590 668176 669596 668228
rect 669648 668216 669654 668228
rect 676122 668216 676128 668228
rect 669648 668188 676128 668216
rect 669648 668176 669654 668188
rect 676122 668176 676128 668188
rect 676180 668176 676186 668228
rect 670418 668108 670424 668160
rect 670476 668148 670482 668160
rect 676214 668148 676220 668160
rect 670476 668120 676220 668148
rect 670476 668108 670482 668120
rect 676214 668108 676220 668120
rect 676272 668108 676278 668160
rect 655514 668040 655520 668092
rect 655572 668080 655578 668092
rect 678974 668080 678980 668092
rect 655572 668052 678980 668080
rect 655572 668040 655578 668052
rect 678974 668040 678980 668052
rect 679032 668040 679038 668092
rect 670602 667972 670608 668024
rect 670660 668012 670666 668024
rect 676306 668012 676312 668024
rect 670660 667984 676312 668012
rect 670660 667972 670666 667984
rect 676306 667972 676312 667984
rect 676364 667972 676370 668024
rect 42242 667836 42248 667888
rect 42300 667876 42306 667888
rect 43162 667876 43168 667888
rect 42300 667848 43168 667876
rect 42300 667836 42306 667848
rect 43162 667836 43168 667848
rect 43220 667836 43226 667888
rect 675202 667836 675208 667888
rect 675260 667876 675266 667888
rect 676030 667876 676036 667888
rect 675260 667848 676036 667876
rect 675260 667836 675266 667848
rect 676030 667836 676036 667848
rect 676088 667836 676094 667888
rect 42150 667700 42156 667752
rect 42208 667740 42214 667752
rect 42334 667740 42340 667752
rect 42208 667712 42340 667740
rect 42208 667700 42214 667712
rect 42334 667700 42340 667712
rect 42392 667700 42398 667752
rect 43162 667700 43168 667752
rect 43220 667740 43226 667752
rect 44174 667740 44180 667752
rect 43220 667712 44180 667740
rect 43220 667700 43226 667712
rect 44174 667700 44180 667712
rect 44232 667700 44238 667752
rect 42150 666680 42156 666732
rect 42208 666720 42214 666732
rect 43622 666720 43628 666732
rect 42208 666692 43628 666720
rect 42208 666680 42214 666692
rect 43622 666680 43628 666692
rect 43680 666680 43686 666732
rect 674558 665932 674564 665984
rect 674616 665972 674622 665984
rect 676030 665972 676036 665984
rect 674616 665944 676036 665972
rect 674616 665932 674622 665944
rect 676030 665932 676036 665944
rect 676088 665932 676094 665984
rect 670234 665252 670240 665304
rect 670292 665292 670298 665304
rect 676214 665292 676220 665304
rect 670292 665264 676220 665292
rect 670292 665252 670298 665264
rect 676214 665252 676220 665264
rect 676272 665252 676278 665304
rect 42150 665184 42156 665236
rect 42208 665224 42214 665236
rect 43254 665224 43260 665236
rect 42208 665196 43260 665224
rect 42208 665184 42214 665196
rect 43254 665184 43260 665196
rect 43312 665184 43318 665236
rect 670326 665224 670332 665236
rect 670322 665196 670332 665224
rect 670326 665184 670332 665196
rect 670384 665224 670390 665236
rect 678974 665224 678980 665236
rect 670384 665196 678980 665224
rect 670384 665184 670390 665196
rect 678974 665184 678980 665196
rect 679032 665184 679038 665236
rect 675018 665116 675024 665168
rect 675076 665156 675082 665168
rect 676030 665156 676036 665168
rect 675076 665128 676036 665156
rect 675076 665116 675082 665128
rect 676030 665116 676036 665128
rect 676088 665116 676094 665168
rect 674742 665048 674748 665100
rect 674800 665088 674806 665100
rect 676122 665088 676128 665100
rect 674800 665060 676128 665088
rect 674800 665048 674806 665060
rect 676122 665048 676128 665060
rect 676180 665048 676186 665100
rect 42150 664640 42156 664692
rect 42208 664680 42214 664692
rect 43530 664680 43536 664692
rect 42208 664652 43536 664680
rect 42208 664640 42214 664652
rect 43530 664640 43536 664652
rect 43588 664640 43594 664692
rect 43622 664504 43628 664556
rect 43680 664544 43686 664556
rect 44266 664544 44272 664556
rect 43680 664516 44272 664544
rect 43680 664504 43686 664516
rect 44266 664504 44272 664516
rect 44324 664504 44330 664556
rect 674650 664300 674656 664352
rect 674708 664340 674714 664352
rect 676030 664340 676036 664352
rect 674708 664312 676036 664340
rect 674708 664300 674714 664312
rect 676030 664300 676036 664312
rect 676088 664300 676094 664352
rect 42150 664164 42156 664216
rect 42208 664204 42214 664216
rect 43162 664204 43168 664216
rect 42208 664176 43168 664204
rect 42208 664164 42214 664176
rect 43162 664164 43168 664176
rect 43220 664164 43226 664216
rect 42150 663348 42156 663400
rect 42208 663388 42214 663400
rect 43070 663388 43076 663400
rect 42208 663360 43076 663388
rect 42208 663348 42214 663360
rect 43070 663348 43076 663360
rect 43128 663348 43134 663400
rect 673822 663076 673828 663128
rect 673880 663116 673886 663128
rect 676030 663116 676036 663128
rect 673880 663088 676036 663116
rect 673880 663076 673886 663088
rect 676030 663076 676036 663088
rect 676088 663076 676094 663128
rect 42150 661036 42156 661088
rect 42208 661076 42214 661088
rect 43346 661076 43352 661088
rect 42208 661048 43352 661076
rect 42208 661036 42214 661048
rect 43346 661036 43352 661048
rect 43404 661036 43410 661088
rect 42150 660492 42156 660544
rect 42208 660532 42214 660544
rect 43254 660532 43260 660544
rect 42208 660504 43260 660532
rect 42208 660492 42214 660504
rect 43254 660492 43260 660504
rect 43312 660492 43318 660544
rect 42426 659676 42432 659728
rect 42484 659716 42490 659728
rect 58434 659716 58440 659728
rect 42484 659688 58440 659716
rect 42484 659676 42490 659688
rect 58434 659676 58440 659688
rect 58492 659676 58498 659728
rect 672166 659676 672172 659728
rect 672224 659716 672230 659728
rect 678974 659716 678980 659728
rect 672224 659688 678980 659716
rect 672224 659676 672230 659688
rect 678974 659676 678980 659688
rect 679032 659676 679038 659728
rect 42242 659608 42248 659660
rect 42300 659648 42306 659660
rect 58526 659648 58532 659660
rect 42300 659620 58532 659648
rect 42300 659608 42306 659620
rect 58526 659608 58532 659620
rect 58584 659608 58590 659660
rect 45738 659540 45744 659592
rect 45796 659580 45802 659592
rect 58618 659580 58624 659592
rect 45796 659552 58624 659580
rect 45796 659540 45802 659552
rect 58618 659540 58624 659552
rect 58676 659540 58682 659592
rect 42242 659472 42248 659524
rect 42300 659512 42306 659524
rect 43622 659512 43628 659524
rect 42300 659484 43628 659512
rect 42300 659472 42306 659484
rect 43622 659472 43628 659484
rect 43680 659472 43686 659524
rect 42150 659200 42156 659252
rect 42208 659240 42214 659252
rect 44082 659240 44088 659252
rect 42208 659212 44088 659240
rect 42208 659200 42214 659212
rect 44082 659200 44088 659212
rect 44140 659200 44146 659252
rect 42150 657364 42156 657416
rect 42208 657404 42214 657416
rect 43530 657404 43536 657416
rect 42208 657376 43536 657404
rect 42208 657364 42214 657376
rect 43530 657364 43536 657376
rect 43588 657364 43594 657416
rect 655698 656888 655704 656940
rect 655756 656928 655762 656940
rect 675386 656928 675392 656940
rect 655756 656900 675392 656928
rect 655756 656888 655762 656900
rect 675386 656888 675392 656900
rect 675444 656888 675450 656940
rect 50982 656820 50988 656872
rect 51040 656860 51046 656872
rect 58434 656860 58440 656872
rect 51040 656832 58440 656860
rect 51040 656820 51046 656832
rect 58434 656820 58440 656832
rect 58492 656820 58498 656872
rect 53834 656752 53840 656804
rect 53892 656792 53898 656804
rect 58986 656792 58992 656804
rect 53892 656764 58992 656792
rect 53892 656752 53898 656764
rect 58986 656752 58992 656764
rect 59044 656752 59050 656804
rect 42150 656004 42156 656056
rect 42208 656044 42214 656056
rect 43898 656044 43904 656056
rect 42208 656016 43904 656044
rect 42208 656004 42214 656016
rect 43898 656004 43904 656016
rect 43956 656004 43962 656056
rect 673730 649544 673736 649596
rect 673788 649584 673794 649596
rect 675386 649584 675392 649596
rect 673788 649556 675392 649584
rect 673788 649544 673794 649556
rect 675386 649544 675392 649556
rect 675444 649544 675450 649596
rect 674650 648932 674656 648984
rect 674708 648972 674714 648984
rect 675110 648972 675116 648984
rect 674708 648944 675116 648972
rect 674708 648932 674714 648944
rect 675110 648932 675116 648944
rect 675168 648932 675174 648984
rect 674558 648864 674564 648916
rect 674616 648904 674622 648916
rect 675294 648904 675300 648916
rect 674616 648876 675300 648904
rect 674616 648864 674622 648876
rect 675294 648864 675300 648876
rect 675352 648864 675358 648916
rect 654410 648592 654416 648644
rect 654468 648632 654474 648644
rect 675110 648632 675116 648644
rect 654468 648604 675116 648632
rect 654468 648592 654474 648604
rect 675110 648592 675116 648604
rect 675168 648592 675174 648644
rect 673454 647708 673460 647760
rect 673512 647748 673518 647760
rect 675386 647748 675392 647760
rect 673512 647720 675392 647748
rect 673512 647708 673518 647720
rect 675386 647708 675392 647720
rect 675444 647708 675450 647760
rect 656434 645872 656440 645924
rect 656492 645912 656498 645924
rect 675202 645912 675208 645924
rect 656492 645884 675208 645912
rect 656492 645872 656498 645884
rect 675202 645872 675208 645884
rect 675260 645872 675266 645924
rect 674742 645192 674748 645244
rect 674800 645232 674806 645244
rect 675386 645232 675392 645244
rect 674800 645204 675392 645232
rect 674800 645192 674806 645204
rect 675386 645192 675392 645204
rect 675444 645192 675450 645244
rect 41506 645056 41512 645108
rect 41564 645096 41570 645108
rect 53834 645096 53840 645108
rect 41564 645068 53840 645096
rect 41564 645056 41570 645068
rect 53834 645056 53840 645068
rect 53892 645056 53898 645108
rect 41782 644988 41788 645040
rect 41840 645028 41846 645040
rect 56502 645028 56508 645040
rect 41840 645000 56508 645028
rect 41840 644988 41846 645000
rect 56502 644988 56508 645000
rect 56560 644988 56566 645040
rect 673822 644580 673828 644632
rect 673880 644620 673886 644632
rect 675386 644620 675392 644632
rect 673880 644592 675392 644620
rect 673880 644580 673886 644592
rect 675386 644580 675392 644592
rect 675444 644580 675450 644632
rect 673270 644240 673276 644292
rect 673328 644280 673334 644292
rect 673730 644280 673736 644292
rect 673328 644252 673736 644280
rect 673328 644240 673334 644252
rect 673730 644240 673736 644252
rect 673788 644240 673794 644292
rect 673730 644104 673736 644156
rect 673788 644144 673794 644156
rect 675386 644144 675392 644156
rect 673788 644116 675392 644144
rect 673788 644104 673794 644116
rect 675386 644104 675392 644116
rect 675444 644104 675450 644156
rect 41782 644036 41788 644088
rect 41840 644076 41846 644088
rect 50982 644076 50988 644088
rect 41840 644048 50988 644076
rect 41840 644036 41846 644048
rect 50982 644036 50988 644048
rect 51040 644036 51046 644088
rect 675478 643560 675484 643612
rect 675536 643560 675542 643612
rect 675110 643492 675116 643544
rect 675168 643532 675174 643544
rect 675386 643532 675392 643544
rect 675168 643504 675392 643532
rect 675168 643492 675174 643504
rect 675386 643492 675392 643504
rect 675444 643492 675450 643544
rect 675496 643464 675524 643560
rect 675220 643436 675524 643464
rect 675220 643408 675248 643436
rect 675202 643356 675208 643408
rect 675260 643356 675266 643408
rect 674650 642200 674656 642252
rect 674708 642240 674714 642252
rect 675110 642240 675116 642252
rect 674708 642212 675116 642240
rect 674708 642200 674714 642212
rect 675110 642200 675116 642212
rect 675168 642200 675174 642252
rect 674650 642064 674656 642116
rect 674708 642104 674714 642116
rect 675386 642104 675392 642116
rect 674708 642076 675392 642104
rect 674708 642064 674714 642076
rect 675386 642064 675392 642076
rect 675444 642064 675450 642116
rect 675110 640772 675116 640824
rect 675168 640772 675174 640824
rect 675128 640744 675156 640772
rect 675294 640744 675300 640756
rect 675128 640716 675300 640744
rect 675294 640704 675300 640716
rect 675352 640704 675358 640756
rect 675018 640228 675024 640280
rect 675076 640268 675082 640280
rect 675386 640268 675392 640280
rect 675076 640240 675392 640268
rect 675076 640228 675082 640240
rect 675386 640228 675392 640240
rect 675444 640228 675450 640280
rect 675202 638664 675208 638716
rect 675260 638664 675266 638716
rect 675220 638512 675248 638664
rect 675202 638460 675208 638512
rect 675260 638460 675266 638512
rect 675110 638392 675116 638444
rect 675168 638432 675174 638444
rect 675478 638432 675484 638444
rect 675168 638404 675484 638432
rect 675168 638392 675174 638404
rect 675478 638392 675484 638404
rect 675536 638392 675542 638444
rect 674558 638188 674564 638240
rect 674616 638228 674622 638240
rect 675754 638228 675760 638240
rect 674616 638200 675760 638228
rect 674616 638188 674622 638200
rect 675754 638188 675760 638200
rect 675812 638188 675818 638240
rect 673730 638052 673736 638104
rect 673788 638092 673794 638104
rect 674558 638092 674564 638104
rect 673788 638064 674564 638092
rect 673788 638052 673794 638064
rect 674558 638052 674564 638064
rect 674616 638052 674622 638104
rect 673270 637916 673276 637968
rect 673328 637956 673334 637968
rect 673730 637956 673736 637968
rect 673328 637928 673736 637956
rect 673328 637916 673334 637928
rect 673730 637916 673736 637928
rect 673788 637916 673794 637968
rect 674742 637780 674748 637832
rect 674800 637820 674806 637832
rect 675202 637820 675208 637832
rect 674800 637792 675208 637820
rect 674800 637780 674806 637792
rect 675202 637780 675208 637792
rect 675260 637780 675266 637832
rect 675662 637508 675668 637560
rect 675720 637548 675726 637560
rect 679066 637548 679072 637560
rect 675720 637520 679072 637548
rect 675720 637508 675726 637520
rect 679066 637508 679072 637520
rect 679124 637508 679130 637560
rect 673822 637236 673828 637288
rect 673880 637276 673886 637288
rect 674650 637276 674656 637288
rect 673880 637248 674656 637276
rect 673880 637236 673886 637248
rect 674650 637236 674656 637248
rect 674708 637236 674714 637288
rect 673454 637100 673460 637152
rect 673512 637140 673518 637152
rect 673822 637140 673828 637152
rect 673512 637112 673828 637140
rect 673512 637100 673518 637112
rect 673822 637100 673828 637112
rect 673880 637100 673886 637152
rect 41506 633224 41512 633276
rect 41564 633264 41570 633276
rect 48406 633264 48412 633276
rect 41564 633236 48412 633264
rect 41564 633224 41570 633236
rect 48406 633224 48412 633236
rect 48464 633224 48470 633276
rect 20622 632612 20628 632664
rect 20680 632652 20686 632664
rect 30190 632652 30196 632664
rect 20680 632624 30196 632652
rect 20680 632612 20686 632624
rect 30190 632612 30196 632624
rect 30248 632612 30254 632664
rect 42426 630912 42432 630964
rect 42484 630952 42490 630964
rect 43714 630952 43720 630964
rect 42484 630924 43720 630952
rect 42484 630912 42490 630924
rect 43714 630912 43720 630924
rect 43772 630912 43778 630964
rect 43162 630844 43168 630896
rect 43220 630884 43226 630896
rect 43806 630884 43812 630896
rect 43220 630856 43812 630884
rect 43220 630844 43226 630856
rect 43806 630844 43812 630856
rect 43864 630844 43870 630896
rect 20622 630776 20628 630828
rect 20680 630816 20686 630828
rect 43714 630816 43720 630828
rect 20680 630788 43720 630816
rect 20680 630776 20686 630788
rect 43714 630776 43720 630788
rect 43772 630776 43778 630828
rect 24762 630708 24768 630760
rect 24820 630748 24826 630760
rect 43162 630748 43168 630760
rect 24820 630720 43168 630748
rect 24820 630708 24826 630720
rect 43162 630708 43168 630720
rect 43220 630708 43226 630760
rect 43070 629348 43076 629400
rect 43128 629388 43134 629400
rect 43990 629388 43996 629400
rect 43128 629360 43996 629388
rect 43128 629348 43134 629360
rect 43990 629348 43996 629360
rect 44048 629348 44054 629400
rect 38470 629212 38476 629264
rect 38528 629252 38534 629264
rect 43070 629252 43076 629264
rect 38528 629224 43076 629252
rect 38528 629212 38534 629224
rect 43070 629212 43076 629224
rect 43128 629212 43134 629264
rect 43346 626832 43352 626884
rect 43404 626872 43410 626884
rect 43622 626872 43628 626884
rect 43404 626844 43628 626872
rect 43404 626832 43410 626844
rect 43622 626832 43628 626844
rect 43680 626832 43686 626884
rect 42702 626696 42708 626748
rect 42760 626736 42766 626748
rect 43346 626736 43352 626748
rect 42760 626708 43352 626736
rect 42760 626696 42766 626708
rect 43346 626696 43352 626708
rect 43404 626696 43410 626748
rect 42702 626560 42708 626612
rect 42760 626600 42766 626612
rect 58526 626600 58532 626612
rect 42760 626572 58532 626600
rect 42760 626560 42766 626572
rect 58526 626560 58532 626572
rect 58584 626560 58590 626612
rect 42150 625268 42156 625320
rect 42208 625308 42214 625320
rect 42334 625308 42340 625320
rect 42208 625280 42340 625308
rect 42208 625268 42214 625280
rect 42334 625268 42340 625280
rect 42392 625268 42398 625320
rect 42334 624452 42340 624504
rect 42392 624492 42398 624504
rect 42702 624492 42708 624504
rect 42392 624464 42708 624492
rect 42392 624452 42398 624464
rect 42702 624452 42708 624464
rect 42760 624452 42766 624504
rect 655790 624112 655796 624164
rect 655848 624152 655854 624164
rect 678974 624152 678980 624164
rect 655848 624124 678980 624152
rect 655848 624112 655854 624124
rect 678974 624112 678980 624124
rect 679032 624112 679038 624164
rect 670602 624084 670608 624096
rect 670600 624056 670608 624084
rect 670602 624044 670608 624056
rect 670660 624084 670666 624096
rect 676214 624084 676220 624096
rect 670660 624056 676220 624084
rect 670660 624044 670666 624056
rect 676214 624044 676220 624056
rect 676272 624044 676278 624096
rect 655606 623976 655612 624028
rect 655664 624016 655670 624028
rect 676306 624016 676312 624028
rect 655664 623988 676312 624016
rect 655664 623976 655670 623988
rect 676306 623976 676312 623988
rect 676364 623976 676370 624028
rect 670510 623908 670516 623960
rect 670568 623948 670574 623960
rect 676122 623948 676128 623960
rect 670568 623920 676128 623948
rect 670568 623908 670574 623920
rect 676122 623908 676128 623920
rect 676180 623908 676186 623960
rect 655422 623840 655428 623892
rect 655480 623880 655486 623892
rect 676030 623880 676036 623892
rect 655480 623852 676036 623880
rect 655480 623840 655486 623852
rect 676030 623840 676036 623852
rect 676088 623840 676094 623892
rect 673270 623772 673276 623824
rect 673328 623812 673334 623824
rect 675938 623812 675944 623824
rect 673328 623784 675944 623812
rect 673328 623772 673334 623784
rect 675938 623772 675944 623784
rect 675996 623772 676002 623824
rect 674926 623704 674932 623756
rect 674984 623744 674990 623756
rect 676030 623744 676036 623756
rect 674984 623716 676036 623744
rect 674984 623704 674990 623716
rect 676030 623704 676036 623716
rect 676088 623704 676094 623756
rect 42150 623432 42156 623484
rect 42208 623472 42214 623484
rect 43254 623472 43260 623484
rect 42208 623444 43260 623472
rect 42208 623432 42214 623444
rect 43254 623432 43260 623444
rect 43312 623432 43318 623484
rect 42242 622412 42248 622464
rect 42300 622452 42306 622464
rect 42702 622452 42708 622464
rect 42300 622424 42708 622452
rect 42300 622412 42306 622424
rect 42702 622412 42708 622424
rect 42760 622412 42766 622464
rect 42334 622208 42340 622260
rect 42392 622248 42398 622260
rect 43070 622248 43076 622260
rect 42392 622220 43076 622248
rect 42392 622208 42398 622220
rect 43070 622208 43076 622220
rect 43128 622208 43134 622260
rect 42334 621664 42340 621716
rect 42392 621704 42398 621716
rect 43438 621704 43444 621716
rect 42392 621676 43444 621704
rect 42392 621664 42398 621676
rect 43438 621664 43444 621676
rect 43496 621664 43502 621716
rect 670602 621120 670608 621172
rect 670660 621160 670666 621172
rect 676122 621160 676128 621172
rect 670660 621132 676128 621160
rect 670660 621120 670666 621132
rect 676122 621120 676128 621132
rect 676180 621120 676186 621172
rect 670418 621052 670424 621104
rect 670476 621092 670482 621104
rect 676214 621092 676220 621104
rect 670476 621064 676220 621092
rect 670476 621052 670482 621064
rect 676214 621052 676220 621064
rect 676272 621052 676278 621104
rect 670234 621024 670240 621036
rect 670224 620996 670240 621024
rect 670234 620984 670240 620996
rect 670292 621024 670298 621036
rect 676306 621024 676312 621036
rect 670292 620996 676312 621024
rect 670292 620984 670298 620996
rect 676306 620984 676312 620996
rect 676364 620984 676370 621036
rect 674282 620916 674288 620968
rect 674340 620956 674346 620968
rect 676030 620956 676036 620968
rect 674340 620928 676036 620956
rect 674340 620916 674346 620928
rect 676030 620916 676036 620928
rect 676088 620916 676094 620968
rect 42058 620780 42064 620832
rect 42116 620820 42122 620832
rect 43622 620820 43628 620832
rect 42116 620792 43628 620820
rect 42116 620780 42122 620792
rect 43622 620780 43628 620792
rect 43680 620780 43686 620832
rect 42058 620168 42064 620220
rect 42116 620208 42122 620220
rect 43070 620208 43076 620220
rect 42116 620180 43076 620208
rect 42116 620168 42122 620180
rect 43070 620168 43076 620180
rect 43128 620168 43134 620220
rect 673546 620100 673552 620152
rect 673604 620140 673610 620152
rect 676030 620140 676036 620152
rect 673604 620112 676036 620140
rect 673604 620100 673610 620112
rect 676030 620100 676036 620112
rect 676088 620100 676094 620152
rect 42426 619148 42432 619200
rect 42484 619188 42490 619200
rect 43162 619188 43168 619200
rect 42484 619160 43168 619188
rect 42484 619148 42490 619160
rect 43162 619148 43168 619160
rect 43220 619148 43226 619200
rect 42702 618196 42708 618248
rect 42760 618236 42766 618248
rect 58158 618236 58164 618248
rect 42760 618208 58164 618236
rect 42760 618196 42766 618208
rect 58158 618196 58164 618208
rect 58216 618196 58222 618248
rect 674466 618196 674472 618248
rect 674524 618236 674530 618248
rect 676030 618236 676036 618248
rect 674524 618208 676036 618236
rect 674524 618196 674530 618208
rect 676030 618196 676036 618208
rect 676088 618196 676094 618248
rect 673638 618060 673644 618112
rect 673696 618100 673702 618112
rect 676030 618100 676036 618112
rect 673696 618072 676036 618100
rect 673696 618060 673702 618072
rect 676030 618060 676036 618072
rect 676088 618060 676094 618112
rect 42058 617312 42064 617364
rect 42116 617352 42122 617364
rect 43346 617352 43352 617364
rect 42116 617324 43352 617352
rect 42116 617312 42122 617324
rect 43346 617312 43352 617324
rect 43404 617312 43410 617364
rect 673362 616700 673368 616752
rect 673420 616740 673426 616752
rect 676214 616740 676220 616752
rect 673420 616712 676220 616740
rect 673420 616700 673426 616712
rect 676214 616700 676220 616712
rect 676272 616700 676278 616752
rect 42334 616020 42340 616072
rect 42392 616060 42398 616072
rect 44082 616060 44088 616072
rect 42392 616032 44088 616060
rect 42392 616020 42398 616032
rect 44082 616020 44088 616032
rect 44140 616020 44146 616072
rect 42242 615952 42248 616004
rect 42300 615992 42306 616004
rect 43714 615992 43720 616004
rect 42300 615964 43720 615992
rect 42300 615952 42306 615964
rect 43714 615952 43720 615964
rect 43772 615952 43778 616004
rect 42150 615816 42156 615868
rect 42208 615856 42214 615868
rect 43806 615856 43812 615868
rect 42208 615828 43812 615856
rect 42208 615816 42214 615828
rect 43806 615816 43812 615828
rect 43864 615816 43870 615868
rect 42426 615476 42432 615528
rect 42484 615516 42490 615528
rect 58526 615516 58532 615528
rect 42484 615488 58532 615516
rect 42484 615476 42490 615488
rect 58526 615476 58532 615488
rect 58584 615476 58590 615528
rect 50982 615408 50988 615460
rect 51040 615448 51046 615460
rect 58158 615448 58164 615460
rect 51040 615420 58164 615448
rect 51040 615408 51046 615420
rect 58158 615408 58164 615420
rect 58216 615408 58222 615460
rect 672258 614592 672264 614644
rect 672316 614632 672322 614644
rect 679066 614632 679072 614644
rect 672316 614604 679072 614632
rect 672316 614592 672322 614604
rect 679066 614592 679072 614604
rect 679124 614592 679130 614644
rect 42150 614184 42156 614236
rect 42208 614224 42214 614236
rect 43990 614224 43996 614236
rect 42208 614196 43996 614224
rect 42208 614184 42214 614196
rect 43990 614184 43996 614196
rect 44048 614184 44054 614236
rect 655422 612824 655428 612876
rect 655480 612864 655486 612876
rect 675662 612864 675668 612876
rect 655480 612836 675668 612864
rect 655480 612824 655486 612836
rect 675662 612824 675668 612836
rect 675720 612824 675726 612876
rect 56502 612688 56508 612740
rect 56560 612728 56566 612740
rect 57974 612728 57980 612740
rect 56560 612700 57980 612728
rect 56560 612688 56566 612700
rect 57974 612688 57980 612700
rect 58032 612688 58038 612740
rect 53834 612076 53840 612128
rect 53892 612116 53898 612128
rect 57974 612116 57980 612128
rect 53892 612088 57980 612116
rect 53892 612076 53898 612088
rect 57974 612076 57980 612088
rect 58032 612076 58038 612128
rect 674282 608948 674288 609000
rect 674340 608988 674346 609000
rect 675570 608988 675576 609000
rect 674340 608960 675576 608988
rect 674340 608948 674346 608960
rect 675570 608948 675576 608960
rect 675628 608948 675634 609000
rect 674466 605072 674472 605124
rect 674524 605112 674530 605124
rect 675202 605112 675208 605124
rect 674524 605084 675208 605112
rect 674524 605072 674530 605084
rect 675202 605072 675208 605084
rect 675260 605072 675266 605124
rect 673638 603440 673644 603492
rect 673696 603480 673702 603492
rect 675478 603480 675484 603492
rect 673696 603452 675484 603480
rect 673696 603440 673702 603452
rect 675478 603440 675484 603452
rect 675536 603440 675542 603492
rect 656802 601740 656808 601792
rect 656860 601780 656866 601792
rect 675202 601780 675208 601792
rect 656860 601752 675208 601780
rect 656860 601740 656866 601752
rect 675202 601740 675208 601752
rect 675260 601740 675266 601792
rect 41782 601672 41788 601724
rect 41840 601712 41846 601724
rect 56502 601712 56508 601724
rect 41840 601684 56508 601712
rect 41840 601672 41846 601684
rect 56502 601672 56508 601684
rect 56560 601672 56566 601724
rect 655606 601672 655612 601724
rect 655664 601712 655670 601724
rect 675294 601712 675300 601724
rect 655664 601684 675300 601712
rect 655664 601672 655670 601684
rect 675294 601672 675300 601684
rect 675352 601672 675358 601724
rect 673546 600380 673552 600432
rect 673604 600420 673610 600432
rect 674466 600420 674472 600432
rect 673604 600392 674472 600420
rect 673604 600380 673610 600392
rect 674466 600380 674472 600392
rect 674524 600380 674530 600432
rect 674466 600244 674472 600296
rect 674524 600284 674530 600296
rect 675478 600284 675484 600296
rect 674524 600256 675484 600284
rect 674524 600244 674530 600256
rect 675478 600244 675484 600256
rect 675536 600244 675542 600296
rect 674282 599904 674288 599956
rect 674340 599944 674346 599956
rect 674650 599944 674656 599956
rect 674340 599916 674656 599944
rect 674340 599904 674346 599916
rect 674650 599904 674656 599916
rect 674708 599904 674714 599956
rect 674282 599768 674288 599820
rect 674340 599808 674346 599820
rect 675478 599808 675484 599820
rect 674340 599780 675484 599808
rect 674340 599768 674346 599780
rect 675478 599768 675484 599780
rect 675536 599768 675542 599820
rect 674926 598952 674932 599004
rect 674984 598992 674990 599004
rect 675386 598992 675392 599004
rect 674984 598964 675392 598992
rect 674984 598952 674990 598964
rect 675386 598952 675392 598964
rect 675444 598952 675450 599004
rect 675202 598884 675208 598936
rect 675260 598924 675266 598936
rect 675260 598896 675432 598924
rect 675260 598884 675266 598896
rect 675294 598816 675300 598868
rect 675352 598816 675358 598868
rect 675312 598664 675340 598816
rect 675404 598732 675432 598896
rect 675386 598680 675392 598732
rect 675444 598680 675450 598732
rect 675294 598612 675300 598664
rect 675352 598612 675358 598664
rect 673454 598544 673460 598596
rect 673512 598584 673518 598596
rect 675478 598584 675484 598596
rect 673512 598556 675484 598584
rect 673512 598544 673518 598556
rect 675478 598544 675484 598556
rect 675536 598544 675542 598596
rect 673546 597252 673552 597304
rect 673604 597292 673610 597304
rect 675202 597292 675208 597304
rect 673604 597264 675208 597292
rect 673604 597252 673610 597264
rect 675202 597252 675208 597264
rect 675260 597252 675266 597304
rect 673546 597116 673552 597168
rect 673604 597156 673610 597168
rect 675386 597156 675392 597168
rect 673604 597128 675392 597156
rect 673604 597116 673610 597128
rect 675386 597116 675392 597128
rect 675444 597116 675450 597168
rect 674650 595416 674656 595468
rect 674708 595456 674714 595468
rect 675202 595456 675208 595468
rect 674708 595428 675208 595456
rect 674708 595416 674714 595428
rect 675202 595416 675208 595428
rect 675260 595416 675266 595468
rect 674650 595280 674656 595332
rect 674708 595320 674714 595332
rect 675386 595320 675392 595332
rect 674708 595292 675392 595320
rect 674708 595280 674714 595292
rect 675386 595280 675392 595292
rect 675444 595280 675450 595332
rect 675294 593512 675300 593564
rect 675352 593552 675358 593564
rect 675352 593524 675708 593552
rect 675352 593512 675358 593524
rect 675202 593172 675208 593224
rect 675260 593212 675266 593224
rect 675570 593212 675576 593224
rect 675260 593184 675576 593212
rect 675260 593172 675266 593184
rect 675570 593172 675576 593184
rect 675628 593172 675634 593224
rect 43070 592968 43076 593020
rect 43128 593008 43134 593020
rect 43346 593008 43352 593020
rect 43128 592980 43352 593008
rect 43128 592968 43134 592980
rect 43346 592968 43352 592980
rect 43404 592968 43410 593020
rect 43346 592832 43352 592884
rect 43404 592872 43410 592884
rect 44082 592872 44088 592884
rect 43404 592844 44088 592872
rect 43404 592832 43410 592844
rect 44082 592832 44088 592844
rect 44140 592832 44146 592884
rect 675680 592860 675708 593524
rect 675680 592832 679020 592860
rect 678992 592804 679020 592832
rect 678974 592752 678980 592804
rect 679032 592752 679038 592804
rect 674926 589364 674932 589416
rect 674984 589404 674990 589416
rect 675294 589404 675300 589416
rect 674984 589376 675300 589404
rect 674984 589364 674990 589376
rect 675294 589364 675300 589376
rect 675352 589364 675358 589416
rect 41506 589228 41512 589280
rect 41564 589268 41570 589280
rect 53834 589268 53840 589280
rect 41564 589240 53840 589268
rect 41564 589228 41570 589240
rect 53834 589228 53840 589240
rect 53892 589228 53898 589280
rect 674466 589228 674472 589280
rect 674524 589268 674530 589280
rect 674926 589268 674932 589280
rect 674524 589240 674932 589268
rect 674524 589228 674530 589240
rect 674926 589228 674932 589240
rect 674984 589228 674990 589280
rect 38562 587800 38568 587852
rect 38620 587840 38626 587852
rect 42334 587840 42340 587852
rect 38620 587812 42340 587840
rect 38620 587800 38626 587812
rect 42334 587800 42340 587812
rect 42392 587800 42398 587852
rect 43070 585148 43076 585200
rect 43128 585188 43134 585200
rect 58526 585188 58532 585200
rect 43128 585160 58532 585188
rect 43128 585148 43134 585160
rect 58526 585148 58532 585160
rect 58584 585148 58590 585200
rect 42426 584196 42432 584248
rect 42484 584236 42490 584248
rect 44266 584236 44272 584248
rect 42484 584208 44272 584236
rect 42484 584196 42490 584208
rect 44266 584196 44272 584208
rect 44324 584196 44330 584248
rect 43346 583856 43352 583908
rect 43404 583896 43410 583908
rect 43404 583868 43576 583896
rect 43404 583856 43410 583868
rect 43548 583704 43576 583868
rect 673454 583720 673460 583772
rect 673512 583760 673518 583772
rect 674466 583760 674472 583772
rect 673512 583732 674472 583760
rect 673512 583720 673518 583732
rect 674466 583720 674472 583732
rect 674524 583720 674530 583772
rect 674650 583720 674656 583772
rect 674708 583760 674714 583772
rect 675202 583760 675208 583772
rect 674708 583732 675208 583760
rect 674708 583720 674714 583732
rect 675202 583720 675208 583732
rect 675260 583720 675266 583772
rect 43530 583652 43536 583704
rect 43588 583652 43594 583704
rect 673546 583584 673552 583636
rect 673604 583624 673610 583636
rect 674650 583624 674656 583636
rect 673604 583596 674656 583624
rect 673604 583584 673610 583596
rect 674650 583584 674656 583596
rect 674708 583584 674714 583636
rect 42242 582564 42248 582616
rect 42300 582604 42306 582616
rect 59354 582604 59360 582616
rect 42300 582576 59360 582604
rect 42300 582564 42306 582576
rect 59354 582564 59360 582576
rect 59412 582564 59418 582616
rect 42150 582088 42156 582140
rect 42208 582128 42214 582140
rect 43254 582128 43260 582140
rect 42208 582100 43260 582128
rect 42208 582088 42214 582100
rect 43254 582088 43260 582100
rect 43312 582088 43318 582140
rect 43254 581952 43260 582004
rect 43312 581992 43318 582004
rect 43530 581992 43536 582004
rect 43312 581964 43536 581992
rect 43312 581952 43318 581964
rect 43530 581952 43536 581964
rect 43588 581952 43594 582004
rect 42150 581476 42156 581528
rect 42208 581516 42214 581528
rect 43070 581516 43076 581528
rect 42208 581488 43076 581516
rect 42208 581476 42214 581488
rect 43070 581476 43076 581488
rect 43128 581476 43134 581528
rect 43438 580388 43444 580440
rect 43496 580428 43502 580440
rect 43990 580428 43996 580440
rect 43496 580400 43996 580428
rect 43496 580388 43502 580400
rect 43990 580388 43996 580400
rect 44048 580388 44054 580440
rect 42242 580320 42248 580372
rect 42300 580320 42306 580372
rect 44082 580320 44088 580372
rect 44140 580320 44146 580372
rect 42260 580168 42288 580320
rect 44100 580168 44128 580320
rect 42242 580116 42248 580168
rect 42300 580116 42306 580168
rect 44082 580116 44088 580168
rect 44140 580116 44146 580168
rect 656158 580048 656164 580100
rect 656216 580088 656222 580100
rect 676214 580088 676220 580100
rect 656216 580060 676220 580088
rect 656216 580048 656222 580060
rect 676214 580048 676220 580060
rect 676272 580048 676278 580100
rect 655974 579912 655980 579964
rect 656032 579952 656038 579964
rect 676122 579952 676128 579964
rect 656032 579924 676128 579952
rect 656032 579912 656038 579924
rect 676122 579912 676128 579924
rect 676180 579912 676186 579964
rect 655514 579776 655520 579828
rect 655572 579816 655578 579828
rect 676306 579816 676312 579828
rect 655572 579788 676312 579816
rect 655572 579776 655578 579788
rect 676306 579776 676312 579788
rect 676364 579776 676370 579828
rect 670510 579680 670516 579692
rect 670504 579652 670516 579680
rect 670510 579640 670516 579652
rect 670568 579680 670574 579692
rect 676214 579680 676220 579692
rect 670568 579652 676220 579680
rect 670568 579640 670574 579652
rect 676214 579640 676220 579652
rect 676272 579640 676278 579692
rect 673270 579028 673276 579080
rect 673328 579068 673334 579080
rect 676030 579068 676036 579080
rect 673328 579040 676036 579068
rect 673328 579028 673334 579040
rect 676030 579028 676036 579040
rect 676088 579028 676094 579080
rect 42242 578960 42248 579012
rect 42300 579000 42306 579012
rect 43622 579000 43628 579012
rect 42300 578972 43628 579000
rect 42300 578960 42306 578972
rect 43622 578960 43628 578972
rect 43680 578960 43686 579012
rect 42150 578756 42156 578808
rect 42208 578796 42214 578808
rect 43162 578796 43168 578808
rect 42208 578768 43168 578796
rect 42208 578756 42214 578768
rect 43162 578756 43168 578768
rect 43220 578756 43226 578808
rect 42150 578416 42156 578468
rect 42208 578456 42214 578468
rect 43806 578456 43812 578468
rect 42208 578428 43812 578456
rect 42208 578416 42214 578428
rect 43806 578416 43812 578428
rect 43864 578416 43870 578468
rect 43898 578416 43904 578468
rect 43956 578416 43962 578468
rect 673362 578416 673368 578468
rect 673420 578456 673426 578468
rect 676214 578456 676220 578468
rect 673420 578428 676220 578456
rect 673420 578416 673426 578428
rect 676214 578416 676220 578428
rect 676272 578416 676278 578468
rect 43916 578264 43944 578416
rect 43898 578212 43904 578264
rect 43956 578212 43962 578264
rect 42242 577124 42248 577176
rect 42300 577164 42306 577176
rect 44082 577164 44088 577176
rect 42300 577136 44088 577164
rect 42300 577124 42306 577136
rect 44082 577124 44088 577136
rect 44140 577124 44146 577176
rect 42150 576920 42156 576972
rect 42208 576960 42214 576972
rect 43070 576960 43076 576972
rect 42208 576932 43076 576960
rect 42208 576920 42214 576932
rect 43070 576920 43076 576932
rect 43128 576920 43134 576972
rect 670418 576960 670424 576972
rect 670406 576932 670424 576960
rect 670418 576920 670424 576932
rect 670476 576960 670482 576972
rect 676214 576960 676220 576972
rect 670476 576932 676220 576960
rect 670476 576920 670482 576932
rect 676214 576920 676220 576932
rect 676272 576920 676278 576972
rect 670602 576892 670608 576904
rect 670588 576864 670608 576892
rect 670602 576852 670608 576864
rect 670660 576892 670666 576904
rect 676122 576892 676128 576904
rect 670660 576864 676128 576892
rect 670660 576852 670666 576864
rect 676122 576852 676128 576864
rect 676180 576852 676186 576904
rect 675018 576784 675024 576836
rect 675076 576824 675082 576836
rect 676030 576824 676036 576836
rect 675076 576796 676036 576824
rect 675076 576784 675082 576796
rect 676030 576784 676036 576796
rect 676088 576784 676094 576836
rect 673730 576716 673736 576768
rect 673788 576756 673794 576768
rect 675938 576756 675944 576768
rect 673788 576728 675944 576756
rect 673788 576716 673794 576728
rect 675938 576716 675944 576728
rect 675996 576716 676002 576768
rect 675110 576036 675116 576088
rect 675168 576076 675174 576088
rect 676030 576076 676036 576088
rect 675168 576048 676036 576076
rect 675168 576036 675174 576048
rect 676030 576036 676036 576048
rect 676088 576036 676094 576088
rect 42334 575968 42340 576020
rect 42392 576008 42398 576020
rect 43530 576008 43536 576020
rect 42392 575980 43536 576008
rect 42392 575968 42398 575980
rect 43530 575968 43536 575980
rect 43588 575968 43594 576020
rect 42426 574064 42432 574116
rect 42484 574104 42490 574116
rect 60642 574104 60648 574116
rect 42484 574076 60648 574104
rect 42484 574064 42490 574076
rect 60642 574064 60648 574076
rect 60700 574064 60706 574116
rect 42150 573792 42156 573844
rect 42208 573832 42214 573844
rect 43346 573832 43352 573844
rect 42208 573804 43352 573832
rect 42208 573792 42214 573804
rect 43346 573792 43352 573804
rect 43404 573792 43410 573844
rect 674742 573656 674748 573708
rect 674800 573696 674806 573708
rect 676030 573696 676036 573708
rect 674800 573668 676036 573696
rect 674800 573656 674806 573668
rect 676030 573656 676036 573668
rect 676088 573656 676094 573708
rect 42334 572840 42340 572892
rect 42392 572880 42398 572892
rect 43438 572880 43444 572892
rect 42392 572852 43444 572880
rect 42392 572840 42398 572852
rect 43438 572840 43444 572852
rect 43496 572840 43502 572892
rect 674558 572772 674564 572824
rect 674616 572812 674622 572824
rect 676030 572812 676036 572824
rect 674616 572784 676036 572812
rect 674616 572772 674622 572784
rect 676030 572772 676036 572784
rect 676088 572772 676094 572824
rect 673822 572364 673828 572416
rect 673880 572404 673886 572416
rect 676030 572404 676036 572416
rect 673880 572376 676036 572404
rect 673880 572364 673886 572376
rect 676030 572364 676036 572376
rect 676088 572364 676094 572416
rect 42242 571956 42248 572008
rect 42300 571996 42306 572008
rect 44082 571996 44088 572008
rect 42300 571968 44088 571996
rect 42300 571956 42306 571968
rect 44082 571956 44088 571968
rect 44140 571956 44146 572008
rect 42334 571616 42340 571668
rect 42392 571656 42398 571668
rect 43714 571656 43720 571668
rect 42392 571628 43720 571656
rect 42392 571616 42398 571628
rect 43714 571616 43720 571628
rect 43772 571616 43778 571668
rect 56502 571276 56508 571328
rect 56560 571316 56566 571328
rect 58710 571316 58716 571328
rect 56560 571288 58716 571316
rect 56560 571276 56566 571288
rect 58710 571276 58716 571288
rect 58768 571276 58774 571328
rect 42058 570936 42064 570988
rect 42116 570976 42122 570988
rect 43254 570976 43260 570988
rect 42116 570948 43260 570976
rect 42116 570936 42122 570948
rect 43254 570936 43260 570948
rect 43312 570936 43318 570988
rect 673454 568760 673460 568812
rect 673512 568800 673518 568812
rect 675386 568800 675392 568812
rect 673512 568772 675392 568800
rect 673512 568760 673518 568772
rect 675386 568760 675392 568772
rect 675444 568760 675450 568812
rect 655974 568624 655980 568676
rect 656032 568664 656038 568676
rect 675386 568664 675392 568676
rect 656032 568636 675392 568664
rect 656032 568624 656038 568636
rect 675386 568624 675392 568636
rect 675444 568624 675450 568676
rect 672350 568556 672356 568608
rect 672408 568596 672414 568608
rect 678974 568596 678980 568608
rect 672408 568568 678980 568596
rect 672408 568556 672414 568568
rect 678974 568556 678980 568568
rect 679032 568556 679038 568608
rect 673822 564408 673828 564460
rect 673880 564448 673886 564460
rect 675294 564448 675300 564460
rect 673880 564420 675300 564448
rect 673880 564408 673886 564420
rect 675294 564408 675300 564420
rect 675352 564408 675358 564460
rect 675018 559512 675024 559564
rect 675076 559552 675082 559564
rect 675478 559552 675484 559564
rect 675076 559524 675484 559552
rect 675076 559512 675082 559524
rect 675478 559512 675484 559524
rect 675536 559512 675542 559564
rect 41506 558764 41512 558816
rect 41564 558804 41570 558816
rect 56502 558804 56508 558816
rect 41564 558776 56508 558804
rect 41564 558764 41570 558776
rect 56502 558764 56508 558776
rect 56560 558764 56566 558816
rect 41506 558628 41512 558680
rect 41564 558668 41570 558680
rect 53926 558668 53932 558680
rect 41564 558640 53932 558668
rect 41564 558628 41570 558640
rect 53926 558628 53932 558640
rect 53984 558628 53990 558680
rect 674282 558220 674288 558272
rect 674340 558260 674346 558272
rect 675386 558260 675392 558272
rect 674340 558232 675392 558260
rect 674340 558220 674346 558232
rect 675386 558220 675392 558232
rect 675444 558220 675450 558272
rect 674558 558016 674564 558068
rect 674616 558056 674622 558068
rect 675294 558056 675300 558068
rect 674616 558028 675300 558056
rect 674616 558016 674622 558028
rect 675294 558016 675300 558028
rect 675352 558016 675358 558068
rect 41506 557540 41512 557592
rect 41564 557580 41570 557592
rect 50982 557580 50988 557592
rect 41564 557552 50988 557580
rect 41564 557540 41570 557552
rect 50982 557540 50988 557552
rect 51040 557540 51046 557592
rect 654226 557540 654232 557592
rect 654284 557580 654290 557592
rect 675110 557580 675116 557592
rect 654284 557552 675116 557580
rect 654284 557540 654290 557552
rect 675110 557540 675116 557552
rect 675168 557540 675174 557592
rect 674742 555228 674748 555280
rect 674800 555268 674806 555280
rect 675386 555268 675392 555280
rect 674800 555240 675392 555268
rect 674800 555228 674806 555240
rect 675386 555228 675392 555240
rect 675444 555228 675450 555280
rect 654134 554752 654140 554804
rect 654192 554792 654198 554804
rect 675294 554792 675300 554804
rect 654192 554764 675300 554792
rect 654192 554752 654198 554764
rect 675294 554752 675300 554764
rect 675352 554752 675358 554804
rect 673086 554684 673092 554736
rect 673144 554724 673150 554736
rect 673454 554724 673460 554736
rect 673144 554696 673460 554724
rect 673144 554684 673150 554696
rect 673454 554684 673460 554696
rect 673512 554684 673518 554736
rect 673454 554548 673460 554600
rect 673512 554588 673518 554600
rect 675386 554588 675392 554600
rect 673512 554560 675392 554588
rect 673512 554548 673518 554560
rect 675386 554548 675392 554560
rect 675444 554548 675450 554600
rect 673730 553800 673736 553852
rect 673788 553840 673794 553852
rect 675570 553840 675576 553852
rect 673788 553812 675576 553840
rect 673788 553800 673794 553812
rect 675570 553800 675576 553812
rect 675628 553800 675634 553852
rect 675478 553732 675484 553784
rect 675536 553732 675542 553784
rect 675110 553460 675116 553512
rect 675168 553500 675174 553512
rect 675386 553500 675392 553512
rect 675168 553472 675392 553500
rect 675168 553460 675174 553472
rect 675386 553460 675392 553472
rect 675444 553460 675450 553512
rect 675110 553324 675116 553376
rect 675168 553364 675174 553376
rect 675496 553364 675524 553732
rect 675168 553336 675524 553364
rect 675168 553324 675174 553336
rect 673178 552168 673184 552220
rect 673236 552208 673242 552220
rect 673822 552208 673828 552220
rect 673236 552180 673828 552208
rect 673236 552168 673242 552180
rect 673822 552168 673828 552180
rect 673880 552168 673886 552220
rect 673822 552032 673828 552084
rect 673880 552072 673886 552084
rect 674558 552072 674564 552084
rect 673880 552044 674564 552072
rect 673880 552032 673886 552044
rect 674558 552032 674564 552044
rect 674616 552032 674622 552084
rect 674558 551896 674564 551948
rect 674616 551936 674622 551948
rect 675386 551936 675392 551948
rect 674616 551908 675392 551936
rect 674616 551896 674622 551908
rect 675386 551896 675392 551908
rect 675444 551896 675450 551948
rect 673270 548972 673276 549024
rect 673328 549012 673334 549024
rect 673454 549012 673460 549024
rect 673328 548984 673460 549012
rect 673328 548972 673334 548984
rect 673454 548972 673460 548984
rect 673512 548972 673518 549024
rect 673454 548836 673460 548888
rect 673512 548876 673518 548888
rect 675294 548876 675300 548888
rect 673512 548848 675300 548876
rect 673512 548836 673518 548848
rect 675294 548836 675300 548848
rect 675352 548836 675358 548888
rect 41506 548632 41512 548684
rect 41564 548672 41570 548684
rect 43622 548672 43628 548684
rect 41564 548644 43628 548672
rect 41564 548632 41570 548644
rect 43622 548632 43628 548644
rect 43680 548632 43686 548684
rect 41506 548428 41512 548480
rect 41564 548468 41570 548480
rect 43254 548468 43260 548480
rect 41564 548440 43260 548468
rect 41564 548428 41570 548440
rect 43254 548428 43260 548440
rect 43312 548428 43318 548480
rect 673086 547952 673092 548004
rect 673144 547992 673150 548004
rect 675386 547992 675392 548004
rect 673144 547964 675392 547992
rect 673144 547952 673150 547964
rect 675386 547952 675392 547964
rect 675444 547952 675450 548004
rect 673178 547612 673184 547664
rect 673236 547652 673242 547664
rect 677594 547652 677600 547664
rect 673236 547624 677600 547652
rect 673236 547612 673242 547624
rect 677594 547612 677600 547624
rect 677652 547612 677658 547664
rect 41506 546864 41512 546916
rect 41564 546904 41570 546916
rect 45738 546904 45744 546916
rect 41564 546876 45744 546904
rect 41564 546864 41570 546876
rect 45738 546864 45744 546876
rect 45796 546864 45802 546916
rect 41598 546388 41604 546440
rect 41656 546428 41662 546440
rect 43714 546428 43720 546440
rect 41656 546400 43720 546428
rect 41656 546388 41662 546400
rect 43714 546388 43720 546400
rect 43772 546388 43778 546440
rect 41414 546320 41420 546372
rect 41472 546360 41478 546372
rect 43438 546360 43444 546372
rect 41472 546332 43444 546360
rect 41472 546320 41478 546332
rect 43438 546320 43444 546332
rect 43496 546320 43502 546372
rect 673822 545232 673828 545284
rect 673880 545272 673886 545284
rect 675570 545272 675576 545284
rect 673880 545244 675576 545272
rect 673880 545232 673886 545244
rect 675570 545232 675576 545244
rect 675628 545232 675634 545284
rect 673822 545096 673828 545148
rect 673880 545136 673886 545148
rect 674282 545136 674288 545148
rect 673880 545108 674288 545136
rect 673880 545096 673886 545108
rect 674282 545096 674288 545108
rect 674340 545096 674346 545148
rect 674742 545096 674748 545148
rect 674800 545136 674806 545148
rect 675018 545136 675024 545148
rect 674800 545108 675024 545136
rect 674800 545096 674806 545108
rect 675018 545096 675024 545108
rect 675076 545096 675082 545148
rect 674834 544756 674840 544808
rect 674892 544796 674898 544808
rect 675110 544796 675116 544808
rect 674892 544768 675116 544796
rect 674892 544756 674898 544768
rect 675110 544756 675116 544768
rect 675168 544756 675174 544808
rect 673730 544552 673736 544604
rect 673788 544592 673794 544604
rect 674282 544592 674288 544604
rect 673788 544564 674288 544592
rect 673788 544552 673794 544564
rect 674282 544552 674288 544564
rect 674340 544552 674346 544604
rect 673270 544416 673276 544468
rect 673328 544456 673334 544468
rect 673730 544456 673736 544468
rect 673328 544428 673736 544456
rect 673328 544416 673334 544428
rect 673730 544416 673736 544428
rect 673788 544416 673794 544468
rect 675386 543668 675392 543720
rect 675444 543708 675450 543720
rect 679434 543708 679440 543720
rect 675444 543680 679440 543708
rect 675444 543668 675450 543680
rect 679434 543668 679440 543680
rect 679492 543668 679498 543720
rect 674834 542104 674840 542156
rect 674892 542144 674898 542156
rect 675294 542144 675300 542156
rect 674892 542116 675300 542144
rect 674892 542104 674898 542116
rect 675294 542104 675300 542116
rect 675352 542104 675358 542156
rect 41782 541016 41788 541068
rect 41840 541016 41846 541068
rect 42242 541016 42248 541068
rect 42300 541016 42306 541068
rect 43070 541016 43076 541068
rect 43128 541056 43134 541068
rect 59262 541056 59268 541068
rect 43128 541028 59268 541056
rect 43128 541016 43134 541028
rect 59262 541016 59268 541028
rect 59320 541016 59326 541068
rect 41800 540796 41828 541016
rect 42260 540988 42288 541016
rect 59446 540988 59452 541000
rect 42260 540960 59452 540988
rect 59446 540948 59452 540960
rect 59504 540948 59510 541000
rect 41782 540744 41788 540796
rect 41840 540744 41846 540796
rect 42058 538908 42064 538960
rect 42116 538948 42122 538960
rect 43346 538948 43352 538960
rect 42116 538920 43352 538948
rect 42116 538908 42122 538920
rect 43346 538908 43352 538920
rect 43404 538908 43410 538960
rect 42242 538092 42248 538144
rect 42300 538132 42306 538144
rect 43070 538132 43076 538144
rect 42300 538104 43076 538132
rect 42300 538092 42306 538104
rect 43070 538092 43076 538104
rect 43128 538092 43134 538144
rect 42058 537072 42064 537124
rect 42116 537112 42122 537124
rect 43162 537112 43168 537124
rect 42116 537084 43168 537112
rect 42116 537072 42122 537084
rect 43162 537072 43168 537084
rect 43220 537072 43226 537124
rect 655882 535712 655888 535764
rect 655940 535752 655946 535764
rect 676030 535752 676036 535764
rect 655940 535724 676036 535752
rect 655940 535712 655946 535724
rect 676030 535712 676036 535724
rect 676088 535712 676094 535764
rect 42150 535576 42156 535628
rect 42208 535616 42214 535628
rect 43254 535616 43260 535628
rect 42208 535588 43260 535616
rect 42208 535576 42214 535588
rect 43254 535576 43260 535588
rect 43312 535576 43318 535628
rect 655698 535576 655704 535628
rect 655756 535616 655762 535628
rect 676214 535616 676220 535628
rect 655756 535588 676220 535616
rect 655756 535576 655762 535588
rect 676214 535576 676220 535588
rect 676272 535576 676278 535628
rect 42058 535032 42064 535084
rect 42116 535072 42122 535084
rect 43714 535072 43720 535084
rect 42116 535044 43720 535072
rect 42116 535032 42122 535044
rect 43714 535032 43720 535044
rect 43772 535032 43778 535084
rect 42150 534420 42156 534472
rect 42208 534460 42214 534472
rect 43622 534460 43628 534472
rect 42208 534432 43628 534460
rect 42208 534420 42214 534432
rect 43622 534420 43628 534432
rect 43680 534420 43686 534472
rect 673362 534080 673368 534132
rect 673420 534120 673426 534132
rect 676030 534120 676036 534132
rect 673420 534092 676036 534120
rect 673420 534080 673426 534092
rect 676030 534080 676036 534092
rect 676088 534080 676094 534132
rect 42150 533944 42156 533996
rect 42208 533984 42214 533996
rect 43346 533984 43352 533996
rect 42208 533956 43352 533984
rect 42208 533944 42214 533956
rect 43346 533944 43352 533956
rect 43404 533944 43410 533996
rect 655790 532856 655796 532908
rect 655848 532896 655854 532908
rect 678974 532896 678980 532908
rect 655848 532868 678980 532896
rect 655848 532856 655854 532868
rect 678974 532856 678980 532868
rect 679032 532856 679038 532908
rect 674926 532788 674932 532840
rect 674984 532828 674990 532840
rect 674984 532800 679020 532828
rect 674984 532788 674990 532800
rect 678992 532772 679020 532800
rect 675202 532720 675208 532772
rect 675260 532760 675266 532772
rect 676214 532760 676220 532772
rect 675260 532732 676220 532760
rect 675260 532720 675266 532732
rect 676214 532720 676220 532732
rect 676272 532720 676278 532772
rect 678974 532720 678980 532772
rect 679032 532720 679038 532772
rect 42150 531428 42156 531480
rect 42208 531468 42214 531480
rect 43438 531468 43444 531480
rect 42208 531440 43444 531468
rect 42208 531428 42214 531440
rect 43438 531428 43444 531440
rect 43496 531428 43502 531480
rect 42150 530680 42156 530732
rect 42208 530720 42214 530732
rect 42334 530720 42340 530732
rect 42208 530692 42340 530720
rect 42208 530680 42214 530692
rect 42334 530680 42340 530692
rect 42392 530680 42398 530732
rect 43254 529932 43260 529984
rect 43312 529972 43318 529984
rect 58526 529972 58532 529984
rect 43312 529944 58532 529972
rect 43312 529932 43318 529944
rect 58526 529932 58532 529944
rect 58584 529932 58590 529984
rect 50982 529864 50988 529916
rect 51040 529904 51046 529916
rect 58342 529904 58348 529916
rect 51040 529876 58348 529904
rect 51040 529864 51046 529876
rect 58342 529864 58348 529876
rect 58400 529864 58406 529916
rect 674650 529864 674656 529916
rect 674708 529904 674714 529916
rect 676030 529904 676036 529916
rect 674708 529876 676036 529904
rect 674708 529864 674714 529876
rect 676030 529864 676036 529876
rect 676088 529864 676094 529916
rect 673638 529796 673644 529848
rect 673696 529836 673702 529848
rect 675754 529836 675760 529848
rect 673696 529808 675760 529836
rect 673696 529796 673702 529808
rect 675754 529796 675760 529808
rect 675812 529796 675818 529848
rect 42150 529456 42156 529508
rect 42208 529496 42214 529508
rect 43070 529496 43076 529508
rect 42208 529468 43076 529496
rect 42208 529456 42214 529468
rect 43070 529456 43076 529468
rect 43128 529456 43134 529508
rect 42150 527756 42156 527808
rect 42208 527796 42214 527808
rect 42426 527796 42432 527808
rect 42208 527768 42432 527796
rect 42208 527756 42214 527768
rect 42426 527756 42432 527768
rect 42484 527756 42490 527808
rect 56502 527076 56508 527128
rect 56560 527116 56566 527128
rect 60642 527116 60648 527128
rect 56560 527088 60648 527116
rect 56560 527076 56566 527088
rect 60642 527076 60648 527088
rect 60700 527076 60706 527128
rect 674466 527076 674472 527128
rect 674524 527116 674530 527128
rect 676030 527116 676036 527128
rect 674524 527088 676036 527116
rect 674524 527076 674530 527088
rect 676030 527076 676036 527088
rect 676088 527076 676094 527128
rect 53926 527008 53932 527060
rect 53984 527048 53990 527060
rect 59354 527048 59360 527060
rect 53984 527020 59360 527048
rect 53984 527008 53990 527020
rect 59354 527008 59360 527020
rect 59412 527008 59418 527060
rect 42150 526396 42156 526448
rect 42208 526436 42214 526448
rect 43162 526436 43168 526448
rect 42208 526408 43168 526436
rect 42208 526396 42214 526408
rect 43162 526396 43168 526408
rect 43220 526396 43226 526448
rect 42150 525716 42156 525768
rect 42208 525756 42214 525768
rect 43254 525756 43260 525768
rect 42208 525728 43260 525756
rect 42208 525716 42214 525728
rect 43254 525716 43260 525728
rect 43312 525716 43318 525768
rect 672442 524424 672448 524476
rect 672500 524464 672506 524476
rect 678974 524464 678980 524476
rect 672500 524436 678980 524464
rect 672500 524424 672506 524436
rect 678974 524424 678980 524436
rect 679032 524424 679038 524476
rect 674742 493348 674748 493400
rect 674800 493388 674806 493400
rect 675846 493388 675852 493400
rect 674800 493360 675852 493388
rect 674800 493348 674806 493360
rect 675846 493348 675852 493360
rect 675904 493348 675910 493400
rect 673454 492532 673460 492584
rect 673512 492572 673518 492584
rect 675478 492572 675484 492584
rect 673512 492544 675484 492572
rect 673512 492532 673518 492544
rect 675478 492532 675484 492544
rect 675536 492532 675542 492584
rect 675386 492328 675392 492380
rect 675444 492368 675450 492380
rect 676030 492368 676036 492380
rect 675444 492340 676036 492368
rect 675444 492328 675450 492340
rect 676030 492328 676036 492340
rect 676088 492328 676094 492380
rect 655606 491648 655612 491700
rect 655664 491688 655670 491700
rect 676030 491688 676036 491700
rect 655664 491660 676036 491688
rect 655664 491648 655670 491660
rect 676030 491648 676036 491660
rect 676088 491648 676094 491700
rect 655514 491512 655520 491564
rect 655572 491552 655578 491564
rect 676030 491552 676036 491564
rect 655572 491524 676036 491552
rect 655572 491512 655578 491524
rect 676030 491512 676036 491524
rect 676088 491512 676094 491564
rect 655422 491376 655428 491428
rect 655480 491416 655486 491428
rect 675938 491416 675944 491428
rect 655480 491388 675944 491416
rect 655480 491376 655486 491388
rect 675938 491376 675944 491388
rect 675996 491376 676002 491428
rect 676214 491240 676220 491292
rect 676272 491280 676278 491292
rect 677410 491280 677416 491292
rect 676272 491252 677416 491280
rect 676272 491240 676278 491252
rect 677410 491240 677416 491252
rect 677468 491240 677474 491292
rect 676214 488520 676220 488572
rect 676272 488560 676278 488572
rect 677482 488560 677488 488572
rect 676272 488532 677488 488560
rect 676272 488520 676278 488532
rect 677482 488520 677488 488532
rect 677540 488520 677546 488572
rect 674834 485732 674840 485784
rect 674892 485772 674898 485784
rect 676030 485772 676036 485784
rect 674892 485744 676036 485772
rect 674892 485732 674898 485744
rect 676030 485732 676036 485744
rect 676088 485732 676094 485784
rect 674558 485664 674564 485716
rect 674616 485704 674622 485716
rect 675938 485704 675944 485716
rect 674616 485676 675944 485704
rect 674616 485664 674622 485676
rect 675938 485664 675944 485676
rect 675996 485664 676002 485716
rect 673822 485596 673828 485648
rect 673880 485636 673886 485648
rect 675846 485636 675852 485648
rect 673880 485608 675852 485636
rect 673880 485596 673886 485608
rect 675846 485596 675852 485608
rect 675904 485596 675910 485648
rect 675018 485460 675024 485512
rect 675076 485500 675082 485512
rect 676030 485500 676036 485512
rect 675076 485472 676036 485500
rect 675076 485460 675082 485472
rect 676030 485460 676036 485472
rect 676088 485460 676094 485512
rect 673546 483420 673552 483472
rect 673604 483460 673610 483472
rect 676030 483460 676036 483472
rect 673604 483432 676036 483460
rect 673604 483420 673610 483432
rect 676030 483420 676036 483432
rect 676088 483420 676094 483472
rect 674282 482944 674288 482996
rect 674340 482984 674346 482996
rect 676030 482984 676036 482996
rect 674340 482956 676036 482984
rect 674340 482944 674346 482956
rect 676030 482944 676036 482956
rect 676088 482944 676094 482996
rect 673730 482876 673736 482928
rect 673788 482916 673794 482928
rect 675938 482916 675944 482928
rect 673788 482888 675944 482916
rect 673788 482876 673794 482888
rect 675938 482876 675944 482888
rect 675996 482876 676002 482928
rect 672534 480700 672540 480752
rect 672592 480740 672598 480752
rect 676030 480740 676036 480752
rect 672592 480712 676036 480740
rect 672592 480700 672598 480712
rect 676030 480700 676036 480712
rect 676088 480700 676094 480752
rect 676122 475396 676128 475448
rect 676180 475436 676186 475448
rect 679160 475436 679166 475448
rect 676180 475408 679166 475436
rect 676180 475396 676186 475408
rect 679160 475396 679166 475408
rect 679218 475396 679224 475448
rect 676030 475208 676036 475260
rect 676088 475248 676094 475260
rect 679618 475248 679624 475260
rect 676088 475220 679624 475248
rect 676088 475208 676094 475220
rect 679618 475208 679624 475220
rect 679676 475208 679682 475260
rect 675938 475016 675944 475068
rect 675996 475056 676002 475068
rect 679434 475056 679440 475068
rect 675996 475028 679440 475056
rect 675996 475016 676002 475028
rect 679434 475016 679440 475028
rect 679492 475016 679498 475068
rect 41782 430856 41788 430908
rect 41840 430896 41846 430908
rect 56502 430896 56508 430908
rect 41840 430868 56508 430896
rect 41840 430856 41846 430868
rect 56502 430856 56508 430868
rect 56560 430856 56566 430908
rect 41782 419432 41788 419484
rect 41840 419472 41846 419484
rect 45922 419472 45928 419484
rect 41840 419444 45928 419472
rect 41840 419432 41846 419444
rect 45922 419432 45928 419444
rect 45980 419432 45986 419484
rect 41966 416644 41972 416696
rect 42024 416684 42030 416696
rect 43162 416684 43168 416696
rect 42024 416656 43168 416684
rect 42024 416644 42030 416656
rect 43162 416644 43168 416656
rect 43220 416644 43226 416696
rect 41874 416576 41880 416628
rect 41932 416616 41938 416628
rect 43070 416616 43076 416628
rect 41932 416588 43076 416616
rect 41932 416576 41938 416588
rect 43070 416576 43076 416588
rect 43128 416576 43134 416628
rect 42334 411204 42340 411256
rect 42392 411244 42398 411256
rect 43070 411244 43076 411256
rect 42392 411216 43076 411244
rect 42392 411204 42398 411216
rect 43070 411204 43076 411216
rect 43128 411204 43134 411256
rect 43070 410796 43076 410848
rect 43128 410836 43134 410848
rect 43806 410836 43812 410848
rect 43128 410808 43812 410836
rect 43128 410796 43134 410808
rect 43806 410796 43812 410808
rect 43864 410796 43870 410848
rect 43806 409844 43812 409896
rect 43864 409884 43870 409896
rect 43990 409884 43996 409896
rect 43864 409856 43996 409884
rect 43864 409844 43870 409856
rect 43990 409844 43996 409856
rect 44048 409844 44054 409896
rect 43990 409708 43996 409760
rect 44048 409748 44054 409760
rect 44174 409748 44180 409760
rect 44048 409720 44180 409748
rect 44048 409708 44054 409720
rect 44174 409708 44180 409720
rect 44232 409708 44238 409760
rect 42242 409504 42248 409556
rect 42300 409544 42306 409556
rect 42300 409516 42380 409544
rect 42300 409504 42306 409516
rect 42352 409352 42380 409516
rect 42334 409300 42340 409352
rect 42392 409300 42398 409352
rect 42058 408008 42064 408060
rect 42116 408048 42122 408060
rect 43254 408048 43260 408060
rect 42116 408020 43260 408048
rect 42116 408008 42122 408020
rect 43254 408008 43260 408020
rect 43312 408008 43318 408060
rect 42150 407872 42156 407924
rect 42208 407912 42214 407924
rect 42334 407912 42340 407924
rect 42208 407884 42340 407912
rect 42208 407872 42214 407884
rect 42334 407872 42340 407884
rect 42392 407872 42398 407924
rect 42150 407600 42156 407652
rect 42208 407640 42214 407652
rect 43162 407640 43168 407652
rect 42208 407612 43168 407640
rect 42208 407600 42214 407612
rect 43162 407600 43168 407612
rect 43220 407600 43226 407652
rect 42058 406784 42064 406836
rect 42116 406824 42122 406836
rect 43346 406824 43352 406836
rect 42116 406796 43352 406824
rect 42116 406784 42122 406796
rect 43346 406784 43352 406796
rect 43404 406784 43410 406836
rect 42150 406172 42156 406224
rect 42208 406212 42214 406224
rect 43622 406212 43628 406224
rect 42208 406184 43628 406212
rect 42208 406172 42214 406184
rect 43622 406172 43628 406184
rect 43680 406172 43686 406224
rect 42242 405628 42248 405680
rect 42300 405668 42306 405680
rect 58158 405668 58164 405680
rect 42300 405640 58164 405668
rect 42300 405628 42306 405640
rect 58158 405628 58164 405640
rect 58216 405628 58222 405680
rect 42242 405492 42248 405544
rect 42300 405532 42306 405544
rect 43070 405532 43076 405544
rect 42300 405504 43076 405532
rect 42300 405492 42306 405504
rect 43070 405492 43076 405504
rect 43128 405492 43134 405544
rect 42426 405152 42432 405204
rect 42484 405192 42490 405204
rect 42702 405192 42708 405204
rect 42484 405164 42708 405192
rect 42484 405152 42490 405164
rect 42702 405152 42708 405164
rect 42760 405152 42766 405204
rect 42150 403860 42156 403912
rect 42208 403900 42214 403912
rect 43990 403900 43996 403912
rect 42208 403872 43996 403900
rect 42208 403860 42214 403872
rect 43990 403860 43996 403872
rect 44048 403860 44054 403912
rect 42150 403316 42156 403368
rect 42208 403356 42214 403368
rect 44082 403356 44088 403368
rect 42208 403328 44088 403356
rect 42208 403316 42214 403328
rect 44082 403316 44088 403328
rect 44140 403316 44146 403368
rect 655698 403112 655704 403164
rect 655756 403152 655762 403164
rect 676214 403152 676220 403164
rect 655756 403124 676220 403152
rect 655756 403112 655762 403124
rect 676214 403112 676220 403124
rect 676272 403112 676278 403164
rect 655514 403044 655520 403096
rect 655572 403084 655578 403096
rect 676306 403084 676312 403096
rect 655572 403056 676312 403084
rect 655572 403044 655578 403056
rect 676306 403044 676312 403056
rect 676364 403044 676370 403096
rect 655422 402976 655428 403028
rect 655480 403016 655486 403028
rect 675846 403016 675852 403028
rect 655480 402988 675852 403016
rect 655480 402976 655486 402988
rect 675846 402976 675852 402988
rect 675904 402976 675910 403028
rect 42334 402908 42340 402960
rect 42392 402948 42398 402960
rect 58158 402948 58164 402960
rect 42392 402920 58164 402948
rect 42392 402908 42398 402920
rect 58158 402908 58164 402920
rect 58216 402908 58222 402960
rect 42334 402772 42340 402824
rect 42392 402812 42398 402824
rect 43530 402812 43536 402824
rect 42392 402784 43536 402812
rect 42392 402772 42398 402784
rect 43530 402772 43536 402784
rect 43588 402772 43594 402824
rect 42334 400596 42340 400648
rect 42392 400636 42398 400648
rect 43438 400636 43444 400648
rect 42392 400608 43444 400636
rect 42392 400596 42398 400608
rect 43438 400596 43444 400608
rect 43496 400596 43502 400648
rect 42334 399644 42340 399696
rect 42392 399684 42398 399696
rect 43806 399684 43812 399696
rect 42392 399656 43812 399684
rect 42392 399644 42398 399656
rect 43806 399644 43812 399656
rect 43864 399644 43870 399696
rect 56502 399644 56508 399696
rect 56560 399684 56566 399696
rect 58158 399684 58164 399696
rect 56560 399656 58164 399684
rect 56560 399644 56566 399656
rect 58158 399644 58164 399656
rect 58216 399644 58222 399696
rect 674466 398216 674472 398268
rect 674524 398256 674530 398268
rect 676030 398256 676036 398268
rect 674524 398228 676036 398256
rect 674524 398216 674530 398228
rect 676030 398216 676036 398228
rect 676088 398216 676094 398268
rect 674558 397604 674564 397656
rect 674616 397644 674622 397656
rect 675938 397644 675944 397656
rect 674616 397616 675944 397644
rect 674616 397604 674622 397616
rect 675938 397604 675944 397616
rect 675996 397604 676002 397656
rect 673730 397536 673736 397588
rect 673788 397576 673794 397588
rect 676122 397576 676128 397588
rect 673788 397548 676128 397576
rect 673788 397536 673794 397548
rect 676122 397536 676128 397548
rect 676180 397536 676186 397588
rect 674650 397468 674656 397520
rect 674708 397508 674714 397520
rect 676030 397508 676036 397520
rect 674708 397480 676036 397508
rect 674708 397468 674714 397480
rect 676030 397468 676036 397480
rect 676088 397468 676094 397520
rect 674282 396992 674288 397044
rect 674340 397032 674346 397044
rect 676030 397032 676036 397044
rect 674340 397004 676036 397032
rect 674340 396992 674346 397004
rect 676030 396992 676036 397004
rect 676088 396992 676094 397044
rect 673454 395360 673460 395412
rect 673512 395400 673518 395412
rect 675846 395400 675852 395412
rect 673512 395372 675852 395400
rect 673512 395360 673518 395372
rect 675846 395360 675852 395372
rect 675904 395360 675910 395412
rect 674834 394952 674840 395004
rect 674892 394992 674898 395004
rect 675938 394992 675944 395004
rect 674892 394964 675944 394992
rect 674892 394952 674898 394964
rect 675938 394952 675944 394964
rect 675996 394952 676002 395004
rect 673546 394884 673552 394936
rect 673604 394924 673610 394936
rect 675846 394924 675852 394936
rect 673604 394896 675852 394924
rect 673604 394884 673610 394896
rect 675846 394884 675852 394896
rect 675904 394884 675910 394936
rect 675018 394816 675024 394868
rect 675076 394856 675082 394868
rect 676122 394856 676128 394868
rect 675076 394828 676128 394856
rect 675076 394816 675082 394828
rect 676122 394816 676128 394828
rect 676180 394816 676186 394868
rect 675110 394748 675116 394800
rect 675168 394788 675174 394800
rect 675938 394788 675944 394800
rect 675168 394760 675944 394788
rect 675168 394748 675174 394760
rect 675938 394748 675944 394760
rect 675996 394748 676002 394800
rect 675202 394680 675208 394732
rect 675260 394720 675266 394732
rect 676030 394720 676036 394732
rect 675260 394692 676036 394720
rect 675260 394680 675266 394692
rect 676030 394680 676036 394692
rect 676088 394680 676094 394732
rect 42150 394612 42156 394664
rect 42208 394652 42214 394664
rect 58894 394652 58900 394664
rect 42208 394624 58900 394652
rect 42208 394612 42214 394624
rect 58894 394612 58900 394624
rect 58952 394612 58958 394664
rect 673638 394136 673644 394188
rect 673696 394176 673702 394188
rect 676030 394176 676036 394188
rect 673696 394148 676036 394176
rect 673696 394136 673702 394148
rect 676030 394136 676036 394148
rect 676088 394136 676094 394188
rect 672810 392028 672816 392080
rect 672868 392068 672874 392080
rect 678974 392068 678980 392080
rect 672868 392040 678980 392068
rect 672868 392028 672874 392040
rect 678974 392028 678980 392040
rect 679032 392028 679038 392080
rect 673822 391960 673828 392012
rect 673880 392000 673886 392012
rect 676030 392000 676036 392012
rect 673880 391972 676036 392000
rect 673880 391960 673886 391972
rect 676030 391960 676036 391972
rect 676088 391960 676094 392012
rect 41506 387812 41512 387864
rect 41564 387852 41570 387864
rect 53926 387852 53932 387864
rect 41564 387824 53932 387852
rect 41564 387812 41570 387824
rect 53926 387812 53932 387824
rect 53984 387812 53990 387864
rect 41782 387744 41788 387796
rect 41840 387784 41846 387796
rect 56502 387784 56508 387796
rect 41840 387756 56508 387784
rect 41840 387744 41846 387756
rect 56502 387744 56508 387756
rect 56560 387744 56566 387796
rect 41506 386656 41512 386708
rect 41564 386696 41570 386708
rect 50982 386696 50988 386708
rect 41564 386668 50988 386696
rect 41564 386656 41570 386668
rect 50982 386656 50988 386668
rect 51040 386656 51046 386708
rect 675754 386588 675760 386640
rect 675812 386588 675818 386640
rect 675772 386028 675800 386588
rect 673362 385976 673368 386028
rect 673420 386016 673426 386028
rect 674558 386016 674564 386028
rect 673420 385988 674564 386016
rect 673420 385976 673426 385988
rect 674558 385976 674564 385988
rect 674616 385976 674622 386028
rect 675386 385976 675392 386028
rect 675444 385976 675450 386028
rect 675754 385976 675760 386028
rect 675812 385976 675818 386028
rect 674558 385840 674564 385892
rect 674616 385880 674622 385892
rect 675404 385880 675432 385976
rect 674616 385852 675432 385880
rect 674616 385840 674622 385852
rect 675202 385568 675208 385620
rect 675260 385608 675266 385620
rect 675386 385608 675392 385620
rect 675260 385580 675392 385608
rect 675260 385568 675266 385580
rect 675386 385568 675392 385580
rect 675444 385568 675450 385620
rect 673730 384956 673736 385008
rect 673788 384996 673794 385008
rect 675202 384996 675208 385008
rect 673788 384968 675208 384996
rect 673788 384956 673794 384968
rect 675202 384956 675208 384968
rect 675260 384956 675266 385008
rect 674466 384752 674472 384804
rect 674524 384792 674530 384804
rect 675386 384792 675392 384804
rect 674524 384764 675392 384792
rect 674524 384752 674530 384764
rect 675386 384752 675392 384764
rect 675444 384752 675450 384804
rect 673362 384684 673368 384736
rect 673420 384724 673426 384736
rect 673638 384724 673644 384736
rect 673420 384696 673644 384724
rect 673420 384684 673426 384696
rect 673638 384684 673644 384696
rect 673696 384684 673702 384736
rect 674650 383120 674656 383172
rect 674708 383160 674714 383172
rect 675386 383160 675392 383172
rect 674708 383132 675392 383160
rect 674708 383120 674714 383132
rect 675386 383120 675392 383132
rect 675444 383120 675450 383172
rect 675018 382440 675024 382492
rect 675076 382480 675082 382492
rect 675386 382480 675392 382492
rect 675076 382452 675392 382480
rect 675076 382440 675082 382452
rect 675386 382440 675392 382452
rect 675444 382440 675450 382492
rect 674834 381896 674840 381948
rect 674892 381936 674898 381948
rect 675386 381936 675392 381948
rect 674892 381908 675392 381936
rect 674892 381896 674898 381908
rect 675386 381896 675392 381908
rect 675444 381896 675450 381948
rect 675110 381284 675116 381336
rect 675168 381324 675174 381336
rect 675386 381324 675392 381336
rect 675168 381296 675392 381324
rect 675168 381284 675174 381296
rect 675386 381284 675392 381296
rect 675444 381284 675450 381336
rect 674282 381148 674288 381200
rect 674340 381188 674346 381200
rect 675110 381188 675116 381200
rect 674340 381160 675116 381188
rect 674340 381148 674346 381160
rect 675110 381148 675116 381160
rect 675168 381148 675174 381200
rect 43438 379448 43444 379500
rect 43496 379448 43502 379500
rect 43346 379176 43352 379228
rect 43404 379216 43410 379228
rect 43456 379216 43484 379448
rect 43530 379312 43536 379364
rect 43588 379352 43594 379364
rect 44082 379352 44088 379364
rect 43588 379324 44088 379352
rect 43588 379312 43594 379324
rect 44082 379312 44088 379324
rect 44140 379312 44146 379364
rect 43404 379188 43484 379216
rect 43404 379176 43410 379188
rect 673638 378768 673644 378820
rect 673696 378808 673702 378820
rect 675386 378808 675392 378820
rect 673696 378780 675392 378808
rect 673696 378768 673702 378780
rect 675386 378768 675392 378780
rect 675444 378768 675450 378820
rect 673730 378156 673736 378208
rect 673788 378196 673794 378208
rect 675478 378196 675484 378208
rect 673788 378168 675484 378196
rect 673788 378156 673794 378168
rect 675478 378156 675484 378168
rect 675536 378156 675542 378208
rect 673546 377408 673552 377460
rect 673604 377448 673610 377460
rect 675386 377448 675392 377460
rect 673604 377420 675392 377448
rect 673604 377408 673610 377420
rect 675386 377408 675392 377420
rect 675444 377408 675450 377460
rect 673822 376932 673828 376984
rect 673880 376972 673886 376984
rect 675478 376972 675484 376984
rect 673880 376944 675484 376972
rect 673880 376932 673886 376944
rect 675478 376932 675484 376944
rect 675536 376932 675542 376984
rect 41782 376184 41788 376236
rect 41840 376224 41846 376236
rect 46014 376224 46020 376236
rect 41840 376196 46020 376224
rect 41840 376184 41846 376196
rect 46014 376184 46020 376196
rect 46072 376184 46078 376236
rect 673454 375708 673460 375760
rect 673512 375748 673518 375760
rect 675386 375748 675392 375760
rect 673512 375720 675392 375748
rect 673512 375708 673518 375720
rect 675386 375708 675392 375720
rect 675444 375708 675450 375760
rect 38194 375300 38200 375352
rect 38252 375340 38258 375352
rect 42242 375340 42248 375352
rect 38252 375312 42248 375340
rect 38252 375300 38258 375312
rect 42242 375300 42248 375312
rect 42300 375300 42306 375352
rect 41414 375232 41420 375284
rect 41472 375272 41478 375284
rect 43254 375272 43260 375284
rect 41472 375244 43260 375272
rect 41472 375232 41478 375244
rect 43254 375232 43260 375244
rect 43312 375232 43318 375284
rect 42334 374212 42340 374264
rect 42392 374252 42398 374264
rect 42702 374252 42708 374264
rect 42392 374224 42708 374252
rect 42392 374212 42398 374224
rect 42702 374212 42708 374224
rect 42760 374212 42766 374264
rect 675018 373464 675024 373516
rect 675076 373504 675082 373516
rect 675294 373504 675300 373516
rect 675076 373476 675300 373504
rect 675076 373464 675082 373476
rect 675294 373464 675300 373476
rect 675352 373464 675358 373516
rect 41598 372784 41604 372836
rect 41656 372824 41662 372836
rect 43990 372824 43996 372836
rect 41656 372796 43996 372824
rect 41656 372784 41662 372796
rect 43990 372784 43996 372796
rect 44048 372784 44054 372836
rect 654502 372512 654508 372564
rect 654560 372552 654566 372564
rect 674558 372552 674564 372564
rect 654560 372524 674564 372552
rect 654560 372512 654566 372524
rect 674558 372512 674564 372524
rect 674616 372512 674622 372564
rect 41506 371424 41512 371476
rect 41564 371464 41570 371476
rect 42702 371464 42708 371476
rect 41564 371436 42708 371464
rect 41564 371424 41570 371436
rect 42702 371424 42708 371436
rect 42760 371424 42766 371476
rect 43714 371288 43720 371340
rect 43772 371328 43778 371340
rect 43772 371300 43852 371328
rect 43772 371288 43778 371300
rect 43824 371136 43852 371300
rect 43806 371084 43812 371136
rect 43864 371084 43870 371136
rect 41966 370200 41972 370252
rect 42024 370200 42030 370252
rect 41984 370036 42012 370200
rect 41984 370008 42288 370036
rect 42260 369368 42288 370008
rect 42242 369316 42248 369368
rect 42300 369316 42306 369368
rect 42150 368092 42156 368144
rect 42208 368132 42214 368144
rect 42334 368132 42340 368144
rect 42208 368104 42340 368132
rect 42208 368092 42214 368104
rect 42334 368092 42340 368104
rect 42392 368092 42398 368144
rect 42150 366256 42156 366308
rect 42208 366296 42214 366308
rect 43162 366296 43168 366308
rect 42208 366268 43168 366296
rect 42208 366256 42214 366268
rect 43162 366256 43168 366268
rect 43220 366256 43226 366308
rect 42334 366120 42340 366172
rect 42392 366160 42398 366172
rect 43162 366160 43168 366172
rect 42392 366132 43168 366160
rect 42392 366120 42398 366132
rect 43162 366120 43168 366132
rect 43220 366120 43226 366172
rect 42334 365032 42340 365084
rect 42392 365072 42398 365084
rect 42392 365044 42840 365072
rect 42392 365032 42398 365044
rect 42150 364760 42156 364812
rect 42208 364800 42214 364812
rect 42702 364800 42708 364812
rect 42208 364772 42708 364800
rect 42208 364760 42214 364772
rect 42702 364760 42708 364772
rect 42760 364760 42766 364812
rect 42702 364624 42708 364676
rect 42760 364664 42766 364676
rect 42812 364664 42840 365044
rect 42760 364636 42840 364664
rect 42760 364624 42766 364636
rect 42242 364080 42248 364132
rect 42300 364120 42306 364132
rect 43438 364120 43444 364132
rect 42300 364092 43444 364120
rect 42300 364080 42306 364092
rect 43438 364080 43444 364092
rect 43496 364080 43502 364132
rect 43438 363944 43444 363996
rect 43496 363984 43502 363996
rect 43898 363984 43904 363996
rect 43496 363956 43904 363984
rect 43496 363944 43502 363956
rect 43898 363944 43904 363956
rect 43956 363944 43962 363996
rect 42150 363808 42156 363860
rect 42208 363848 42214 363860
rect 43254 363848 43260 363860
rect 42208 363820 43260 363848
rect 42208 363808 42214 363820
rect 43254 363808 43260 363820
rect 43312 363808 43318 363860
rect 43162 363740 43168 363792
rect 43220 363780 43226 363792
rect 43990 363780 43996 363792
rect 43220 363752 43996 363780
rect 43220 363740 43226 363752
rect 43990 363740 43996 363752
rect 44048 363740 44054 363792
rect 42150 363128 42156 363180
rect 42208 363168 42214 363180
rect 43530 363168 43536 363180
rect 42208 363140 43536 363168
rect 42208 363128 42214 363140
rect 43530 363128 43536 363140
rect 43588 363128 43594 363180
rect 42426 361904 42432 361956
rect 42484 361944 42490 361956
rect 43070 361944 43076 361956
rect 42484 361916 43076 361944
rect 42484 361904 42490 361916
rect 43070 361904 43076 361916
rect 43128 361904 43134 361956
rect 42334 361564 42340 361616
rect 42392 361564 42398 361616
rect 42352 361536 42380 361564
rect 58342 361536 58348 361548
rect 42352 361508 58348 361536
rect 58342 361496 58348 361508
rect 58400 361496 58406 361548
rect 42702 361292 42708 361344
rect 42760 361332 42766 361344
rect 58158 361332 58164 361344
rect 42760 361304 58164 361332
rect 42760 361292 42766 361304
rect 58158 361292 58164 361304
rect 58216 361292 58222 361344
rect 42058 360612 42064 360664
rect 42116 360652 42122 360664
rect 43898 360652 43904 360664
rect 42116 360624 43904 360652
rect 42116 360612 42122 360624
rect 43898 360612 43904 360624
rect 43956 360612 43962 360664
rect 42334 360272 42340 360324
rect 42392 360312 42398 360324
rect 43438 360312 43444 360324
rect 42392 360284 43444 360312
rect 42392 360272 42398 360284
rect 43438 360272 43444 360284
rect 43496 360272 43502 360324
rect 42150 359932 42156 359984
rect 42208 359972 42214 359984
rect 43990 359972 43996 359984
rect 42208 359944 43996 359972
rect 42208 359932 42214 359944
rect 43990 359932 43996 359944
rect 44048 359932 44054 359984
rect 50982 358708 50988 358760
rect 51040 358748 51046 358760
rect 58526 358748 58532 358760
rect 51040 358720 58532 358748
rect 51040 358708 51046 358720
rect 58526 358708 58532 358720
rect 58584 358708 58590 358760
rect 42426 358300 42432 358352
rect 42484 358340 42490 358352
rect 43346 358340 43352 358352
rect 42484 358312 43352 358340
rect 42484 358300 42490 358312
rect 43346 358300 43352 358312
rect 43404 358300 43410 358352
rect 673086 357008 673092 357060
rect 673144 357048 673150 357060
rect 675662 357048 675668 357060
rect 673144 357020 675668 357048
rect 673144 357008 673150 357020
rect 675662 357008 675668 357020
rect 675720 357008 675726 357060
rect 42426 356464 42432 356516
rect 42484 356504 42490 356516
rect 43622 356504 43628 356516
rect 42484 356476 43628 356504
rect 42484 356464 42490 356476
rect 43622 356464 43628 356476
rect 43680 356464 43686 356516
rect 655514 356464 655520 356516
rect 655572 356504 655578 356516
rect 675938 356504 675944 356516
rect 655572 356476 675944 356504
rect 655572 356464 655578 356476
rect 675938 356464 675944 356476
rect 675996 356464 676002 356516
rect 42334 356396 42340 356448
rect 42392 356436 42398 356448
rect 43806 356436 43812 356448
rect 42392 356408 43812 356436
rect 42392 356396 42398 356408
rect 43806 356396 43812 356408
rect 43864 356396 43870 356448
rect 655422 356328 655428 356380
rect 655480 356368 655486 356380
rect 676030 356368 676036 356380
rect 655480 356340 676036 356368
rect 655480 356328 655486 356340
rect 676030 356328 676036 356340
rect 676088 356328 676094 356380
rect 655606 356192 655612 356244
rect 655664 356232 655670 356244
rect 675846 356232 675852 356244
rect 655664 356204 675852 356232
rect 655664 356192 655670 356204
rect 675846 356192 675852 356204
rect 675904 356192 675910 356244
rect 673362 356124 673368 356176
rect 673420 356164 673426 356176
rect 676030 356164 676036 356176
rect 673420 356136 676036 356164
rect 673420 356124 673426 356136
rect 676030 356124 676036 356136
rect 676088 356124 676094 356176
rect 56502 355988 56508 356040
rect 56560 356028 56566 356040
rect 58066 356028 58072 356040
rect 56560 356000 58072 356028
rect 56560 355988 56566 356000
rect 58066 355988 58072 356000
rect 58124 355988 58130 356040
rect 53926 355920 53932 355972
rect 53984 355960 53990 355972
rect 59354 355960 59360 355972
rect 53984 355932 59360 355960
rect 53984 355920 53990 355932
rect 59354 355920 59360 355932
rect 59412 355920 59418 355972
rect 673178 355376 673184 355428
rect 673236 355416 673242 355428
rect 676030 355416 676036 355428
rect 673236 355388 676036 355416
rect 673236 355376 673242 355388
rect 676030 355376 676036 355388
rect 676088 355376 676094 355428
rect 673270 354560 673276 354612
rect 673328 354600 673334 354612
rect 676030 354600 676036 354612
rect 673328 354572 676036 354600
rect 673328 354560 673334 354572
rect 676030 354560 676036 354572
rect 676088 354560 676094 354612
rect 674650 353472 674656 353524
rect 674708 353512 674714 353524
rect 676030 353512 676036 353524
rect 674708 353484 676036 353512
rect 674708 353472 674714 353484
rect 676030 353472 676036 353484
rect 676088 353472 676094 353524
rect 675110 353268 675116 353320
rect 675168 353308 675174 353320
rect 676030 353308 676036 353320
rect 675168 353280 676036 353308
rect 675168 353268 675174 353280
rect 676030 353268 676036 353280
rect 676088 353268 676094 353320
rect 674834 351432 674840 351484
rect 674892 351472 674898 351484
rect 676030 351472 676036 351484
rect 674892 351444 676036 351472
rect 674892 351432 674898 351444
rect 676030 351432 676036 351444
rect 676088 351432 676094 351484
rect 673730 351024 673736 351076
rect 673788 351064 673794 351076
rect 675938 351064 675944 351076
rect 673788 351036 675944 351064
rect 673788 351024 673794 351036
rect 675938 351024 675944 351036
rect 675996 351024 676002 351076
rect 673546 350820 673552 350872
rect 673604 350860 673610 350872
rect 675846 350860 675852 350872
rect 673604 350832 675852 350860
rect 673604 350820 673610 350832
rect 675846 350820 675852 350832
rect 675904 350820 675910 350872
rect 673454 350684 673460 350736
rect 673512 350724 673518 350736
rect 675846 350724 675852 350736
rect 673512 350696 675852 350724
rect 673512 350684 673518 350696
rect 675846 350684 675852 350696
rect 675904 350684 675910 350736
rect 674558 350616 674564 350668
rect 674616 350656 674622 350668
rect 675938 350656 675944 350668
rect 674616 350628 675944 350656
rect 674616 350616 674622 350628
rect 675938 350616 675944 350628
rect 675996 350616 676002 350668
rect 675202 350548 675208 350600
rect 675260 350588 675266 350600
rect 676030 350588 676036 350600
rect 675260 350560 676036 350588
rect 675260 350548 675266 350560
rect 676030 350548 676036 350560
rect 676088 350548 676094 350600
rect 42150 350480 42156 350532
rect 42208 350520 42214 350532
rect 58618 350520 58624 350532
rect 42208 350492 58624 350520
rect 42208 350480 42214 350492
rect 58618 350480 58624 350492
rect 58676 350480 58682 350532
rect 674282 349800 674288 349852
rect 674340 349840 674346 349852
rect 676030 349840 676036 349852
rect 674340 349812 676036 349840
rect 674340 349800 674346 349812
rect 676030 349800 676036 349812
rect 676088 349800 676094 349852
rect 673638 347896 673644 347948
rect 673696 347936 673702 347948
rect 675846 347936 675852 347948
rect 673696 347908 675852 347936
rect 673696 347896 673702 347908
rect 675846 347896 675852 347908
rect 675904 347896 675910 347948
rect 674466 347828 674472 347880
rect 674524 347868 674530 347880
rect 675938 347868 675944 347880
rect 674524 347840 675944 347868
rect 674524 347828 674530 347840
rect 675938 347828 675944 347840
rect 675996 347828 676002 347880
rect 675018 347760 675024 347812
rect 675076 347800 675082 347812
rect 676030 347800 676036 347812
rect 675076 347772 676036 347800
rect 675076 347760 675082 347772
rect 676030 347760 676036 347772
rect 676088 347760 676094 347812
rect 672902 347216 672908 347268
rect 672960 347256 672966 347268
rect 676030 347256 676036 347268
rect 672960 347228 676036 347256
rect 672960 347216 672966 347228
rect 676030 347216 676036 347228
rect 676088 347216 676094 347268
rect 41506 344224 41512 344276
rect 41564 344264 41570 344276
rect 46566 344264 46572 344276
rect 41564 344236 46572 344264
rect 41564 344224 41570 344236
rect 46566 344224 46572 344236
rect 46624 344224 46630 344276
rect 41506 343816 41512 343868
rect 41564 343856 41570 343868
rect 46382 343856 46388 343868
rect 41564 343828 46388 343856
rect 41564 343816 41570 343828
rect 46382 343816 46388 343828
rect 46440 343816 46446 343868
rect 41506 343408 41512 343460
rect 41564 343448 41570 343460
rect 46474 343448 46480 343460
rect 41564 343420 46480 343448
rect 41564 343408 41570 343420
rect 46474 343408 46480 343420
rect 46532 343408 46538 343460
rect 41506 342864 41512 342916
rect 41564 342904 41570 342916
rect 44082 342904 44088 342916
rect 41564 342876 44088 342904
rect 41564 342864 41570 342876
rect 44082 342864 44088 342876
rect 44140 342864 44146 342916
rect 673822 341776 673828 341828
rect 673880 341816 673886 341828
rect 674282 341816 674288 341828
rect 673880 341788 674288 341816
rect 673880 341776 673886 341788
rect 674282 341776 674288 341788
rect 674340 341776 674346 341828
rect 674282 341640 674288 341692
rect 674340 341680 674346 341692
rect 674466 341680 674472 341692
rect 674340 341652 674472 341680
rect 674340 341640 674346 341652
rect 674466 341640 674472 341652
rect 674524 341640 674530 341692
rect 674558 341368 674564 341420
rect 674616 341408 674622 341420
rect 675386 341408 675392 341420
rect 674616 341380 675392 341408
rect 674616 341368 674622 341380
rect 675386 341368 675392 341380
rect 675444 341368 675450 341420
rect 675110 340824 675116 340876
rect 675168 340824 675174 340876
rect 675018 340796 675024 340808
rect 674944 340768 675024 340796
rect 674944 340456 674972 340768
rect 675018 340756 675024 340768
rect 675076 340756 675082 340808
rect 675128 340796 675156 340824
rect 675478 340796 675484 340808
rect 675128 340768 675484 340796
rect 675478 340756 675484 340768
rect 675536 340756 675542 340808
rect 675018 340620 675024 340672
rect 675076 340660 675082 340672
rect 675386 340660 675392 340672
rect 675076 340632 675392 340660
rect 675076 340620 675082 340632
rect 675386 340620 675392 340632
rect 675444 340620 675450 340672
rect 675110 340456 675116 340468
rect 674944 340428 675116 340456
rect 675110 340416 675116 340428
rect 675168 340416 675174 340468
rect 674650 339532 674656 339584
rect 674708 339572 674714 339584
rect 675478 339572 675484 339584
rect 674708 339544 675484 339572
rect 674708 339532 674714 339544
rect 675478 339532 675484 339544
rect 675536 339532 675542 339584
rect 674834 337900 674840 337952
rect 674892 337940 674898 337952
rect 675478 337940 675484 337952
rect 674892 337912 675484 337940
rect 674892 337900 674898 337912
rect 675478 337900 675484 337912
rect 675536 337900 675542 337952
rect 674466 336676 674472 336728
rect 674524 336716 674530 336728
rect 675202 336716 675208 336728
rect 674524 336688 675208 336716
rect 674524 336676 674530 336688
rect 675202 336676 675208 336688
rect 675260 336676 675266 336728
rect 674282 335452 674288 335504
rect 674340 335492 674346 335504
rect 675110 335492 675116 335504
rect 674340 335464 675116 335492
rect 674340 335452 674346 335464
rect 675110 335452 675116 335464
rect 675168 335452 675174 335504
rect 673730 335384 673736 335436
rect 673788 335424 673794 335436
rect 675202 335424 675208 335436
rect 673788 335396 675208 335424
rect 673788 335384 673794 335396
rect 675202 335384 675208 335396
rect 675260 335384 675266 335436
rect 655974 335316 655980 335368
rect 656032 335356 656038 335368
rect 675018 335356 675024 335368
rect 656032 335328 675024 335356
rect 656032 335316 656038 335328
rect 675018 335316 675024 335328
rect 675076 335316 675082 335368
rect 41598 332800 41604 332852
rect 41656 332840 41662 332852
rect 46198 332840 46204 332852
rect 41656 332812 46204 332840
rect 41656 332800 41662 332812
rect 46198 332800 46204 332812
rect 46256 332800 46262 332852
rect 673822 332392 673828 332444
rect 673880 332432 673886 332444
rect 675110 332432 675116 332444
rect 673880 332404 675116 332432
rect 673880 332392 673886 332404
rect 675110 332392 675116 332404
rect 675168 332392 675174 332444
rect 673638 331712 673644 331764
rect 673696 331752 673702 331764
rect 675110 331752 675116 331764
rect 673696 331724 675116 331752
rect 673696 331712 673702 331724
rect 675110 331712 675116 331724
rect 675168 331712 675174 331764
rect 41414 331168 41420 331220
rect 41472 331208 41478 331220
rect 43530 331208 43536 331220
rect 41472 331180 43536 331208
rect 41472 331168 41478 331180
rect 43530 331168 43536 331180
rect 43588 331168 43594 331220
rect 673454 331100 673460 331152
rect 673512 331140 673518 331152
rect 675110 331140 675116 331152
rect 673512 331112 675116 331140
rect 673512 331100 673518 331112
rect 675110 331100 675116 331112
rect 675168 331100 675174 331152
rect 41506 330080 41512 330132
rect 41564 330120 41570 330132
rect 43070 330120 43076 330132
rect 41564 330092 43076 330120
rect 41564 330080 41570 330092
rect 43070 330080 43076 330092
rect 43128 330080 43134 330132
rect 33042 329944 33048 329996
rect 33100 329984 33106 329996
rect 42242 329984 42248 329996
rect 33100 329956 42248 329984
rect 33100 329944 33106 329956
rect 42242 329944 42248 329956
rect 42300 329944 42306 329996
rect 674558 328720 674564 328772
rect 674616 328760 674622 328772
rect 675386 328760 675392 328772
rect 674616 328732 675392 328760
rect 674616 328720 674622 328732
rect 675386 328720 675392 328732
rect 675444 328720 675450 328772
rect 41782 326952 41788 327004
rect 41840 326952 41846 327004
rect 41800 326800 41828 326952
rect 673546 326884 673552 326936
rect 673604 326924 673610 326936
rect 675386 326924 675392 326936
rect 673604 326896 675392 326924
rect 673604 326884 673610 326896
rect 675386 326884 675392 326896
rect 675444 326884 675450 326936
rect 41782 326748 41788 326800
rect 41840 326748 41846 326800
rect 42242 323144 42248 323196
rect 42300 323144 42306 323196
rect 42260 322992 42288 323144
rect 42242 322940 42248 322992
rect 42300 322940 42306 322992
rect 42242 321988 42248 322040
rect 42300 322028 42306 322040
rect 43714 322028 43720 322040
rect 42300 322000 43720 322028
rect 42300 321988 42306 322000
rect 43714 321988 43720 322000
rect 43772 321988 43778 322040
rect 42242 321784 42248 321836
rect 42300 321824 42306 321836
rect 43254 321824 43260 321836
rect 42300 321796 43260 321824
rect 42300 321784 42306 321796
rect 43254 321784 43260 321796
rect 43312 321784 43318 321836
rect 42150 321580 42156 321632
rect 42208 321620 42214 321632
rect 43438 321620 43444 321632
rect 42208 321592 43444 321620
rect 42208 321580 42214 321592
rect 43438 321580 43444 321592
rect 43496 321580 43502 321632
rect 42242 320560 42248 320612
rect 42300 320600 42306 320612
rect 43162 320600 43168 320612
rect 42300 320572 43168 320600
rect 42300 320560 42306 320572
rect 43162 320560 43168 320572
rect 43220 320560 43226 320612
rect 42150 320424 42156 320476
rect 42208 320464 42214 320476
rect 43622 320464 43628 320476
rect 42208 320436 43628 320464
rect 42208 320424 42214 320436
rect 43622 320424 43628 320436
rect 43680 320424 43686 320476
rect 42426 318724 42432 318776
rect 42484 318764 42490 318776
rect 42702 318764 42708 318776
rect 42484 318736 42708 318764
rect 42484 318724 42490 318736
rect 42702 318724 42708 318736
rect 42760 318724 42766 318776
rect 43714 318724 43720 318776
rect 43772 318764 43778 318776
rect 58434 318764 58440 318776
rect 43772 318736 58440 318764
rect 43772 318724 43778 318736
rect 58434 318724 58440 318736
rect 58492 318724 58498 318776
rect 42334 317364 42340 317416
rect 42392 317404 42398 317416
rect 58158 317404 58164 317416
rect 42392 317376 58164 317404
rect 42392 317364 42398 317376
rect 58158 317364 58164 317376
rect 58216 317364 58222 317416
rect 42426 316888 42432 316940
rect 42484 316928 42490 316940
rect 43070 316928 43076 316940
rect 42484 316900 43076 316928
rect 42484 316888 42490 316900
rect 43070 316888 43076 316900
rect 43128 316888 43134 316940
rect 42334 316820 42340 316872
rect 42392 316860 42398 316872
rect 43530 316860 43536 316872
rect 42392 316832 43536 316860
rect 42392 316820 42398 316832
rect 43530 316820 43536 316832
rect 43588 316820 43594 316872
rect 46474 314576 46480 314628
rect 46532 314616 46538 314628
rect 58526 314616 58532 314628
rect 46532 314588 58532 314616
rect 46532 314576 46538 314588
rect 58526 314576 58532 314588
rect 58584 314576 58590 314628
rect 46566 314508 46572 314560
rect 46624 314548 46630 314560
rect 58158 314548 58164 314560
rect 46624 314520 58164 314548
rect 46624 314508 46630 314520
rect 58158 314508 58164 314520
rect 58216 314508 58222 314560
rect 673086 312400 673092 312452
rect 673144 312440 673150 312452
rect 676030 312440 676036 312452
rect 673144 312412 676036 312440
rect 673144 312400 673150 312412
rect 676030 312400 676036 312412
rect 676088 312400 676094 312452
rect 655422 312128 655428 312180
rect 655480 312168 655486 312180
rect 676214 312168 676220 312180
rect 655480 312140 676220 312168
rect 655480 312128 655486 312140
rect 676214 312128 676220 312140
rect 676272 312128 676278 312180
rect 655698 311992 655704 312044
rect 655756 312032 655762 312044
rect 676306 312032 676312 312044
rect 655756 312004 676312 312032
rect 655756 311992 655762 312004
rect 676306 311992 676312 312004
rect 676364 311992 676370 312044
rect 655514 311924 655520 311976
rect 655572 311964 655578 311976
rect 676122 311964 676128 311976
rect 655572 311936 676128 311964
rect 655572 311924 655578 311936
rect 676122 311924 676128 311936
rect 676180 311924 676186 311976
rect 671614 311856 671620 311908
rect 671672 311896 671678 311908
rect 676214 311896 676220 311908
rect 671672 311868 676220 311896
rect 671672 311856 671678 311868
rect 676214 311856 676220 311868
rect 676272 311856 676278 311908
rect 46382 311788 46388 311840
rect 46440 311828 46446 311840
rect 58526 311828 58532 311840
rect 46440 311800 58532 311828
rect 46440 311788 46446 311800
rect 58526 311788 58532 311800
rect 58584 311788 58590 311840
rect 673362 311652 673368 311704
rect 673420 311692 673426 311704
rect 676030 311692 676036 311704
rect 673420 311664 676036 311692
rect 673420 311652 673426 311664
rect 676030 311652 676036 311664
rect 676088 311652 676094 311704
rect 673362 311040 673368 311092
rect 673420 311080 673426 311092
rect 676214 311080 676220 311092
rect 673420 311052 676220 311080
rect 673420 311040 673426 311052
rect 676214 311040 676220 311052
rect 676272 311040 676278 311092
rect 673178 310632 673184 310684
rect 673236 310672 673242 310684
rect 676214 310672 676220 310684
rect 673236 310644 676220 310672
rect 673236 310632 673242 310644
rect 676214 310632 676220 310644
rect 676272 310632 676278 310684
rect 671706 310224 671712 310276
rect 671764 310264 671770 310276
rect 676214 310264 676220 310276
rect 671764 310236 676220 310264
rect 671764 310224 671770 310236
rect 676214 310224 676220 310236
rect 676272 310224 676278 310276
rect 673270 309856 673276 309868
rect 673268 309828 673276 309856
rect 673270 309816 673276 309828
rect 673328 309856 673334 309868
rect 676214 309856 676220 309868
rect 673328 309828 676220 309856
rect 673328 309816 673334 309828
rect 676214 309816 676220 309828
rect 676272 309816 676278 309868
rect 671798 309408 671804 309460
rect 671856 309448 671862 309460
rect 676214 309448 676220 309460
rect 671856 309420 676220 309448
rect 671856 309408 671862 309420
rect 676214 309408 676220 309420
rect 676272 309408 676278 309460
rect 674650 309136 674656 309188
rect 674708 309176 674714 309188
rect 676030 309176 676036 309188
rect 674708 309148 676036 309176
rect 674708 309136 674714 309148
rect 676030 309136 676036 309148
rect 676088 309136 676094 309188
rect 673454 308048 673460 308100
rect 673512 308088 673518 308100
rect 676030 308088 676036 308100
rect 673512 308060 676036 308088
rect 673512 308048 673518 308060
rect 676030 308048 676036 308060
rect 676088 308048 676094 308100
rect 674466 306824 674472 306876
rect 674524 306864 674530 306876
rect 676030 306864 676036 306876
rect 674524 306836 676036 306864
rect 674524 306824 674530 306836
rect 676030 306824 676036 306836
rect 676088 306824 676094 306876
rect 674558 306416 674564 306468
rect 674616 306456 674622 306468
rect 676030 306456 676036 306468
rect 674616 306428 676036 306456
rect 674616 306416 674622 306428
rect 676030 306416 676036 306428
rect 676088 306416 676094 306468
rect 673546 306348 673552 306400
rect 673604 306388 673610 306400
rect 676122 306388 676128 306400
rect 673604 306360 676128 306388
rect 673604 306348 673610 306360
rect 676122 306348 676128 306360
rect 676180 306348 676186 306400
rect 42058 306280 42064 306332
rect 42116 306320 42122 306332
rect 58342 306320 58348 306332
rect 42116 306292 58348 306320
rect 42116 306280 42122 306292
rect 58342 306280 58348 306292
rect 58400 306280 58406 306332
rect 675202 306008 675208 306060
rect 675260 306048 675266 306060
rect 676030 306048 676036 306060
rect 675260 306020 676036 306048
rect 675260 306008 675266 306020
rect 676030 306008 676036 306020
rect 676088 306008 676094 306060
rect 673638 305056 673644 305108
rect 673696 305096 673702 305108
rect 676122 305096 676128 305108
rect 673696 305068 676128 305096
rect 673696 305056 673702 305068
rect 676122 305056 676128 305068
rect 676180 305056 676186 305108
rect 675018 304784 675024 304836
rect 675076 304824 675082 304836
rect 676030 304824 676036 304836
rect 675076 304796 676036 304824
rect 675076 304784 675082 304796
rect 676030 304784 676036 304796
rect 676088 304784 676094 304836
rect 673822 304308 673828 304360
rect 673880 304348 673886 304360
rect 676122 304348 676128 304360
rect 673880 304320 676128 304348
rect 673880 304308 673886 304320
rect 676122 304308 676128 304320
rect 676180 304308 676186 304360
rect 674834 304172 674840 304224
rect 674892 304212 674898 304224
rect 676030 304212 676036 304224
rect 674892 304184 676036 304212
rect 674892 304172 674898 304184
rect 676030 304172 676036 304184
rect 676088 304172 676094 304224
rect 674282 303900 674288 303952
rect 674340 303940 674346 303952
rect 676122 303940 676128 303952
rect 674340 303912 676128 303940
rect 674340 303900 674346 303912
rect 676122 303900 676128 303912
rect 676180 303900 676186 303952
rect 673730 303696 673736 303748
rect 673788 303736 673794 303748
rect 676030 303736 676036 303748
rect 673788 303708 676036 303736
rect 673788 303696 673794 303708
rect 676030 303696 676036 303708
rect 676088 303696 676094 303748
rect 41874 301384 41880 301436
rect 41932 301424 41938 301436
rect 54018 301424 54024 301436
rect 41932 301396 54024 301424
rect 41932 301384 41938 301396
rect 54018 301384 54024 301396
rect 54076 301384 54082 301436
rect 41782 301316 41788 301368
rect 41840 301356 41846 301368
rect 57882 301356 57888 301368
rect 41840 301328 57888 301356
rect 41840 301316 41846 301328
rect 57882 301316 57888 301328
rect 57940 301316 57946 301368
rect 41782 301180 41788 301232
rect 41840 301220 41846 301232
rect 43346 301220 43352 301232
rect 41840 301192 43352 301220
rect 41840 301180 41846 301192
rect 43346 301180 43352 301192
rect 43404 301180 43410 301232
rect 672994 300840 673000 300892
rect 673052 300880 673058 300892
rect 678974 300880 678980 300892
rect 673052 300852 678980 300880
rect 673052 300840 673058 300852
rect 678974 300840 678980 300852
rect 679032 300840 679038 300892
rect 675110 298256 675116 298308
rect 675168 298296 675174 298308
rect 675386 298296 675392 298308
rect 675168 298268 675392 298296
rect 675168 298256 675174 298268
rect 675386 298256 675392 298268
rect 675444 298256 675450 298308
rect 655054 298120 655060 298172
rect 655112 298160 655118 298172
rect 675386 298160 675392 298172
rect 655112 298132 675392 298160
rect 655112 298120 655118 298132
rect 675386 298120 675392 298132
rect 675444 298120 675450 298172
rect 674650 295400 674656 295452
rect 674708 295440 674714 295452
rect 675294 295440 675300 295452
rect 674708 295412 675300 295440
rect 674708 295400 674714 295412
rect 675294 295400 675300 295412
rect 675352 295400 675358 295452
rect 42334 295332 42340 295384
rect 42392 295372 42398 295384
rect 58526 295372 58532 295384
rect 42392 295344 58532 295372
rect 42392 295332 42398 295344
rect 58526 295332 58532 295344
rect 58584 295332 58590 295384
rect 674558 295196 674564 295248
rect 674616 295236 674622 295248
rect 675386 295236 675392 295248
rect 674616 295208 675392 295236
rect 674616 295196 674622 295208
rect 675386 295196 675392 295208
rect 675444 295196 675450 295248
rect 674466 294108 674472 294160
rect 674524 294148 674530 294160
rect 675294 294148 675300 294160
rect 674524 294120 675300 294148
rect 674524 294108 674530 294120
rect 675294 294108 675300 294120
rect 675352 294108 675358 294160
rect 674558 293904 674564 293956
rect 674616 293944 674622 293956
rect 675110 293944 675116 293956
rect 674616 293916 675116 293944
rect 674616 293904 674622 293916
rect 675110 293904 675116 293916
rect 675168 293904 675174 293956
rect 43346 292544 43352 292596
rect 43404 292584 43410 292596
rect 58342 292584 58348 292596
rect 43404 292556 58348 292584
rect 43404 292544 43410 292556
rect 58342 292544 58348 292556
rect 58400 292544 58406 292596
rect 41782 291864 41788 291916
rect 41840 291904 41846 291916
rect 43438 291904 43444 291916
rect 41840 291876 43444 291904
rect 41840 291864 41846 291876
rect 43438 291864 43444 291876
rect 43496 291864 43502 291916
rect 674834 291252 674840 291304
rect 674892 291252 674898 291304
rect 674852 291088 674880 291252
rect 675110 291088 675116 291100
rect 674852 291060 675116 291088
rect 675110 291048 675116 291060
rect 675168 291048 675174 291100
rect 674282 290436 674288 290488
rect 674340 290476 674346 290488
rect 675110 290476 675116 290488
rect 674340 290448 675116 290476
rect 674340 290436 674346 290448
rect 675110 290436 675116 290448
rect 675168 290436 675174 290488
rect 41782 289824 41788 289876
rect 41840 289864 41846 289876
rect 42702 289864 42708 289876
rect 41840 289836 42708 289864
rect 41840 289824 41846 289836
rect 42702 289824 42708 289836
rect 42760 289824 42766 289876
rect 54018 289756 54024 289808
rect 54076 289796 54082 289808
rect 58526 289796 58532 289808
rect 54076 289768 58532 289796
rect 54076 289756 54082 289768
rect 58526 289756 58532 289768
rect 58584 289756 58590 289808
rect 654134 289076 654140 289128
rect 654192 289116 654198 289128
rect 667014 289116 667020 289128
rect 654192 289088 667020 289116
rect 654192 289076 654198 289088
rect 667014 289076 667020 289088
rect 667072 289076 667078 289128
rect 30006 288844 30012 288856
rect 24826 288816 30012 288844
rect 24826 288436 24854 288816
rect 30006 288804 30012 288816
rect 30064 288804 30070 288856
rect 673546 288600 673552 288652
rect 673604 288640 673610 288652
rect 675386 288640 675392 288652
rect 673604 288612 675392 288640
rect 673604 288600 673610 288612
rect 675386 288600 675392 288612
rect 675444 288600 675450 288652
rect 42242 288436 42248 288448
rect 24826 288408 42248 288436
rect 42242 288396 42248 288408
rect 42300 288396 42306 288448
rect 673822 287376 673828 287428
rect 673880 287416 673886 287428
rect 675110 287416 675116 287428
rect 673880 287388 675116 287416
rect 673880 287376 673886 287388
rect 675110 287376 675116 287388
rect 675168 287376 675174 287428
rect 656802 287240 656808 287292
rect 656860 287280 656866 287292
rect 666830 287280 666836 287292
rect 656860 287252 666836 287280
rect 656860 287240 656866 287252
rect 666830 287240 666836 287252
rect 666888 287240 666894 287292
rect 56502 287104 56508 287156
rect 56560 287144 56566 287156
rect 57974 287144 57980 287156
rect 56560 287116 57980 287144
rect 56560 287104 56566 287116
rect 57974 287104 57980 287116
rect 58032 287104 58038 287156
rect 46106 287036 46112 287088
rect 46164 287076 46170 287088
rect 58526 287076 58532 287088
rect 46164 287048 58532 287076
rect 46164 287036 46170 287048
rect 58526 287036 58532 287048
rect 58584 287036 58590 287088
rect 654134 287036 654140 287088
rect 654192 287076 654198 287088
rect 670234 287076 670240 287088
rect 654192 287048 670240 287076
rect 654192 287036 654198 287048
rect 670234 287036 670240 287048
rect 670292 287036 670298 287088
rect 673454 286764 673460 286816
rect 673512 286804 673518 286816
rect 675110 286804 675116 286816
rect 673512 286776 675116 286804
rect 673512 286764 673518 286776
rect 675110 286764 675116 286776
rect 675168 286764 675174 286816
rect 673638 286696 673644 286748
rect 673696 286736 673702 286748
rect 675202 286736 675208 286748
rect 673696 286708 675208 286736
rect 673696 286696 673702 286708
rect 675202 286696 675208 286708
rect 675260 286696 675266 286748
rect 673454 286628 673460 286680
rect 673512 286668 673518 286680
rect 674558 286668 674564 286680
rect 673512 286640 674564 286668
rect 673512 286628 673518 286640
rect 674558 286628 674564 286640
rect 674616 286628 674622 286680
rect 673730 286560 673736 286612
rect 673788 286600 673794 286612
rect 675386 286600 675392 286612
rect 673788 286572 675392 286600
rect 673788 286560 673794 286572
rect 675386 286560 675392 286572
rect 675444 286560 675450 286612
rect 43070 285608 43076 285660
rect 43128 285648 43134 285660
rect 43714 285648 43720 285660
rect 43128 285620 43720 285648
rect 43128 285608 43134 285620
rect 43714 285608 43720 285620
rect 43772 285608 43778 285660
rect 42426 285472 42432 285524
rect 42484 285512 42490 285524
rect 43070 285512 43076 285524
rect 42484 285484 43076 285512
rect 42484 285472 42490 285484
rect 43070 285472 43076 285484
rect 43128 285472 43134 285524
rect 53926 285132 53932 285184
rect 53984 285172 53990 285184
rect 57974 285172 57980 285184
rect 53984 285144 57980 285172
rect 53984 285132 53990 285144
rect 57974 285132 57980 285144
rect 58032 285132 58038 285184
rect 655238 284928 655244 284980
rect 655296 284968 655302 284980
rect 670326 284968 670332 284980
rect 655296 284940 670332 284968
rect 655296 284928 655302 284940
rect 670326 284928 670332 284940
rect 670384 284928 670390 284980
rect 654502 284656 654508 284708
rect 654560 284696 654566 284708
rect 666738 284696 666744 284708
rect 654560 284668 666744 284696
rect 654560 284656 654566 284668
rect 666738 284656 666744 284668
rect 666796 284656 666802 284708
rect 51074 284316 51080 284368
rect 51132 284356 51138 284368
rect 58526 284356 58532 284368
rect 51132 284328 58532 284356
rect 51132 284316 51138 284328
rect 58526 284316 58532 284328
rect 58584 284316 58590 284368
rect 43990 284248 43996 284300
rect 44048 284288 44054 284300
rect 44266 284288 44272 284300
rect 44048 284260 44272 284288
rect 44048 284248 44054 284260
rect 44266 284248 44272 284260
rect 44324 284248 44330 284300
rect 41874 283772 41880 283824
rect 41932 283772 41938 283824
rect 41892 283620 41920 283772
rect 41874 283568 41880 283620
rect 41932 283568 41938 283620
rect 654226 283160 654232 283212
rect 654284 283200 654290 283212
rect 669958 283200 669964 283212
rect 654284 283172 669964 283200
rect 654284 283160 654290 283172
rect 669958 283160 669964 283172
rect 670016 283160 670022 283212
rect 673454 282820 673460 282872
rect 673512 282860 673518 282872
rect 675110 282860 675116 282872
rect 673512 282832 675116 282860
rect 673512 282820 673518 282832
rect 675110 282820 675116 282832
rect 675168 282820 675174 282872
rect 42150 281732 42156 281784
rect 42208 281772 42214 281784
rect 43622 281772 43628 281784
rect 42208 281744 43628 281772
rect 42208 281732 42214 281744
rect 43622 281732 43628 281744
rect 43680 281732 43686 281784
rect 43622 281596 43628 281648
rect 43680 281636 43686 281648
rect 44266 281636 44272 281648
rect 43680 281608 44272 281636
rect 43680 281596 43686 281608
rect 44266 281596 44272 281608
rect 44324 281596 44330 281648
rect 48498 281528 48504 281580
rect 48556 281568 48562 281580
rect 57974 281568 57980 281580
rect 48556 281540 57980 281568
rect 48556 281528 48562 281540
rect 57974 281528 57980 281540
rect 58032 281528 58038 281580
rect 655238 281528 655244 281580
rect 655296 281568 655302 281580
rect 670050 281568 670056 281580
rect 655296 281540 670056 281568
rect 655296 281528 655302 281540
rect 670050 281528 670056 281540
rect 670108 281528 670114 281580
rect 42150 281052 42156 281104
rect 42208 281092 42214 281104
rect 42334 281092 42340 281104
rect 42208 281064 42340 281092
rect 42208 281052 42214 281064
rect 42334 281052 42340 281064
rect 42392 281052 42398 281104
rect 42334 280440 42340 280492
rect 42392 280480 42398 280492
rect 43438 280480 43444 280492
rect 42392 280452 43444 280480
rect 42392 280440 42398 280452
rect 43438 280440 43444 280452
rect 43496 280440 43502 280492
rect 654134 280372 654140 280424
rect 654192 280412 654198 280424
rect 670142 280412 670148 280424
rect 654192 280384 670148 280412
rect 654192 280372 654198 280384
rect 670142 280372 670148 280384
rect 670200 280372 670206 280424
rect 42150 279828 42156 279880
rect 42208 279868 42214 279880
rect 43162 279868 43168 279880
rect 42208 279840 43168 279868
rect 42208 279828 42214 279840
rect 43162 279828 43168 279840
rect 43220 279828 43226 279880
rect 42150 279216 42156 279268
rect 42208 279256 42214 279268
rect 43346 279256 43352 279268
rect 42208 279228 43352 279256
rect 42208 279216 42214 279228
rect 43346 279216 43352 279228
rect 43404 279216 43410 279268
rect 654870 278740 654876 278792
rect 654928 278780 654934 278792
rect 666646 278780 666652 278792
rect 654928 278752 666652 278780
rect 654928 278740 654934 278752
rect 666646 278740 666652 278752
rect 666704 278740 666710 278792
rect 42058 278604 42064 278656
rect 42116 278644 42122 278656
rect 42702 278644 42708 278656
rect 42116 278616 42708 278644
rect 42116 278604 42122 278616
rect 42702 278604 42708 278616
rect 42760 278604 42766 278656
rect 42702 278468 42708 278520
rect 42760 278508 42766 278520
rect 43898 278508 43904 278520
rect 42760 278480 43904 278508
rect 42760 278468 42766 278480
rect 43898 278468 43904 278480
rect 43956 278468 43962 278520
rect 671614 278372 671620 278384
rect 671606 278344 671620 278372
rect 671614 278332 671620 278344
rect 671672 278372 671678 278384
rect 678974 278372 678980 278384
rect 671672 278344 678980 278372
rect 671672 278332 671678 278344
rect 678974 278332 678980 278344
rect 679032 278332 679038 278384
rect 671706 278304 671712 278316
rect 671694 278276 671712 278304
rect 671706 278264 671712 278276
rect 671764 278304 671770 278316
rect 679066 278304 679072 278316
rect 671764 278276 679072 278304
rect 671764 278264 671770 278276
rect 679066 278264 679072 278276
rect 679124 278264 679130 278316
rect 671798 278100 671804 278112
rect 671792 278072 671804 278100
rect 671798 278060 671804 278072
rect 671856 278100 671862 278112
rect 679158 278100 679164 278112
rect 671856 278072 679164 278100
rect 671856 278060 671862 278072
rect 679158 278060 679164 278072
rect 679216 278060 679222 278112
rect 48314 277584 48320 277636
rect 48372 277624 48378 277636
rect 648614 277624 648620 277636
rect 48372 277596 648620 277624
rect 48372 277584 48378 277596
rect 648614 277584 648620 277596
rect 648672 277584 648678 277636
rect 48406 277516 48412 277568
rect 48464 277556 48470 277568
rect 654134 277556 654140 277568
rect 48464 277528 654140 277556
rect 48464 277516 48470 277528
rect 654134 277516 654140 277528
rect 654192 277516 654198 277568
rect 48222 277380 48228 277432
rect 48280 277420 48286 277432
rect 666554 277420 666560 277432
rect 48280 277392 666560 277420
rect 48280 277380 48286 277392
rect 666554 277380 666560 277392
rect 666612 277380 666618 277432
rect 42334 276768 42340 276820
rect 42392 276808 42398 276820
rect 43806 276808 43812 276820
rect 42392 276780 43812 276808
rect 42392 276768 42398 276780
rect 43806 276768 43812 276780
rect 43864 276768 43870 276820
rect 42242 276700 42248 276752
rect 42300 276740 42306 276752
rect 43070 276740 43076 276752
rect 42300 276712 43076 276740
rect 42300 276700 42306 276712
rect 43070 276700 43076 276712
rect 43128 276700 43134 276752
rect 42058 276564 42064 276616
rect 42116 276604 42122 276616
rect 43530 276604 43536 276616
rect 42116 276576 43536 276604
rect 42116 276564 42122 276576
rect 43530 276564 43536 276576
rect 43588 276564 43594 276616
rect 387242 276020 387248 276072
rect 387300 276060 387306 276072
rect 405090 276060 405096 276072
rect 387300 276032 405096 276060
rect 387300 276020 387306 276032
rect 405090 276020 405096 276032
rect 405148 276020 405154 276072
rect 347774 275952 347780 276004
rect 347832 275992 347838 276004
rect 478322 275992 478328 276004
rect 347832 275964 478328 275992
rect 347832 275952 347838 275964
rect 478322 275952 478328 275964
rect 478380 275952 478386 276004
rect 350166 275884 350172 275936
rect 350224 275924 350230 275936
rect 485498 275924 485504 275936
rect 350224 275896 485504 275924
rect 350224 275884 350230 275896
rect 485498 275884 485504 275896
rect 485556 275884 485562 275936
rect 353202 275816 353208 275868
rect 353260 275856 353266 275868
rect 492582 275856 492588 275868
rect 353260 275828 492588 275856
rect 353260 275816 353266 275828
rect 492582 275816 492588 275828
rect 492640 275816 492646 275868
rect 355778 275748 355784 275800
rect 355836 275788 355842 275800
rect 499666 275788 499672 275800
rect 355836 275760 499672 275788
rect 355836 275748 355842 275760
rect 499666 275748 499672 275760
rect 499724 275748 499730 275800
rect 358538 275680 358544 275732
rect 358596 275720 358602 275732
rect 506750 275720 506756 275732
rect 358596 275692 506756 275720
rect 358596 275680 358602 275692
rect 506750 275680 506756 275692
rect 506808 275680 506814 275732
rect 361482 275612 361488 275664
rect 361540 275652 361546 275664
rect 513834 275652 513840 275664
rect 361540 275624 513840 275652
rect 361540 275612 361546 275624
rect 513834 275612 513840 275624
rect 513892 275612 513898 275664
rect 42426 275544 42432 275596
rect 42484 275584 42490 275596
rect 42702 275584 42708 275596
rect 42484 275556 42708 275584
rect 42484 275544 42490 275556
rect 42702 275544 42708 275556
rect 42760 275544 42766 275596
rect 363966 275544 363972 275596
rect 364024 275584 364030 275596
rect 520918 275584 520924 275596
rect 364024 275556 520924 275584
rect 364024 275544 364030 275556
rect 520918 275544 520924 275556
rect 520976 275544 520982 275596
rect 366450 275476 366456 275528
rect 366508 275516 366514 275528
rect 528002 275516 528008 275528
rect 366508 275488 528008 275516
rect 366508 275476 366514 275488
rect 528002 275476 528008 275488
rect 528060 275476 528066 275528
rect 369118 275408 369124 275460
rect 369176 275448 369182 275460
rect 535086 275448 535092 275460
rect 369176 275420 535092 275448
rect 369176 275408 369182 275420
rect 535086 275408 535092 275420
rect 535144 275408 535150 275460
rect 371786 275340 371792 275392
rect 371844 275380 371850 275392
rect 542170 275380 542176 275392
rect 371844 275352 542176 275380
rect 371844 275340 371850 275352
rect 542170 275340 542176 275352
rect 542228 275340 542234 275392
rect 375282 275272 375288 275324
rect 375340 275312 375346 275324
rect 550450 275312 550456 275324
rect 375340 275284 550456 275312
rect 375340 275272 375346 275284
rect 550450 275272 550456 275284
rect 550508 275272 550514 275324
rect 377950 275204 377956 275256
rect 378008 275244 378014 275256
rect 557534 275244 557540 275256
rect 378008 275216 557540 275244
rect 378008 275204 378014 275216
rect 557534 275204 557540 275216
rect 557592 275204 557598 275256
rect 380342 275136 380348 275188
rect 380400 275176 380406 275188
rect 564618 275176 564624 275188
rect 380400 275148 564624 275176
rect 380400 275136 380406 275148
rect 564618 275136 564624 275148
rect 564676 275136 564682 275188
rect 382918 275068 382924 275120
rect 382976 275108 382982 275120
rect 571702 275108 571708 275120
rect 382976 275080 571708 275108
rect 382976 275068 382982 275080
rect 571702 275068 571708 275080
rect 571760 275068 571766 275120
rect 385586 275000 385592 275052
rect 385644 275040 385650 275052
rect 578878 275040 578884 275052
rect 385644 275012 578884 275040
rect 385644 275000 385650 275012
rect 578878 275000 578884 275012
rect 578936 275000 578942 275052
rect 401594 274932 401600 274984
rect 401652 274972 401658 274984
rect 585962 274972 585968 274984
rect 401652 274944 585968 274972
rect 401652 274932 401658 274944
rect 585962 274932 585968 274944
rect 586020 274932 586026 274984
rect 320266 274864 320272 274916
rect 320324 274904 320330 274916
rect 387242 274904 387248 274916
rect 320324 274876 387248 274904
rect 320324 274864 320330 274876
rect 387242 274864 387248 274876
rect 387300 274864 387306 274916
rect 405366 274864 405372 274916
rect 405424 274904 405430 274916
rect 627270 274904 627276 274916
rect 405424 274876 627276 274904
rect 405424 274864 405430 274876
rect 627270 274864 627276 274876
rect 627328 274864 627334 274916
rect 361546 274808 391934 274836
rect 319898 274728 319904 274780
rect 319956 274768 319962 274780
rect 361546 274768 361574 274808
rect 319956 274740 361574 274768
rect 391906 274768 391934 274808
rect 401686 274796 401692 274848
rect 401744 274836 401750 274848
rect 593046 274836 593052 274848
rect 401744 274808 593052 274836
rect 401744 274796 401750 274808
rect 593046 274796 593052 274808
rect 593104 274796 593110 274848
rect 403894 274768 403900 274780
rect 391906 274740 403900 274768
rect 319956 274728 319962 274740
rect 403894 274728 403900 274740
rect 403952 274728 403958 274780
rect 404262 274728 404268 274780
rect 404320 274768 404326 274780
rect 628466 274768 628472 274780
rect 404320 274740 628472 274768
rect 404320 274728 404326 274740
rect 628466 274728 628472 274740
rect 628524 274728 628530 274780
rect 321002 274660 321008 274712
rect 321060 274700 321066 274712
rect 407482 274700 407488 274712
rect 321060 274672 407488 274700
rect 321060 274660 321066 274672
rect 407482 274660 407488 274672
rect 407540 274660 407546 274712
rect 409230 274660 409236 274712
rect 409288 274700 409294 274712
rect 409288 274672 419534 274700
rect 409288 274660 409294 274672
rect 322750 274592 322756 274644
rect 322808 274632 322814 274644
rect 410978 274632 410984 274644
rect 322808 274604 410984 274632
rect 322808 274592 322814 274604
rect 410978 274592 410984 274604
rect 411036 274592 411042 274644
rect 419506 274632 419534 274672
rect 429102 274660 429108 274712
rect 429160 274700 429166 274712
rect 634354 274700 634360 274712
rect 429160 274672 634360 274700
rect 429160 274660 429166 274672
rect 634354 274660 634360 274672
rect 634412 274660 634418 274712
rect 641438 274632 641444 274644
rect 419506 274604 641444 274632
rect 641438 274592 641444 274604
rect 641496 274592 641502 274644
rect 343726 274524 343732 274576
rect 343784 274564 343790 274576
rect 467742 274564 467748 274576
rect 343784 274536 467748 274564
rect 343784 274524 343790 274536
rect 467742 274524 467748 274536
rect 467800 274524 467806 274576
rect 345106 274456 345112 274508
rect 345164 274496 345170 274508
rect 471238 274496 471244 274508
rect 345164 274468 471244 274496
rect 345164 274456 345170 274468
rect 471238 274456 471244 274468
rect 471296 274456 471302 274508
rect 342530 274388 342536 274440
rect 342588 274428 342594 274440
rect 464154 274428 464160 274440
rect 342588 274400 464160 274428
rect 342588 274388 342594 274400
rect 464154 274388 464160 274400
rect 464212 274388 464218 274440
rect 339770 274320 339776 274372
rect 339828 274360 339834 274372
rect 457070 274360 457076 274372
rect 339828 274332 457076 274360
rect 339828 274320 339834 274332
rect 457070 274320 457076 274332
rect 457128 274320 457134 274372
rect 42150 274252 42156 274304
rect 42208 274292 42214 274304
rect 44082 274292 44088 274304
rect 42208 274264 44088 274292
rect 42208 274252 42214 274264
rect 44082 274252 44088 274264
rect 44140 274252 44146 274304
rect 337102 274252 337108 274304
rect 337160 274292 337166 274304
rect 449986 274292 449992 274304
rect 337160 274264 449992 274292
rect 337160 274252 337166 274264
rect 449986 274252 449992 274264
rect 450044 274252 450050 274304
rect 335722 274184 335728 274236
rect 335780 274224 335786 274236
rect 446490 274224 446496 274236
rect 335780 274196 446496 274224
rect 335780 274184 335786 274196
rect 446490 274184 446496 274196
rect 446548 274184 446554 274236
rect 334342 274116 334348 274168
rect 334400 274156 334406 274168
rect 442902 274156 442908 274168
rect 334400 274128 442908 274156
rect 334400 274116 334406 274128
rect 442902 274116 442908 274128
rect 442960 274116 442966 274168
rect 333422 274048 333428 274100
rect 333480 274088 333486 274100
rect 439314 274088 439320 274100
rect 333480 274060 439320 274088
rect 333480 274048 333486 274060
rect 439314 274048 439320 274060
rect 439372 274048 439378 274100
rect 331674 273980 331680 274032
rect 331732 274020 331738 274032
rect 435818 274020 435824 274032
rect 331732 273992 435824 274020
rect 331732 273980 331738 273992
rect 435818 273980 435824 273992
rect 435876 273980 435882 274032
rect 330754 273912 330760 273964
rect 330812 273952 330818 273964
rect 432230 273952 432236 273964
rect 330812 273924 432236 273952
rect 330812 273912 330818 273924
rect 432230 273912 432236 273924
rect 432288 273912 432294 273964
rect 329006 273844 329012 273896
rect 329064 273884 329070 273896
rect 428734 273884 428740 273896
rect 329064 273856 428740 273884
rect 329064 273844 329070 273856
rect 428734 273844 428740 273856
rect 428792 273844 428798 273896
rect 327718 273776 327724 273828
rect 327776 273816 327782 273828
rect 425146 273816 425152 273828
rect 327776 273788 425152 273816
rect 327776 273776 327782 273788
rect 425146 273776 425152 273788
rect 425204 273776 425210 273828
rect 325510 273708 325516 273760
rect 325568 273748 325574 273760
rect 418062 273748 418068 273760
rect 325568 273720 418068 273748
rect 325568 273708 325574 273720
rect 418062 273708 418068 273720
rect 418120 273708 418126 273760
rect 326338 273640 326344 273692
rect 326396 273680 326402 273692
rect 421650 273680 421656 273692
rect 326396 273652 421656 273680
rect 326396 273640 326402 273652
rect 421650 273640 421656 273652
rect 421708 273640 421714 273692
rect 323670 273572 323676 273624
rect 323728 273612 323734 273624
rect 414566 273612 414572 273624
rect 323728 273584 414572 273612
rect 323728 273572 323734 273584
rect 414566 273572 414572 273584
rect 414624 273572 414630 273624
rect 42058 273504 42064 273556
rect 42116 273544 42122 273556
rect 43622 273544 43628 273556
rect 42116 273516 43628 273544
rect 42116 273504 42122 273516
rect 43622 273504 43628 273516
rect 43680 273504 43686 273556
rect 388254 273504 388260 273556
rect 388312 273544 388318 273556
rect 401594 273544 401600 273556
rect 388312 273516 401600 273544
rect 388312 273504 388318 273516
rect 401594 273504 401600 273516
rect 401652 273504 401658 273556
rect 429102 273544 429108 273556
rect 419506 273516 429108 273544
rect 406562 273436 406568 273488
rect 406620 273476 406626 273488
rect 419506 273476 419534 273516
rect 429102 273504 429108 273516
rect 429160 273504 429166 273556
rect 406620 273448 419534 273476
rect 406620 273436 406626 273448
rect 391014 273232 391020 273284
rect 391072 273272 391078 273284
rect 401686 273272 401692 273284
rect 391072 273244 401692 273272
rect 391072 273232 391078 273244
rect 401686 273232 401692 273244
rect 401744 273232 401750 273284
rect 154482 273164 154488 273216
rect 154540 273204 154546 273216
rect 225322 273204 225328 273216
rect 154540 273176 225328 273204
rect 154540 273164 154546 273176
rect 225322 273164 225328 273176
rect 225380 273164 225386 273216
rect 263226 273164 263232 273216
rect 263284 273204 263290 273216
rect 266722 273204 266728 273216
rect 263284 273176 266728 273204
rect 263284 273164 263290 273176
rect 266722 273164 266728 273176
rect 266780 273164 266786 273216
rect 291194 273164 291200 273216
rect 291252 273204 291258 273216
rect 328270 273204 328276 273216
rect 291252 273176 328276 273204
rect 291252 273164 291258 273176
rect 328270 273164 328276 273176
rect 328328 273164 328334 273216
rect 345474 273164 345480 273216
rect 345532 273204 345538 273216
rect 472434 273204 472440 273216
rect 345532 273176 472440 273204
rect 345532 273164 345538 273176
rect 472434 273164 472440 273176
rect 472492 273164 472498 273216
rect 472526 273164 472532 273216
rect 472584 273204 472590 273216
rect 610710 273204 610716 273216
rect 472584 273176 610716 273204
rect 472584 273164 472590 273176
rect 610710 273164 610716 273176
rect 610768 273164 610774 273216
rect 156874 273096 156880 273148
rect 156932 273136 156938 273148
rect 208302 273136 208308 273148
rect 156932 273108 208308 273136
rect 156932 273096 156938 273108
rect 208302 273096 208308 273108
rect 208360 273096 208366 273148
rect 260926 273096 260932 273148
rect 260984 273136 260990 273148
rect 265802 273136 265808 273148
rect 260984 273108 265808 273136
rect 260984 273096 260990 273108
rect 265802 273096 265808 273108
rect 265860 273096 265866 273148
rect 292114 273096 292120 273148
rect 292172 273136 292178 273148
rect 330570 273136 330576 273148
rect 292172 273108 330576 273136
rect 292172 273096 292178 273108
rect 330570 273096 330576 273108
rect 330628 273096 330634 273148
rect 356238 273096 356244 273148
rect 356296 273136 356302 273148
rect 500862 273136 500868 273148
rect 356296 273108 500868 273136
rect 356296 273096 356302 273108
rect 500862 273096 500868 273108
rect 500920 273096 500926 273148
rect 149790 273028 149796 273080
rect 149848 273068 149854 273080
rect 224402 273068 224408 273080
rect 149848 273040 224408 273068
rect 149848 273028 149854 273040
rect 224402 273028 224408 273040
rect 224460 273028 224466 273080
rect 243170 273028 243176 273080
rect 243228 273068 243234 273080
rect 259178 273068 259184 273080
rect 243228 273040 259184 273068
rect 243228 273028 243234 273040
rect 259178 273028 259184 273040
rect 259236 273028 259242 273080
rect 259730 273028 259736 273080
rect 259788 273068 259794 273080
rect 265342 273068 265348 273080
rect 259788 273040 265348 273068
rect 259788 273028 259794 273040
rect 265342 273028 265348 273040
rect 265400 273028 265406 273080
rect 293862 273028 293868 273080
rect 293920 273068 293926 273080
rect 335354 273068 335360 273080
rect 293920 273040 335360 273068
rect 293920 273028 293926 273040
rect 335354 273028 335360 273040
rect 335412 273028 335418 273080
rect 342806 273028 342812 273080
rect 342864 273068 342870 273080
rect 465350 273068 465356 273080
rect 342864 273040 465356 273068
rect 342864 273028 342870 273040
rect 465350 273028 465356 273040
rect 465408 273028 465414 273080
rect 467742 273028 467748 273080
rect 467800 273068 467806 273080
rect 617794 273068 617800 273080
rect 467800 273040 617800 273068
rect 467800 273028 467806 273040
rect 617794 273028 617800 273040
rect 617852 273028 617858 273080
rect 143902 272960 143908 273012
rect 143960 273000 143966 273012
rect 221274 273000 221280 273012
rect 143960 272972 221280 273000
rect 143960 272960 143966 272972
rect 221274 272960 221280 272972
rect 221332 272960 221338 273012
rect 241974 272960 241980 273012
rect 242032 273000 242038 273012
rect 258718 273000 258724 273012
rect 242032 272972 258724 273000
rect 242032 272960 242038 272972
rect 258718 272960 258724 272972
rect 258776 272960 258782 273012
rect 296070 272960 296076 273012
rect 296128 273000 296134 273012
rect 341242 273000 341248 273012
rect 296128 272972 341248 273000
rect 296128 272960 296134 272972
rect 341242 272960 341248 272972
rect 341300 272960 341306 273012
rect 347866 272960 347872 273012
rect 347924 273000 347930 273012
rect 351914 273000 351920 273012
rect 347924 272972 351920 273000
rect 347924 272960 347930 272972
rect 351914 272960 351920 272972
rect 351972 272960 351978 273012
rect 361574 272960 361580 273012
rect 361632 273000 361638 273012
rect 515030 273000 515036 273012
rect 361632 272972 515036 273000
rect 361632 272960 361638 272972
rect 515030 272960 515036 272972
rect 515088 272960 515094 273012
rect 148594 272892 148600 272944
rect 148652 272932 148658 272944
rect 223206 272932 223212 272944
rect 148652 272904 223212 272932
rect 148652 272892 148658 272904
rect 223206 272892 223212 272904
rect 223264 272892 223270 272944
rect 236086 272892 236092 272944
rect 236144 272932 236150 272944
rect 256418 272932 256424 272944
rect 236144 272904 256424 272932
rect 236144 272892 236150 272904
rect 256418 272892 256424 272904
rect 256476 272892 256482 272944
rect 294874 272892 294880 272944
rect 294932 272932 294938 272944
rect 337746 272932 337752 272944
rect 294932 272904 337752 272932
rect 294932 272892 294938 272904
rect 337746 272892 337752 272904
rect 337804 272892 337810 272944
rect 350074 272892 350080 272944
rect 350132 272932 350138 272944
rect 484302 272932 484308 272944
rect 350132 272904 484308 272932
rect 350132 272892 350138 272904
rect 484302 272892 484308 272904
rect 484360 272892 484366 272944
rect 485038 272892 485044 272944
rect 485096 272932 485102 272944
rect 635550 272932 635556 272944
rect 485096 272904 635556 272932
rect 485096 272892 485102 272904
rect 635550 272892 635556 272904
rect 635608 272892 635614 272944
rect 145098 272824 145104 272876
rect 145156 272864 145162 272876
rect 222194 272864 222200 272876
rect 145156 272836 222200 272864
rect 145156 272824 145162 272836
rect 222194 272824 222200 272836
rect 222252 272824 222258 272876
rect 234890 272824 234896 272876
rect 234948 272864 234954 272876
rect 256050 272864 256056 272876
rect 234948 272836 256056 272864
rect 234948 272824 234954 272836
rect 256050 272824 256056 272836
rect 256108 272824 256114 272876
rect 301406 272824 301412 272876
rect 301464 272864 301470 272876
rect 355410 272864 355416 272876
rect 301464 272836 355416 272864
rect 301464 272824 301470 272836
rect 355410 272824 355416 272836
rect 355468 272824 355474 272876
rect 372798 272824 372804 272876
rect 372856 272864 372862 272876
rect 381446 272864 381452 272876
rect 372856 272836 381452 272864
rect 372856 272824 372862 272836
rect 381446 272824 381452 272836
rect 381504 272824 381510 272876
rect 383654 272824 383660 272876
rect 383712 272864 383718 272876
rect 388530 272864 388536 272876
rect 383712 272836 388536 272864
rect 383712 272824 383718 272836
rect 388530 272824 388536 272836
rect 388588 272824 388594 272876
rect 390462 272824 390468 272876
rect 390520 272864 390526 272876
rect 526806 272864 526812 272876
rect 390520 272836 526812 272864
rect 390520 272824 390526 272836
rect 526806 272824 526812 272836
rect 526864 272824 526870 272876
rect 146202 272756 146208 272808
rect 146260 272796 146266 272808
rect 223022 272796 223028 272808
rect 146260 272768 223028 272796
rect 146260 272756 146266 272768
rect 223022 272756 223028 272768
rect 223080 272756 223086 272808
rect 238478 272756 238484 272808
rect 238536 272796 238542 272808
rect 257430 272796 257436 272808
rect 238536 272768 257436 272796
rect 238536 272756 238542 272768
rect 257430 272756 257436 272768
rect 257488 272756 257494 272808
rect 301866 272756 301872 272808
rect 301924 272796 301930 272808
rect 356606 272796 356612 272808
rect 301924 272768 356612 272796
rect 301924 272756 301930 272768
rect 356606 272756 356612 272768
rect 356664 272756 356670 272808
rect 363874 272756 363880 272808
rect 363932 272796 363938 272808
rect 519722 272796 519728 272808
rect 363932 272768 519728 272796
rect 363932 272756 363938 272768
rect 519722 272756 519728 272768
rect 519780 272756 519786 272808
rect 139118 272688 139124 272740
rect 139176 272728 139182 272740
rect 220354 272728 220360 272740
rect 139176 272700 220360 272728
rect 139176 272688 139182 272700
rect 220354 272688 220360 272700
rect 220412 272688 220418 272740
rect 239582 272688 239588 272740
rect 239640 272728 239646 272740
rect 257798 272728 257804 272740
rect 239640 272700 257804 272728
rect 239640 272688 239646 272700
rect 257798 272688 257804 272700
rect 257856 272688 257862 272740
rect 295242 272688 295248 272740
rect 295300 272728 295306 272740
rect 338850 272728 338856 272740
rect 295300 272700 338856 272728
rect 295300 272688 295306 272700
rect 338850 272688 338856 272700
rect 338908 272688 338914 272740
rect 339402 272688 339408 272740
rect 339460 272728 339466 272740
rect 455874 272728 455880 272740
rect 339460 272700 455880 272728
rect 339460 272688 339466 272700
rect 455874 272688 455880 272700
rect 455932 272688 455938 272740
rect 455966 272688 455972 272740
rect 456024 272728 456030 272740
rect 624970 272728 624976 272740
rect 456024 272700 624976 272728
rect 456024 272688 456030 272700
rect 624970 272688 624976 272700
rect 625028 272688 625034 272740
rect 137922 272620 137928 272672
rect 137980 272660 137986 272672
rect 219434 272660 219440 272672
rect 137980 272632 219440 272660
rect 137980 272620 137986 272632
rect 219434 272620 219440 272632
rect 219492 272620 219498 272672
rect 232498 272620 232504 272672
rect 232556 272660 232562 272672
rect 255130 272660 255136 272672
rect 232556 272632 255136 272660
rect 232556 272620 232562 272632
rect 255130 272620 255136 272632
rect 255188 272620 255194 272672
rect 304074 272620 304080 272672
rect 304132 272660 304138 272672
rect 362494 272660 362500 272672
rect 304132 272632 362500 272660
rect 304132 272620 304138 272632
rect 362494 272620 362500 272632
rect 362552 272620 362558 272672
rect 375374 272620 375380 272672
rect 375432 272660 375438 272672
rect 551646 272660 551652 272672
rect 375432 272632 551652 272660
rect 375432 272620 375438 272632
rect 551646 272620 551652 272632
rect 551704 272620 551710 272672
rect 136818 272552 136824 272604
rect 136876 272592 136882 272604
rect 218606 272592 218612 272604
rect 136876 272564 218612 272592
rect 136876 272552 136882 272564
rect 218606 272552 218612 272564
rect 218664 272552 218670 272604
rect 237282 272552 237288 272604
rect 237340 272592 237346 272604
rect 257246 272592 257252 272604
rect 237340 272564 257252 272592
rect 237340 272552 237346 272564
rect 257246 272552 257252 272564
rect 257304 272552 257310 272604
rect 304534 272552 304540 272604
rect 304592 272592 304598 272604
rect 363690 272592 363696 272604
rect 304592 272564 363696 272592
rect 304592 272552 304598 272564
rect 363690 272552 363696 272564
rect 363748 272552 363754 272604
rect 378042 272552 378048 272604
rect 378100 272592 378106 272604
rect 558730 272592 558736 272604
rect 378100 272564 558736 272592
rect 378100 272552 378106 272564
rect 558730 272552 558736 272564
rect 558788 272552 558794 272604
rect 130838 272484 130844 272536
rect 130896 272524 130902 272536
rect 216858 272524 216864 272536
rect 130896 272496 216864 272524
rect 130896 272484 130902 272496
rect 216858 272484 216864 272496
rect 216916 272484 216922 272536
rect 233694 272484 233700 272536
rect 233752 272524 233758 272536
rect 255590 272524 255596 272536
rect 233752 272496 255596 272524
rect 233752 272484 233758 272496
rect 255590 272484 255596 272496
rect 255648 272484 255654 272536
rect 288158 272484 288164 272536
rect 288216 272524 288222 272536
rect 319990 272524 319996 272536
rect 288216 272496 319996 272524
rect 288216 272484 288222 272496
rect 319990 272484 319996 272496
rect 320048 272484 320054 272536
rect 320082 272484 320088 272536
rect 320140 272524 320146 272536
rect 377858 272524 377864 272536
rect 320140 272496 377864 272524
rect 320140 272484 320146 272496
rect 377858 272484 377864 272496
rect 377916 272484 377922 272536
rect 390480 272496 391244 272524
rect 132034 272416 132040 272468
rect 132092 272456 132098 272468
rect 217686 272456 217692 272468
rect 132092 272428 217692 272456
rect 132092 272416 132098 272428
rect 217686 272416 217692 272428
rect 217744 272416 217750 272468
rect 227806 272416 227812 272468
rect 227864 272456 227870 272468
rect 253382 272456 253388 272468
rect 227864 272428 253388 272456
rect 227864 272416 227870 272428
rect 253382 272416 253388 272428
rect 253440 272416 253446 272468
rect 293402 272416 293408 272468
rect 293460 272456 293466 272468
rect 334158 272456 334164 272468
rect 293460 272428 334164 272456
rect 293460 272416 293466 272428
rect 334158 272416 334164 272428
rect 334216 272416 334222 272468
rect 334250 272416 334256 272468
rect 334308 272456 334314 272468
rect 390480 272456 390508 272496
rect 334308 272428 390508 272456
rect 391216 272456 391244 272496
rect 391566 272484 391572 272536
rect 391624 272524 391630 272536
rect 572898 272524 572904 272536
rect 391624 272496 572904 272524
rect 391624 272484 391630 272496
rect 572898 272484 572904 272496
rect 572956 272484 572962 272536
rect 441706 272456 441712 272468
rect 391216 272428 441712 272456
rect 334308 272416 334314 272428
rect 441706 272416 441712 272428
rect 441764 272416 441770 272468
rect 441798 272416 441804 272468
rect 441856 272456 441862 272468
rect 632054 272456 632060 272468
rect 441856 272428 632060 272456
rect 441856 272416 441862 272428
rect 632054 272416 632060 272428
rect 632112 272416 632118 272468
rect 129642 272348 129648 272400
rect 129700 272388 129706 272400
rect 215662 272388 215668 272400
rect 129700 272360 215668 272388
rect 129700 272348 129706 272360
rect 215662 272348 215668 272360
rect 215720 272348 215726 272400
rect 231302 272348 231308 272400
rect 231360 272388 231366 272400
rect 254670 272388 254676 272400
rect 231360 272360 254676 272388
rect 231360 272348 231366 272360
rect 254670 272348 254676 272360
rect 254728 272348 254734 272400
rect 307202 272348 307208 272400
rect 307260 272388 307266 272400
rect 370774 272388 370780 272400
rect 307260 272360 370780 272388
rect 307260 272348 307266 272360
rect 370774 272348 370780 272360
rect 370832 272348 370838 272400
rect 372062 272348 372068 272400
rect 372120 272388 372126 272400
rect 390462 272388 390468 272400
rect 372120 272360 390468 272388
rect 372120 272348 372126 272360
rect 390462 272348 390468 272360
rect 390520 272348 390526 272400
rect 391198 272348 391204 272400
rect 391256 272388 391262 272400
rect 579982 272388 579988 272400
rect 391256 272360 579988 272388
rect 391256 272348 391262 272360
rect 579982 272348 579988 272360
rect 580040 272348 580046 272400
rect 124950 272280 124956 272332
rect 125008 272320 125014 272332
rect 215018 272320 215024 272332
rect 125008 272292 215024 272320
rect 125008 272280 125014 272292
rect 215018 272280 215024 272292
rect 215076 272280 215082 272332
rect 229002 272280 229008 272332
rect 229060 272320 229066 272332
rect 253750 272320 253756 272332
rect 229060 272292 253756 272320
rect 229060 272280 229066 272292
rect 253750 272280 253756 272292
rect 253808 272280 253814 272332
rect 287606 272280 287612 272332
rect 287664 272320 287670 272332
rect 318794 272320 318800 272332
rect 287664 272292 318800 272320
rect 287664 272280 287670 272292
rect 318794 272280 318800 272292
rect 318852 272280 318858 272332
rect 318886 272280 318892 272332
rect 318944 272320 318950 272332
rect 384942 272320 384948 272332
rect 318944 272292 384948 272320
rect 318944 272280 318950 272292
rect 384942 272280 384948 272292
rect 385000 272280 385006 272332
rect 390002 272280 390008 272332
rect 390060 272320 390066 272332
rect 390060 272292 391060 272320
rect 390060 272280 390066 272292
rect 123754 272212 123760 272264
rect 123812 272252 123818 272264
rect 214190 272252 214196 272264
rect 123812 272224 214196 272252
rect 123812 272212 123818 272224
rect 214190 272212 214196 272224
rect 214248 272212 214254 272264
rect 230198 272212 230204 272264
rect 230256 272252 230262 272264
rect 254210 272252 254216 272264
rect 230256 272224 254216 272252
rect 230256 272212 230262 272224
rect 254210 272212 254216 272224
rect 254268 272212 254274 272264
rect 288894 272212 288900 272264
rect 288952 272252 288958 272264
rect 321186 272252 321192 272264
rect 288952 272224 321192 272252
rect 288952 272212 288958 272224
rect 321186 272212 321192 272224
rect 321244 272212 321250 272264
rect 325326 272212 325332 272264
rect 325384 272252 325390 272264
rect 390922 272252 390928 272264
rect 325384 272224 390928 272252
rect 325384 272212 325390 272224
rect 390922 272212 390928 272224
rect 390980 272212 390986 272264
rect 391032 272252 391060 272292
rect 391106 272280 391112 272332
rect 391164 272320 391170 272332
rect 587066 272320 587072 272332
rect 391164 272292 587072 272320
rect 391164 272280 391170 272292
rect 587066 272280 587072 272292
rect 587124 272280 587130 272332
rect 590654 272252 590660 272264
rect 391032 272224 590660 272252
rect 590654 272212 590660 272224
rect 590712 272212 590718 272264
rect 104894 272144 104900 272196
rect 104952 272184 104958 272196
rect 206278 272184 206284 272196
rect 104952 272156 206284 272184
rect 104952 272144 104958 272156
rect 206278 272144 206284 272156
rect 206336 272144 206342 272196
rect 226610 272144 226616 272196
rect 226668 272184 226674 272196
rect 252922 272184 252928 272196
rect 226668 272156 252928 272184
rect 226668 272144 226674 272156
rect 252922 272144 252928 272156
rect 252980 272144 252986 272196
rect 286686 272144 286692 272196
rect 286744 272184 286750 272196
rect 315206 272184 315212 272196
rect 286744 272156 315212 272184
rect 286744 272144 286750 272156
rect 315206 272144 315212 272156
rect 315264 272144 315270 272196
rect 315298 272144 315304 272196
rect 315356 272184 315362 272196
rect 392118 272184 392124 272196
rect 315356 272156 392124 272184
rect 315356 272144 315362 272156
rect 392118 272144 392124 272156
rect 392176 272144 392182 272196
rect 394050 272144 394056 272196
rect 394108 272184 394114 272196
rect 601326 272184 601332 272196
rect 394108 272156 601332 272184
rect 394108 272144 394114 272156
rect 601326 272144 601332 272156
rect 601384 272144 601390 272196
rect 97810 272076 97816 272128
rect 97868 272116 97874 272128
rect 203886 272116 203892 272128
rect 97868 272088 203892 272116
rect 97868 272076 97874 272088
rect 203886 272076 203892 272088
rect 203944 272076 203950 272128
rect 205358 272076 205364 272128
rect 205416 272116 205422 272128
rect 244918 272116 244924 272128
rect 205416 272088 244924 272116
rect 205416 272076 205422 272088
rect 244918 272076 244924 272088
rect 244976 272076 244982 272128
rect 258258 272116 258264 272128
rect 245626 272088 258264 272116
rect 91830 272008 91836 272060
rect 91888 272048 91894 272060
rect 195974 272048 195980 272060
rect 91888 272020 195980 272048
rect 91888 272008 91894 272020
rect 195974 272008 195980 272020
rect 196032 272008 196038 272060
rect 201770 272008 201776 272060
rect 201828 272048 201834 272060
rect 240134 272048 240140 272060
rect 201828 272020 240140 272048
rect 201828 272008 201834 272020
rect 240134 272008 240140 272020
rect 240192 272008 240198 272060
rect 89530 271940 89536 271992
rect 89588 271980 89594 271992
rect 200758 271980 200764 271992
rect 89588 271952 200764 271980
rect 89588 271940 89594 271952
rect 200758 271940 200764 271952
rect 200816 271940 200822 271992
rect 208302 271940 208308 271992
rect 208360 271980 208366 271992
rect 227070 271980 227076 271992
rect 208360 271952 227076 271980
rect 208360 271940 208366 271952
rect 227070 271940 227076 271952
rect 227128 271940 227134 271992
rect 240778 271940 240784 271992
rect 240836 271980 240842 271992
rect 245626 271980 245654 272088
rect 258258 272076 258264 272088
rect 258316 272076 258322 272128
rect 292574 272076 292580 272128
rect 292632 272116 292638 272128
rect 331766 272116 331772 272128
rect 292632 272088 331772 272116
rect 292632 272076 292638 272088
rect 331766 272076 331772 272088
rect 331824 272076 331830 272128
rect 331858 272076 331864 272128
rect 331916 272116 331922 272128
rect 434622 272116 434628 272128
rect 331916 272088 434628 272116
rect 331916 272076 331922 272088
rect 434622 272076 434628 272088
rect 434680 272076 434686 272128
rect 435726 272076 435732 272128
rect 435784 272116 435790 272128
rect 642634 272116 642640 272128
rect 435784 272088 642640 272116
rect 435784 272076 435790 272088
rect 642634 272076 642640 272088
rect 642692 272076 642698 272128
rect 260006 272048 260012 272060
rect 240836 271952 245654 271980
rect 246500 272020 260012 272048
rect 240836 271940 240842 271952
rect 82446 271872 82452 271924
rect 82504 271912 82510 271924
rect 198550 271912 198556 271924
rect 82504 271884 198556 271912
rect 82504 271872 82510 271884
rect 198550 271872 198556 271884
rect 198608 271872 198614 271924
rect 245562 271872 245568 271924
rect 245620 271912 245626 271924
rect 246500 271912 246528 272020
rect 260006 272008 260012 272020
rect 260064 272008 260070 272060
rect 287146 272008 287152 272060
rect 287204 272048 287210 272060
rect 317598 272048 317604 272060
rect 287204 272020 317604 272048
rect 287204 272008 287210 272020
rect 317598 272008 317604 272020
rect 317656 272008 317662 272060
rect 317874 272008 317880 272060
rect 317932 272048 317938 272060
rect 399202 272048 399208 272060
rect 317932 272020 399208 272048
rect 317932 272008 317938 272020
rect 399202 272008 399208 272020
rect 399260 272008 399266 272060
rect 399570 272008 399576 272060
rect 399628 272048 399634 272060
rect 611906 272048 611912 272060
rect 399628 272020 611912 272048
rect 399628 272008 399634 272020
rect 611906 272008 611912 272020
rect 611964 272008 611970 272060
rect 262122 271940 262128 271992
rect 262180 271980 262186 271992
rect 266262 271980 266268 271992
rect 262180 271952 266268 271980
rect 262180 271940 262186 271952
rect 266262 271940 266268 271952
rect 266320 271940 266326 271992
rect 286962 271940 286968 271992
rect 287020 271980 287026 271992
rect 316402 271980 316408 271992
rect 287020 271952 316408 271980
rect 287020 271940 287026 271952
rect 316402 271940 316408 271952
rect 316460 271940 316466 271992
rect 318794 271940 318800 271992
rect 318852 271980 318858 271992
rect 401502 271980 401508 271992
rect 318852 271952 401508 271980
rect 318852 271940 318858 271952
rect 401502 271940 401508 271952
rect 401560 271940 401566 271992
rect 407390 271940 407396 271992
rect 407448 271980 407454 271992
rect 407448 271952 413600 271980
rect 407448 271940 407454 271952
rect 259546 271912 259552 271924
rect 245620 271884 246528 271912
rect 246684 271884 259552 271912
rect 245620 271872 245626 271884
rect 65886 271804 65892 271856
rect 65944 271844 65950 271856
rect 176838 271844 176844 271856
rect 65944 271816 176844 271844
rect 65944 271804 65950 271816
rect 176838 271804 176844 271816
rect 176896 271804 176902 271856
rect 194686 271804 194692 271856
rect 194744 271844 194750 271856
rect 240870 271844 240876 271856
rect 194744 271816 240876 271844
rect 194744 271804 194750 271816
rect 240870 271804 240876 271816
rect 240928 271804 240934 271856
rect 244366 271804 244372 271856
rect 244424 271844 244430 271856
rect 246684 271844 246712 271884
rect 259546 271872 259552 271884
rect 259604 271872 259610 271924
rect 289538 271872 289544 271924
rect 289596 271912 289602 271924
rect 322382 271912 322388 271924
rect 289596 271884 322388 271912
rect 289596 271872 289602 271884
rect 322382 271872 322388 271884
rect 322440 271872 322446 271924
rect 406286 271912 406292 271924
rect 322906 271884 406292 271912
rect 244424 271816 246712 271844
rect 244424 271804 244430 271816
rect 246758 271804 246764 271856
rect 246816 271844 246822 271856
rect 260466 271844 260472 271856
rect 246816 271816 260472 271844
rect 246816 271804 246822 271816
rect 260466 271804 260472 271816
rect 260524 271804 260530 271856
rect 264422 271804 264428 271856
rect 264480 271844 264486 271856
rect 267182 271844 267188 271856
rect 264480 271816 267188 271844
rect 264480 271804 264486 271816
rect 267182 271804 267188 271816
rect 267240 271804 267246 271856
rect 289630 271804 289636 271856
rect 289688 271844 289694 271856
rect 289688 271816 313504 271844
rect 289688 271804 289694 271816
rect 155678 271736 155684 271788
rect 155736 271776 155742 271788
rect 225874 271776 225880 271788
rect 155736 271748 225880 271776
rect 155736 271736 155742 271748
rect 225874 271736 225880 271748
rect 225932 271736 225938 271788
rect 249058 271736 249064 271788
rect 249116 271776 249122 271788
rect 261386 271776 261392 271788
rect 249116 271748 261392 271776
rect 249116 271736 249122 271748
rect 261386 271736 261392 271748
rect 261444 271736 261450 271788
rect 291654 271736 291660 271788
rect 291712 271776 291718 271788
rect 313366 271776 313372 271788
rect 291712 271748 313372 271776
rect 291712 271736 291718 271748
rect 313366 271736 313372 271748
rect 313424 271736 313430 271788
rect 161566 271668 161572 271720
rect 161624 271708 161630 271720
rect 227990 271708 227996 271720
rect 161624 271680 227996 271708
rect 161624 271668 161630 271680
rect 227990 271668 227996 271680
rect 228048 271668 228054 271720
rect 251450 271668 251456 271720
rect 251508 271708 251514 271720
rect 262214 271708 262220 271720
rect 251508 271680 262220 271708
rect 251508 271668 251514 271680
rect 262214 271668 262220 271680
rect 262272 271668 262278 271720
rect 285398 271668 285404 271720
rect 285456 271708 285462 271720
rect 312906 271708 312912 271720
rect 285456 271680 312912 271708
rect 285456 271668 285462 271680
rect 312906 271668 312912 271680
rect 312964 271668 312970 271720
rect 163958 271600 163964 271652
rect 164016 271640 164022 271652
rect 229738 271640 229744 271652
rect 164016 271612 229744 271640
rect 164016 271600 164022 271612
rect 229738 271600 229744 271612
rect 229796 271600 229802 271652
rect 253842 271600 253848 271652
rect 253900 271640 253906 271652
rect 263134 271640 263140 271652
rect 253900 271612 263140 271640
rect 253900 271600 253906 271612
rect 263134 271600 263140 271612
rect 263192 271600 263198 271652
rect 290734 271600 290740 271652
rect 290792 271640 290798 271652
rect 313274 271640 313280 271652
rect 290792 271612 313280 271640
rect 290792 271600 290798 271612
rect 313274 271600 313280 271612
rect 313332 271600 313338 271652
rect 313476 271640 313504 271816
rect 313550 271804 313556 271856
rect 313608 271804 313614 271856
rect 320542 271804 320548 271856
rect 320600 271844 320606 271856
rect 322906 271844 322934 271884
rect 406286 271872 406292 271884
rect 406344 271872 406350 271924
rect 411438 271872 411444 271924
rect 411496 271912 411502 271924
rect 413572 271912 413600 271952
rect 413646 271940 413652 271992
rect 413704 271980 413710 271992
rect 622578 271980 622584 271992
rect 413704 271952 622584 271980
rect 413704 271940 413710 271952
rect 622578 271940 622584 271952
rect 622636 271940 622642 271992
rect 636746 271912 636752 271924
rect 411496 271884 413508 271912
rect 413572 271884 636752 271912
rect 411496 271872 411502 271884
rect 320600 271816 322934 271844
rect 320600 271804 320606 271816
rect 323210 271804 323216 271856
rect 323268 271844 323274 271856
rect 413370 271844 413376 271856
rect 323268 271816 413376 271844
rect 323268 271804 323274 271816
rect 413370 271804 413376 271816
rect 413428 271804 413434 271856
rect 413480 271844 413508 271884
rect 636746 271872 636752 271884
rect 636804 271872 636810 271924
rect 647418 271844 647424 271856
rect 413480 271816 647424 271844
rect 647418 271804 647424 271816
rect 647476 271804 647482 271856
rect 313568 271776 313596 271804
rect 329466 271776 329472 271788
rect 313568 271748 329472 271776
rect 329466 271736 329472 271748
rect 329524 271736 329530 271788
rect 353570 271736 353576 271788
rect 353628 271776 353634 271788
rect 493686 271776 493692 271788
rect 353628 271748 493692 271776
rect 353628 271736 353634 271748
rect 493686 271736 493692 271748
rect 493744 271736 493750 271788
rect 498654 271736 498660 271788
rect 498712 271776 498718 271788
rect 603626 271776 603632 271788
rect 498712 271748 603632 271776
rect 498712 271736 498718 271748
rect 603626 271736 603632 271748
rect 603684 271736 603690 271788
rect 313550 271668 313556 271720
rect 313608 271708 313614 271720
rect 349522 271708 349528 271720
rect 313608 271680 349528 271708
rect 313608 271668 313614 271680
rect 349522 271668 349528 271680
rect 349580 271668 349586 271720
rect 350902 271668 350908 271720
rect 350960 271708 350966 271720
rect 486602 271708 486608 271720
rect 350960 271680 486608 271708
rect 350960 271668 350966 271680
rect 486602 271668 486608 271680
rect 486660 271668 486666 271720
rect 323486 271640 323492 271652
rect 313476 271612 323492 271640
rect 323486 271600 323492 271612
rect 323544 271600 323550 271652
rect 348234 271600 348240 271652
rect 348292 271640 348298 271652
rect 479518 271640 479524 271652
rect 348292 271612 479524 271640
rect 348292 271600 348298 271612
rect 479518 271600 479524 271612
rect 479576 271600 479582 271652
rect 162762 271532 162768 271584
rect 162820 271572 162826 271584
rect 228818 271572 228824 271584
rect 162820 271544 228824 271572
rect 162820 271532 162826 271544
rect 228818 271532 228824 271544
rect 228876 271532 228882 271584
rect 257338 271532 257344 271584
rect 257396 271572 257402 271584
rect 264514 271572 264520 271584
rect 257396 271544 264520 271572
rect 257396 271532 257402 271544
rect 264514 271532 264520 271544
rect 264572 271532 264578 271584
rect 289814 271532 289820 271584
rect 289872 271572 289878 271584
rect 324682 271572 324688 271584
rect 289872 271544 324688 271572
rect 289872 271532 289878 271544
rect 324682 271532 324688 271544
rect 324740 271532 324746 271584
rect 347590 271532 347596 271584
rect 347648 271572 347654 271584
rect 477218 271572 477224 271584
rect 347648 271544 477224 271572
rect 347648 271532 347654 271544
rect 477218 271532 477224 271544
rect 477276 271532 477282 271584
rect 171042 271464 171048 271516
rect 171100 271504 171106 271516
rect 232406 271504 232412 271516
rect 171100 271476 232412 271504
rect 171100 271464 171106 271476
rect 232406 271464 232412 271476
rect 232464 271464 232470 271516
rect 258534 271464 258540 271516
rect 258592 271504 258598 271516
rect 264882 271504 264888 271516
rect 258592 271476 264888 271504
rect 258592 271464 258598 271476
rect 264882 271464 264888 271476
rect 264940 271464 264946 271516
rect 266814 271464 266820 271516
rect 266872 271504 266878 271516
rect 268010 271504 268016 271516
rect 266872 271476 268016 271504
rect 266872 271464 266878 271476
rect 268010 271464 268016 271476
rect 268068 271464 268074 271516
rect 290274 271464 290280 271516
rect 290332 271504 290338 271516
rect 290332 271476 313228 271504
rect 290332 271464 290338 271476
rect 134426 271396 134432 271448
rect 134484 271436 134490 271448
rect 195790 271436 195796 271448
rect 134484 271408 195796 271436
rect 134484 271396 134490 271408
rect 195790 271396 195796 271408
rect 195848 271396 195854 271448
rect 197078 271396 197084 271448
rect 197136 271436 197142 271448
rect 241790 271436 241796 271448
rect 197136 271408 241796 271436
rect 197136 271396 197142 271408
rect 241790 271396 241796 271408
rect 241848 271396 241854 271448
rect 254946 271396 254952 271448
rect 255004 271436 255010 271448
rect 263594 271436 263600 271448
rect 255004 271408 263600 271436
rect 255004 271396 255010 271408
rect 263594 271396 263600 271408
rect 263652 271396 263658 271448
rect 285858 271396 285864 271448
rect 285916 271436 285922 271448
rect 285916 271408 309456 271436
rect 285916 271396 285922 271408
rect 168742 271328 168748 271380
rect 168800 271368 168806 271380
rect 230658 271368 230664 271380
rect 168800 271340 230664 271368
rect 168800 271328 168806 271340
rect 230658 271328 230664 271340
rect 230716 271328 230722 271380
rect 252646 271328 252652 271380
rect 252704 271368 252710 271380
rect 262858 271368 262864 271380
rect 252704 271340 262864 271368
rect 252704 271328 252710 271340
rect 262858 271328 262864 271340
rect 262916 271328 262922 271380
rect 284202 271328 284208 271380
rect 284260 271368 284266 271380
rect 309318 271368 309324 271380
rect 284260 271340 309324 271368
rect 284260 271328 284266 271340
rect 309318 271328 309324 271340
rect 309376 271328 309382 271380
rect 169846 271260 169852 271312
rect 169904 271300 169910 271312
rect 231486 271300 231492 271312
rect 169904 271272 231492 271300
rect 169904 271260 169910 271272
rect 231486 271260 231492 271272
rect 231544 271260 231550 271312
rect 250254 271260 250260 271312
rect 250312 271300 250318 271312
rect 261846 271300 261852 271312
rect 250312 271272 261852 271300
rect 250312 271260 250318 271272
rect 261846 271260 261852 271272
rect 261904 271260 261910 271312
rect 309428 271300 309456 271408
rect 313200 271368 313228 271476
rect 313274 271464 313280 271516
rect 313332 271504 313338 271516
rect 327074 271504 327080 271516
rect 313332 271476 327080 271504
rect 313332 271464 313338 271476
rect 327074 271464 327080 271476
rect 327132 271464 327138 271516
rect 344830 271504 344836 271516
rect 332520 271476 344836 271504
rect 314654 271396 314660 271448
rect 314712 271436 314718 271448
rect 332520 271436 332548 271476
rect 344830 271464 344836 271476
rect 344888 271464 344894 271516
rect 344922 271464 344928 271516
rect 344980 271504 344986 271516
rect 470134 271504 470140 271516
rect 344980 271476 470140 271504
rect 344980 271464 344986 271476
rect 470134 271464 470140 271476
rect 470192 271464 470198 271516
rect 314712 271408 332548 271436
rect 314712 271396 314718 271408
rect 342162 271396 342168 271448
rect 342220 271436 342226 271448
rect 462958 271436 462964 271448
rect 342220 271408 462964 271436
rect 342220 271396 342226 271408
rect 462958 271396 462964 271408
rect 463016 271396 463022 271448
rect 325878 271368 325884 271380
rect 313200 271340 325884 271368
rect 325878 271328 325884 271340
rect 325936 271328 325942 271380
rect 340138 271328 340144 271380
rect 340196 271368 340202 271380
rect 458266 271368 458272 271380
rect 340196 271340 458272 271368
rect 340196 271328 340202 271340
rect 458266 271328 458272 271340
rect 458324 271328 458330 271380
rect 314102 271300 314108 271312
rect 309428 271272 314108 271300
rect 314102 271260 314108 271272
rect 314160 271260 314166 271312
rect 336458 271260 336464 271312
rect 336516 271300 336522 271312
rect 448790 271300 448796 271312
rect 336516 271272 448796 271300
rect 336516 271260 336522 271272
rect 448790 271260 448796 271272
rect 448848 271260 448854 271312
rect 176838 271192 176844 271244
rect 176896 271232 176902 271244
rect 192110 271232 192116 271244
rect 176896 271204 192116 271232
rect 176896 271192 176902 271204
rect 192110 271192 192116 271204
rect 192168 271192 192174 271244
rect 193876 271204 197308 271232
rect 178126 271124 178132 271176
rect 178184 271164 178190 271176
rect 193876 271164 193904 271204
rect 178184 271136 193904 271164
rect 197280 271164 197308 271204
rect 197354 271192 197360 271244
rect 197412 271232 197418 271244
rect 233326 271232 233332 271244
rect 197412 271204 233332 271232
rect 197412 271192 197418 271204
rect 233326 271192 233332 271204
rect 233384 271192 233390 271244
rect 337470 271192 337476 271244
rect 337528 271232 337534 271244
rect 451182 271232 451188 271244
rect 337528 271204 451188 271232
rect 337528 271192 337534 271204
rect 451182 271192 451188 271204
rect 451240 271192 451246 271244
rect 231854 271164 231860 271176
rect 197280 271136 231860 271164
rect 178184 271124 178190 271136
rect 231854 271124 231860 271136
rect 231912 271124 231918 271176
rect 334802 271124 334808 271176
rect 334860 271164 334866 271176
rect 444098 271164 444104 271176
rect 334860 271136 444104 271164
rect 334860 271124 334866 271136
rect 444098 271124 444104 271136
rect 444156 271124 444162 271176
rect 175826 271056 175832 271108
rect 175884 271096 175890 271108
rect 197170 271096 197176 271108
rect 175884 271068 197176 271096
rect 175884 271056 175890 271068
rect 197170 271056 197176 271068
rect 197228 271056 197234 271108
rect 197262 271056 197268 271108
rect 197320 271096 197326 271108
rect 234154 271096 234160 271108
rect 197320 271068 234160 271096
rect 197320 271056 197326 271068
rect 234154 271056 234160 271068
rect 234212 271056 234218 271108
rect 247862 271056 247868 271108
rect 247920 271096 247926 271108
rect 260926 271096 260932 271108
rect 247920 271068 260932 271096
rect 247920 271056 247926 271068
rect 260926 271056 260932 271068
rect 260984 271056 260990 271108
rect 332134 271056 332140 271108
rect 332192 271096 332198 271108
rect 437014 271096 437020 271108
rect 332192 271068 437020 271096
rect 332192 271056 332198 271068
rect 437014 271056 437020 271068
rect 437072 271056 437078 271108
rect 182910 270988 182916 271040
rect 182968 271028 182974 271040
rect 235994 271028 236000 271040
rect 182968 271000 236000 271028
rect 182968 270988 182974 271000
rect 235994 270988 236000 271000
rect 236052 270988 236058 271040
rect 332410 270988 332416 271040
rect 332468 271028 332474 271040
rect 429930 271028 429936 271040
rect 332468 271000 429936 271028
rect 332468 270988 332474 271000
rect 429930 270988 429936 271000
rect 429988 270988 429994 271040
rect 187602 270920 187608 270972
rect 187660 270960 187666 270972
rect 238202 270960 238208 270972
rect 187660 270932 238208 270960
rect 187660 270920 187666 270932
rect 238202 270920 238208 270932
rect 238260 270920 238266 270972
rect 328638 270920 328644 270972
rect 328696 270960 328702 270972
rect 427538 270960 427544 270972
rect 328696 270932 427544 270960
rect 328696 270920 328702 270932
rect 427538 270920 427544 270932
rect 427596 270920 427602 270972
rect 186406 270852 186412 270904
rect 186464 270892 186470 270904
rect 237282 270892 237288 270904
rect 186464 270864 237288 270892
rect 186464 270852 186470 270864
rect 237282 270852 237288 270864
rect 237340 270852 237346 270904
rect 325970 270852 325976 270904
rect 326028 270892 326034 270904
rect 420454 270892 420460 270904
rect 326028 270864 420460 270892
rect 326028 270852 326034 270864
rect 420454 270852 420460 270864
rect 420512 270852 420518 270904
rect 142706 270784 142712 270836
rect 142764 270824 142770 270836
rect 146202 270824 146208 270836
rect 142764 270796 146208 270824
rect 142764 270784 142770 270796
rect 146202 270784 146208 270796
rect 146260 270784 146266 270836
rect 188798 270784 188804 270836
rect 188856 270824 188862 270836
rect 239122 270824 239128 270836
rect 188856 270796 239128 270824
rect 188856 270784 188862 270796
rect 239122 270784 239128 270796
rect 239180 270784 239186 270836
rect 324130 270784 324136 270836
rect 324188 270824 324194 270836
rect 415762 270824 415768 270836
rect 324188 270796 415768 270824
rect 324188 270784 324194 270796
rect 415762 270784 415768 270796
rect 415820 270784 415826 270836
rect 176930 270716 176936 270768
rect 176988 270756 176994 270768
rect 197262 270756 197268 270768
rect 176988 270728 197268 270756
rect 176988 270716 176994 270728
rect 197262 270716 197268 270728
rect 197320 270716 197326 270768
rect 234614 270756 234620 270768
rect 198200 270728 234620 270756
rect 133230 270512 133236 270564
rect 133288 270552 133294 270564
rect 133288 270524 137968 270552
rect 133288 270512 133294 270524
rect 137940 270280 137968 270524
rect 191190 270512 191196 270564
rect 191248 270552 191254 270564
rect 198200 270552 198228 270728
rect 234614 270716 234620 270728
rect 234672 270716 234678 270768
rect 327166 270716 327172 270768
rect 327224 270756 327230 270768
rect 383838 270756 383844 270768
rect 327224 270728 383844 270756
rect 327224 270716 327230 270728
rect 383838 270716 383844 270728
rect 383896 270716 383902 270768
rect 386230 270716 386236 270768
rect 386288 270756 386294 270768
rect 391198 270756 391204 270768
rect 386288 270728 391204 270756
rect 386288 270716 386294 270728
rect 391198 270716 391204 270728
rect 391256 270716 391262 270768
rect 402054 270716 402060 270768
rect 402112 270756 402118 270768
rect 413646 270756 413652 270768
rect 402112 270728 413652 270756
rect 402112 270716 402118 270728
rect 413646 270716 413652 270728
rect 413704 270716 413710 270768
rect 199562 270648 199568 270700
rect 199620 270688 199626 270700
rect 242618 270688 242624 270700
rect 199620 270660 242624 270688
rect 199620 270648 199626 270660
rect 242618 270648 242624 270660
rect 242676 270648 242682 270700
rect 256142 270648 256148 270700
rect 256200 270688 256206 270700
rect 264054 270688 264060 270700
rect 256200 270660 264060 270688
rect 256200 270648 256206 270660
rect 264054 270648 264060 270660
rect 264112 270648 264118 270700
rect 320174 270648 320180 270700
rect 320232 270688 320238 270700
rect 374362 270688 374368 270700
rect 320232 270660 374368 270688
rect 320232 270648 320238 270660
rect 374362 270648 374368 270660
rect 374420 270648 374426 270700
rect 383470 270648 383476 270700
rect 383528 270688 383534 270700
rect 391566 270688 391572 270700
rect 383528 270660 391572 270688
rect 383528 270648 383534 270660
rect 391566 270648 391572 270660
rect 391624 270648 391630 270700
rect 198274 270580 198280 270632
rect 198332 270620 198338 270632
rect 242250 270620 242256 270632
rect 198332 270592 242256 270620
rect 198332 270580 198338 270592
rect 242250 270580 242256 270592
rect 242308 270580 242314 270632
rect 327534 270580 327540 270632
rect 327592 270620 327598 270632
rect 376754 270620 376760 270632
rect 327592 270592 376760 270620
rect 327592 270580 327598 270592
rect 376754 270580 376760 270592
rect 376812 270580 376818 270632
rect 388990 270580 388996 270632
rect 389048 270620 389054 270632
rect 391106 270620 391112 270632
rect 389048 270592 391112 270620
rect 389048 270580 389054 270592
rect 391106 270580 391112 270592
rect 391164 270580 391170 270632
rect 191248 270524 198228 270552
rect 191248 270512 191254 270524
rect 312538 270512 312544 270564
rect 312596 270552 312602 270564
rect 342438 270552 342444 270564
rect 312596 270524 342444 270552
rect 312596 270512 312602 270524
rect 342438 270512 342444 270524
rect 342496 270512 342502 270564
rect 347130 270552 347136 270564
rect 344664 270524 347136 270552
rect 147398 270444 147404 270496
rect 147456 270484 147462 270496
rect 208118 270484 208124 270496
rect 147456 270456 208124 270484
rect 147456 270444 147462 270456
rect 208118 270444 208124 270456
rect 208176 270444 208182 270496
rect 220814 270484 220820 270496
rect 208228 270456 220820 270484
rect 141510 270376 141516 270428
rect 141568 270416 141574 270428
rect 208228 270416 208256 270456
rect 220814 270444 220820 270456
rect 220872 270444 220878 270496
rect 225414 270444 225420 270496
rect 225472 270484 225478 270496
rect 252462 270484 252468 270496
rect 225472 270456 252468 270484
rect 225472 270444 225478 270456
rect 252462 270444 252468 270456
rect 252520 270444 252526 270496
rect 265618 270444 265624 270496
rect 265676 270484 265682 270496
rect 267550 270484 267556 270496
rect 265676 270456 267556 270484
rect 265676 270444 265682 270456
rect 267550 270444 267556 270456
rect 267608 270444 267614 270496
rect 269390 270444 269396 270496
rect 269448 270484 269454 270496
rect 270310 270484 270316 270496
rect 269448 270456 270316 270484
rect 269448 270444 269454 270456
rect 270310 270444 270316 270456
rect 270368 270444 270374 270496
rect 271138 270444 271144 270496
rect 271196 270484 271202 270496
rect 275094 270484 275100 270496
rect 271196 270456 275100 270484
rect 271196 270444 271202 270456
rect 275094 270444 275100 270456
rect 275152 270444 275158 270496
rect 276934 270444 276940 270496
rect 276992 270484 276998 270496
rect 290458 270484 290464 270496
rect 276992 270456 290464 270484
rect 276992 270444 276998 270456
rect 290458 270444 290464 270456
rect 290516 270444 290522 270496
rect 295610 270444 295616 270496
rect 295668 270484 295674 270496
rect 340046 270484 340052 270496
rect 295668 270456 340052 270484
rect 295668 270444 295674 270456
rect 340046 270444 340052 270456
rect 340104 270444 340110 270496
rect 219986 270416 219992 270428
rect 141568 270388 208256 270416
rect 208320 270388 219992 270416
rect 141568 270376 141574 270388
rect 140314 270308 140320 270360
rect 140372 270348 140378 270360
rect 208320 270348 208348 270388
rect 219986 270376 219992 270388
rect 220044 270376 220050 270428
rect 224218 270376 224224 270428
rect 224276 270416 224282 270428
rect 252002 270416 252008 270428
rect 224276 270388 252008 270416
rect 224276 270376 224282 270388
rect 252002 270376 252008 270388
rect 252060 270376 252066 270428
rect 269850 270376 269856 270428
rect 269908 270416 269914 270428
rect 271506 270416 271512 270428
rect 269908 270388 271512 270416
rect 269908 270376 269914 270388
rect 271506 270376 271512 270388
rect 271564 270376 271570 270428
rect 271598 270376 271604 270428
rect 271656 270416 271662 270428
rect 276198 270416 276204 270428
rect 271656 270388 276204 270416
rect 271656 270376 271662 270388
rect 276198 270376 276204 270388
rect 276256 270376 276262 270428
rect 277486 270376 277492 270428
rect 277544 270416 277550 270428
rect 277544 270388 281672 270416
rect 277544 270376 277550 270388
rect 219066 270348 219072 270360
rect 140372 270320 208348 270348
rect 218026 270320 219072 270348
rect 140372 270308 140378 270320
rect 207842 270280 207848 270292
rect 137940 270252 207848 270280
rect 207842 270240 207848 270252
rect 207900 270240 207906 270292
rect 207934 270240 207940 270292
rect 207992 270280 207998 270292
rect 215478 270280 215484 270292
rect 207992 270252 215484 270280
rect 207992 270240 207998 270252
rect 215478 270240 215484 270252
rect 215536 270240 215542 270292
rect 135622 270172 135628 270224
rect 135680 270212 135686 270224
rect 218026 270212 218054 270320
rect 219066 270308 219072 270320
rect 219124 270308 219130 270360
rect 221918 270308 221924 270360
rect 221976 270348 221982 270360
rect 251082 270348 251088 270360
rect 221976 270320 251088 270348
rect 221976 270308 221982 270320
rect 251082 270308 251088 270320
rect 251140 270308 251146 270360
rect 272058 270308 272064 270360
rect 272116 270348 272122 270360
rect 277394 270348 277400 270360
rect 272116 270320 277400 270348
rect 272116 270308 272122 270320
rect 277394 270308 277400 270320
rect 277452 270308 277458 270360
rect 277854 270308 277860 270360
rect 277912 270348 277918 270360
rect 281644 270348 281672 270388
rect 296990 270376 296996 270428
rect 297048 270416 297054 270428
rect 343634 270416 343640 270428
rect 297048 270388 343640 270416
rect 297048 270376 297054 270388
rect 343634 270376 343640 270388
rect 343692 270376 343698 270428
rect 291562 270348 291568 270360
rect 277912 270320 281580 270348
rect 281644 270320 291568 270348
rect 277912 270308 277918 270320
rect 218330 270240 218336 270292
rect 218388 270280 218394 270292
rect 249794 270280 249800 270292
rect 218388 270252 249800 270280
rect 218388 270240 218394 270252
rect 249794 270240 249800 270252
rect 249852 270240 249858 270292
rect 135680 270184 218054 270212
rect 135680 270172 135686 270184
rect 220722 270172 220728 270224
rect 220780 270212 220786 270224
rect 250714 270212 250720 270224
rect 220780 270184 250720 270212
rect 220780 270172 220786 270184
rect 250714 270172 250720 270184
rect 250772 270172 250778 270224
rect 270678 270172 270684 270224
rect 270736 270212 270742 270224
rect 273898 270212 273904 270224
rect 270736 270184 273904 270212
rect 270736 270172 270742 270184
rect 273898 270172 273904 270184
rect 273956 270172 273962 270224
rect 278682 270172 278688 270224
rect 278740 270212 278746 270224
rect 281552 270212 281580 270320
rect 291562 270308 291568 270320
rect 291620 270308 291626 270360
rect 298278 270308 298284 270360
rect 298336 270348 298342 270360
rect 344664 270348 344692 270524
rect 347130 270512 347136 270524
rect 347188 270512 347194 270564
rect 346026 270444 346032 270496
rect 346084 270484 346090 270496
rect 473630 270484 473636 270496
rect 346084 270456 473636 270484
rect 346084 270444 346090 270456
rect 473630 270444 473636 270456
rect 473688 270444 473694 270496
rect 346854 270376 346860 270428
rect 346912 270416 346918 270428
rect 476022 270416 476028 270428
rect 346912 270388 476028 270416
rect 346912 270376 346918 270388
rect 476022 270376 476028 270388
rect 476080 270376 476086 270428
rect 298336 270320 344692 270348
rect 298336 270308 298342 270320
rect 348602 270308 348608 270360
rect 348660 270348 348666 270360
rect 480714 270348 480720 270360
rect 348660 270320 480720 270348
rect 348660 270308 348666 270320
rect 480714 270308 480720 270320
rect 480772 270308 480778 270360
rect 297910 270240 297916 270292
rect 297968 270280 297974 270292
rect 345934 270280 345940 270292
rect 297968 270252 345940 270280
rect 297968 270240 297974 270252
rect 345934 270240 345940 270252
rect 345992 270240 345998 270292
rect 349522 270240 349528 270292
rect 349580 270280 349586 270292
rect 483106 270280 483112 270292
rect 349580 270252 483112 270280
rect 349580 270240 349586 270252
rect 483106 270240 483112 270252
rect 483164 270240 483170 270292
rect 292758 270212 292764 270224
rect 278740 270184 281488 270212
rect 281552 270184 292764 270212
rect 278740 270172 278746 270184
rect 126146 270104 126152 270156
rect 126204 270144 126210 270156
rect 213454 270144 213460 270156
rect 126204 270116 213460 270144
rect 126204 270104 126210 270116
rect 213454 270104 213460 270116
rect 213512 270104 213518 270156
rect 213638 270104 213644 270156
rect 213696 270144 213702 270156
rect 248046 270144 248052 270156
rect 213696 270116 248052 270144
rect 213696 270104 213702 270116
rect 248046 270104 248052 270116
rect 248104 270104 248110 270156
rect 272978 270104 272984 270156
rect 273036 270144 273042 270156
rect 279786 270144 279792 270156
rect 273036 270116 279792 270144
rect 273036 270104 273042 270116
rect 279786 270104 279792 270116
rect 279844 270104 279850 270156
rect 281460 270144 281488 270184
rect 292758 270172 292764 270184
rect 292816 270172 292822 270224
rect 300118 270172 300124 270224
rect 300176 270212 300182 270224
rect 347866 270212 347872 270224
rect 300176 270184 347872 270212
rect 300176 270172 300182 270184
rect 347866 270172 347872 270184
rect 347924 270172 347930 270224
rect 351270 270172 351276 270224
rect 351328 270212 351334 270224
rect 487798 270212 487804 270224
rect 351328 270184 487804 270212
rect 351328 270172 351334 270184
rect 487798 270172 487804 270184
rect 487856 270172 487862 270224
rect 295150 270144 295156 270156
rect 281460 270116 295156 270144
rect 295150 270104 295156 270116
rect 295208 270104 295214 270156
rect 298738 270104 298744 270156
rect 298796 270144 298802 270156
rect 348326 270144 348332 270156
rect 298796 270116 348332 270144
rect 298796 270104 298802 270116
rect 348326 270104 348332 270116
rect 348384 270104 348390 270156
rect 359366 270104 359372 270156
rect 359424 270144 359430 270156
rect 509050 270144 509056 270156
rect 359424 270116 509056 270144
rect 359424 270104 359430 270116
rect 509050 270104 509056 270116
rect 509108 270104 509114 270156
rect 127342 270036 127348 270088
rect 127400 270076 127406 270088
rect 207934 270076 207940 270088
rect 127400 270048 207940 270076
rect 127400 270036 127406 270048
rect 207934 270036 207940 270048
rect 207992 270036 207998 270088
rect 208118 270036 208124 270088
rect 208176 270076 208182 270088
rect 222654 270076 222660 270088
rect 208176 270048 222660 270076
rect 208176 270036 208182 270048
rect 222654 270036 222660 270048
rect 222712 270036 222718 270088
rect 223114 270036 223120 270088
rect 223172 270076 223178 270088
rect 251542 270076 251548 270088
rect 223172 270048 251548 270076
rect 223172 270036 223178 270048
rect 251542 270036 251548 270048
rect 251600 270036 251606 270088
rect 273714 270036 273720 270088
rect 273772 270076 273778 270088
rect 280982 270076 280988 270088
rect 273772 270048 280988 270076
rect 273772 270036 273778 270048
rect 280982 270036 280988 270048
rect 281040 270036 281046 270088
rect 281074 270036 281080 270088
rect 281132 270076 281138 270088
rect 293954 270076 293960 270088
rect 281132 270048 293960 270076
rect 281132 270036 281138 270048
rect 293954 270036 293960 270048
rect 294012 270036 294018 270088
rect 300578 270036 300584 270088
rect 300636 270076 300642 270088
rect 353110 270076 353116 270088
rect 300636 270048 353116 270076
rect 300636 270036 300642 270048
rect 353110 270036 353116 270048
rect 353168 270036 353174 270088
rect 360194 270036 360200 270088
rect 360252 270076 360258 270088
rect 511442 270076 511448 270088
rect 360252 270048 511448 270076
rect 360252 270036 360258 270048
rect 511442 270036 511448 270048
rect 511500 270036 511506 270088
rect 121454 269968 121460 270020
rect 121512 270008 121518 270020
rect 213730 270008 213736 270020
rect 121512 269980 213736 270008
rect 121512 269968 121518 269980
rect 213730 269968 213736 269980
rect 213788 269968 213794 270020
rect 215938 269968 215944 270020
rect 215996 270008 216002 270020
rect 248874 270008 248880 270020
rect 215996 269980 248880 270008
rect 215996 269968 216002 269980
rect 248874 269968 248880 269980
rect 248932 269968 248938 270020
rect 272518 269968 272524 270020
rect 272576 270008 272582 270020
rect 278590 270008 278596 270020
rect 272576 269980 278596 270008
rect 272576 269968 272582 269980
rect 278590 269968 278596 269980
rect 278648 269968 278654 270020
rect 279142 269968 279148 270020
rect 279200 270008 279206 270020
rect 296346 270008 296352 270020
rect 279200 269980 296352 270008
rect 279200 269968 279206 269980
rect 296346 269968 296352 269980
rect 296404 269968 296410 270020
rect 303246 269968 303252 270020
rect 303304 270008 303310 270020
rect 359918 270008 359924 270020
rect 303304 269980 359924 270008
rect 303304 269968 303310 269980
rect 359918 269968 359924 269980
rect 359976 269968 359982 270020
rect 364702 269968 364708 270020
rect 364760 270008 364766 270020
rect 523310 270008 523316 270020
rect 364760 269980 523316 270008
rect 364760 269968 364766 269980
rect 523310 269968 523316 269980
rect 523368 269968 523374 270020
rect 119062 269900 119068 269952
rect 119120 269940 119126 269952
rect 211890 269940 211896 269952
rect 119120 269912 211896 269940
rect 119120 269900 119126 269912
rect 211890 269900 211896 269912
rect 211948 269900 211954 269952
rect 217134 269900 217140 269952
rect 217192 269940 217198 269952
rect 249334 269940 249340 269952
rect 217192 269912 249340 269940
rect 217192 269900 217198 269912
rect 249334 269900 249340 269912
rect 249392 269900 249398 269952
rect 279602 269900 279608 269952
rect 279660 269940 279666 269952
rect 297542 269940 297548 269952
rect 279660 269912 297548 269940
rect 279660 269900 279666 269912
rect 297542 269900 297548 269912
rect 297600 269900 297606 269952
rect 302786 269900 302792 269952
rect 302844 269940 302850 269952
rect 358998 269940 359004 269952
rect 302844 269912 359004 269940
rect 302844 269900 302850 269912
rect 358998 269900 359004 269912
rect 359056 269900 359062 269952
rect 367370 269900 367376 269952
rect 367428 269940 367434 269952
rect 530394 269940 530400 269952
rect 367428 269912 530400 269940
rect 367428 269900 367434 269912
rect 530394 269900 530400 269912
rect 530452 269900 530458 269952
rect 114370 269832 114376 269884
rect 114428 269872 114434 269884
rect 211062 269872 211068 269884
rect 114428 269844 211068 269872
rect 114428 269832 114434 269844
rect 211062 269832 211068 269844
rect 211120 269832 211126 269884
rect 212442 269832 212448 269884
rect 212500 269872 212506 269884
rect 247586 269872 247592 269884
rect 212500 269844 247592 269872
rect 212500 269832 212506 269844
rect 247586 269832 247592 269844
rect 247644 269832 247650 269884
rect 280062 269832 280068 269884
rect 280120 269872 280126 269884
rect 298462 269872 298468 269884
rect 280120 269844 298468 269872
rect 280120 269832 280126 269844
rect 298462 269832 298468 269844
rect 298520 269832 298526 269884
rect 305454 269832 305460 269884
rect 305512 269872 305518 269884
rect 366082 269872 366088 269884
rect 305512 269844 366088 269872
rect 305512 269832 305518 269844
rect 366082 269832 366088 269844
rect 366140 269832 366146 269884
rect 368198 269832 368204 269884
rect 368256 269872 368262 269884
rect 532694 269872 532700 269884
rect 368256 269844 532700 269872
rect 368256 269832 368262 269844
rect 532694 269832 532700 269844
rect 532752 269832 532758 269884
rect 113174 269764 113180 269816
rect 113232 269804 113238 269816
rect 210142 269804 210148 269816
rect 113232 269776 210148 269804
rect 113232 269764 113238 269776
rect 210142 269764 210148 269776
rect 210200 269764 210206 269816
rect 214834 269764 214840 269816
rect 214892 269804 214898 269816
rect 248414 269804 248420 269816
rect 214892 269776 248420 269804
rect 214892 269764 214898 269776
rect 248414 269764 248420 269776
rect 248472 269764 248478 269816
rect 280522 269764 280528 269816
rect 280580 269804 280586 269816
rect 299842 269804 299848 269816
rect 280580 269776 299848 269804
rect 280580 269764 280586 269776
rect 299842 269764 299848 269776
rect 299900 269764 299906 269816
rect 306742 269764 306748 269816
rect 306800 269804 306806 269816
rect 369578 269804 369584 269816
rect 306800 269776 369584 269804
rect 306800 269764 306806 269776
rect 369578 269764 369584 269776
rect 369636 269764 369642 269816
rect 372706 269764 372712 269816
rect 372764 269804 372770 269816
rect 544562 269804 544568 269816
rect 372764 269776 544568 269804
rect 372764 269764 372770 269776
rect 544562 269764 544568 269776
rect 544620 269764 544626 269816
rect 109586 269696 109592 269748
rect 109644 269736 109650 269748
rect 208854 269736 208860 269748
rect 109644 269708 208860 269736
rect 109644 269696 109650 269708
rect 208854 269696 208860 269708
rect 208912 269696 208918 269748
rect 211246 269696 211252 269748
rect 211304 269736 211310 269748
rect 247126 269736 247132 269748
rect 211304 269708 247132 269736
rect 211304 269696 211310 269708
rect 247126 269696 247132 269708
rect 247184 269696 247190 269748
rect 278314 269696 278320 269748
rect 278372 269736 278378 269748
rect 281074 269736 281080 269748
rect 278372 269708 281080 269736
rect 278372 269696 278378 269708
rect 281074 269696 281080 269708
rect 281132 269696 281138 269748
rect 284478 269736 284484 269748
rect 281184 269708 284484 269736
rect 108390 269628 108396 269680
rect 108448 269668 108454 269680
rect 207934 269668 207940 269680
rect 108448 269640 207940 269668
rect 108448 269628 108454 269640
rect 207934 269628 207940 269640
rect 207992 269628 207998 269680
rect 208026 269628 208032 269680
rect 208084 269668 208090 269680
rect 245746 269668 245752 269680
rect 208084 269640 245752 269668
rect 208084 269628 208090 269640
rect 245746 269628 245752 269640
rect 245804 269628 245810 269680
rect 274726 269628 274732 269680
rect 274784 269668 274790 269680
rect 281184 269668 281212 269708
rect 284478 269696 284484 269708
rect 284536 269696 284542 269748
rect 305914 269696 305920 269748
rect 305972 269736 305978 269748
rect 367278 269736 367284 269748
rect 305972 269708 367284 269736
rect 305972 269696 305978 269708
rect 367278 269696 367284 269708
rect 367336 269696 367342 269748
rect 373994 269696 374000 269748
rect 374052 269736 374058 269748
rect 548058 269736 548064 269748
rect 374052 269708 548064 269736
rect 374052 269696 374058 269708
rect 548058 269696 548064 269708
rect 548116 269696 548122 269748
rect 274784 269640 281212 269668
rect 274784 269628 274790 269640
rect 281810 269628 281816 269680
rect 281868 269668 281874 269680
rect 303430 269668 303436 269680
rect 281868 269640 303436 269668
rect 281868 269628 281874 269640
rect 303430 269628 303436 269640
rect 303488 269628 303494 269680
rect 308214 269628 308220 269680
rect 308272 269668 308278 269680
rect 373166 269668 373172 269680
rect 308272 269640 373172 269668
rect 308272 269628 308278 269640
rect 373166 269628 373172 269640
rect 373224 269628 373230 269680
rect 379330 269628 379336 269680
rect 379388 269668 379394 269680
rect 562318 269668 562324 269680
rect 379388 269640 562324 269668
rect 379388 269628 379394 269640
rect 562318 269628 562324 269640
rect 562376 269628 562382 269680
rect 102502 269560 102508 269612
rect 102560 269600 102566 269612
rect 206186 269600 206192 269612
rect 102560 269572 206192 269600
rect 102560 269560 102566 269572
rect 206186 269560 206192 269572
rect 206244 269560 206250 269612
rect 210050 269560 210056 269612
rect 210108 269600 210114 269612
rect 246666 269600 246672 269612
rect 210108 269572 246672 269600
rect 210108 269560 210114 269572
rect 246666 269560 246672 269572
rect 246724 269560 246730 269612
rect 281442 269560 281448 269612
rect 281500 269600 281506 269612
rect 302234 269600 302240 269612
rect 281500 269572 302240 269600
rect 281500 269560 281506 269572
rect 302234 269560 302240 269572
rect 302292 269560 302298 269612
rect 310790 269560 310796 269612
rect 310848 269600 310854 269612
rect 380250 269600 380256 269612
rect 310848 269572 380256 269600
rect 310848 269560 310854 269572
rect 380250 269560 380256 269572
rect 380308 269560 380314 269612
rect 384666 269560 384672 269612
rect 384724 269600 384730 269612
rect 576486 269600 576492 269612
rect 384724 269572 576492 269600
rect 384724 269560 384730 269572
rect 576486 269560 576492 269572
rect 576544 269560 576550 269612
rect 94222 269492 94228 269544
rect 94280 269532 94286 269544
rect 202598 269532 202604 269544
rect 94280 269504 202604 269532
rect 94280 269492 94286 269504
rect 202598 269492 202604 269504
rect 202656 269492 202662 269544
rect 209130 269492 209136 269544
rect 209188 269532 209194 269544
rect 246206 269532 246212 269544
rect 209188 269504 246212 269532
rect 209188 269492 209194 269504
rect 246206 269492 246212 269504
rect 246264 269492 246270 269544
rect 280982 269492 280988 269544
rect 281040 269532 281046 269544
rect 301038 269532 301044 269544
rect 281040 269504 301044 269532
rect 281040 269492 281046 269504
rect 301038 269492 301044 269504
rect 301096 269492 301102 269544
rect 313458 269492 313464 269544
rect 313516 269532 313522 269544
rect 386966 269532 386972 269544
rect 313516 269504 386972 269532
rect 313516 269492 313522 269504
rect 386966 269492 386972 269504
rect 387024 269492 387030 269544
rect 387334 269492 387340 269544
rect 387392 269532 387398 269544
rect 583570 269532 583576 269544
rect 387392 269504 583576 269532
rect 387392 269492 387398 269504
rect 583570 269492 583576 269504
rect 583628 269492 583634 269544
rect 95418 269424 95424 269476
rect 95476 269464 95482 269476
rect 203518 269464 203524 269476
rect 95476 269436 203524 269464
rect 95476 269424 95482 269436
rect 203518 269424 203524 269436
rect 203576 269424 203582 269476
rect 206554 269424 206560 269476
rect 206612 269464 206618 269476
rect 245286 269464 245292 269476
rect 206612 269436 245292 269464
rect 206612 269424 206618 269436
rect 245286 269424 245292 269436
rect 245344 269424 245350 269476
rect 282730 269424 282736 269476
rect 282788 269464 282794 269476
rect 305822 269464 305828 269476
rect 282788 269436 305828 269464
rect 282788 269424 282794 269436
rect 305822 269424 305828 269436
rect 305880 269424 305886 269476
rect 316126 269424 316132 269476
rect 316184 269464 316190 269476
rect 316184 269436 387656 269464
rect 316184 269424 316190 269436
rect 42426 269356 42432 269408
rect 42484 269396 42490 269408
rect 43254 269396 43260 269408
rect 42484 269368 43260 269396
rect 42484 269356 42490 269368
rect 43254 269356 43260 269368
rect 43312 269356 43318 269408
rect 87138 269356 87144 269408
rect 87196 269396 87202 269408
rect 200390 269396 200396 269408
rect 87196 269368 200396 269396
rect 87196 269356 87202 269368
rect 200390 269356 200396 269368
rect 200448 269356 200454 269408
rect 202966 269356 202972 269408
rect 203024 269396 203030 269408
rect 243998 269396 244004 269408
rect 203024 269368 244004 269396
rect 203024 269356 203030 269368
rect 243998 269356 244004 269368
rect 244056 269356 244062 269408
rect 282270 269356 282276 269408
rect 282328 269396 282334 269408
rect 304626 269396 304632 269408
rect 282328 269368 304632 269396
rect 282328 269356 282334 269368
rect 304626 269356 304632 269368
rect 304684 269356 304690 269408
rect 316586 269356 316592 269408
rect 316644 269396 316650 269408
rect 387628 269396 387656 269436
rect 392762 269424 392768 269476
rect 392820 269464 392826 269476
rect 597738 269464 597744 269476
rect 392820 269436 597744 269464
rect 392820 269424 392826 269436
rect 597738 269424 597744 269436
rect 597796 269424 597802 269476
rect 394418 269396 394424 269408
rect 316644 269368 387564 269396
rect 387628 269368 394424 269396
rect 316644 269356 316650 269368
rect 75362 269288 75368 269340
rect 75420 269328 75426 269340
rect 195422 269328 195428 269340
rect 75420 269300 195428 269328
rect 75420 269288 75426 269300
rect 195422 269288 195428 269300
rect 195480 269288 195486 269340
rect 204162 269288 204168 269340
rect 204220 269328 204226 269340
rect 244458 269328 244464 269340
rect 204220 269300 244464 269328
rect 204220 269288 204226 269300
rect 244458 269288 244464 269300
rect 244516 269288 244522 269340
rect 283650 269288 283656 269340
rect 283708 269328 283714 269340
rect 308122 269328 308128 269340
rect 283708 269300 308128 269328
rect 283708 269288 283714 269300
rect 308122 269288 308128 269300
rect 308180 269288 308186 269340
rect 317506 269288 317512 269340
rect 317564 269328 317570 269340
rect 387426 269328 387432 269340
rect 317564 269300 387432 269328
rect 317564 269288 317570 269300
rect 387426 269288 387432 269300
rect 387484 269288 387490 269340
rect 387536 269328 387564 269368
rect 394418 269356 394424 269368
rect 394476 269356 394482 269408
rect 396718 269356 396724 269408
rect 396776 269396 396782 269408
rect 608410 269396 608416 269408
rect 396776 269368 608416 269396
rect 396776 269356 396782 269368
rect 608410 269356 608416 269368
rect 608468 269356 608474 269408
rect 395614 269328 395620 269340
rect 387536 269300 395620 269328
rect 395614 269288 395620 269300
rect 395672 269288 395678 269340
rect 399386 269288 399392 269340
rect 399444 269328 399450 269340
rect 615494 269328 615500 269340
rect 399444 269300 615500 269328
rect 399444 269288 399450 269300
rect 615494 269288 615500 269300
rect 615552 269288 615558 269340
rect 72970 269220 72976 269272
rect 73028 269260 73034 269272
rect 195054 269260 195060 269272
rect 73028 269232 195060 269260
rect 73028 269220 73034 269232
rect 195054 269220 195060 269232
rect 195112 269220 195118 269272
rect 200574 269220 200580 269272
rect 200632 269260 200638 269272
rect 243078 269260 243084 269272
rect 200632 269232 243084 269260
rect 200632 269220 200638 269232
rect 243078 269220 243084 269232
rect 243136 269220 243142 269272
rect 283190 269220 283196 269272
rect 283248 269260 283254 269272
rect 307018 269260 307024 269272
rect 283248 269232 307024 269260
rect 283248 269220 283254 269232
rect 307018 269220 307024 269232
rect 307076 269220 307082 269272
rect 319254 269220 319260 269272
rect 319312 269260 319318 269272
rect 319312 269232 397316 269260
rect 319312 269220 319318 269232
rect 195882 269152 195888 269204
rect 195940 269192 195946 269204
rect 241330 269192 241336 269204
rect 195940 269164 241336 269192
rect 195940 269152 195946 269164
rect 241330 269152 241336 269164
rect 241388 269152 241394 269204
rect 284938 269152 284944 269204
rect 284996 269192 285002 269204
rect 311710 269192 311716 269204
rect 284996 269164 311716 269192
rect 284996 269152 285002 269164
rect 311710 269152 311716 269164
rect 311768 269152 311774 269204
rect 321922 269152 321928 269204
rect 321980 269192 321986 269204
rect 397178 269192 397184 269204
rect 321980 269164 397184 269192
rect 321980 269152 321986 269164
rect 397178 269152 397184 269164
rect 397236 269152 397242 269204
rect 397288 269192 397316 269232
rect 400766 269220 400772 269272
rect 400824 269260 400830 269272
rect 618990 269260 618996 269272
rect 400824 269232 618996 269260
rect 400824 269220 400830 269232
rect 618990 269220 618996 269232
rect 619048 269220 619054 269272
rect 402698 269192 402704 269204
rect 397288 269164 402704 269192
rect 402698 269152 402704 269164
rect 402756 269152 402762 269204
rect 408770 269152 408776 269204
rect 408828 269192 408834 269204
rect 640334 269192 640340 269204
rect 408828 269164 640340 269192
rect 408828 269152 408834 269164
rect 640334 269152 640340 269164
rect 640392 269152 640398 269204
rect 67082 269084 67088 269136
rect 67140 269124 67146 269136
rect 192754 269124 192760 269136
rect 67140 269096 192760 269124
rect 67140 269084 67146 269096
rect 192754 269084 192760 269096
rect 192812 269084 192818 269136
rect 193490 269084 193496 269136
rect 193548 269124 193554 269136
rect 240410 269124 240416 269136
rect 193548 269096 240416 269124
rect 193548 269084 193554 269096
rect 240410 269084 240416 269096
rect 240468 269084 240474 269136
rect 270310 269084 270316 269136
rect 270368 269124 270374 269136
rect 272702 269124 272708 269136
rect 270368 269096 272708 269124
rect 270368 269084 270374 269096
rect 272702 269084 272708 269096
rect 272760 269084 272766 269136
rect 284478 269084 284484 269136
rect 284536 269124 284542 269136
rect 310514 269124 310520 269136
rect 284536 269096 310520 269124
rect 284536 269084 284542 269096
rect 310514 269084 310520 269096
rect 310572 269084 310578 269136
rect 322842 269084 322848 269136
rect 322900 269124 322906 269136
rect 401594 269124 401600 269136
rect 322900 269096 401600 269124
rect 322900 269084 322906 269096
rect 401594 269084 401600 269096
rect 401652 269084 401658 269136
rect 403894 269084 403900 269136
rect 403952 269124 403958 269136
rect 405366 269124 405372 269136
rect 403952 269096 405372 269124
rect 403952 269084 403958 269096
rect 405366 269084 405372 269096
rect 405424 269084 405430 269136
rect 411898 269084 411904 269136
rect 411956 269124 411962 269136
rect 648706 269124 648712 269136
rect 411956 269096 648712 269124
rect 411956 269084 411962 269096
rect 648706 269084 648712 269096
rect 648764 269084 648770 269136
rect 153378 269016 153384 269068
rect 153436 269056 153442 269068
rect 225782 269056 225788 269068
rect 153436 269028 225788 269056
rect 153436 269016 153442 269028
rect 225782 269016 225788 269028
rect 225840 269016 225846 269068
rect 234614 269016 234620 269068
rect 234672 269056 234678 269068
rect 239582 269056 239588 269068
rect 234672 269028 239588 269056
rect 234672 269016 234678 269028
rect 239582 269016 239588 269028
rect 239640 269016 239646 269068
rect 294322 269016 294328 269068
rect 294380 269056 294386 269068
rect 336550 269056 336556 269068
rect 294380 269028 336556 269056
rect 294380 269016 294386 269028
rect 336550 269016 336556 269028
rect 336608 269016 336614 269068
rect 343266 269016 343272 269068
rect 343324 269056 343330 269068
rect 466546 269056 466552 269068
rect 343324 269028 466552 269056
rect 343324 269016 343330 269028
rect 466546 269016 466552 269028
rect 466604 269016 466610 269068
rect 152182 268948 152188 269000
rect 152240 268988 152246 269000
rect 224862 268988 224868 269000
rect 152240 268960 224868 268988
rect 152240 268948 152246 268960
rect 224862 268948 224868 268960
rect 224920 268948 224926 269000
rect 292942 268948 292948 269000
rect 293000 268988 293006 269000
rect 332962 268988 332968 269000
rect 293000 268960 332968 268988
rect 293000 268948 293006 268960
rect 332962 268948 332968 268960
rect 333020 268948 333026 269000
rect 344186 268948 344192 269000
rect 344244 268988 344250 269000
rect 468938 268988 468944 269000
rect 344244 268960 468944 268988
rect 344244 268948 344250 268960
rect 468938 268948 468944 268960
rect 468996 268948 469002 269000
rect 165154 268880 165160 268932
rect 165212 268920 165218 268932
rect 229278 268920 229284 268932
rect 165212 268892 229284 268920
rect 165212 268880 165218 268892
rect 229278 268880 229284 268892
rect 229336 268880 229342 268932
rect 297450 268880 297456 268932
rect 297508 268920 297514 268932
rect 314654 268920 314660 268932
rect 297508 268892 314660 268920
rect 297508 268880 297514 268892
rect 314654 268880 314660 268892
rect 314712 268880 314718 268932
rect 341518 268880 341524 268932
rect 341576 268920 341582 268932
rect 461854 268920 461860 268932
rect 341576 268892 461860 268920
rect 341576 268880 341582 268892
rect 461854 268880 461860 268892
rect 461912 268880 461918 268932
rect 160462 268812 160468 268864
rect 160520 268852 160526 268864
rect 228450 268852 228456 268864
rect 160520 268824 228456 268852
rect 160520 268812 160526 268824
rect 228450 268812 228456 268824
rect 228508 268812 228514 268864
rect 340598 268812 340604 268864
rect 340656 268852 340662 268864
rect 459462 268852 459468 268864
rect 340656 268824 459468 268852
rect 340656 268812 340662 268824
rect 459462 268812 459468 268824
rect 459520 268812 459526 268864
rect 167546 268744 167552 268796
rect 167604 268784 167610 268796
rect 231118 268784 231124 268796
rect 167604 268756 231124 268784
rect 167604 268744 167610 268756
rect 231118 268744 231124 268756
rect 231176 268744 231182 268796
rect 296530 268744 296536 268796
rect 296588 268784 296594 268796
rect 312538 268784 312544 268796
rect 296588 268756 312544 268784
rect 296588 268744 296594 268756
rect 312538 268744 312544 268756
rect 312596 268744 312602 268796
rect 338850 268744 338856 268796
rect 338908 268784 338914 268796
rect 454678 268784 454684 268796
rect 338908 268756 454684 268784
rect 338908 268744 338914 268756
rect 454678 268744 454684 268756
rect 454736 268744 454742 268796
rect 166350 268676 166356 268728
rect 166408 268716 166414 268728
rect 230198 268716 230204 268728
rect 166408 268688 230204 268716
rect 166408 268676 166414 268688
rect 230198 268676 230204 268688
rect 230256 268676 230262 268728
rect 273806 268676 273812 268728
rect 273864 268716 273870 268728
rect 282178 268716 282184 268728
rect 273864 268688 282184 268716
rect 273864 268676 273870 268688
rect 282178 268676 282184 268688
rect 282236 268676 282242 268728
rect 309870 268676 309876 268728
rect 309928 268716 309934 268728
rect 320082 268716 320088 268728
rect 309928 268688 320088 268716
rect 309928 268676 309934 268688
rect 320082 268676 320088 268688
rect 320140 268676 320146 268728
rect 337930 268676 337936 268728
rect 337988 268716 337994 268728
rect 452378 268716 452384 268728
rect 337988 268688 452384 268716
rect 337988 268676 337994 268688
rect 452378 268676 452384 268688
rect 452436 268676 452442 268728
rect 172238 268608 172244 268660
rect 172296 268648 172302 268660
rect 231946 268648 231952 268660
rect 172296 268620 231952 268648
rect 172296 268608 172302 268620
rect 231946 268608 231952 268620
rect 232004 268608 232010 268660
rect 274266 268608 274272 268660
rect 274324 268648 274330 268660
rect 283374 268648 283380 268660
rect 274324 268620 283380 268648
rect 274324 268608 274330 268620
rect 283374 268608 283380 268620
rect 283432 268608 283438 268660
rect 299198 268608 299204 268660
rect 299256 268648 299262 268660
rect 313550 268648 313556 268660
rect 299256 268620 313556 268648
rect 299256 268608 299262 268620
rect 313550 268608 313556 268620
rect 313608 268608 313614 268660
rect 336182 268608 336188 268660
rect 336240 268648 336246 268660
rect 447594 268648 447600 268660
rect 336240 268620 447600 268648
rect 336240 268608 336246 268620
rect 447594 268608 447600 268620
rect 447652 268608 447658 268660
rect 173434 268540 173440 268592
rect 173492 268580 173498 268592
rect 232866 268580 232872 268592
rect 173492 268552 232872 268580
rect 173492 268540 173498 268552
rect 232866 268540 232872 268552
rect 232924 268540 232930 268592
rect 312538 268540 312544 268592
rect 312596 268580 312602 268592
rect 318886 268580 318892 268592
rect 312596 268552 318892 268580
rect 312596 268540 312602 268552
rect 318886 268540 318892 268552
rect 318944 268540 318950 268592
rect 335262 268540 335268 268592
rect 335320 268580 335326 268592
rect 445294 268580 445300 268592
rect 335320 268552 445300 268580
rect 335320 268540 335326 268552
rect 445294 268540 445300 268552
rect 445352 268540 445358 268592
rect 174630 268472 174636 268524
rect 174688 268512 174694 268524
rect 233786 268512 233792 268524
rect 174688 268484 233792 268512
rect 174688 268472 174694 268484
rect 233786 268472 233792 268484
rect 233844 268472 233850 268524
rect 240134 268472 240140 268524
rect 240192 268512 240198 268524
rect 243538 268512 243544 268524
rect 240192 268484 243544 268512
rect 240192 268472 240198 268484
rect 243538 268472 243544 268484
rect 243596 268472 243602 268524
rect 331306 268472 331312 268524
rect 331364 268512 331370 268524
rect 331858 268512 331864 268524
rect 331364 268484 331864 268512
rect 331364 268472 331370 268484
rect 331858 268472 331864 268484
rect 331916 268472 331922 268524
rect 333514 268472 333520 268524
rect 333572 268512 333578 268524
rect 440510 268512 440516 268524
rect 333572 268484 440516 268512
rect 333572 268472 333578 268484
rect 440510 268472 440516 268484
rect 440568 268472 440574 268524
rect 179322 268404 179328 268456
rect 179380 268444 179386 268456
rect 234614 268444 234620 268456
rect 179380 268416 234620 268444
rect 179380 268404 179386 268416
rect 234614 268404 234620 268416
rect 234672 268404 234678 268456
rect 332594 268404 332600 268456
rect 332652 268444 332658 268456
rect 438210 268444 438216 268456
rect 332652 268416 438216 268444
rect 332652 268404 332658 268416
rect 438210 268404 438216 268416
rect 438268 268404 438274 268456
rect 181714 268336 181720 268388
rect 181772 268376 181778 268388
rect 236454 268376 236460 268388
rect 181772 268348 236460 268376
rect 181772 268336 181778 268348
rect 236454 268336 236460 268348
rect 236512 268336 236518 268388
rect 330846 268336 330852 268388
rect 330904 268376 330910 268388
rect 433426 268376 433432 268388
rect 330904 268348 433432 268376
rect 330904 268336 330910 268348
rect 433426 268336 433432 268348
rect 433484 268336 433490 268388
rect 180518 268268 180524 268320
rect 180576 268308 180582 268320
rect 235534 268308 235540 268320
rect 180576 268280 235540 268308
rect 180576 268268 180582 268280
rect 235534 268268 235540 268280
rect 235592 268268 235598 268320
rect 275186 268268 275192 268320
rect 275244 268308 275250 268320
rect 285674 268308 285680 268320
rect 275244 268280 285680 268308
rect 275244 268268 275250 268280
rect 285674 268268 285680 268280
rect 285732 268268 285738 268320
rect 329926 268268 329932 268320
rect 329984 268308 329990 268320
rect 431126 268308 431132 268320
rect 329984 268280 431132 268308
rect 329984 268268 329990 268280
rect 431126 268268 431132 268280
rect 431184 268268 431190 268320
rect 184106 268200 184112 268252
rect 184164 268240 184170 268252
rect 236914 268240 236920 268252
rect 184164 268212 236920 268240
rect 184164 268200 184170 268212
rect 236914 268200 236920 268212
rect 236972 268200 236978 268252
rect 275646 268200 275652 268252
rect 275704 268240 275710 268252
rect 286870 268240 286876 268252
rect 275704 268212 286876 268240
rect 275704 268200 275710 268212
rect 286870 268200 286876 268212
rect 286928 268200 286934 268252
rect 309410 268200 309416 268252
rect 309468 268240 309474 268252
rect 327534 268240 327540 268252
rect 309468 268212 327540 268240
rect 309468 268200 309474 268212
rect 327534 268200 327540 268212
rect 327592 268200 327598 268252
rect 328178 268200 328184 268252
rect 328236 268240 328242 268252
rect 426342 268240 426348 268252
rect 328236 268212 426348 268240
rect 328236 268200 328242 268212
rect 426342 268200 426348 268212
rect 426400 268200 426406 268252
rect 185210 268132 185216 268184
rect 185268 268172 185274 268184
rect 237742 268172 237748 268184
rect 185268 268144 237748 268172
rect 185268 268132 185274 268144
rect 237742 268132 237748 268144
rect 237800 268132 237806 268184
rect 312078 268132 312084 268184
rect 312136 268172 312142 268184
rect 327166 268172 327172 268184
rect 312136 268144 327172 268172
rect 312136 268132 312142 268144
rect 327166 268132 327172 268144
rect 327224 268132 327230 268184
rect 327258 268132 327264 268184
rect 327316 268172 327322 268184
rect 423950 268172 423956 268184
rect 327316 268144 423956 268172
rect 327316 268132 327322 268144
rect 423950 268132 423956 268144
rect 424008 268132 424014 268184
rect 189994 268064 190000 268116
rect 190052 268104 190058 268116
rect 238662 268104 238668 268116
rect 190052 268076 238668 268104
rect 190052 268064 190058 268076
rect 238662 268064 238668 268076
rect 238720 268064 238726 268116
rect 313918 268064 313924 268116
rect 313976 268104 313982 268116
rect 313976 268076 332548 268104
rect 313976 268064 313982 268076
rect 192386 267996 192392 268048
rect 192444 268036 192450 268048
rect 239950 268036 239956 268048
rect 192444 268008 239956 268036
rect 192444 267996 192450 268008
rect 239950 267996 239956 268008
rect 240008 267996 240014 268048
rect 314838 267996 314844 268048
rect 314896 268036 314902 268048
rect 325326 268036 325332 268048
rect 314896 268008 325332 268036
rect 314896 267996 314902 268008
rect 325326 267996 325332 268008
rect 325384 267996 325390 268048
rect 329466 267996 329472 268048
rect 329524 268036 329530 268048
rect 332410 268036 332416 268048
rect 329524 268008 332416 268036
rect 329524 267996 329530 268008
rect 332410 267996 332416 268008
rect 332468 267996 332474 268048
rect 332520 268036 332548 268076
rect 332686 268064 332692 268116
rect 332744 268104 332750 268116
rect 332744 268076 401548 268104
rect 332744 268064 332750 268076
rect 383654 268036 383660 268048
rect 332520 268008 383660 268036
rect 383654 267996 383660 268008
rect 383712 267996 383718 268048
rect 387426 267996 387432 268048
rect 387484 268036 387490 268048
rect 398006 268036 398012 268048
rect 387484 268008 398012 268036
rect 387484 267996 387490 268008
rect 398006 267996 398012 268008
rect 398064 267996 398070 268048
rect 401520 268036 401548 268076
rect 401594 268064 401600 268116
rect 401652 268104 401658 268116
rect 412174 268104 412180 268116
rect 401652 268076 412180 268104
rect 401652 268064 401658 268076
rect 412174 268064 412180 268076
rect 412232 268064 412238 268116
rect 656158 268064 656164 268116
rect 656216 268104 656222 268116
rect 676214 268104 676220 268116
rect 656216 268076 676220 268104
rect 656216 268064 656222 268076
rect 676214 268064 676220 268076
rect 676272 268064 676278 268116
rect 416866 268036 416872 268048
rect 401520 268008 416872 268036
rect 416866 267996 416872 268008
rect 416924 267996 416930 268048
rect 195790 267928 195796 267980
rect 195848 267968 195854 267980
rect 218146 267968 218152 267980
rect 195848 267940 218152 267968
rect 195848 267928 195854 267940
rect 218146 267928 218152 267940
rect 218204 267928 218210 267980
rect 219526 267928 219532 267980
rect 219584 267968 219590 267980
rect 250254 267968 250260 267980
rect 219584 267940 250260 267968
rect 219584 267928 219590 267940
rect 250254 267928 250260 267940
rect 250312 267928 250318 267980
rect 276474 267928 276480 267980
rect 276532 267968 276538 267980
rect 289262 267968 289268 267980
rect 276532 267940 289268 267968
rect 276532 267928 276538 267940
rect 289262 267928 289268 267940
rect 289320 267928 289326 267980
rect 311250 267928 311256 267980
rect 311308 267968 311314 267980
rect 311308 267940 361574 267968
rect 311308 267928 311314 267940
rect 74166 267860 74172 267912
rect 74224 267900 74230 267912
rect 195882 267900 195888 267912
rect 74224 267872 195888 267900
rect 74224 267860 74230 267872
rect 195882 267860 195888 267872
rect 195940 267860 195946 267912
rect 207842 267860 207848 267912
rect 207900 267900 207906 267912
rect 217318 267900 217324 267912
rect 207900 267872 217324 267900
rect 207900 267860 207906 267872
rect 217318 267860 217324 267872
rect 217376 267860 217382 267912
rect 231854 267860 231860 267912
rect 231912 267900 231918 267912
rect 235074 267900 235080 267912
rect 231912 267872 235080 267900
rect 231912 267860 231918 267872
rect 235074 267860 235080 267872
rect 235132 267860 235138 267912
rect 276290 267860 276296 267912
rect 276348 267900 276354 267912
rect 288066 267900 288072 267912
rect 276348 267872 288072 267900
rect 276348 267860 276354 267872
rect 288066 267860 288072 267872
rect 288124 267860 288130 267912
rect 324590 267860 324596 267912
rect 324648 267900 324654 267912
rect 332686 267900 332692 267912
rect 324648 267872 332692 267900
rect 324648 267860 324654 267872
rect 332686 267860 332692 267872
rect 332744 267860 332750 267912
rect 361546 267900 361574 267940
rect 371326 267928 371332 267980
rect 371384 267968 371390 267980
rect 372522 267968 372528 267980
rect 371384 267940 372528 267968
rect 371384 267928 371390 267940
rect 372522 267928 372528 267940
rect 372580 267928 372586 267980
rect 397178 267928 397184 267980
rect 397236 267968 397242 267980
rect 409782 267968 409788 267980
rect 397236 267940 409788 267968
rect 397236 267928 397242 267940
rect 409782 267928 409788 267940
rect 409840 267928 409846 267980
rect 655974 267928 655980 267980
rect 656032 267968 656038 267980
rect 676030 267968 676036 267980
rect 656032 267940 676036 267968
rect 656032 267928 656038 267940
rect 676030 267928 676036 267940
rect 676088 267928 676094 267980
rect 372798 267900 372804 267912
rect 361546 267872 372804 267900
rect 372798 267860 372804 267872
rect 372856 267860 372862 267912
rect 308582 267792 308588 267844
rect 308640 267832 308646 267844
rect 320174 267832 320180 267844
rect 308640 267804 320180 267832
rect 308640 267792 308646 267804
rect 320174 267792 320180 267804
rect 320232 267792 320238 267844
rect 213454 267724 213460 267776
rect 213512 267764 213518 267776
rect 214650 267764 214656 267776
rect 213512 267736 214656 267764
rect 213512 267724 213518 267736
rect 214650 267724 214656 267736
rect 214708 267724 214714 267776
rect 398098 267724 398104 267776
rect 398156 267764 398162 267776
rect 399570 267764 399576 267776
rect 398156 267736 399576 267764
rect 398156 267724 398162 267736
rect 399570 267724 399576 267736
rect 399628 267724 399634 267776
rect 655790 267724 655796 267776
rect 655848 267764 655854 267776
rect 676122 267764 676128 267776
rect 655848 267736 676128 267764
rect 655848 267724 655854 267736
rect 676122 267724 676128 267736
rect 676180 267724 676186 267776
rect 367738 267656 367744 267708
rect 367796 267696 367802 267708
rect 531590 267696 531596 267708
rect 367796 267668 531596 267696
rect 367796 267656 367802 267668
rect 531590 267656 531596 267668
rect 531648 267656 531654 267708
rect 370498 267588 370504 267640
rect 370556 267628 370562 267640
rect 538674 267628 538680 267640
rect 370556 267600 538680 267628
rect 370556 267588 370562 267600
rect 538674 267588 538680 267600
rect 538732 267588 538738 267640
rect 373166 267520 373172 267572
rect 373224 267560 373230 267572
rect 545758 267560 545764 267572
rect 373224 267532 545764 267560
rect 373224 267520 373230 267532
rect 545758 267520 545764 267532
rect 545816 267520 545822 267572
rect 373534 267452 373540 267504
rect 373592 267492 373598 267504
rect 546954 267492 546960 267504
rect 373592 267464 546960 267492
rect 373592 267452 373598 267464
rect 546954 267452 546960 267464
rect 547012 267452 547018 267504
rect 374454 267384 374460 267436
rect 374512 267424 374518 267436
rect 549254 267424 549260 267436
rect 374512 267396 549260 267424
rect 374512 267384 374518 267396
rect 549254 267384 549260 267396
rect 549312 267384 549318 267436
rect 376202 267316 376208 267368
rect 376260 267356 376266 267368
rect 554038 267356 554044 267368
rect 376260 267328 554044 267356
rect 376260 267316 376266 267328
rect 554038 267316 554044 267328
rect 554096 267316 554102 267368
rect 375834 267248 375840 267300
rect 375892 267288 375898 267300
rect 552842 267288 552848 267300
rect 375892 267260 552848 267288
rect 375892 267248 375898 267260
rect 552842 267248 552848 267260
rect 552900 267248 552906 267300
rect 377122 267180 377128 267232
rect 377180 267220 377186 267232
rect 556338 267220 556344 267232
rect 377180 267192 556344 267220
rect 377180 267180 377186 267192
rect 556338 267180 556344 267192
rect 556396 267180 556402 267232
rect 299658 267112 299664 267164
rect 299716 267152 299722 267164
rect 350718 267152 350724 267164
rect 299716 267124 350724 267152
rect 299716 267112 299722 267124
rect 350718 267112 350724 267124
rect 350776 267112 350782 267164
rect 378502 267112 378508 267164
rect 378560 267152 378566 267164
rect 559926 267152 559932 267164
rect 378560 267124 559932 267152
rect 378560 267112 378566 267124
rect 559926 267112 559932 267124
rect 559984 267112 559990 267164
rect 300946 267044 300952 267096
rect 301004 267084 301010 267096
rect 354214 267084 354220 267096
rect 301004 267056 354220 267084
rect 301004 267044 301010 267056
rect 354214 267044 354220 267056
rect 354272 267044 354278 267096
rect 378870 267044 378876 267096
rect 378928 267084 378934 267096
rect 561122 267084 561128 267096
rect 378928 267056 561128 267084
rect 378928 267044 378934 267056
rect 561122 267044 561128 267056
rect 561180 267044 561186 267096
rect 302326 266976 302332 267028
rect 302384 267016 302390 267028
rect 357802 267016 357808 267028
rect 302384 266988 357808 267016
rect 302384 266976 302390 266988
rect 357802 266976 357808 266988
rect 357860 266976 357866 267028
rect 379790 266976 379796 267028
rect 379848 267016 379854 267028
rect 563422 267016 563428 267028
rect 379848 266988 563428 267016
rect 379848 266976 379854 266988
rect 563422 266976 563428 266988
rect 563480 266976 563486 267028
rect 303706 266908 303712 266960
rect 303764 266948 303770 266960
rect 361390 266948 361396 266960
rect 303764 266920 361396 266948
rect 303764 266908 303770 266920
rect 361390 266908 361396 266920
rect 361448 266908 361454 266960
rect 381630 266908 381636 266960
rect 381688 266948 381694 266960
rect 568206 266948 568212 266960
rect 381688 266920 568212 266948
rect 381688 266908 381694 266920
rect 568206 266908 568212 266920
rect 568264 266908 568270 266960
rect 304994 266840 305000 266892
rect 305052 266880 305058 266892
rect 364886 266880 364892 266892
rect 305052 266852 364892 266880
rect 305052 266840 305058 266852
rect 364886 266840 364892 266852
rect 364944 266840 364950 266892
rect 381170 266840 381176 266892
rect 381228 266880 381234 266892
rect 567010 266880 567016 266892
rect 381228 266852 567016 266880
rect 381228 266840 381234 266852
rect 567010 266840 567016 266852
rect 567068 266840 567074 266892
rect 306374 266772 306380 266824
rect 306432 266812 306438 266824
rect 368474 266812 368480 266824
rect 306432 266784 368480 266812
rect 306432 266772 306438 266784
rect 368474 266772 368480 266784
rect 368532 266772 368538 266824
rect 382458 266772 382464 266824
rect 382516 266812 382522 266824
rect 570598 266812 570604 266824
rect 382516 266784 570604 266812
rect 382516 266772 382522 266784
rect 570598 266772 570604 266784
rect 570656 266772 570662 266824
rect 307662 266704 307668 266756
rect 307720 266744 307726 266756
rect 371970 266744 371976 266756
rect 307720 266716 371976 266744
rect 307720 266704 307726 266716
rect 371970 266704 371976 266716
rect 372028 266704 372034 266756
rect 384298 266704 384304 266756
rect 384356 266744 384362 266756
rect 575290 266744 575296 266756
rect 384356 266716 575296 266744
rect 384356 266704 384362 266716
rect 575290 266704 575296 266716
rect 575348 266704 575354 266756
rect 309042 266636 309048 266688
rect 309100 266676 309106 266688
rect 375558 266676 375564 266688
rect 309100 266648 375564 266676
rect 309100 266636 309106 266648
rect 375558 266636 375564 266648
rect 375616 266636 375622 266688
rect 383838 266636 383844 266688
rect 383896 266676 383902 266688
rect 574094 266676 574100 266688
rect 383896 266648 574100 266676
rect 383896 266636 383902 266648
rect 574094 266636 574100 266648
rect 574152 266636 574158 266688
rect 673362 266636 673368 266688
rect 673420 266676 673426 266688
rect 676030 266676 676036 266688
rect 673420 266648 676036 266676
rect 673420 266636 673426 266648
rect 676030 266636 676036 266648
rect 676088 266636 676094 266688
rect 310330 266568 310336 266620
rect 310388 266608 310394 266620
rect 379054 266608 379060 266620
rect 310388 266580 379060 266608
rect 310388 266568 310394 266580
rect 379054 266568 379060 266580
rect 379112 266568 379118 266620
rect 385126 266568 385132 266620
rect 385184 266608 385190 266620
rect 577682 266608 577688 266620
rect 385184 266580 577688 266608
rect 385184 266568 385190 266580
rect 577682 266568 577688 266580
rect 577740 266568 577746 266620
rect 311710 266500 311716 266552
rect 311768 266540 311774 266552
rect 382642 266540 382648 266552
rect 311768 266512 382648 266540
rect 311768 266500 311774 266512
rect 382642 266500 382648 266512
rect 382700 266500 382706 266552
rect 386506 266500 386512 266552
rect 386564 266540 386570 266552
rect 581178 266540 581184 266552
rect 386564 266512 581184 266540
rect 386564 266500 386570 266512
rect 581178 266500 581184 266512
rect 581236 266500 581242 266552
rect 312998 266432 313004 266484
rect 313056 266472 313062 266484
rect 386138 266472 386144 266484
rect 313056 266444 386144 266472
rect 313056 266432 313062 266444
rect 386138 266432 386144 266444
rect 386196 266432 386202 266484
rect 387794 266432 387800 266484
rect 387852 266472 387858 266484
rect 584766 266472 584772 266484
rect 387852 266444 584772 266472
rect 387852 266432 387858 266444
rect 584766 266432 584772 266444
rect 584824 266432 584830 266484
rect 116670 266364 116676 266416
rect 116728 266404 116734 266416
rect 211522 266404 211528 266416
rect 116728 266376 211528 266404
rect 116728 266364 116734 266376
rect 211522 266364 211528 266376
rect 211580 266364 211586 266416
rect 389174 266364 389180 266416
rect 389232 266404 389238 266416
rect 588262 266404 588268 266416
rect 389232 266376 588268 266404
rect 389232 266364 389238 266376
rect 588262 266364 588268 266376
rect 588320 266364 588326 266416
rect 68186 266296 68192 266348
rect 68244 266336 68250 266348
rect 193214 266336 193220 266348
rect 68244 266308 193220 266336
rect 68244 266296 68250 266308
rect 193214 266296 193220 266308
rect 193272 266296 193278 266348
rect 315666 266296 315672 266348
rect 315724 266336 315730 266348
rect 392210 266336 392216 266348
rect 315724 266308 392216 266336
rect 315724 266296 315730 266308
rect 392210 266296 392216 266308
rect 392268 266296 392274 266348
rect 392302 266296 392308 266348
rect 392360 266336 392366 266348
rect 596542 266336 596548 266348
rect 392360 266308 596548 266336
rect 392360 266296 392366 266308
rect 596542 266296 596548 266308
rect 596600 266296 596606 266348
rect 365070 266228 365076 266280
rect 365128 266268 365134 266280
rect 524506 266268 524512 266280
rect 365128 266240 524512 266268
rect 365128 266228 365134 266240
rect 524506 266228 524512 266240
rect 524564 266228 524570 266280
rect 362402 266160 362408 266212
rect 362460 266200 362466 266212
rect 517330 266200 517336 266212
rect 362460 266172 517336 266200
rect 362460 266160 362466 266172
rect 517330 266160 517336 266172
rect 517388 266160 517394 266212
rect 359734 266092 359740 266144
rect 359792 266132 359798 266144
rect 510246 266132 510252 266144
rect 359792 266104 510252 266132
rect 359792 266092 359798 266104
rect 510246 266092 510252 266104
rect 510304 266092 510310 266144
rect 357066 266024 357072 266076
rect 357124 266064 357130 266076
rect 503162 266064 503168 266076
rect 357124 266036 503168 266064
rect 357124 266024 357130 266036
rect 503162 266024 503168 266036
rect 503220 266024 503226 266076
rect 354398 265956 354404 266008
rect 354456 265996 354462 266008
rect 496078 265996 496084 266008
rect 354456 265968 496084 265996
rect 354456 265956 354462 265968
rect 496078 265956 496084 265968
rect 496136 265956 496142 266008
rect 351730 265888 351736 265940
rect 351788 265928 351794 265940
rect 488994 265928 489000 265940
rect 351788 265900 489000 265928
rect 351788 265888 351794 265900
rect 488994 265888 489000 265900
rect 489052 265888 489058 265940
rect 349062 265820 349068 265872
rect 349120 265860 349126 265872
rect 481910 265860 481916 265872
rect 349120 265832 481916 265860
rect 349120 265820 349126 265832
rect 481910 265820 481916 265832
rect 481968 265820 481974 265872
rect 346394 265752 346400 265804
rect 346452 265792 346458 265804
rect 474826 265792 474832 265804
rect 346452 265764 474832 265792
rect 346452 265752 346458 265764
rect 474826 265752 474832 265764
rect 474884 265752 474890 265804
rect 341058 265684 341064 265736
rect 341116 265724 341122 265736
rect 460658 265724 460664 265736
rect 341116 265696 460664 265724
rect 341116 265684 341122 265696
rect 460658 265684 460664 265696
rect 460716 265684 460722 265736
rect 338390 265616 338396 265668
rect 338448 265656 338454 265668
rect 453574 265656 453580 265668
rect 338448 265628 453580 265656
rect 338448 265616 338454 265628
rect 453574 265616 453580 265628
rect 453632 265616 453638 265668
rect 317046 265548 317052 265600
rect 317104 265588 317110 265600
rect 394694 265588 394700 265600
rect 317104 265560 394700 265588
rect 317104 265548 317110 265560
rect 394694 265548 394700 265560
rect 394752 265548 394758 265600
rect 394970 265548 394976 265600
rect 395028 265588 395034 265600
rect 498654 265588 498660 265600
rect 395028 265560 498660 265588
rect 395028 265548 395034 265560
rect 498654 265548 498660 265560
rect 498712 265548 498718 265600
rect 675202 265548 675208 265600
rect 675260 265588 675266 265600
rect 676030 265588 676036 265600
rect 675260 265560 676036 265588
rect 675260 265548 675266 265560
rect 676030 265548 676036 265560
rect 676088 265548 676094 265600
rect 326798 265480 326804 265532
rect 326856 265520 326862 265532
rect 422846 265520 422852 265532
rect 326856 265492 422852 265520
rect 326856 265480 326862 265492
rect 422846 265480 422852 265492
rect 422904 265480 422910 265532
rect 325602 265412 325608 265464
rect 325660 265452 325666 265464
rect 419258 265452 419264 265464
rect 325660 265424 419264 265452
rect 325660 265412 325666 265424
rect 419258 265412 419264 265424
rect 419316 265412 419322 265464
rect 321462 265344 321468 265396
rect 321520 265384 321526 265396
rect 321520 265356 391934 265384
rect 321520 265344 321526 265356
rect 314378 265276 314384 265328
rect 314436 265316 314442 265328
rect 389726 265316 389732 265328
rect 314436 265288 389732 265316
rect 314436 265276 314442 265288
rect 389726 265276 389732 265288
rect 389784 265276 389790 265328
rect 391906 265316 391934 265356
rect 394694 265344 394700 265396
rect 394752 265384 394758 265396
rect 396810 265384 396816 265396
rect 394752 265356 396816 265384
rect 394752 265344 394758 265356
rect 396810 265344 396816 265356
rect 396868 265344 396874 265396
rect 408586 265384 408592 265396
rect 396920 265356 408592 265384
rect 396920 265316 396948 265356
rect 408586 265344 408592 265356
rect 408644 265344 408650 265396
rect 409598 265344 409604 265396
rect 409656 265384 409662 265396
rect 435726 265384 435732 265396
rect 409656 265356 435732 265384
rect 409656 265344 409662 265356
rect 435726 265344 435732 265356
rect 435784 265344 435790 265396
rect 391906 265288 396948 265316
rect 400306 265276 400312 265328
rect 400364 265316 400370 265328
rect 467742 265316 467748 265328
rect 400364 265288 467748 265316
rect 400364 265276 400370 265288
rect 467742 265276 467748 265288
rect 467800 265276 467806 265328
rect 318334 265208 318340 265260
rect 318392 265248 318398 265260
rect 400214 265248 400220 265260
rect 318392 265220 400220 265248
rect 318392 265208 318398 265220
rect 400214 265208 400220 265220
rect 400272 265208 400278 265260
rect 42150 264732 42156 264784
rect 42208 264772 42214 264784
rect 59446 264772 59452 264784
rect 42208 264744 59452 264772
rect 42208 264732 42214 264744
rect 59446 264732 59452 264744
rect 59504 264732 59510 264784
rect 673822 263032 673828 263084
rect 673880 263072 673886 263084
rect 676030 263072 676036 263084
rect 673880 263044 676036 263072
rect 673880 263032 673886 263044
rect 676030 263032 676036 263044
rect 676088 263032 676094 263084
rect 673454 262488 673460 262540
rect 673512 262528 673518 262540
rect 676122 262528 676128 262540
rect 673512 262500 676128 262528
rect 673512 262488 673518 262500
rect 676122 262488 676128 262500
rect 676180 262488 676186 262540
rect 673546 262284 673552 262336
rect 673604 262324 673610 262336
rect 676122 262324 676128 262336
rect 673604 262296 676128 262324
rect 673604 262284 673610 262296
rect 676122 262284 676128 262296
rect 676180 262284 676186 262336
rect 674466 262216 674472 262268
rect 674524 262256 674530 262268
rect 676030 262256 676036 262268
rect 674524 262228 676036 262256
rect 674524 262216 674530 262228
rect 676030 262216 676036 262228
rect 676088 262216 676094 262268
rect 674926 261808 674932 261860
rect 674984 261848 674990 261860
rect 676030 261848 676036 261860
rect 674984 261820 676036 261848
rect 674984 261808 674990 261820
rect 676030 261808 676036 261820
rect 676088 261808 676094 261860
rect 673638 260176 673644 260228
rect 673696 260216 673702 260228
rect 675662 260216 675668 260228
rect 673696 260188 675668 260216
rect 673696 260176 673702 260188
rect 675662 260176 675668 260188
rect 675720 260176 675726 260228
rect 673730 259700 673736 259752
rect 673788 259740 673794 259752
rect 675662 259740 675668 259752
rect 673788 259712 675668 259740
rect 673788 259700 673794 259712
rect 675662 259700 675668 259712
rect 675720 259700 675726 259752
rect 674742 259632 674748 259684
rect 674800 259672 674806 259684
rect 676122 259672 676128 259684
rect 674800 259644 676128 259672
rect 674800 259632 674806 259644
rect 676122 259632 676128 259644
rect 676180 259632 676186 259684
rect 674650 259564 674656 259616
rect 674708 259604 674714 259616
rect 675938 259604 675944 259616
rect 674708 259576 675944 259604
rect 674708 259564 674714 259576
rect 675938 259564 675944 259576
rect 675996 259564 676002 259616
rect 674834 259496 674840 259548
rect 674892 259536 674898 259548
rect 676122 259536 676128 259548
rect 674892 259508 676128 259536
rect 674892 259496 674898 259508
rect 676122 259496 676128 259508
rect 676180 259496 676186 259548
rect 675018 259428 675024 259480
rect 675076 259468 675082 259480
rect 676030 259468 676036 259480
rect 675076 259440 676036 259468
rect 675076 259428 675082 259440
rect 676030 259428 676036 259440
rect 676088 259428 676094 259480
rect 674282 258952 674288 259004
rect 674340 258992 674346 259004
rect 676030 258992 676036 259004
rect 674340 258964 676036 258992
rect 674340 258952 674346 258964
rect 676030 258952 676036 258964
rect 676088 258952 676094 259004
rect 41782 258068 41788 258120
rect 41840 258108 41846 258120
rect 53926 258108 53932 258120
rect 41840 258080 53932 258108
rect 41840 258068 41846 258080
rect 53926 258068 53932 258080
rect 53984 258068 53990 258120
rect 41506 257932 41512 257984
rect 41564 257972 41570 257984
rect 51074 257972 51080 257984
rect 41564 257944 51080 257972
rect 41564 257932 41570 257944
rect 51074 257932 51080 257944
rect 51132 257932 51138 257984
rect 41506 257524 41512 257576
rect 41564 257564 41570 257576
rect 46106 257564 46112 257576
rect 41564 257536 46112 257564
rect 41564 257524 41570 257536
rect 46106 257524 46112 257536
rect 46164 257524 46170 257576
rect 672626 256776 672632 256828
rect 672684 256816 672690 256828
rect 678974 256816 678980 256828
rect 672684 256788 678980 256816
rect 672684 256776 672690 256788
rect 678974 256776 678980 256788
rect 679032 256776 679038 256828
rect 52270 256708 52276 256760
rect 52328 256748 52334 256760
rect 184934 256748 184940 256760
rect 52328 256720 184940 256748
rect 52328 256708 52334 256720
rect 184934 256708 184940 256720
rect 184992 256708 184998 256760
rect 674558 256708 674564 256760
rect 674616 256748 674622 256760
rect 676030 256748 676036 256760
rect 674616 256720 676036 256748
rect 674616 256708 674622 256720
rect 676030 256708 676036 256720
rect 676088 256708 676094 256760
rect 673546 252696 673552 252748
rect 673604 252696 673610 252748
rect 673564 252544 673592 252696
rect 673546 252492 673552 252544
rect 673604 252492 673610 252544
rect 673730 252288 673736 252340
rect 673788 252328 673794 252340
rect 674282 252328 674288 252340
rect 673788 252300 674288 252328
rect 673788 252288 673794 252300
rect 674282 252288 674288 252300
rect 674340 252288 674346 252340
rect 674282 252152 674288 252204
rect 674340 252192 674346 252204
rect 674558 252192 674564 252204
rect 674340 252164 674564 252192
rect 674340 252152 674346 252164
rect 674558 252152 674564 252164
rect 674616 252152 674622 252204
rect 674650 251880 674656 251932
rect 674708 251920 674714 251932
rect 674834 251920 674840 251932
rect 674708 251892 674840 251920
rect 674708 251880 674714 251892
rect 674834 251880 674840 251892
rect 674892 251880 674898 251932
rect 675662 251336 675668 251388
rect 675720 251336 675726 251388
rect 675754 251336 675760 251388
rect 675812 251336 675818 251388
rect 416774 251200 416780 251252
rect 416832 251240 416838 251252
rect 567102 251240 567108 251252
rect 416832 251212 567108 251240
rect 416832 251200 416838 251212
rect 567102 251200 567108 251212
rect 567160 251200 567166 251252
rect 674742 251200 674748 251252
rect 674800 251240 674806 251252
rect 675294 251240 675300 251252
rect 674800 251212 675300 251240
rect 674800 251200 674806 251212
rect 675294 251200 675300 251212
rect 675352 251200 675358 251252
rect 675294 250928 675300 250980
rect 675352 250968 675358 250980
rect 675680 250968 675708 251336
rect 675352 250940 675708 250968
rect 675352 250928 675358 250940
rect 675772 250776 675800 251336
rect 675754 250724 675760 250776
rect 675812 250724 675818 250776
rect 675018 250180 675024 250232
rect 675076 250220 675082 250232
rect 675478 250220 675484 250232
rect 675076 250192 675484 250220
rect 675076 250180 675082 250192
rect 675478 250180 675484 250192
rect 675536 250180 675542 250232
rect 675018 249772 675024 249824
rect 675076 249812 675082 249824
rect 675294 249812 675300 249824
rect 675076 249784 675300 249812
rect 675076 249772 675082 249784
rect 675294 249772 675300 249784
rect 675352 249772 675358 249824
rect 674466 249636 674472 249688
rect 674524 249676 674530 249688
rect 675294 249676 675300 249688
rect 674524 249648 675300 249676
rect 674524 249636 674530 249648
rect 675294 249636 675300 249648
rect 675352 249636 675358 249688
rect 673822 249568 673828 249620
rect 673880 249608 673886 249620
rect 675386 249608 675392 249620
rect 673880 249580 675392 249608
rect 673880 249568 673886 249580
rect 675386 249568 675392 249580
rect 675444 249568 675450 249620
rect 673362 249500 673368 249552
rect 673420 249540 673426 249552
rect 674466 249540 674472 249552
rect 673420 249512 674472 249540
rect 673420 249500 673426 249512
rect 674466 249500 674472 249512
rect 674524 249500 674530 249552
rect 416774 248412 416780 248464
rect 416832 248452 416838 248464
rect 564342 248452 564348 248464
rect 416832 248424 564348 248452
rect 416832 248412 416838 248424
rect 564342 248412 564348 248424
rect 564400 248412 564406 248464
rect 41414 247664 41420 247716
rect 41472 247704 41478 247716
rect 45646 247704 45652 247716
rect 41472 247676 45652 247704
rect 41472 247664 41478 247676
rect 45646 247664 45652 247676
rect 45704 247664 45710 247716
rect 674834 247256 674840 247308
rect 674892 247296 674898 247308
rect 675386 247296 675392 247308
rect 674892 247268 675392 247296
rect 674892 247256 674898 247268
rect 675386 247256 675392 247268
rect 675444 247256 675450 247308
rect 674926 246984 674932 247036
rect 674984 247024 674990 247036
rect 675202 247024 675208 247036
rect 674984 246996 675208 247024
rect 674984 246984 674990 246996
rect 675202 246984 675208 246996
rect 675260 246984 675266 247036
rect 41506 246916 41512 246968
rect 41564 246956 41570 246968
rect 43346 246956 43352 246968
rect 41564 246928 43352 246956
rect 41564 246916 41570 246928
rect 43346 246916 43352 246928
rect 43404 246916 43410 246968
rect 674558 246508 674564 246560
rect 674616 246548 674622 246560
rect 675386 246548 675392 246560
rect 674616 246520 675392 246548
rect 674616 246508 674622 246520
rect 675386 246508 675392 246520
rect 675444 246508 675450 246560
rect 674650 246032 674656 246084
rect 674708 246072 674714 246084
rect 675386 246072 675392 246084
rect 674708 246044 675392 246072
rect 674708 246032 674714 246044
rect 675386 246032 675392 246044
rect 675444 246032 675450 246084
rect 20714 245828 20720 245880
rect 20772 245868 20778 245880
rect 30098 245868 30104 245880
rect 20772 245840 30104 245868
rect 20772 245828 20778 245840
rect 30098 245828 30104 245840
rect 30156 245828 30162 245880
rect 52178 245760 52184 245812
rect 52236 245800 52242 245812
rect 184934 245800 184940 245812
rect 52236 245772 184940 245800
rect 52236 245760 52242 245772
rect 184934 245760 184940 245772
rect 184992 245760 184998 245812
rect 41506 245692 41512 245744
rect 41564 245732 41570 245744
rect 56686 245732 56692 245744
rect 41564 245704 56692 245732
rect 41564 245692 41570 245704
rect 56686 245692 56692 245704
rect 56744 245692 56750 245744
rect 41414 245624 41420 245676
rect 41472 245664 41478 245676
rect 56594 245664 56600 245676
rect 41472 245636 56600 245664
rect 41472 245624 41478 245636
rect 56594 245624 56600 245636
rect 56652 245624 56658 245676
rect 416774 245624 416780 245676
rect 416832 245664 416838 245676
rect 564526 245664 564532 245676
rect 416832 245636 564532 245664
rect 416832 245624 416838 245636
rect 564526 245624 564532 245636
rect 564584 245624 564590 245676
rect 43254 245556 43260 245608
rect 43312 245596 43318 245608
rect 43312 245568 43484 245596
rect 43312 245556 43318 245568
rect 43456 245540 43484 245568
rect 655606 245556 655612 245608
rect 655664 245596 655670 245608
rect 675294 245596 675300 245608
rect 655664 245568 675300 245596
rect 655664 245556 655670 245568
rect 675294 245556 675300 245568
rect 675352 245556 675358 245608
rect 43438 245488 43444 245540
rect 43496 245488 43502 245540
rect 38102 245420 38108 245472
rect 38160 245460 38166 245472
rect 43254 245460 43260 245472
rect 38160 245432 43260 245460
rect 38160 245420 38166 245432
rect 43254 245420 43260 245432
rect 43312 245420 43318 245472
rect 674282 245420 674288 245472
rect 674340 245460 674346 245472
rect 675294 245460 675300 245472
rect 674340 245432 675300 245460
rect 674340 245420 674346 245432
rect 675294 245420 675300 245432
rect 675352 245420 675358 245472
rect 38194 245352 38200 245404
rect 38252 245392 38258 245404
rect 43070 245392 43076 245404
rect 38252 245364 43076 245392
rect 38252 245352 38258 245364
rect 43070 245352 43076 245364
rect 43128 245352 43134 245404
rect 43714 244808 43720 244860
rect 43772 244848 43778 244860
rect 43898 244848 43904 244860
rect 43772 244820 43904 244848
rect 43772 244808 43778 244820
rect 43898 244808 43904 244820
rect 43956 244808 43962 244860
rect 43438 244672 43444 244724
rect 43496 244712 43502 244724
rect 43714 244712 43720 244724
rect 43496 244684 43720 244712
rect 43496 244672 43502 244684
rect 43714 244672 43720 244684
rect 43772 244672 43778 244724
rect 42334 244536 42340 244588
rect 42392 244576 42398 244588
rect 43438 244576 43444 244588
rect 42392 244548 43444 244576
rect 42392 244536 42398 244548
rect 43438 244536 43444 244548
rect 43496 244536 43502 244588
rect 20714 244332 20720 244384
rect 20772 244372 20778 244384
rect 42242 244372 42248 244384
rect 20772 244344 42248 244372
rect 20772 244332 20778 244344
rect 42242 244332 42248 244344
rect 42300 244332 42306 244384
rect 673546 243584 673552 243636
rect 673604 243624 673610 243636
rect 675386 243624 675392 243636
rect 673604 243596 675392 243624
rect 673604 243584 673610 243596
rect 675386 243584 675392 243596
rect 675444 243584 675450 243636
rect 673730 242904 673736 242956
rect 673788 242944 673794 242956
rect 675386 242944 675392 242956
rect 673788 242916 675392 242944
rect 673788 242904 673794 242916
rect 675386 242904 675392 242916
rect 675444 242904 675450 242956
rect 673638 242156 673644 242208
rect 673696 242196 673702 242208
rect 675386 242196 675392 242208
rect 673696 242168 675392 242196
rect 673696 242156 673702 242168
rect 675386 242156 675392 242168
rect 675444 242156 675450 242208
rect 673454 241068 673460 241120
rect 673512 241108 673518 241120
rect 675294 241108 675300 241120
rect 673512 241080 675300 241108
rect 673512 241068 673518 241080
rect 675294 241068 675300 241080
rect 675352 241068 675358 241120
rect 674466 239912 674472 239964
rect 674524 239952 674530 239964
rect 675294 239952 675300 239964
rect 674524 239924 675300 239952
rect 674524 239912 674530 239924
rect 675294 239912 675300 239924
rect 675352 239912 675358 239964
rect 42242 239708 42248 239760
rect 42300 239748 42306 239760
rect 42702 239748 42708 239760
rect 42300 239720 42708 239748
rect 42300 239708 42306 239720
rect 42702 239708 42708 239720
rect 42760 239708 42766 239760
rect 42150 238484 42156 238536
rect 42208 238524 42214 238536
rect 43806 238524 43812 238536
rect 42208 238496 43812 238524
rect 42208 238484 42214 238496
rect 43806 238484 43812 238496
rect 43864 238484 43870 238536
rect 184934 237436 184940 237448
rect 184806 237408 184940 237436
rect 42242 236036 42248 236088
rect 42300 236076 42306 236088
rect 43070 236076 43076 236088
rect 42300 236048 43076 236076
rect 42300 236036 42306 236048
rect 43070 236036 43076 236048
rect 43128 236036 43134 236088
rect 42150 235356 42156 235408
rect 42208 235396 42214 235408
rect 43346 235396 43352 235408
rect 42208 235368 43352 235396
rect 42208 235356 42214 235368
rect 43346 235356 43352 235368
rect 43404 235356 43410 235408
rect 42150 234608 42156 234660
rect 42208 234648 42214 234660
rect 43162 234648 43168 234660
rect 42208 234620 43168 234648
rect 42208 234608 42214 234620
rect 43162 234608 43168 234620
rect 43220 234608 43226 234660
rect 42242 233520 42248 233572
rect 42300 233560 42306 233572
rect 43254 233560 43260 233572
rect 42300 233532 43260 233560
rect 42300 233520 42306 233532
rect 43254 233520 43260 233532
rect 43312 233520 43318 233572
rect 42150 233316 42156 233368
rect 42208 233356 42214 233368
rect 43530 233356 43536 233368
rect 42208 233328 43536 233356
rect 42208 233316 42214 233328
rect 43530 233316 43536 233328
rect 43588 233316 43594 233368
rect 52086 230796 52092 230848
rect 52144 230836 52150 230848
rect 184806 230836 184834 237408
rect 184934 237396 184940 237408
rect 184992 237396 184998 237448
rect 674926 235560 674932 235612
rect 674984 235600 674990 235612
rect 675754 235600 675760 235612
rect 674984 235572 675760 235600
rect 674984 235560 674990 235572
rect 675754 235560 675760 235572
rect 675812 235560 675818 235612
rect 674742 235492 674748 235544
rect 674800 235532 674806 235544
rect 675662 235532 675668 235544
rect 674800 235504 675668 235532
rect 674800 235492 674806 235504
rect 675662 235492 675668 235504
rect 675720 235492 675726 235544
rect 345934 231140 345940 231192
rect 345992 231180 345998 231192
rect 414014 231180 414020 231192
rect 345992 231152 414020 231180
rect 345992 231140 345998 231152
rect 414014 231140 414020 231152
rect 414072 231140 414078 231192
rect 355870 231072 355876 231124
rect 355928 231112 355934 231124
rect 437290 231112 437296 231124
rect 355928 231084 437296 231112
rect 355928 231072 355934 231084
rect 437290 231072 437296 231084
rect 437348 231072 437354 231124
rect 347314 231004 347320 231056
rect 347372 231044 347378 231056
rect 417142 231044 417148 231056
rect 347372 231016 417148 231044
rect 347372 231004 347378 231016
rect 417142 231004 417148 231016
rect 417200 231004 417206 231056
rect 356238 230936 356244 230988
rect 356296 230976 356302 230988
rect 439774 230976 439780 230988
rect 356296 230948 439780 230976
rect 356296 230936 356302 230948
rect 439774 230936 439780 230948
rect 439832 230936 439838 230988
rect 348786 230868 348792 230920
rect 348844 230908 348850 230920
rect 420454 230908 420460 230920
rect 348844 230880 420460 230908
rect 348844 230868 348850 230880
rect 420454 230868 420460 230880
rect 420512 230868 420518 230920
rect 52144 230808 184834 230836
rect 52144 230796 52150 230808
rect 351638 230800 351644 230852
rect 351696 230840 351702 230852
rect 427170 230840 427176 230852
rect 351696 230812 427176 230840
rect 351696 230800 351702 230812
rect 427170 230800 427176 230812
rect 427228 230800 427234 230852
rect 354490 230732 354496 230784
rect 354548 230772 354554 230784
rect 433886 230772 433892 230784
rect 354548 230744 433892 230772
rect 354548 230732 354554 230744
rect 433886 230732 433892 230744
rect 433944 230732 433950 230784
rect 45922 230664 45928 230716
rect 45980 230704 45986 230716
rect 656894 230704 656900 230716
rect 45980 230676 656900 230704
rect 45980 230664 45986 230676
rect 656894 230664 656900 230676
rect 656952 230664 656958 230716
rect 46198 230596 46204 230648
rect 46256 230636 46262 230648
rect 659746 230636 659752 230648
rect 46256 230608 659752 230636
rect 46256 230596 46262 230608
rect 659746 230596 659752 230608
rect 659804 230596 659810 230648
rect 42242 230528 42248 230580
rect 42300 230568 42306 230580
rect 43714 230568 43720 230580
rect 42300 230540 43720 230568
rect 42300 230528 42306 230540
rect 43714 230528 43720 230540
rect 43772 230528 43778 230580
rect 46014 230528 46020 230580
rect 46072 230568 46078 230580
rect 659654 230568 659660 230580
rect 46072 230540 659660 230568
rect 46072 230528 46078 230540
rect 659654 230528 659660 230540
rect 659712 230528 659718 230580
rect 45646 230460 45652 230512
rect 45704 230500 45710 230512
rect 662782 230500 662788 230512
rect 45704 230472 662788 230500
rect 45704 230460 45710 230472
rect 662782 230460 662788 230472
rect 662840 230460 662846 230512
rect 42150 230324 42156 230376
rect 42208 230364 42214 230376
rect 43990 230364 43996 230376
rect 42208 230336 43996 230364
rect 42208 230324 42214 230336
rect 43990 230324 43996 230336
rect 44048 230324 44054 230376
rect 359090 230324 359096 230376
rect 359148 230364 359154 230376
rect 446582 230364 446588 230376
rect 359148 230336 446588 230364
rect 359148 230324 359154 230336
rect 446582 230324 446588 230336
rect 446640 230324 446646 230376
rect 357710 230256 357716 230308
rect 357768 230296 357774 230308
rect 443178 230296 443184 230308
rect 357768 230268 443184 230296
rect 357768 230256 357774 230268
rect 443178 230256 443184 230268
rect 443236 230256 443242 230308
rect 363046 230188 363052 230240
rect 363104 230228 363110 230240
rect 454126 230228 454132 230240
rect 363104 230200 454132 230228
rect 363104 230188 363110 230200
rect 454126 230188 454132 230200
rect 454184 230188 454190 230240
rect 361942 230120 361948 230172
rect 362000 230160 362006 230172
rect 453298 230160 453304 230172
rect 362000 230132 453304 230160
rect 362000 230120 362006 230132
rect 453298 230120 453304 230132
rect 453356 230120 453362 230172
rect 360562 230052 360568 230104
rect 360620 230092 360626 230104
rect 449894 230092 449900 230104
rect 360620 230064 449900 230092
rect 360620 230052 360626 230064
rect 449894 230052 449900 230064
rect 449952 230052 449958 230104
rect 364794 229984 364800 230036
rect 364852 230024 364858 230036
rect 460014 230024 460020 230036
rect 364852 229996 460020 230024
rect 364852 229984 364858 229996
rect 460014 229984 460020 229996
rect 460072 229984 460078 230036
rect 363414 229916 363420 229968
rect 363472 229956 363478 229968
rect 456610 229956 456616 229968
rect 363472 229928 456616 229956
rect 363472 229916 363478 229928
rect 456610 229916 456616 229928
rect 456668 229916 456674 229968
rect 42150 229848 42156 229900
rect 42208 229888 42214 229900
rect 43898 229888 43904 229900
rect 42208 229860 43904 229888
rect 42208 229848 42214 229860
rect 43898 229848 43904 229860
rect 43956 229848 43962 229900
rect 364058 229848 364064 229900
rect 364116 229888 364122 229900
rect 455782 229888 455788 229900
rect 364116 229860 455788 229888
rect 364116 229848 364122 229860
rect 455782 229848 455788 229860
rect 455840 229848 455846 229900
rect 366910 229780 366916 229832
rect 366968 229820 366974 229832
rect 462498 229820 462504 229832
rect 366968 229792 462504 229820
rect 366968 229780 366974 229792
rect 462498 229780 462504 229792
rect 462556 229780 462562 229832
rect 366266 229712 366272 229764
rect 366324 229752 366330 229764
rect 463694 229752 463700 229764
rect 366324 229724 463700 229752
rect 366324 229712 366330 229724
rect 463694 229712 463700 229724
rect 463752 229712 463758 229764
rect 372614 229644 372620 229696
rect 372672 229684 372678 229696
rect 476022 229684 476028 229696
rect 372672 229656 476028 229684
rect 372672 229644 372678 229656
rect 476022 229644 476028 229656
rect 476080 229644 476086 229696
rect 370498 229576 370504 229628
rect 370556 229616 370562 229628
rect 473446 229616 473452 229628
rect 370556 229588 473452 229616
rect 370556 229576 370562 229588
rect 473446 229576 473452 229588
rect 473504 229576 473510 229628
rect 369118 229508 369124 229560
rect 369176 229548 369182 229560
rect 470134 229548 470140 229560
rect 369176 229520 470140 229548
rect 369176 229508 369182 229520
rect 470134 229508 470140 229520
rect 470192 229508 470198 229560
rect 371234 229440 371240 229492
rect 371292 229480 371298 229492
rect 472618 229480 472624 229492
rect 371292 229452 472624 229480
rect 371292 229440 371298 229452
rect 472618 229440 472624 229452
rect 472676 229440 472682 229492
rect 373350 229372 373356 229424
rect 373408 229412 373414 229424
rect 480346 229412 480352 229424
rect 373408 229384 480352 229412
rect 373408 229372 373414 229384
rect 480346 229372 480352 229384
rect 480404 229372 480410 229424
rect 374822 229304 374828 229356
rect 374880 229344 374886 229356
rect 483014 229344 483020 229356
rect 374880 229316 483020 229344
rect 374880 229304 374886 229316
rect 483014 229304 483020 229316
rect 483072 229304 483078 229356
rect 376202 229236 376208 229288
rect 376260 229276 376266 229288
rect 487154 229276 487160 229288
rect 376260 229248 487160 229276
rect 376260 229236 376266 229248
rect 487154 229236 487160 229248
rect 487212 229236 487218 229288
rect 393682 229168 393688 229220
rect 393740 229208 393746 229220
rect 528370 229208 528376 229220
rect 393740 229180 528376 229208
rect 393740 229168 393746 229180
rect 528370 229168 528376 229180
rect 528428 229168 528434 229220
rect 396902 229100 396908 229152
rect 396960 229140 396966 229152
rect 536650 229140 536656 229152
rect 396960 229112 536656 229140
rect 396960 229100 396966 229112
rect 536650 229100 536656 229112
rect 536708 229100 536714 229152
rect 158714 229032 158720 229084
rect 158772 229072 158778 229084
rect 237558 229072 237564 229084
rect 158772 229044 237564 229072
rect 158772 229032 158778 229044
rect 237558 229032 237564 229044
rect 237616 229032 237622 229084
rect 246206 229032 246212 229084
rect 246264 229072 246270 229084
rect 258534 229072 258540 229084
rect 246264 229044 258540 229072
rect 246264 229032 246270 229044
rect 258534 229032 258540 229044
rect 258592 229032 258598 229084
rect 296346 229032 296352 229084
rect 296404 229072 296410 229084
rect 298462 229072 298468 229084
rect 296404 229044 298468 229072
rect 296404 229032 296410 229044
rect 298462 229032 298468 229044
rect 298520 229032 298526 229084
rect 298830 229032 298836 229084
rect 298888 229072 298894 229084
rect 302694 229072 302700 229084
rect 298888 229044 302700 229072
rect 298888 229032 298894 229044
rect 302694 229032 302700 229044
rect 302752 229032 302758 229084
rect 304166 229032 304172 229084
rect 304224 229072 304230 229084
rect 314654 229072 314660 229084
rect 304224 229044 314660 229072
rect 304224 229032 304230 229044
rect 314654 229032 314660 229044
rect 314712 229032 314718 229084
rect 339126 229032 339132 229084
rect 339184 229072 339190 229084
rect 377030 229072 377036 229084
rect 339184 229044 377036 229072
rect 339184 229032 339190 229044
rect 377030 229032 377036 229044
rect 377088 229032 377094 229084
rect 397362 229072 397368 229084
rect 391906 229044 397368 229072
rect 152826 228964 152832 229016
rect 152884 229004 152890 229016
rect 233970 229004 233976 229016
rect 152884 228976 233976 229004
rect 152884 228964 152890 228976
rect 233970 228964 233976 228976
rect 234028 228964 234034 229016
rect 243538 228964 243544 229016
rect 243596 229004 243602 229016
rect 272426 229004 272432 229016
rect 243596 228976 272432 229004
rect 243596 228964 243602 228976
rect 272426 228964 272432 228976
rect 272484 228964 272490 229016
rect 293218 228964 293224 229016
rect 293276 229004 293282 229016
rect 294598 229004 294604 229016
rect 293276 228976 294604 229004
rect 293276 228964 293282 228976
rect 294598 228964 294604 228976
rect 294656 228964 294662 229016
rect 297450 228964 297456 229016
rect 297508 229004 297514 229016
rect 299382 229004 299388 229016
rect 297508 228976 299388 229004
rect 297508 228964 297514 228976
rect 299382 228964 299388 228976
rect 299440 228964 299446 229016
rect 303522 228964 303528 229016
rect 303580 229004 303586 229016
rect 315298 229004 315304 229016
rect 303580 228976 315304 229004
rect 303580 228964 303586 228976
rect 315298 228964 315304 228976
rect 315356 228964 315362 229016
rect 318794 228964 318800 229016
rect 318852 229004 318858 229016
rect 340966 229004 340972 229016
rect 318852 228976 340972 229004
rect 318852 228964 318858 228976
rect 340966 228964 340972 228976
rect 341024 228964 341030 229016
rect 342346 228964 342352 229016
rect 342404 229004 342410 229016
rect 380894 229004 380900 229016
rect 342404 228976 380900 229004
rect 342404 228964 342410 228976
rect 380894 228964 380900 228976
rect 380952 228964 380958 229016
rect 388346 228964 388352 229016
rect 388404 229004 388410 229016
rect 391906 229004 391934 229044
rect 397362 229032 397368 229044
rect 397420 229032 397426 229084
rect 401502 229032 401508 229084
rect 401560 229072 401566 229084
rect 458174 229072 458180 229084
rect 401560 229044 458180 229072
rect 401560 229032 401566 229044
rect 458174 229032 458180 229044
rect 458232 229032 458238 229084
rect 388404 228976 391934 229004
rect 388404 228964 388410 228976
rect 392118 228964 392124 229016
rect 392176 229004 392182 229016
rect 467006 229004 467012 229016
rect 392176 228976 467012 229004
rect 392176 228964 392182 228976
rect 467006 228964 467012 228976
rect 467064 228964 467070 229016
rect 156966 228896 156972 228948
rect 157024 228936 157030 228948
rect 237190 228936 237196 228948
rect 157024 228908 237196 228936
rect 157024 228896 157030 228908
rect 237190 228896 237196 228908
rect 237248 228896 237254 228948
rect 241238 228896 241244 228948
rect 241296 228936 241302 228948
rect 269574 228936 269580 228948
rect 241296 228908 269580 228936
rect 241296 228896 241302 228908
rect 269574 228896 269580 228908
rect 269632 228896 269638 228948
rect 296714 228896 296720 228948
rect 296772 228936 296778 228948
rect 300210 228936 300216 228948
rect 296772 228908 300216 228936
rect 296772 228896 296778 228908
rect 300210 228896 300216 228908
rect 300268 228896 300274 228948
rect 304534 228896 304540 228948
rect 304592 228936 304598 228948
rect 316126 228936 316132 228948
rect 304592 228908 316132 228936
rect 304592 228896 304598 228908
rect 316126 228896 316132 228908
rect 316184 228896 316190 228948
rect 336274 228896 336280 228948
rect 336332 228936 336338 228948
rect 378502 228936 378508 228948
rect 336332 228908 378508 228936
rect 336332 228896 336338 228908
rect 378502 228896 378508 228908
rect 378560 228896 378566 228948
rect 389726 228896 389732 228948
rect 389784 228936 389790 228948
rect 464430 228936 464436 228948
rect 389784 228908 464436 228936
rect 389784 228896 389790 228908
rect 464430 228896 464436 228908
rect 464488 228896 464494 228948
rect 150250 228828 150256 228880
rect 150308 228868 150314 228880
rect 234338 228868 234344 228880
rect 150308 228840 234344 228868
rect 150308 228828 150314 228840
rect 234338 228828 234344 228840
rect 234396 228828 234402 228880
rect 239766 228828 239772 228880
rect 239824 228868 239830 228880
rect 266722 228868 266728 228880
rect 239824 228840 266728 228868
rect 239824 228828 239830 228840
rect 266722 228828 266728 228840
rect 266780 228828 266786 228880
rect 308490 228828 308496 228880
rect 308548 228868 308554 228880
rect 324590 228868 324596 228880
rect 308548 228840 324596 228868
rect 308548 228828 308554 228840
rect 324590 228828 324596 228840
rect 324648 228828 324654 228880
rect 340874 228828 340880 228880
rect 340932 228868 340938 228880
rect 383746 228868 383752 228880
rect 340932 228840 383752 228868
rect 340932 228828 340938 228840
rect 383746 228828 383752 228840
rect 383804 228828 383810 228880
rect 387242 228828 387248 228880
rect 387300 228868 387306 228880
rect 401502 228868 401508 228880
rect 387300 228840 401508 228868
rect 387300 228828 387306 228840
rect 401502 228828 401508 228840
rect 401560 228828 401566 228880
rect 469950 228868 469956 228880
rect 402624 228840 469956 228868
rect 151722 228760 151728 228812
rect 151780 228800 151786 228812
rect 234706 228800 234712 228812
rect 151780 228772 234712 228800
rect 151780 228760 151786 228772
rect 234706 228760 234712 228772
rect 234764 228760 234770 228812
rect 239950 228760 239956 228812
rect 240008 228800 240014 228812
rect 265342 228800 265348 228812
rect 240008 228772 265348 228800
rect 240008 228760 240014 228772
rect 265342 228760 265348 228772
rect 265400 228760 265406 228812
rect 305638 228760 305644 228812
rect 305696 228800 305702 228812
rect 317874 228800 317880 228812
rect 305696 228772 317880 228800
rect 305696 228760 305702 228772
rect 317874 228760 317880 228772
rect 317932 228760 317938 228812
rect 340598 228760 340604 228812
rect 340656 228800 340662 228812
rect 391750 228800 391756 228812
rect 340656 228772 391756 228800
rect 340656 228760 340662 228772
rect 391750 228760 391756 228772
rect 391808 228760 391814 228812
rect 394050 228760 394056 228812
rect 394108 228800 394114 228812
rect 402624 228800 402652 228840
rect 469950 228828 469956 228840
rect 470008 228828 470014 228880
rect 394108 228772 402652 228800
rect 394108 228760 394114 228772
rect 403342 228760 403348 228812
rect 403400 228800 403406 228812
rect 416774 228800 416780 228812
rect 403400 228772 416780 228800
rect 403400 228760 403406 228772
rect 416774 228760 416780 228772
rect 416832 228760 416838 228812
rect 416866 228760 416872 228812
rect 416924 228800 416930 228812
rect 477494 228800 477500 228812
rect 416924 228772 477500 228800
rect 416924 228760 416930 228772
rect 477494 228760 477500 228772
rect 477552 228760 477558 228812
rect 146018 228692 146024 228744
rect 146076 228732 146082 228744
rect 231118 228732 231124 228744
rect 146076 228704 231124 228732
rect 146076 228692 146082 228704
rect 231118 228692 231124 228704
rect 231176 228692 231182 228744
rect 241974 228692 241980 228744
rect 242032 228732 242038 228744
rect 272150 228732 272156 228744
rect 242032 228704 272156 228732
rect 242032 228692 242038 228704
rect 272150 228692 272156 228704
rect 272208 228692 272214 228744
rect 306650 228692 306656 228744
rect 306708 228732 306714 228744
rect 323854 228732 323860 228744
rect 306708 228704 323860 228732
rect 306708 228692 306714 228704
rect 323854 228692 323860 228704
rect 323912 228692 323918 228744
rect 337746 228692 337752 228744
rect 337804 228732 337810 228744
rect 389082 228732 389088 228744
rect 337804 228704 389088 228732
rect 337804 228692 337810 228704
rect 389082 228692 389088 228704
rect 389140 228692 389146 228744
rect 396166 228692 396172 228744
rect 396224 228732 396230 228744
rect 473262 228732 473268 228744
rect 396224 228704 473268 228732
rect 396224 228692 396230 228704
rect 473262 228692 473268 228704
rect 473320 228692 473326 228744
rect 138474 228624 138480 228676
rect 138532 228664 138538 228676
rect 229002 228664 229008 228676
rect 138532 228636 229008 228664
rect 138532 228624 138538 228636
rect 229002 228624 229008 228636
rect 229060 228624 229066 228676
rect 245286 228624 245292 228676
rect 245344 228664 245350 228676
rect 273530 228664 273536 228676
rect 245344 228636 273536 228664
rect 245344 228624 245350 228636
rect 273530 228624 273536 228636
rect 273588 228624 273594 228676
rect 304902 228624 304908 228676
rect 304960 228664 304966 228676
rect 318702 228664 318708 228676
rect 304960 228636 318708 228664
rect 304960 228624 304966 228636
rect 318702 228624 318708 228636
rect 318760 228624 318766 228676
rect 323486 228624 323492 228676
rect 323544 228664 323550 228676
rect 362402 228664 362408 228676
rect 323544 228636 362408 228664
rect 323544 228624 323550 228636
rect 362402 228624 362408 228636
rect 362460 228624 362466 228676
rect 376570 228624 376576 228676
rect 376628 228664 376634 228676
rect 460934 228664 460940 228676
rect 376628 228636 460940 228664
rect 376628 228624 376634 228636
rect 460934 228624 460940 228636
rect 460992 228624 460998 228676
rect 143442 228556 143448 228608
rect 143500 228596 143506 228608
rect 231486 228596 231492 228608
rect 143500 228568 231492 228596
rect 143500 228556 143506 228568
rect 231486 228556 231492 228568
rect 231544 228556 231550 228608
rect 239858 228556 239864 228608
rect 239916 228596 239922 228608
rect 268194 228596 268200 228608
rect 239916 228568 268200 228596
rect 239916 228556 239922 228568
rect 268194 228556 268200 228568
rect 268252 228556 268258 228608
rect 307386 228556 307392 228608
rect 307444 228596 307450 228608
rect 322934 228596 322940 228608
rect 307444 228568 322940 228596
rect 307444 228556 307450 228568
rect 322934 228556 322940 228568
rect 322992 228556 322998 228608
rect 336642 228556 336648 228608
rect 336700 228596 336706 228608
rect 375282 228596 375288 228608
rect 336700 228568 375288 228596
rect 336700 228556 336706 228568
rect 375282 228556 375288 228568
rect 375340 228556 375346 228608
rect 377950 228556 377956 228608
rect 378008 228596 378014 228608
rect 474734 228596 474740 228608
rect 378008 228568 474740 228596
rect 378008 228556 378014 228568
rect 474734 228556 474740 228568
rect 474792 228556 474798 228608
rect 145190 228488 145196 228540
rect 145248 228528 145254 228540
rect 231854 228528 231860 228540
rect 145248 228500 231860 228528
rect 145248 228488 145254 228500
rect 231854 228488 231860 228500
rect 231912 228488 231918 228540
rect 240134 228488 240140 228540
rect 240192 228528 240198 228540
rect 271046 228528 271052 228540
rect 240192 228500 271052 228528
rect 240192 228488 240198 228500
rect 271046 228488 271052 228500
rect 271104 228488 271110 228540
rect 308858 228488 308864 228540
rect 308916 228528 308922 228540
rect 326246 228528 326252 228540
rect 308916 228500 326252 228528
rect 308916 228488 308922 228500
rect 326246 228488 326252 228500
rect 326304 228488 326310 228540
rect 335170 228488 335176 228540
rect 335228 228528 335234 228540
rect 373994 228528 374000 228540
rect 335228 228500 374000 228528
rect 335228 228488 335234 228500
rect 373994 228488 374000 228500
rect 374052 228488 374058 228540
rect 375466 228488 375472 228540
rect 375524 228528 375530 228540
rect 480254 228528 480260 228540
rect 375524 228500 480260 228528
rect 375524 228488 375530 228500
rect 480254 228488 480260 228500
rect 480312 228488 480318 228540
rect 136818 228420 136824 228472
rect 136876 228460 136882 228472
rect 228634 228460 228640 228472
rect 136876 228432 228640 228460
rect 136876 228420 136882 228432
rect 228634 228420 228640 228432
rect 228692 228420 228698 228472
rect 238570 228420 238576 228472
rect 238628 228460 238634 228472
rect 270678 228460 270684 228472
rect 238628 228432 270684 228460
rect 238628 228420 238634 228432
rect 270678 228420 270684 228432
rect 270736 228420 270742 228472
rect 307754 228420 307760 228472
rect 307812 228460 307818 228472
rect 325694 228460 325700 228472
rect 307812 228432 325700 228460
rect 307812 228420 307818 228432
rect 325694 228420 325700 228432
rect 325752 228420 325758 228472
rect 332042 228420 332048 228472
rect 332100 228460 332106 228472
rect 376846 228460 376852 228472
rect 332100 228432 376852 228460
rect 332100 228420 332106 228432
rect 376846 228420 376852 228432
rect 376904 228420 376910 228472
rect 379422 228420 379428 228472
rect 379480 228460 379486 228472
rect 494514 228460 494520 228472
rect 379480 228432 494520 228460
rect 379480 228420 379486 228432
rect 494514 228420 494520 228432
rect 494572 228420 494578 228472
rect 131758 228352 131764 228404
rect 131816 228392 131822 228404
rect 226150 228392 226156 228404
rect 131816 228364 226156 228392
rect 131816 228352 131822 228364
rect 226150 228352 226156 228364
rect 226208 228352 226214 228404
rect 235258 228352 235264 228404
rect 235316 228392 235322 228404
rect 269298 228392 269304 228404
rect 235316 228364 269304 228392
rect 235316 228352 235322 228364
rect 269298 228352 269304 228364
rect 269356 228352 269362 228404
rect 302786 228352 302792 228404
rect 302844 228392 302850 228404
rect 311158 228392 311164 228404
rect 302844 228364 311164 228392
rect 302844 228352 302850 228364
rect 311158 228352 311164 228364
rect 311216 228352 311222 228404
rect 317414 228352 317420 228404
rect 317472 228392 317478 228404
rect 317472 228364 329144 228392
rect 317472 228352 317478 228364
rect 125042 228284 125048 228336
rect 125100 228324 125106 228336
rect 223298 228324 223304 228336
rect 125100 228296 223304 228324
rect 125100 228284 125106 228296
rect 223298 228284 223304 228296
rect 223356 228284 223362 228336
rect 229278 228284 229284 228336
rect 229336 228324 229342 228336
rect 267458 228324 267464 228336
rect 229336 228296 267464 228324
rect 229336 228284 229342 228296
rect 267458 228284 267464 228296
rect 267516 228284 267522 228336
rect 308122 228284 308128 228336
rect 308180 228324 308186 228336
rect 327074 228324 327080 228336
rect 308180 228296 327080 228324
rect 308180 228284 308186 228296
rect 327074 228284 327080 228296
rect 327132 228284 327138 228336
rect 130102 228216 130108 228268
rect 130160 228256 130166 228268
rect 225782 228256 225788 228268
rect 130160 228228 225788 228256
rect 130160 228216 130166 228228
rect 225782 228216 225788 228228
rect 225840 228216 225846 228268
rect 227622 228216 227628 228268
rect 227680 228256 227686 228268
rect 267090 228256 267096 228268
rect 227680 228228 267096 228256
rect 227680 228216 227686 228228
rect 267090 228216 267096 228228
rect 267148 228216 267154 228268
rect 300946 228216 300952 228268
rect 301004 228256 301010 228268
rect 310238 228256 310244 228268
rect 301004 228228 310244 228256
rect 301004 228216 301010 228228
rect 310238 228216 310244 228228
rect 310296 228216 310302 228268
rect 123386 228148 123392 228200
rect 123444 228188 123450 228200
rect 222930 228188 222936 228200
rect 123444 228160 222936 228188
rect 123444 228148 123450 228160
rect 222930 228148 222936 228160
rect 222988 228148 222994 228200
rect 231670 228148 231676 228200
rect 231728 228188 231734 228200
rect 267826 228188 267832 228200
rect 231728 228160 267832 228188
rect 231728 228148 231734 228160
rect 267826 228148 267832 228160
rect 267884 228148 267890 228200
rect 307018 228148 307024 228200
rect 307076 228188 307082 228200
rect 321186 228188 321192 228200
rect 307076 228160 321192 228188
rect 307076 228148 307082 228160
rect 321186 228148 321192 228160
rect 321244 228148 321250 228200
rect 329116 228188 329144 228364
rect 329190 228352 329196 228404
rect 329248 228392 329254 228404
rect 375926 228392 375932 228404
rect 329248 228364 375932 228392
rect 329248 228352 329254 228364
rect 375926 228352 375932 228364
rect 375984 228352 375990 228404
rect 382274 228352 382280 228404
rect 382332 228392 382338 228404
rect 501230 228392 501236 228404
rect 382332 228364 501236 228392
rect 382332 228352 382338 228364
rect 501230 228352 501236 228364
rect 501288 228352 501294 228404
rect 334894 228284 334900 228336
rect 334952 228324 334958 228336
rect 381998 228324 382004 228336
rect 334952 228296 382004 228324
rect 334952 228284 334958 228296
rect 381998 228284 382004 228296
rect 382056 228284 382062 228336
rect 384390 228284 384396 228336
rect 384448 228324 384454 228336
rect 506290 228324 506296 228336
rect 384448 228296 506296 228324
rect 384448 228284 384454 228296
rect 506290 228284 506296 228296
rect 506348 228284 506354 228336
rect 330570 228216 330576 228268
rect 330628 228256 330634 228268
rect 379238 228256 379244 228268
rect 330628 228228 379244 228256
rect 330628 228216 330634 228228
rect 379238 228216 379244 228228
rect 379296 228216 379302 228268
rect 386506 228216 386512 228268
rect 386564 228256 386570 228268
rect 511350 228256 511356 228268
rect 386564 228228 511356 228256
rect 386564 228216 386570 228228
rect 511350 228216 511356 228228
rect 511408 228216 511414 228268
rect 337654 228188 337660 228200
rect 329116 228160 337660 228188
rect 337654 228148 337660 228160
rect 337712 228148 337718 228200
rect 339494 228148 339500 228200
rect 339552 228188 339558 228200
rect 391842 228188 391848 228200
rect 339552 228160 391848 228188
rect 339552 228148 339558 228160
rect 391842 228148 391848 228160
rect 391900 228148 391906 228200
rect 400490 228148 400496 228200
rect 400548 228188 400554 228200
rect 416866 228188 416872 228200
rect 400548 228160 416872 228188
rect 400548 228148 400554 228160
rect 416866 228148 416872 228160
rect 416924 228148 416930 228200
rect 416958 228148 416964 228200
rect 417016 228188 417022 228200
rect 550266 228188 550272 228200
rect 417016 228160 550272 228188
rect 417016 228148 417022 228160
rect 550266 228148 550272 228160
rect 550324 228148 550330 228200
rect 114922 228080 114928 228132
rect 114980 228120 114986 228132
rect 218974 228120 218980 228132
rect 114980 228092 218980 228120
rect 114980 228080 114986 228092
rect 218974 228080 218980 228092
rect 219032 228080 219038 228132
rect 223482 228080 223488 228132
rect 223540 228120 223546 228132
rect 263870 228120 263876 228132
rect 223540 228092 263876 228120
rect 223540 228080 223546 228092
rect 263870 228080 263876 228092
rect 263928 228080 263934 228132
rect 309502 228080 309508 228132
rect 309560 228120 309566 228132
rect 330478 228120 330484 228132
rect 309560 228092 330484 228120
rect 309560 228080 309566 228092
rect 330478 228080 330484 228092
rect 330536 228080 330542 228132
rect 333422 228080 333428 228132
rect 333480 228120 333486 228132
rect 385954 228120 385960 228132
rect 333480 228092 385960 228120
rect 333480 228080 333486 228092
rect 385954 228080 385960 228092
rect 386012 228080 386018 228132
rect 403618 228080 403624 228132
rect 403676 228120 403682 228132
rect 552014 228120 552020 228132
rect 403676 228092 552020 228120
rect 403676 228080 403682 228092
rect 552014 228080 552020 228092
rect 552072 228080 552078 228132
rect 108206 228012 108212 228064
rect 108264 228052 108270 228064
rect 216122 228052 216128 228064
rect 108264 228024 216128 228052
rect 108264 228012 108270 228024
rect 216122 228012 216128 228024
rect 216180 228012 216186 228064
rect 216674 228012 216680 228064
rect 216732 228052 216738 228064
rect 261018 228052 261024 228064
rect 216732 228024 261024 228052
rect 216732 228012 216738 228024
rect 261018 228012 261024 228024
rect 261076 228012 261082 228064
rect 311710 228012 311716 228064
rect 311768 228052 311774 228064
rect 332962 228052 332968 228064
rect 311768 228024 332968 228052
rect 311768 228012 311774 228024
rect 332962 228012 332968 228024
rect 333020 228012 333026 228064
rect 337010 228012 337016 228064
rect 337068 228052 337074 228064
rect 391934 228052 391940 228064
rect 337068 228024 391940 228052
rect 337068 228012 337074 228024
rect 391934 228012 391940 228024
rect 391992 228012 391998 228064
rect 402974 228012 402980 228064
rect 403032 228052 403038 228064
rect 416958 228052 416964 228064
rect 403032 228024 416964 228052
rect 403032 228012 403038 228024
rect 416958 228012 416964 228024
rect 417016 228012 417022 228064
rect 417050 228012 417056 228064
rect 417108 228052 417114 228064
rect 549254 228052 549260 228064
rect 417108 228024 549260 228052
rect 417108 228012 417114 228024
rect 549254 228012 549260 228024
rect 549312 228012 549318 228064
rect 72050 227944 72056 227996
rect 72108 227984 72114 227996
rect 199746 227984 199752 227996
rect 72108 227956 199752 227984
rect 72108 227944 72114 227956
rect 199746 227944 199752 227956
rect 199804 227944 199810 227996
rect 203242 227944 203248 227996
rect 203300 227984 203306 227996
rect 255314 227984 255320 227996
rect 203300 227956 255320 227984
rect 203300 227944 203306 227956
rect 255314 227944 255320 227956
rect 255372 227944 255378 227996
rect 255958 227944 255964 227996
rect 256016 227984 256022 227996
rect 275646 227984 275652 227996
rect 256016 227956 275652 227984
rect 256016 227944 256022 227956
rect 275646 227944 275652 227956
rect 275704 227944 275710 227996
rect 311342 227944 311348 227996
rect 311400 227984 311406 227996
rect 331306 227984 331312 227996
rect 311400 227956 331312 227984
rect 311400 227944 311406 227956
rect 331306 227944 331312 227956
rect 331364 227944 331370 227996
rect 341242 227944 341248 227996
rect 341300 227984 341306 227996
rect 396534 227984 396540 227996
rect 341300 227956 396540 227984
rect 341300 227944 341306 227956
rect 396534 227944 396540 227956
rect 396592 227944 396598 227996
rect 406838 227944 406844 227996
rect 406896 227984 406902 227996
rect 559282 227984 559288 227996
rect 406896 227956 559288 227984
rect 406896 227944 406902 227956
rect 559282 227944 559288 227956
rect 559340 227944 559346 227996
rect 78766 227876 78772 227928
rect 78824 227916 78830 227928
rect 193766 227916 193772 227928
rect 78824 227888 193772 227916
rect 78824 227876 78830 227888
rect 193766 227876 193772 227888
rect 193824 227876 193830 227928
rect 200114 227916 200120 227928
rect 193876 227888 200120 227916
rect 69474 227808 69480 227860
rect 69532 227848 69538 227860
rect 193876 227848 193904 227888
rect 200114 227876 200120 227888
rect 200172 227876 200178 227928
rect 209590 227876 209596 227928
rect 209648 227916 209654 227928
rect 258166 227916 258172 227928
rect 209648 227888 258172 227916
rect 209648 227876 209654 227888
rect 258166 227876 258172 227888
rect 258224 227876 258230 227928
rect 258350 227876 258356 227928
rect 258408 227916 258414 227928
rect 277486 227916 277492 227928
rect 258408 227888 277492 227916
rect 258408 227876 258414 227888
rect 277486 227876 277492 227888
rect 277544 227876 277550 227928
rect 301682 227876 301688 227928
rect 301740 227916 301746 227928
rect 309410 227916 309416 227928
rect 301740 227888 309416 227916
rect 301740 227876 301746 227888
rect 309410 227876 309416 227888
rect 309468 227876 309474 227928
rect 310606 227876 310612 227928
rect 310664 227916 310670 227928
rect 332134 227916 332140 227928
rect 310664 227888 332140 227916
rect 310664 227876 310670 227888
rect 332134 227876 332140 227888
rect 332192 227876 332198 227928
rect 338390 227876 338396 227928
rect 338448 227916 338454 227928
rect 392946 227916 392952 227928
rect 338448 227888 392952 227916
rect 338448 227876 338454 227888
rect 392946 227876 392952 227888
rect 393004 227876 393010 227928
rect 409046 227876 409052 227928
rect 409104 227916 409110 227928
rect 564434 227916 564440 227928
rect 409104 227888 564440 227916
rect 409104 227876 409110 227888
rect 564434 227876 564440 227888
rect 564492 227876 564498 227928
rect 69532 227820 193904 227848
rect 69532 227808 69538 227820
rect 198734 227808 198740 227860
rect 198792 227848 198798 227860
rect 203978 227848 203984 227860
rect 198792 227820 203984 227848
rect 198792 227808 198798 227820
rect 203978 227808 203984 227820
rect 204036 227808 204042 227860
rect 254670 227848 254676 227860
rect 204088 227820 254676 227848
rect 65334 227740 65340 227792
rect 65392 227780 65398 227792
rect 196894 227780 196900 227792
rect 65392 227752 196900 227780
rect 65392 227740 65398 227752
rect 196894 227740 196900 227752
rect 196952 227740 196958 227792
rect 198918 227740 198924 227792
rect 198976 227780 198982 227792
rect 204088 227780 204116 227820
rect 254670 227808 254676 227820
rect 254728 227808 254734 227860
rect 259546 227808 259552 227860
rect 259604 227848 259610 227860
rect 278866 227848 278872 227860
rect 259604 227820 278872 227848
rect 259604 227808 259610 227820
rect 278866 227808 278872 227820
rect 278924 227808 278930 227860
rect 312078 227808 312084 227860
rect 312136 227848 312142 227860
rect 335538 227848 335544 227860
rect 312136 227820 335544 227848
rect 312136 227808 312142 227820
rect 335538 227808 335544 227820
rect 335596 227808 335602 227860
rect 341610 227808 341616 227860
rect 341668 227848 341674 227860
rect 403618 227848 403624 227860
rect 341668 227820 403624 227848
rect 341668 227808 341674 227820
rect 403618 227808 403624 227820
rect 403676 227808 403682 227860
rect 409322 227808 409328 227860
rect 409380 227848 409386 227860
rect 565446 227848 565452 227860
rect 409380 227820 565452 227848
rect 409380 227808 409386 227820
rect 565446 227808 565452 227820
rect 565504 227808 565510 227860
rect 254302 227780 254308 227792
rect 198976 227752 204116 227780
rect 204180 227752 254308 227780
rect 198976 227740 198982 227752
rect 52730 227672 52736 227724
rect 52788 227712 52794 227724
rect 192938 227712 192944 227724
rect 52788 227684 192944 227712
rect 52788 227672 52794 227684
rect 192938 227672 192944 227684
rect 192996 227672 193002 227724
rect 197354 227672 197360 227724
rect 197412 227712 197418 227724
rect 204180 227712 204208 227752
rect 254302 227740 254308 227752
rect 254360 227740 254366 227792
rect 256510 227740 256516 227792
rect 256568 227780 256574 227792
rect 277118 227780 277124 227792
rect 256568 227752 277124 227780
rect 256568 227740 256574 227752
rect 277118 227740 277124 227752
rect 277176 227740 277182 227792
rect 312722 227740 312728 227792
rect 312780 227780 312786 227792
rect 334710 227780 334716 227792
rect 312780 227752 334716 227780
rect 312780 227740 312786 227752
rect 334710 227740 334716 227752
rect 334768 227740 334774 227792
rect 341978 227740 341984 227792
rect 342036 227780 342042 227792
rect 402974 227780 402980 227792
rect 342036 227752 402980 227780
rect 342036 227740 342042 227752
rect 402974 227740 402980 227752
rect 403032 227740 403038 227792
rect 407206 227740 407212 227792
rect 407264 227780 407270 227792
rect 560386 227780 560392 227792
rect 407264 227752 560392 227780
rect 407264 227740 407270 227752
rect 560386 227740 560392 227752
rect 560444 227740 560450 227792
rect 197412 227684 204208 227712
rect 197412 227672 197418 227684
rect 204254 227672 204260 227724
rect 204312 227712 204318 227724
rect 251818 227712 251824 227724
rect 204312 227684 251824 227712
rect 204312 227672 204318 227684
rect 251818 227672 251824 227684
rect 251876 227672 251882 227724
rect 253750 227672 253756 227724
rect 253808 227712 253814 227724
rect 276750 227712 276756 227724
rect 253808 227684 276756 227712
rect 253808 227672 253814 227684
rect 276750 227672 276756 227684
rect 276808 227672 276814 227724
rect 315942 227672 315948 227724
rect 316000 227712 316006 227724
rect 338298 227712 338304 227724
rect 316000 227684 338304 227712
rect 316000 227672 316006 227684
rect 338298 227672 338304 227684
rect 338356 227672 338362 227724
rect 344462 227672 344468 227724
rect 344520 227712 344526 227724
rect 410334 227712 410340 227724
rect 344520 227684 410340 227712
rect 344520 227672 344526 227684
rect 410334 227672 410340 227684
rect 410392 227672 410398 227724
rect 411530 227672 411536 227724
rect 411588 227712 411594 227724
rect 570230 227712 570236 227724
rect 411588 227684 570236 227712
rect 411588 227672 411594 227684
rect 570230 227672 570236 227684
rect 570288 227672 570294 227724
rect 156138 227604 156144 227656
rect 156196 227644 156202 227656
rect 235350 227644 235356 227656
rect 156196 227616 235356 227644
rect 156196 227604 156202 227616
rect 235350 227604 235356 227616
rect 235408 227604 235414 227656
rect 248690 227604 248696 227656
rect 248748 227644 248754 227656
rect 275002 227644 275008 227656
rect 248748 227616 275008 227644
rect 248748 227604 248754 227616
rect 275002 227604 275008 227616
rect 275060 227604 275066 227656
rect 306006 227604 306012 227656
rect 306064 227644 306070 227656
rect 319530 227644 319536 227656
rect 306064 227616 319536 227644
rect 306064 227604 306070 227616
rect 319530 227604 319536 227616
rect 319588 227604 319594 227656
rect 322014 227604 322020 227656
rect 322072 227644 322078 227656
rect 359090 227644 359096 227656
rect 322072 227616 359096 227644
rect 322072 227604 322078 227616
rect 359090 227604 359096 227616
rect 359148 227604 359154 227656
rect 385126 227604 385132 227656
rect 385184 227644 385190 227656
rect 453850 227644 453856 227656
rect 385184 227616 453856 227644
rect 385184 227604 385190 227616
rect 453850 227604 453856 227616
rect 453908 227604 453914 227656
rect 162762 227536 162768 227588
rect 162820 227576 162826 227588
rect 238202 227576 238208 227588
rect 162820 227548 238208 227576
rect 162820 227536 162826 227548
rect 238202 227536 238208 227548
rect 238260 227536 238266 227588
rect 250346 227536 250352 227588
rect 250404 227576 250410 227588
rect 275278 227576 275284 227588
rect 250404 227548 275284 227576
rect 250404 227536 250410 227548
rect 275278 227536 275284 227548
rect 275336 227536 275342 227588
rect 320266 227536 320272 227588
rect 320324 227576 320330 227588
rect 342070 227576 342076 227588
rect 320324 227548 342076 227576
rect 320324 227536 320330 227548
rect 342070 227536 342076 227548
rect 342128 227536 342134 227588
rect 343726 227536 343732 227588
rect 343784 227576 343790 227588
rect 378134 227576 378140 227588
rect 343784 227548 378140 227576
rect 343784 227536 343790 227548
rect 378134 227536 378140 227548
rect 378192 227536 378198 227588
rect 383010 227536 383016 227588
rect 383068 227576 383074 227588
rect 452562 227576 452568 227588
rect 383068 227548 452568 227576
rect 383068 227536 383074 227548
rect 452562 227536 452568 227548
rect 452620 227536 452626 227588
rect 165430 227468 165436 227520
rect 165488 227508 165494 227520
rect 240410 227508 240416 227520
rect 165488 227480 240416 227508
rect 165488 227468 165494 227480
rect 240410 227468 240416 227480
rect 240468 227468 240474 227520
rect 252002 227468 252008 227520
rect 252060 227508 252066 227520
rect 276382 227508 276388 227520
rect 252060 227480 276388 227508
rect 252060 227468 252066 227480
rect 276382 227468 276388 227480
rect 276440 227468 276446 227520
rect 305270 227468 305276 227520
rect 305328 227508 305334 227520
rect 320358 227508 320364 227520
rect 305328 227480 320364 227508
rect 305328 227468 305334 227480
rect 320358 227468 320364 227480
rect 320416 227468 320422 227520
rect 320634 227468 320640 227520
rect 320692 227508 320698 227520
rect 356054 227508 356060 227520
rect 320692 227480 356060 227508
rect 320692 227468 320698 227480
rect 356054 227468 356060 227480
rect 356112 227468 356118 227520
rect 374454 227468 374460 227520
rect 374512 227508 374518 227520
rect 435726 227508 435732 227520
rect 374512 227480 435732 227508
rect 374512 227468 374518 227480
rect 435726 227468 435732 227480
rect 435784 227468 435790 227520
rect 163682 227400 163688 227452
rect 163740 227440 163746 227452
rect 240042 227440 240048 227452
rect 163740 227412 240048 227440
rect 163740 227400 163746 227412
rect 240042 227400 240048 227412
rect 240100 227400 240106 227452
rect 258718 227400 258724 227452
rect 258776 227440 258782 227452
rect 274266 227440 274272 227452
rect 258776 227412 274272 227440
rect 258776 227400 258782 227412
rect 274266 227400 274272 227412
rect 274324 227400 274330 227452
rect 303798 227400 303804 227452
rect 303856 227440 303862 227452
rect 317414 227440 317420 227452
rect 303856 227412 317420 227440
rect 303856 227400 303862 227412
rect 317414 227400 317420 227412
rect 317472 227400 317478 227452
rect 321646 227400 321652 227452
rect 321704 227440 321710 227452
rect 342898 227440 342904 227452
rect 321704 227412 342904 227440
rect 321704 227400 321710 227412
rect 342898 227400 342904 227412
rect 342956 227400 342962 227452
rect 371602 227400 371608 227452
rect 371660 227440 371666 227452
rect 433150 227440 433156 227452
rect 371660 227412 433156 227440
rect 371660 227400 371666 227412
rect 433150 227400 433156 227412
rect 433208 227400 433214 227452
rect 42058 227332 42064 227384
rect 42116 227372 42122 227384
rect 43438 227372 43444 227384
rect 42116 227344 43444 227372
rect 42116 227332 42122 227344
rect 43438 227332 43444 227344
rect 43496 227332 43502 227384
rect 167086 227332 167092 227384
rect 167144 227372 167150 227384
rect 241422 227372 241428 227384
rect 167144 227344 241428 227372
rect 167144 227332 167150 227344
rect 241422 227332 241428 227344
rect 241480 227332 241486 227384
rect 253566 227332 253572 227384
rect 253624 227372 253630 227384
rect 272794 227372 272800 227384
rect 253624 227344 272800 227372
rect 253624 227332 253630 227344
rect 272794 227332 272800 227344
rect 272852 227332 272858 227384
rect 303154 227332 303160 227384
rect 303212 227372 303218 227384
rect 312814 227372 312820 227384
rect 303212 227344 312820 227372
rect 303212 227332 303218 227344
rect 312814 227332 312820 227344
rect 312872 227332 312878 227384
rect 323118 227332 323124 227384
rect 323176 227372 323182 227384
rect 342990 227372 342996 227384
rect 323176 227344 342996 227372
rect 323176 227332 323182 227344
rect 342990 227332 342996 227344
rect 343048 227332 343054 227384
rect 365898 227332 365904 227384
rect 365956 227372 365962 227384
rect 425422 227372 425428 227384
rect 365956 227344 425428 227372
rect 365956 227332 365962 227344
rect 425422 227332 425428 227344
rect 425480 227332 425486 227384
rect 173618 227264 173624 227316
rect 173676 227304 173682 227316
rect 244274 227304 244280 227316
rect 173676 227276 244280 227304
rect 173676 227264 173682 227276
rect 244274 227264 244280 227276
rect 244332 227264 244338 227316
rect 253198 227264 253204 227316
rect 253256 227304 253262 227316
rect 271414 227304 271420 227316
rect 253256 227276 271420 227304
rect 253256 227264 253262 227276
rect 271414 227264 271420 227276
rect 271472 227264 271478 227316
rect 295242 227264 295248 227316
rect 295300 227304 295306 227316
rect 296806 227304 296812 227316
rect 295300 227276 296812 227304
rect 295300 227264 295306 227276
rect 296806 227264 296812 227276
rect 296864 227264 296870 227316
rect 298738 227264 298744 227316
rect 298796 227304 298802 227316
rect 301038 227304 301044 227316
rect 298796 227276 301044 227304
rect 298796 227264 298802 227276
rect 301038 227264 301044 227276
rect 301096 227264 301102 227316
rect 302418 227264 302424 227316
rect 302476 227304 302482 227316
rect 313642 227304 313648 227316
rect 302476 227276 313648 227304
rect 302476 227264 302482 227276
rect 313642 227264 313648 227276
rect 313700 227264 313706 227316
rect 325970 227264 325976 227316
rect 326028 227304 326034 227316
rect 345290 227304 345296 227316
rect 326028 227276 345296 227304
rect 326028 227264 326034 227276
rect 345290 227264 345296 227276
rect 345348 227264 345354 227316
rect 350166 227264 350172 227316
rect 350224 227304 350230 227316
rect 408494 227304 408500 227316
rect 350224 227276 408500 227304
rect 350224 227264 350230 227276
rect 408494 227264 408500 227276
rect 408552 227264 408558 227316
rect 169570 227196 169576 227248
rect 169628 227236 169634 227248
rect 241054 227236 241060 227248
rect 169628 227208 241060 227236
rect 169628 227196 169634 227208
rect 241054 227196 241060 227208
rect 241112 227196 241118 227248
rect 248506 227196 248512 227248
rect 248564 227236 248570 227248
rect 268562 227236 268568 227248
rect 248564 227208 268568 227236
rect 248564 227196 248570 227208
rect 268562 227196 268568 227208
rect 268620 227196 268626 227248
rect 302050 227196 302056 227248
rect 302108 227236 302114 227248
rect 311986 227236 311992 227248
rect 302108 227208 311992 227236
rect 302108 227196 302114 227208
rect 311986 227196 311992 227208
rect 312044 227196 312050 227248
rect 368750 227196 368756 227248
rect 368808 227236 368814 227248
rect 430390 227236 430396 227248
rect 368808 227208 430396 227236
rect 368808 227196 368814 227208
rect 430390 227196 430396 227208
rect 430448 227196 430454 227248
rect 172146 227128 172152 227180
rect 172204 227168 172210 227180
rect 243262 227168 243268 227180
rect 172204 227140 243268 227168
rect 172204 227128 172210 227140
rect 243262 227128 243268 227140
rect 243320 227128 243326 227180
rect 256602 227128 256608 227180
rect 256660 227168 256666 227180
rect 258718 227168 258724 227180
rect 256660 227140 258724 227168
rect 256660 227128 256666 227140
rect 258718 227128 258724 227140
rect 258776 227128 258782 227180
rect 273898 227168 273904 227180
rect 258828 227140 273904 227168
rect 181898 227060 181904 227112
rect 181956 227100 181962 227112
rect 246114 227100 246120 227112
rect 181956 227072 246120 227100
rect 181956 227060 181962 227072
rect 246114 227060 246120 227072
rect 246172 227060 246178 227112
rect 247034 227060 247040 227112
rect 247092 227100 247098 227112
rect 258828 227100 258856 227140
rect 273898 227128 273904 227140
rect 273956 227128 273962 227180
rect 309226 227128 309232 227180
rect 309284 227168 309290 227180
rect 328822 227168 328828 227180
rect 309284 227140 328828 227168
rect 309284 227128 309290 227140
rect 328822 227128 328828 227140
rect 328880 227128 328886 227180
rect 331674 227128 331680 227180
rect 331732 227168 331738 227180
rect 347774 227168 347780 227180
rect 331732 227140 347780 227168
rect 331732 227128 331738 227140
rect 347774 227128 347780 227140
rect 347832 227128 347838 227180
rect 353018 227128 353024 227180
rect 353076 227168 353082 227180
rect 413186 227168 413192 227180
rect 353076 227140 413192 227168
rect 353076 227128 353082 227140
rect 413186 227128 413192 227140
rect 413244 227128 413250 227180
rect 247092 227072 258856 227100
rect 247092 227060 247098 227072
rect 258902 227060 258908 227112
rect 258960 227100 258966 227112
rect 276014 227100 276020 227112
rect 258960 227072 276020 227100
rect 258960 227060 258966 227072
rect 276014 227060 276020 227072
rect 276072 227060 276078 227112
rect 306374 227060 306380 227112
rect 306432 227100 306438 227112
rect 322014 227100 322020 227112
rect 306432 227072 322020 227100
rect 306432 227060 306438 227072
rect 322014 227060 322020 227072
rect 322072 227060 322078 227112
rect 358722 227060 358728 227112
rect 358780 227100 358786 227112
rect 415302 227100 415308 227112
rect 358780 227072 415308 227100
rect 358780 227060 358786 227072
rect 415302 227060 415308 227072
rect 415360 227060 415366 227112
rect 176378 226992 176384 227044
rect 176436 227032 176442 227044
rect 243906 227032 243912 227044
rect 176436 227004 243912 227032
rect 176436 226992 176442 227004
rect 243906 226992 243912 227004
rect 243964 226992 243970 227044
rect 255498 226992 255504 227044
rect 255556 227032 255562 227044
rect 271782 227032 271788 227044
rect 255556 227004 271788 227032
rect 255556 226992 255562 227004
rect 271782 226992 271788 227004
rect 271840 226992 271846 227044
rect 338022 226992 338028 227044
rect 338080 227032 338086 227044
rect 372062 227032 372068 227044
rect 338080 227004 372068 227032
rect 338080 226992 338086 227004
rect 372062 226992 372068 227004
rect 372120 226992 372126 227044
rect 372982 226992 372988 227044
rect 373040 227032 373046 227044
rect 433242 227032 433248 227044
rect 373040 227004 433248 227032
rect 373040 226992 373046 227004
rect 433242 226992 433248 227004
rect 433300 226992 433306 227044
rect 180518 226924 180524 226976
rect 180576 226964 180582 226976
rect 247126 226964 247132 226976
rect 180576 226936 247132 226964
rect 180576 226924 180582 226936
rect 247126 226924 247132 226936
rect 247184 226924 247190 226976
rect 251450 226964 251456 226976
rect 248524 226936 251456 226964
rect 190362 226856 190368 226908
rect 190420 226896 190426 226908
rect 248524 226896 248552 226936
rect 251450 226924 251456 226936
rect 251508 226924 251514 226976
rect 258718 226924 258724 226976
rect 258776 226964 258782 226976
rect 274634 226964 274640 226976
rect 258776 226936 274640 226964
rect 258776 226924 258782 226936
rect 274634 226924 274640 226936
rect 274692 226924 274698 226976
rect 298094 226924 298100 226976
rect 298152 226964 298158 226976
rect 301958 226964 301964 226976
rect 298152 226936 301964 226964
rect 298152 226924 298158 226936
rect 301958 226924 301964 226936
rect 302016 226924 302022 226976
rect 310514 226924 310520 226976
rect 310572 226964 310578 226976
rect 329650 226964 329656 226976
rect 310572 226936 329656 226964
rect 310572 226924 310578 226936
rect 329650 226924 329656 226936
rect 329708 226924 329714 226976
rect 364426 226924 364432 226976
rect 364484 226964 364490 226976
rect 422294 226964 422300 226976
rect 364484 226936 422300 226964
rect 364484 226924 364490 226936
rect 422294 226924 422300 226936
rect 422352 226924 422358 226976
rect 190420 226868 248552 226896
rect 190420 226856 190426 226868
rect 248598 226856 248604 226908
rect 248656 226896 248662 226908
rect 269942 226896 269948 226908
rect 248656 226868 269948 226896
rect 248656 226856 248662 226868
rect 269942 226856 269948 226868
rect 270000 226856 270006 226908
rect 290734 226856 290740 226908
rect 290792 226896 290798 226908
rect 292390 226896 292396 226908
rect 290792 226868 292396 226896
rect 290792 226856 290798 226868
rect 292390 226856 292396 226868
rect 292448 226856 292454 226908
rect 300670 226856 300676 226908
rect 300728 226896 300734 226908
rect 308582 226896 308588 226908
rect 300728 226868 308588 226896
rect 300728 226856 300734 226868
rect 308582 226856 308588 226868
rect 308640 226856 308646 226908
rect 361574 226856 361580 226908
rect 361632 226896 361638 226908
rect 416866 226896 416872 226908
rect 361632 226868 416872 226896
rect 361632 226856 361638 226868
rect 416866 226856 416872 226868
rect 416924 226856 416930 226908
rect 42150 226788 42156 226840
rect 42208 226828 42214 226840
rect 43622 226828 43628 226840
rect 42208 226800 43628 226828
rect 42208 226788 42214 226800
rect 43622 226788 43628 226800
rect 43680 226788 43686 226840
rect 189258 226788 189264 226840
rect 189316 226828 189322 226840
rect 248966 226828 248972 226840
rect 189316 226800 248972 226828
rect 189316 226788 189322 226800
rect 248966 226788 248972 226800
rect 249024 226788 249030 226840
rect 265710 226828 265716 226840
rect 249076 226800 265716 226828
rect 186406 226720 186412 226772
rect 186464 226760 186470 226772
rect 248230 226760 248236 226772
rect 186464 226732 248236 226760
rect 186464 226720 186470 226732
rect 248230 226720 248236 226732
rect 248288 226720 248294 226772
rect 248414 226720 248420 226772
rect 248472 226760 248478 226772
rect 249076 226760 249104 226800
rect 265710 226788 265716 226800
rect 265768 226788 265774 226840
rect 299566 226788 299572 226840
rect 299624 226828 299630 226840
rect 306926 226828 306932 226840
rect 299624 226800 306932 226828
rect 299624 226788 299630 226800
rect 306926 226788 306932 226800
rect 306984 226788 306990 226840
rect 359826 226788 359832 226840
rect 359884 226828 359890 226840
rect 404538 226828 404544 226840
rect 359884 226800 404544 226828
rect 359884 226788 359890 226800
rect 404538 226788 404544 226800
rect 404596 226788 404602 226840
rect 409690 226788 409696 226840
rect 409748 226828 409754 226840
rect 447134 226828 447140 226840
rect 409748 226800 447140 226828
rect 409748 226788 409754 226800
rect 447134 226788 447140 226800
rect 447192 226788 447198 226840
rect 248472 226732 249104 226760
rect 248472 226720 248478 226732
rect 255774 226720 255780 226772
rect 255832 226760 255838 226772
rect 268930 226760 268936 226772
rect 255832 226732 268936 226760
rect 255832 226720 255838 226732
rect 268930 226720 268936 226732
rect 268988 226720 268994 226772
rect 299198 226720 299204 226772
rect 299256 226760 299262 226772
rect 305270 226760 305276 226772
rect 299256 226732 305276 226760
rect 299256 226720 299262 226732
rect 305270 226720 305276 226732
rect 305328 226720 305334 226772
rect 368382 226720 368388 226772
rect 368440 226760 368446 226772
rect 408770 226760 408776 226772
rect 368440 226732 408776 226760
rect 368440 226720 368446 226732
rect 408770 226720 408776 226732
rect 408828 226720 408834 226772
rect 195882 226652 195888 226704
rect 195940 226692 195946 226704
rect 251082 226692 251088 226704
rect 195940 226664 251088 226692
rect 195940 226652 195946 226664
rect 251082 226652 251088 226664
rect 251140 226652 251146 226704
rect 258810 226652 258816 226704
rect 258868 226692 258874 226704
rect 273162 226692 273168 226704
rect 258868 226664 273168 226692
rect 258868 226652 258874 226664
rect 273162 226652 273168 226664
rect 273220 226652 273226 226704
rect 297818 226652 297824 226704
rect 297876 226692 297882 226704
rect 301866 226692 301872 226704
rect 297876 226664 301872 226692
rect 297876 226652 297882 226664
rect 301866 226652 301872 226664
rect 301924 226652 301930 226704
rect 301958 226652 301964 226704
rect 302016 226692 302022 226704
rect 303614 226692 303620 226704
rect 302016 226664 303620 226692
rect 302016 226652 302022 226664
rect 303614 226652 303620 226664
rect 303672 226652 303678 226704
rect 329098 226652 329104 226704
rect 329156 226692 329162 226704
rect 345106 226692 345112 226704
rect 329156 226664 345112 226692
rect 329156 226652 329162 226664
rect 345106 226652 345112 226664
rect 345164 226652 345170 226704
rect 365530 226652 365536 226704
rect 365588 226692 365594 226704
rect 405826 226692 405832 226704
rect 365588 226664 405832 226692
rect 365588 226652 365594 226664
rect 405826 226652 405832 226664
rect 405884 226652 405890 226704
rect 408678 226652 408684 226704
rect 408736 226692 408742 226704
rect 444374 226692 444380 226704
rect 408736 226664 444380 226692
rect 408736 226652 408742 226664
rect 444374 226652 444380 226664
rect 444432 226652 444438 226704
rect 193030 226584 193036 226636
rect 193088 226624 193094 226636
rect 204254 226624 204260 226636
rect 193088 226596 204260 226624
rect 193088 226584 193094 226596
rect 204254 226584 204260 226596
rect 204312 226584 204318 226636
rect 236270 226584 236276 226636
rect 236328 226624 236334 226636
rect 256786 226624 256792 226636
rect 236328 226596 256792 226624
rect 236328 226584 236334 226596
rect 256786 226584 256792 226596
rect 256844 226584 256850 226636
rect 300302 226584 300308 226636
rect 300360 226624 300366 226636
rect 306374 226624 306380 226636
rect 300360 226596 306380 226624
rect 300360 226584 300366 226596
rect 306374 226584 306380 226596
rect 306432 226584 306438 226636
rect 395798 226584 395804 226636
rect 395856 226624 395862 226636
rect 438762 226624 438768 226636
rect 395856 226596 438768 226624
rect 395856 226584 395862 226596
rect 438762 226584 438768 226596
rect 438820 226584 438826 226636
rect 193766 226516 193772 226568
rect 193824 226556 193830 226568
rect 202598 226556 202604 226568
rect 193824 226528 202604 226556
rect 193824 226516 193830 226528
rect 202598 226516 202604 226528
rect 202656 226516 202662 226568
rect 301314 226516 301320 226568
rect 301372 226556 301378 226568
rect 307754 226556 307760 226568
rect 301372 226528 307760 226556
rect 301372 226516 301378 226528
rect 307754 226516 307760 226528
rect 307812 226516 307818 226568
rect 402606 226516 402612 226568
rect 402664 226556 402670 226568
rect 417050 226556 417056 226568
rect 402664 226528 417056 226556
rect 402664 226516 402670 226528
rect 417050 226516 417056 226528
rect 417108 226516 417114 226568
rect 441614 226556 441620 226568
rect 419506 226528 441620 226556
rect 255314 226448 255320 226500
rect 255372 226488 255378 226500
rect 270310 226488 270316 226500
rect 255372 226460 270316 226488
rect 255372 226448 255378 226460
rect 270310 226448 270316 226460
rect 270368 226448 270374 226500
rect 374086 226448 374092 226500
rect 374144 226488 374150 226500
rect 405734 226488 405740 226500
rect 374144 226460 405740 226488
rect 374144 226448 374150 226460
rect 405734 226448 405740 226460
rect 405792 226448 405798 226500
rect 201586 226380 201592 226432
rect 201644 226420 201650 226432
rect 209038 226420 209044 226432
rect 201644 226392 209044 226420
rect 201644 226380 201650 226392
rect 209038 226380 209044 226392
rect 209096 226380 209102 226432
rect 233510 226380 233516 226432
rect 233568 226420 233574 226432
rect 247494 226420 247500 226432
rect 233568 226392 247500 226420
rect 233568 226380 233574 226392
rect 247494 226380 247500 226392
rect 247552 226380 247558 226432
rect 404354 226380 404360 226432
rect 404412 226420 404418 226432
rect 419506 226420 419534 226528
rect 441614 226516 441620 226528
rect 441672 226516 441678 226568
rect 404412 226392 419534 226420
rect 404412 226380 404418 226392
rect 183002 226312 183008 226364
rect 183060 226352 183066 226364
rect 192294 226352 192300 226364
rect 183060 226324 192300 226352
rect 183060 226312 183066 226324
rect 192294 226312 192300 226324
rect 192352 226312 192358 226364
rect 258166 226312 258172 226364
rect 258224 226352 258230 226364
rect 264606 226352 264612 226364
rect 258224 226324 264612 226352
rect 258224 226312 258230 226324
rect 264606 226312 264612 226324
rect 264664 226312 264670 226364
rect 299934 226312 299940 226364
rect 299992 226352 299998 226364
rect 304350 226352 304356 226364
rect 299992 226324 304356 226352
rect 299992 226312 299998 226324
rect 304350 226312 304356 226324
rect 304408 226312 304414 226364
rect 309870 226312 309876 226364
rect 309928 226352 309934 226364
rect 327902 226352 327908 226364
rect 309928 226324 327908 226352
rect 309928 226312 309934 226324
rect 327902 226312 327908 226324
rect 327960 226312 327966 226364
rect 144362 226244 144368 226296
rect 144420 226284 144426 226296
rect 230750 226284 230756 226296
rect 144420 226256 230756 226284
rect 144420 226244 144426 226256
rect 230750 226244 230756 226256
rect 230808 226244 230814 226296
rect 349430 226244 349436 226296
rect 349488 226284 349494 226296
rect 425054 226284 425060 226296
rect 349488 226256 425060 226284
rect 349488 226244 349494 226256
rect 425054 226244 425060 226256
rect 425112 226244 425118 226296
rect 430390 226244 430396 226296
rect 430448 226284 430454 226296
rect 467558 226284 467564 226296
rect 430448 226256 467564 226284
rect 430448 226244 430454 226256
rect 467558 226244 467564 226256
rect 467616 226244 467622 226296
rect 147766 226176 147772 226228
rect 147824 226216 147830 226228
rect 232222 226216 232228 226228
rect 147824 226188 232228 226216
rect 147824 226176 147830 226188
rect 232222 226176 232228 226188
rect 232280 226176 232286 226228
rect 352650 226176 352656 226228
rect 352708 226216 352714 226228
rect 428918 226216 428924 226228
rect 352708 226188 428924 226216
rect 352708 226176 352714 226188
rect 428918 226176 428924 226188
rect 428976 226176 428982 226228
rect 433150 226176 433156 226228
rect 433208 226216 433214 226228
rect 474274 226216 474280 226228
rect 433208 226188 474280 226216
rect 433208 226176 433214 226188
rect 474274 226176 474280 226188
rect 474332 226176 474338 226228
rect 141050 226108 141056 226160
rect 141108 226148 141114 226160
rect 229370 226148 229376 226160
rect 141108 226120 229376 226148
rect 141108 226108 141114 226120
rect 229370 226108 229376 226120
rect 229428 226108 229434 226160
rect 353754 226108 353760 226160
rect 353812 226148 353818 226160
rect 434806 226148 434812 226160
rect 353812 226120 434812 226148
rect 353812 226108 353818 226120
rect 434806 226108 434812 226120
rect 434864 226108 434870 226160
rect 137646 226040 137652 226092
rect 137704 226080 137710 226092
rect 227898 226080 227904 226092
rect 137704 226052 227904 226080
rect 137704 226040 137710 226052
rect 227898 226040 227904 226052
rect 227956 226040 227962 226092
rect 352282 226040 352288 226092
rect 352340 226080 352346 226092
rect 431402 226080 431408 226092
rect 352340 226052 431408 226080
rect 352340 226040 352346 226052
rect 431402 226040 431408 226052
rect 431460 226040 431466 226092
rect 433242 226040 433248 226092
rect 433300 226080 433306 226092
rect 477770 226080 477776 226092
rect 433300 226052 477776 226080
rect 433300 226040 433306 226052
rect 477770 226040 477776 226052
rect 477828 226040 477834 226092
rect 134242 225972 134248 226024
rect 134300 226012 134306 226024
rect 226518 226012 226524 226024
rect 134300 225984 226524 226012
rect 134300 225972 134306 225984
rect 226518 225972 226524 225984
rect 226576 225972 226582 226024
rect 356974 225972 356980 226024
rect 357032 226012 357038 226024
rect 439038 226012 439044 226024
rect 357032 225984 439044 226012
rect 357032 225972 357038 225984
rect 439038 225972 439044 225984
rect 439096 225972 439102 226024
rect 480990 226012 480996 226024
rect 458146 225984 480996 226012
rect 130930 225904 130936 225956
rect 130988 225944 130994 225956
rect 225046 225944 225052 225956
rect 130988 225916 225052 225944
rect 130988 225904 130994 225916
rect 225046 225904 225052 225916
rect 225104 225904 225110 225956
rect 243078 225904 243084 225956
rect 243136 225944 243142 225956
rect 252922 225944 252928 225956
rect 243136 225916 252928 225944
rect 243136 225904 243142 225916
rect 252922 225904 252928 225916
rect 252980 225904 252986 225956
rect 355502 225904 355508 225956
rect 355560 225944 355566 225956
rect 435634 225944 435640 225956
rect 355560 225916 435640 225944
rect 355560 225904 355566 225916
rect 435634 225904 435640 225916
rect 435692 225904 435698 225956
rect 435726 225904 435732 225956
rect 435784 225944 435790 225956
rect 458146 225944 458174 225984
rect 480990 225972 480996 225984
rect 481048 225972 481054 226024
rect 435784 225916 458174 225944
rect 435784 225904 435790 225916
rect 127526 225836 127532 225888
rect 127584 225876 127590 225888
rect 223666 225876 223672 225888
rect 127584 225848 223672 225876
rect 127584 225836 127590 225848
rect 223666 225836 223672 225848
rect 223724 225836 223730 225888
rect 242986 225836 242992 225888
rect 243044 225876 243050 225888
rect 252830 225876 252836 225888
rect 243044 225848 252836 225876
rect 243044 225836 243050 225848
rect 252830 225836 252836 225848
rect 252888 225836 252894 225888
rect 356606 225836 356612 225888
rect 356664 225876 356670 225888
rect 429102 225876 429108 225888
rect 356664 225848 429108 225876
rect 356664 225836 356670 225848
rect 429102 225836 429108 225848
rect 429160 225836 429166 225888
rect 448238 225876 448244 225888
rect 430546 225848 448244 225876
rect 119154 225768 119160 225820
rect 119212 225808 119218 225820
rect 219710 225808 219716 225820
rect 119212 225780 219716 225808
rect 119212 225768 119218 225780
rect 219710 225768 219716 225780
rect 219768 225768 219774 225820
rect 231302 225768 231308 225820
rect 231360 225808 231366 225820
rect 249610 225808 249616 225820
rect 231360 225780 249616 225808
rect 231360 225768 231366 225780
rect 249610 225768 249616 225780
rect 249668 225768 249674 225820
rect 359458 225768 359464 225820
rect 359516 225808 359522 225820
rect 430546 225808 430574 225848
rect 448238 225836 448244 225848
rect 448296 225836 448302 225888
rect 474734 225836 474740 225888
rect 474792 225876 474798 225888
rect 491294 225876 491300 225888
rect 474792 225848 491300 225876
rect 474792 225836 474798 225848
rect 491294 225836 491300 225848
rect 491352 225836 491358 225888
rect 359516 225780 430574 225808
rect 440160 225780 452516 225808
rect 359516 225768 359522 225780
rect 124122 225700 124128 225752
rect 124180 225740 124186 225752
rect 222194 225740 222200 225752
rect 124180 225712 222200 225740
rect 124180 225700 124186 225712
rect 222194 225700 222200 225712
rect 222252 225700 222258 225752
rect 232038 225700 232044 225752
rect 232096 225740 232102 225752
rect 253934 225740 253940 225752
rect 232096 225712 253940 225740
rect 232096 225700 232102 225712
rect 253934 225700 253940 225712
rect 253992 225700 253998 225752
rect 362310 225700 362316 225752
rect 362368 225740 362374 225752
rect 440160 225740 440188 225780
rect 451550 225740 451556 225752
rect 362368 225712 440188 225740
rect 440252 225712 451556 225740
rect 362368 225700 362374 225712
rect 114094 225632 114100 225684
rect 114152 225672 114158 225684
rect 217962 225672 217968 225684
rect 114152 225644 217968 225672
rect 114152 225632 114158 225644
rect 217962 225632 217968 225644
rect 218020 225632 218026 225684
rect 252462 225672 252468 225684
rect 226306 225644 252468 225672
rect 110690 225564 110696 225616
rect 110748 225604 110754 225616
rect 216490 225604 216496 225616
rect 110748 225576 216496 225604
rect 110748 225564 110754 225576
rect 216490 225564 216496 225576
rect 216548 225564 216554 225616
rect 216582 225564 216588 225616
rect 216640 225604 216646 225616
rect 226306 225604 226334 225644
rect 252462 225632 252468 225644
rect 252520 225632 252526 225684
rect 360838 225632 360844 225684
rect 360896 225672 360902 225684
rect 440252 225672 440280 225712
rect 451550 225700 451556 225712
rect 451608 225700 451614 225752
rect 452488 225740 452516 225780
rect 452562 225768 452568 225820
rect 452620 225808 452626 225820
rect 503162 225808 503168 225820
rect 452620 225780 503168 225808
rect 452620 225768 452626 225780
rect 503162 225768 503168 225780
rect 503220 225768 503226 225820
rect 454954 225740 454960 225752
rect 452488 225712 454960 225740
rect 454954 225700 454960 225712
rect 455012 225700 455018 225752
rect 460934 225700 460940 225752
rect 460992 225740 460998 225752
rect 487798 225740 487804 225752
rect 460992 225712 487804 225740
rect 460992 225700 460998 225712
rect 487798 225700 487804 225712
rect 487856 225700 487862 225752
rect 461670 225672 461676 225684
rect 360896 225644 440280 225672
rect 440436 225644 461676 225672
rect 360896 225632 360902 225644
rect 216640 225576 226334 225604
rect 216640 225564 216646 225576
rect 228450 225564 228456 225616
rect 228508 225604 228514 225616
rect 266446 225604 266452 225616
rect 228508 225576 266452 225604
rect 228508 225564 228514 225576
rect 266446 225564 266452 225576
rect 266504 225564 266510 225616
rect 362678 225564 362684 225616
rect 362736 225604 362742 225616
rect 440326 225604 440332 225616
rect 362736 225576 440332 225604
rect 362736 225564 362742 225576
rect 440326 225564 440332 225576
rect 440384 225564 440390 225616
rect 105722 225496 105728 225548
rect 105780 225536 105786 225548
rect 214006 225536 214012 225548
rect 105780 225508 214012 225536
rect 105780 225496 105786 225508
rect 214006 225496 214012 225508
rect 214064 225496 214070 225548
rect 218422 225496 218428 225548
rect 218480 225536 218486 225548
rect 262122 225536 262128 225548
rect 218480 225508 262128 225536
rect 218480 225496 218486 225508
rect 262122 225496 262128 225508
rect 262180 225496 262186 225548
rect 365162 225496 365168 225548
rect 365220 225536 365226 225548
rect 440436 225536 440464 225644
rect 461670 225632 461676 225644
rect 461728 225632 461734 225684
rect 467006 225632 467012 225684
rect 467064 225672 467070 225684
rect 523954 225672 523960 225684
rect 467064 225644 523960 225672
rect 467064 225632 467070 225644
rect 523954 225632 523960 225644
rect 524012 225632 524018 225684
rect 440510 225564 440516 225616
rect 440568 225604 440574 225616
rect 452654 225604 452660 225616
rect 440568 225576 452660 225604
rect 440568 225564 440574 225576
rect 452654 225564 452660 225576
rect 452712 225564 452718 225616
rect 453850 225564 453856 225616
rect 453908 225604 453914 225616
rect 507946 225604 507952 225616
rect 453908 225576 507952 225604
rect 453908 225564 453914 225576
rect 507946 225564 507952 225576
rect 508004 225564 508010 225616
rect 458450 225536 458456 225548
rect 365220 225508 440464 225536
rect 449866 225508 458456 225536
rect 365220 225496 365226 225508
rect 107378 225428 107384 225480
rect 107436 225468 107442 225480
rect 215110 225468 215116 225480
rect 107436 225440 215116 225468
rect 107436 225428 107442 225440
rect 215110 225428 215116 225440
rect 215168 225428 215174 225480
rect 221734 225428 221740 225480
rect 221792 225468 221798 225480
rect 263594 225468 263600 225480
rect 221792 225440 263600 225468
rect 221792 225428 221798 225440
rect 263594 225428 263600 225440
rect 263652 225428 263658 225480
rect 363690 225428 363696 225480
rect 363748 225468 363754 225480
rect 449866 225468 449894 225508
rect 458450 225496 458456 225508
rect 458508 225496 458514 225548
rect 464430 225496 464436 225548
rect 464488 225536 464494 225548
rect 518894 225536 518900 225548
rect 464488 225508 518900 225536
rect 464488 225496 464494 225508
rect 518894 225496 518900 225508
rect 518952 225496 518958 225548
rect 363748 225440 449894 225468
rect 363748 225428 363754 225440
rect 458174 225428 458180 225480
rect 458232 225468 458238 225480
rect 513374 225468 513380 225480
rect 458232 225440 513380 225468
rect 458232 225428 458238 225440
rect 513374 225428 513380 225440
rect 513432 225428 513438 225480
rect 100662 225360 100668 225412
rect 100720 225400 100726 225412
rect 192754 225400 192760 225412
rect 100720 225372 192760 225400
rect 100720 225360 100726 225372
rect 192754 225360 192760 225372
rect 192812 225360 192818 225412
rect 207014 225400 207020 225412
rect 192864 225372 207020 225400
rect 97258 225292 97264 225344
rect 97316 225332 97322 225344
rect 192864 225332 192892 225372
rect 207014 225360 207020 225372
rect 207072 225360 207078 225412
rect 225138 225360 225144 225412
rect 225196 225400 225202 225412
rect 264974 225400 264980 225412
rect 225196 225372 264980 225400
rect 225196 225360 225202 225372
rect 264974 225360 264980 225372
rect 265032 225360 265038 225412
rect 355134 225360 355140 225412
rect 355192 225400 355198 225412
rect 438118 225400 438124 225412
rect 355192 225372 438124 225400
rect 355192 225360 355198 225372
rect 438118 225360 438124 225372
rect 438176 225360 438182 225412
rect 438762 225360 438768 225412
rect 438820 225400 438826 225412
rect 532694 225400 532700 225412
rect 438820 225372 532700 225400
rect 438820 225360 438826 225372
rect 532694 225360 532700 225372
rect 532752 225360 532758 225412
rect 209682 225332 209688 225344
rect 97316 225304 192892 225332
rect 197280 225304 209688 225332
rect 97316 225292 97322 225304
rect 95602 225224 95608 225276
rect 95660 225264 95666 225276
rect 197280 225264 197308 225304
rect 209682 225292 209688 225304
rect 209740 225292 209746 225344
rect 215018 225292 215024 225344
rect 215076 225332 215082 225344
rect 260742 225332 260748 225344
rect 215076 225304 260748 225332
rect 215076 225292 215082 225304
rect 260742 225292 260748 225304
rect 260800 225292 260806 225344
rect 366542 225292 366548 225344
rect 366600 225332 366606 225344
rect 465074 225332 465080 225344
rect 366600 225304 465080 225332
rect 366600 225292 366606 225304
rect 465074 225292 465080 225304
rect 465132 225292 465138 225344
rect 469950 225292 469956 225344
rect 470008 225332 470014 225344
rect 529014 225332 529020 225344
rect 470008 225304 529020 225332
rect 470008 225292 470014 225304
rect 529014 225292 529020 225304
rect 529072 225292 529078 225344
rect 95660 225236 197308 225264
rect 95660 225224 95666 225236
rect 211706 225224 211712 225276
rect 211764 225264 211770 225276
rect 259270 225264 259276 225276
rect 211764 225236 259276 225264
rect 211764 225224 211770 225236
rect 259270 225224 259276 225236
rect 259328 225224 259334 225276
rect 343082 225224 343088 225276
rect 343140 225264 343146 225276
rect 365714 225264 365720 225276
rect 343140 225236 365720 225264
rect 343140 225224 343146 225236
rect 365714 225224 365720 225236
rect 365772 225224 365778 225276
rect 368014 225224 368020 225276
rect 368072 225264 368078 225276
rect 468386 225264 468392 225276
rect 368072 225236 468392 225264
rect 368072 225224 368078 225236
rect 468386 225224 468392 225236
rect 468444 225224 468450 225276
rect 473262 225224 473268 225276
rect 473320 225264 473326 225276
rect 533982 225264 533988 225276
rect 473320 225236 533988 225264
rect 473320 225224 473326 225236
rect 533982 225224 533988 225236
rect 534040 225224 534046 225276
rect 88886 225156 88892 225208
rect 88944 225196 88950 225208
rect 192662 225196 192668 225208
rect 88944 225168 192668 225196
rect 88944 225156 88950 225168
rect 192662 225156 192668 225168
rect 192720 225156 192726 225208
rect 192754 225156 192760 225208
rect 192812 225196 192818 225208
rect 197446 225196 197452 225208
rect 192812 225168 197452 225196
rect 192812 225156 192818 225168
rect 197446 225156 197452 225168
rect 197504 225156 197510 225208
rect 208302 225156 208308 225208
rect 208360 225196 208366 225208
rect 257890 225196 257896 225208
rect 208360 225168 257896 225196
rect 208360 225156 208366 225168
rect 257890 225156 257896 225168
rect 257948 225156 257954 225208
rect 313458 225156 313464 225208
rect 313516 225196 313522 225208
rect 338850 225196 338856 225208
rect 313516 225168 338856 225196
rect 313516 225156 313522 225168
rect 338850 225156 338856 225168
rect 338908 225156 338914 225208
rect 339862 225156 339868 225208
rect 339920 225196 339926 225208
rect 368566 225196 368572 225208
rect 339920 225168 368572 225196
rect 339920 225156 339926 225168
rect 368566 225156 368572 225168
rect 368624 225156 368630 225208
rect 369762 225156 369768 225208
rect 369820 225196 369826 225208
rect 469214 225196 469220 225208
rect 369820 225168 469220 225196
rect 369820 225156 369826 225168
rect 469214 225156 469220 225168
rect 469272 225156 469278 225208
rect 477494 225156 477500 225208
rect 477552 225196 477558 225208
rect 544102 225196 544108 225208
rect 477552 225168 544108 225196
rect 477552 225156 477558 225168
rect 544102 225156 544108 225168
rect 544160 225156 544166 225208
rect 92198 225088 92204 225140
rect 92256 225128 92262 225140
rect 208026 225128 208032 225140
rect 92256 225100 208032 225128
rect 92256 225088 92262 225100
rect 208026 225088 208032 225100
rect 208084 225088 208090 225140
rect 209222 225088 209228 225140
rect 209280 225128 209286 225140
rect 257154 225128 257160 225140
rect 209280 225100 257160 225128
rect 209280 225088 209286 225100
rect 257154 225088 257160 225100
rect 257212 225088 257218 225140
rect 314930 225088 314936 225140
rect 314988 225128 314994 225140
rect 342530 225128 342536 225140
rect 314988 225100 342536 225128
rect 314988 225088 314994 225100
rect 342530 225088 342536 225100
rect 342588 225088 342594 225140
rect 358354 225088 358360 225140
rect 358412 225128 358418 225140
rect 358412 225100 436508 225128
rect 358412 225088 358418 225100
rect 73706 225020 73712 225072
rect 73764 225060 73770 225072
rect 200850 225060 200856 225072
rect 73764 225032 200856 225060
rect 73764 225020 73770 225032
rect 200850 225020 200856 225032
rect 200908 225020 200914 225072
rect 201402 225020 201408 225072
rect 201460 225060 201466 225072
rect 255038 225060 255044 225072
rect 201460 225032 255044 225060
rect 201460 225020 201466 225032
rect 255038 225020 255044 225032
rect 255096 225020 255102 225072
rect 317782 225020 317788 225072
rect 317840 225060 317846 225072
rect 348970 225060 348976 225072
rect 317840 225032 348976 225060
rect 317840 225020 317846 225032
rect 348970 225020 348976 225032
rect 349028 225020 349034 225072
rect 357986 225020 357992 225072
rect 358044 225060 358050 225072
rect 436480 225060 436508 225100
rect 441614 225088 441620 225140
rect 441672 225128 441678 225140
rect 554314 225128 554320 225140
rect 441672 225100 554320 225128
rect 441672 225088 441678 225100
rect 554314 225088 554320 225100
rect 554372 225088 554378 225140
rect 442350 225060 442356 225072
rect 358044 225032 436416 225060
rect 436480 225032 442356 225060
rect 358044 225020 358050 225032
rect 60274 224952 60280 225004
rect 60332 224992 60338 225004
rect 195146 224992 195152 225004
rect 60332 224964 195152 224992
rect 60332 224952 60338 224964
rect 195146 224952 195152 224964
rect 195204 224952 195210 225004
rect 195238 224952 195244 225004
rect 195296 224992 195302 225004
rect 252186 224992 252192 225004
rect 195296 224964 252192 224992
rect 195296 224952 195302 224964
rect 252186 224952 252192 224964
rect 252244 224952 252250 225004
rect 319162 224952 319168 225004
rect 319220 224992 319226 225004
rect 352374 224992 352380 225004
rect 319220 224964 352380 224992
rect 319220 224952 319226 224964
rect 352374 224952 352380 224964
rect 352432 224952 352438 225004
rect 361206 224952 361212 225004
rect 361264 224992 361270 225004
rect 434622 224992 434628 225004
rect 361264 224964 434628 224992
rect 361264 224952 361270 224964
rect 434622 224952 434628 224964
rect 434680 224952 434686 225004
rect 436388 224992 436416 225032
rect 442350 225020 442356 225032
rect 442408 225020 442414 225072
rect 444374 225020 444380 225072
rect 444432 225060 444438 225072
rect 563698 225060 563704 225072
rect 444432 225032 563704 225060
rect 444432 225020 444438 225032
rect 563698 225020 563704 225032
rect 563756 225020 563762 225072
rect 444834 224992 444840 225004
rect 434732 224964 436324 224992
rect 436388 224964 444840 224992
rect 55122 224884 55128 224936
rect 55180 224924 55186 224936
rect 192570 224924 192576 224936
rect 55180 224896 192576 224924
rect 55180 224884 55186 224896
rect 192570 224884 192576 224896
rect 192628 224884 192634 224936
rect 192662 224884 192668 224936
rect 192720 224924 192726 224936
rect 206830 224924 206836 224936
rect 192720 224896 206836 224924
rect 192720 224884 192726 224896
rect 206830 224884 206836 224896
rect 206888 224884 206894 224936
rect 206922 224884 206928 224936
rect 206980 224924 206986 224936
rect 250714 224924 250720 224936
rect 206980 224896 250720 224924
rect 206980 224884 206986 224896
rect 250714 224884 250720 224896
rect 250772 224884 250778 224936
rect 316310 224884 316316 224936
rect 316368 224924 316374 224936
rect 345658 224924 345664 224936
rect 316368 224896 345664 224924
rect 316368 224884 316374 224896
rect 345658 224884 345664 224896
rect 345716 224884 345722 224936
rect 346578 224884 346584 224936
rect 346636 224924 346642 224936
rect 416682 224924 416688 224936
rect 346636 224896 416688 224924
rect 346636 224884 346642 224896
rect 416682 224884 416688 224896
rect 416740 224884 416746 224936
rect 416774 224884 416780 224936
rect 416832 224924 416838 224936
rect 434732 224924 434760 224964
rect 416832 224896 434760 224924
rect 436296 224924 436324 224964
rect 444834 224952 444840 224964
rect 444892 224952 444898 225004
rect 447134 224952 447140 225004
rect 447192 224992 447198 225004
rect 565998 224992 566004 225004
rect 447192 224964 566004 224992
rect 447192 224952 447198 224964
rect 565998 224952 566004 224964
rect 566056 224952 566062 225004
rect 549346 224924 549352 224936
rect 436296 224896 549352 224924
rect 416832 224884 416838 224896
rect 549346 224884 549352 224896
rect 549404 224884 549410 224936
rect 114278 224816 114284 224868
rect 114336 224856 114342 224868
rect 197998 224856 198004 224868
rect 114336 224828 198004 224856
rect 114336 224816 114342 224828
rect 197998 224816 198004 224828
rect 198056 224816 198062 224868
rect 198182 224816 198188 224868
rect 198240 224856 198246 224868
rect 253290 224856 253296 224868
rect 198240 224828 253296 224856
rect 198240 224816 198246 224828
rect 253290 224816 253296 224828
rect 253348 224816 253354 224868
rect 350902 224816 350908 224868
rect 350960 224856 350966 224868
rect 427998 224856 428004 224868
rect 350960 224828 428004 224856
rect 350960 224816 350966 224828
rect 427998 224816 428004 224828
rect 428056 224816 428062 224868
rect 434622 224816 434628 224868
rect 434680 224856 434686 224868
rect 449066 224856 449072 224868
rect 434680 224828 449072 224856
rect 434680 224816 434686 224828
rect 449066 224816 449072 224828
rect 449124 224816 449130 224868
rect 154482 224748 154488 224800
rect 154540 224788 154546 224800
rect 235074 224788 235080 224800
rect 154540 224760 235080 224788
rect 154540 224748 154546 224760
rect 235074 224748 235080 224760
rect 235132 224748 235138 224800
rect 354122 224748 354128 224800
rect 354180 224788 354186 224800
rect 425238 224788 425244 224800
rect 354180 224760 425244 224788
rect 354180 224748 354186 224760
rect 425238 224748 425244 224760
rect 425296 224748 425302 224800
rect 425514 224788 425520 224800
rect 425348 224760 425520 224788
rect 151078 224680 151084 224732
rect 151136 224720 151142 224732
rect 233602 224720 233608 224732
rect 151136 224692 233608 224720
rect 151136 224680 151142 224692
rect 233602 224680 233608 224692
rect 233660 224680 233666 224732
rect 351270 224680 351276 224732
rect 351328 224720 351334 224732
rect 425348 224720 425376 224760
rect 425514 224748 425520 224760
rect 425572 224748 425578 224800
rect 429102 224748 429108 224800
rect 429160 224788 429166 224800
rect 441614 224788 441620 224800
rect 429160 224760 441620 224788
rect 429160 224748 429166 224760
rect 441614 224748 441620 224760
rect 441672 224748 441678 224800
rect 351328 224692 425376 224720
rect 351328 224680 351334 224692
rect 425422 224680 425428 224732
rect 425480 224720 425486 224732
rect 460934 224720 460940 224732
rect 425480 224692 460940 224720
rect 425480 224680 425486 224692
rect 460934 224680 460940 224692
rect 460992 224680 460998 224732
rect 161198 224612 161204 224664
rect 161256 224652 161262 224664
rect 237926 224652 237932 224664
rect 161256 224624 237932 224652
rect 161256 224612 161262 224624
rect 237926 224612 237932 224624
rect 237984 224612 237990 224664
rect 349798 224612 349804 224664
rect 349856 224652 349862 224664
rect 401502 224652 401508 224664
rect 349856 224624 401508 224652
rect 349856 224612 349862 224624
rect 401502 224612 401508 224624
rect 401560 224612 401566 224664
rect 416682 224612 416688 224664
rect 416740 224652 416746 224664
rect 417970 224652 417976 224664
rect 416740 224624 417976 224652
rect 416740 224612 416746 224624
rect 417970 224612 417976 224624
rect 418028 224612 418034 224664
rect 422294 224612 422300 224664
rect 422352 224652 422358 224664
rect 457438 224652 457444 224664
rect 422352 224624 457444 224652
rect 422352 224612 422358 224624
rect 457438 224612 457444 224624
rect 457496 224612 457502 224664
rect 157794 224544 157800 224596
rect 157852 224584 157858 224596
rect 236454 224584 236460 224596
rect 157852 224556 236460 224584
rect 157852 224544 157858 224556
rect 236454 224544 236460 224556
rect 236512 224544 236518 224596
rect 342714 224544 342720 224596
rect 342772 224584 342778 224596
rect 405642 224584 405648 224596
rect 342772 224556 405648 224584
rect 342772 224544 342778 224556
rect 405642 224544 405648 224556
rect 405700 224544 405706 224596
rect 405734 224544 405740 224596
rect 405792 224584 405798 224596
rect 479334 224584 479340 224596
rect 405792 224556 479340 224584
rect 405792 224544 405798 224556
rect 479334 224544 479340 224556
rect 479392 224544 479398 224596
rect 169110 224476 169116 224528
rect 169168 224516 169174 224528
rect 240778 224516 240784 224528
rect 169168 224488 240784 224516
rect 169168 224476 169174 224488
rect 240778 224476 240784 224488
rect 240836 224476 240842 224528
rect 348050 224476 348056 224528
rect 348108 224516 348114 224528
rect 421282 224516 421288 224528
rect 348108 224488 421288 224516
rect 348108 224476 348114 224488
rect 421282 224476 421288 224488
rect 421340 224476 421346 224528
rect 425238 224476 425244 224528
rect 425296 224516 425302 224528
rect 432230 224516 432236 224528
rect 425296 224488 432236 224516
rect 425296 224476 425302 224488
rect 432230 224476 432236 224488
rect 432288 224476 432294 224528
rect 166350 224408 166356 224460
rect 166408 224448 166414 224460
rect 239306 224448 239312 224460
rect 166408 224420 239312 224448
rect 166408 224408 166414 224420
rect 239306 224408 239312 224420
rect 239364 224408 239370 224460
rect 346946 224408 346952 224460
rect 347004 224448 347010 224460
rect 415394 224448 415400 224460
rect 347004 224420 415400 224448
rect 347004 224408 347010 224420
rect 415394 224408 415400 224420
rect 415452 224408 415458 224460
rect 416866 224408 416872 224460
rect 416924 224448 416930 224460
rect 450722 224448 450728 224460
rect 416924 224420 450728 224448
rect 416924 224408 416930 224420
rect 450722 224408 450728 224420
rect 450780 224408 450786 224460
rect 171042 224340 171048 224392
rect 171100 224380 171106 224392
rect 242158 224380 242164 224392
rect 171100 224352 242164 224380
rect 171100 224340 171106 224352
rect 242158 224340 242164 224352
rect 242216 224340 242222 224392
rect 348418 224340 348424 224392
rect 348476 224380 348482 224392
rect 418798 224380 418804 224392
rect 348476 224352 418804 224380
rect 348476 224340 348482 224352
rect 418798 224340 418804 224352
rect 418856 224340 418862 224392
rect 176654 224272 176660 224324
rect 176712 224312 176718 224324
rect 243630 224312 243636 224324
rect 176712 224284 243636 224312
rect 176712 224272 176718 224284
rect 243630 224272 243636 224284
rect 243688 224272 243694 224324
rect 345198 224272 345204 224324
rect 345256 224312 345262 224324
rect 414566 224312 414572 224324
rect 345256 224284 414572 224312
rect 345256 224272 345262 224284
rect 414566 224272 414572 224284
rect 414624 224272 414630 224324
rect 415302 224272 415308 224324
rect 415360 224312 415366 224324
rect 444374 224312 444380 224324
rect 415360 224284 444380 224312
rect 415360 224272 415366 224284
rect 444374 224272 444380 224284
rect 444432 224272 444438 224324
rect 181346 224204 181352 224256
rect 181404 224244 181410 224256
rect 246482 224244 246488 224256
rect 181404 224216 246488 224244
rect 181404 224204 181410 224216
rect 246482 224204 246488 224216
rect 246540 224204 246546 224256
rect 345566 224204 345572 224256
rect 345624 224244 345630 224256
rect 412082 224244 412088 224256
rect 345624 224216 412088 224244
rect 345624 224204 345630 224216
rect 412082 224204 412088 224216
rect 412140 224204 412146 224256
rect 413186 224204 413192 224256
rect 413244 224244 413250 224256
rect 430574 224244 430580 224256
rect 413244 224216 430580 224244
rect 413244 224204 413250 224216
rect 430574 224204 430580 224216
rect 430632 224204 430638 224256
rect 178034 224136 178040 224188
rect 178092 224176 178098 224188
rect 245010 224176 245016 224188
rect 178092 224148 245016 224176
rect 178092 224136 178098 224148
rect 245010 224136 245016 224148
rect 245068 224136 245074 224188
rect 344094 224136 344100 224188
rect 344152 224176 344158 224188
rect 408678 224176 408684 224188
rect 344152 224148 408684 224176
rect 344152 224136 344158 224148
rect 408678 224136 408684 224148
rect 408736 224136 408742 224188
rect 408770 224136 408776 224188
rect 408828 224176 408834 224188
rect 465902 224176 465908 224188
rect 408828 224148 465908 224176
rect 408828 224136 408834 224148
rect 465902 224136 465908 224148
rect 465960 224136 465966 224188
rect 184750 224068 184756 224120
rect 184808 224108 184814 224120
rect 247862 224108 247868 224120
rect 184808 224080 247868 224108
rect 184808 224068 184814 224080
rect 247862 224068 247868 224080
rect 247920 224068 247926 224120
rect 340230 224068 340236 224120
rect 340288 224108 340294 224120
rect 400398 224108 400404 224120
rect 340288 224080 400404 224108
rect 340288 224068 340294 224080
rect 400398 224068 400404 224080
rect 400456 224068 400462 224120
rect 405826 224068 405832 224120
rect 405884 224108 405890 224120
rect 459186 224108 459192 224120
rect 405884 224080 459192 224108
rect 405884 224068 405890 224080
rect 459186 224068 459192 224080
rect 459244 224068 459250 224120
rect 146294 224000 146300 224052
rect 146352 224040 146358 224052
rect 146352 224012 168374 224040
rect 146352 224000 146358 224012
rect 168346 223700 168374 224012
rect 197446 224000 197452 224052
rect 197504 224040 197510 224052
rect 212258 224040 212264 224052
rect 197504 224012 212264 224040
rect 197504 224000 197510 224012
rect 212258 224000 212264 224012
rect 212316 224000 212322 224052
rect 216122 224000 216128 224052
rect 216180 224040 216186 224052
rect 246758 224040 246764 224052
rect 216180 224012 246764 224040
rect 216180 224000 216186 224012
rect 246758 224000 246764 224012
rect 246816 224000 246822 224052
rect 383746 224000 383752 224052
rect 383804 224040 383810 224052
rect 404446 224040 404452 224052
rect 383804 224012 404452 224040
rect 383804 224000 383810 224012
rect 404446 224000 404452 224012
rect 404504 224000 404510 224052
rect 404538 224000 404544 224052
rect 404596 224040 404602 224052
rect 445662 224040 445668 224052
rect 404596 224012 445668 224040
rect 404596 224000 404602 224012
rect 445662 224000 445668 224012
rect 445720 224000 445726 224052
rect 188154 223932 188160 223984
rect 188212 223972 188218 223984
rect 249334 223972 249340 223984
rect 188212 223944 249340 223972
rect 188212 223932 188218 223944
rect 249334 223932 249340 223944
rect 249392 223932 249398 223984
rect 378134 223932 378140 223984
rect 378192 223972 378198 223984
rect 378192 223944 399892 223972
rect 378192 223932 378198 223944
rect 204898 223864 204904 223916
rect 204956 223904 204962 223916
rect 256418 223904 256424 223916
rect 204956 223876 256424 223904
rect 204956 223864 204962 223876
rect 256418 223864 256424 223876
rect 256476 223864 256482 223916
rect 380894 223864 380900 223916
rect 380952 223904 380958 223916
rect 399864 223904 399892 223944
rect 401502 223932 401508 223984
rect 401560 223972 401566 223984
rect 422294 223972 422300 223984
rect 401560 223944 422300 223972
rect 401560 223932 401566 223944
rect 422294 223932 422300 223944
rect 422352 223932 422358 223984
rect 380952 223876 391934 223904
rect 399864 223876 411254 223904
rect 380952 223864 380958 223876
rect 188430 223796 188436 223848
rect 188488 223836 188494 223848
rect 232498 223836 232504 223848
rect 188488 223808 232504 223836
rect 188488 223796 188494 223808
rect 232498 223796 232504 223808
rect 232556 223796 232562 223848
rect 391906 223836 391934 223876
rect 411226 223848 411254 223876
rect 407850 223836 407856 223848
rect 391906 223808 407856 223836
rect 407850 223796 407856 223808
rect 407908 223796 407914 223848
rect 411226 223808 411260 223848
rect 411254 223796 411260 223808
rect 411312 223796 411318 223848
rect 191466 223728 191472 223780
rect 191524 223768 191530 223780
rect 206922 223768 206928 223780
rect 191524 223740 206928 223768
rect 191524 223728 191530 223740
rect 206922 223728 206928 223740
rect 206980 223728 206986 223780
rect 208946 223728 208952 223780
rect 209004 223768 209010 223780
rect 239674 223768 239680 223780
rect 209004 223740 239680 223768
rect 209004 223728 209010 223740
rect 239674 223728 239680 223740
rect 239732 223728 239738 223780
rect 168346 223672 189396 223700
rect 185578 223592 185584 223644
rect 185636 223632 185642 223644
rect 189258 223632 189264 223644
rect 185636 223604 189264 223632
rect 185636 223592 185642 223604
rect 189258 223592 189264 223604
rect 189316 223592 189322 223644
rect 189368 223632 189396 223672
rect 209682 223660 209688 223712
rect 209740 223700 209746 223712
rect 236822 223700 236828 223712
rect 209740 223672 236828 223700
rect 209740 223660 209746 223672
rect 236822 223660 236828 223672
rect 236880 223660 236886 223712
rect 209406 223632 209412 223644
rect 189368 223604 209412 223632
rect 209406 223592 209412 223604
rect 209464 223592 209470 223644
rect 214926 223592 214932 223644
rect 214984 223632 214990 223644
rect 242526 223632 242532 223644
rect 214984 223604 242532 223632
rect 214984 223592 214990 223604
rect 242526 223592 242532 223604
rect 242584 223592 242590 223644
rect 408494 223592 408500 223644
rect 408552 223632 408558 223644
rect 423858 223632 423864 223644
rect 408552 223604 423864 223632
rect 408552 223592 408558 223604
rect 423858 223592 423864 223604
rect 423916 223592 423922 223644
rect 480254 223592 480260 223644
rect 480312 223632 480318 223644
rect 484394 223632 484400 223644
rect 480312 223604 484400 223632
rect 480312 223592 480318 223604
rect 484394 223592 484400 223604
rect 484452 223592 484458 223644
rect 155310 223524 155316 223576
rect 155368 223564 155374 223576
rect 236086 223564 236092 223576
rect 155368 223536 236092 223564
rect 155368 223524 155374 223536
rect 236086 223524 236092 223536
rect 236144 223524 236150 223576
rect 278682 223524 278688 223576
rect 278740 223564 278746 223576
rect 287790 223564 287796 223576
rect 278740 223536 287796 223564
rect 278740 223524 278746 223536
rect 287790 223524 287796 223536
rect 287848 223524 287854 223576
rect 324498 223524 324504 223576
rect 324556 223564 324562 223576
rect 363230 223564 363236 223576
rect 324556 223536 363236 223564
rect 324556 223524 324562 223536
rect 363230 223524 363236 223536
rect 363288 223524 363294 223576
rect 392946 223524 392952 223576
rect 393004 223564 393010 223576
rect 395246 223564 395252 223576
rect 393004 223536 395252 223564
rect 393004 223524 393010 223536
rect 395246 223524 395252 223536
rect 395304 223524 395310 223576
rect 402974 223524 402980 223576
rect 403032 223564 403038 223576
rect 406194 223564 406200 223576
rect 403032 223536 406200 223564
rect 403032 223524 403038 223536
rect 406194 223524 406200 223536
rect 406252 223524 406258 223576
rect 503806 223524 503812 223576
rect 503864 223564 503870 223576
rect 623406 223564 623412 223576
rect 503864 223536 623412 223564
rect 503864 223524 503870 223536
rect 623406 223524 623412 223536
rect 623464 223524 623470 223576
rect 93762 223456 93768 223508
rect 93820 223496 93826 223508
rect 146294 223496 146300 223508
rect 93820 223468 146300 223496
rect 93820 223456 93826 223468
rect 146294 223456 146300 223468
rect 146352 223456 146358 223508
rect 153654 223456 153660 223508
rect 153712 223496 153718 223508
rect 235718 223496 235724 223508
rect 153712 223468 235724 223496
rect 153712 223456 153718 223468
rect 235718 223456 235724 223468
rect 235776 223456 235782 223508
rect 241146 223456 241152 223508
rect 241204 223496 241210 223508
rect 253566 223496 253572 223508
rect 241204 223468 253572 223496
rect 241204 223456 241210 223468
rect 253566 223456 253572 223468
rect 253624 223456 253630 223508
rect 322382 223456 322388 223508
rect 322440 223496 322446 223508
rect 360746 223496 360752 223508
rect 322440 223468 360752 223496
rect 322440 223456 322446 223468
rect 360746 223456 360752 223468
rect 360804 223456 360810 223508
rect 494054 223456 494060 223508
rect 494112 223496 494118 223508
rect 607582 223496 607588 223508
rect 494112 223468 607588 223496
rect 494112 223456 494118 223468
rect 607582 223456 607588 223468
rect 607640 223456 607646 223508
rect 146938 223388 146944 223440
rect 146996 223428 147002 223440
rect 232866 223428 232872 223440
rect 146996 223400 232872 223428
rect 146996 223388 147002 223400
rect 232866 223388 232872 223400
rect 232924 223388 232930 223440
rect 324130 223388 324136 223440
rect 324188 223428 324194 223440
rect 361758 223428 361764 223440
rect 324188 223400 361764 223428
rect 324188 223388 324194 223400
rect 361758 223388 361764 223400
rect 361816 223388 361822 223440
rect 397270 223388 397276 223440
rect 397328 223428 397334 223440
rect 406562 223428 406568 223440
rect 397328 223400 406568 223428
rect 397328 223388 397334 223400
rect 406562 223388 406568 223400
rect 406620 223388 406626 223440
rect 499482 223388 499488 223440
rect 499540 223428 499546 223440
rect 608042 223428 608048 223440
rect 499540 223400 608048 223428
rect 499540 223388 499546 223400
rect 608042 223388 608048 223400
rect 608100 223388 608106 223440
rect 148594 223320 148600 223372
rect 148652 223360 148658 223372
rect 233234 223360 233240 223372
rect 148652 223332 233240 223360
rect 148652 223320 148658 223332
rect 233234 223320 233240 223332
rect 233292 223320 233298 223372
rect 237742 223320 237748 223372
rect 237800 223360 237806 223372
rect 253198 223360 253204 223372
rect 237800 223332 253204 223360
rect 237800 223320 237806 223332
rect 253198 223320 253204 223332
rect 253256 223320 253262 223372
rect 324866 223320 324872 223372
rect 324924 223360 324930 223372
rect 365806 223360 365812 223372
rect 324924 223332 365812 223360
rect 324924 223320 324930 223332
rect 365806 223320 365812 223332
rect 365864 223320 365870 223372
rect 398282 223320 398288 223372
rect 398340 223360 398346 223372
rect 539042 223360 539048 223372
rect 398340 223332 539048 223360
rect 398340 223320 398346 223332
rect 539042 223320 539048 223332
rect 539100 223320 539106 223372
rect 87138 223252 87144 223304
rect 87196 223292 87202 223304
rect 172422 223292 172428 223304
rect 87196 223264 172428 223292
rect 87196 223252 87202 223264
rect 172422 223252 172428 223264
rect 172480 223252 172486 223304
rect 175458 223252 175464 223304
rect 175516 223292 175522 223304
rect 244642 223292 244648 223304
rect 175516 223264 244648 223292
rect 175516 223252 175522 223264
rect 244642 223252 244648 223264
rect 244700 223252 244706 223304
rect 326982 223252 326988 223304
rect 327040 223292 327046 223304
rect 368290 223292 368296 223304
rect 327040 223264 368296 223292
rect 327040 223252 327046 223264
rect 368290 223252 368296 223264
rect 368348 223252 368354 223304
rect 399018 223252 399024 223304
rect 399076 223292 399082 223304
rect 536282 223292 536288 223304
rect 399076 223264 536288 223292
rect 399076 223252 399082 223264
rect 536282 223252 536288 223264
rect 536340 223252 536346 223304
rect 536374 223252 536380 223304
rect 536432 223292 536438 223304
rect 536432 223264 536696 223292
rect 536432 223252 536438 223264
rect 536668 223236 536696 223264
rect 141878 223184 141884 223236
rect 141936 223224 141942 223236
rect 230382 223224 230388 223236
rect 141936 223196 230388 223224
rect 141936 223184 141942 223196
rect 230382 223184 230388 223196
rect 230440 223184 230446 223236
rect 239398 223184 239404 223236
rect 239456 223224 239462 223236
rect 255498 223224 255504 223236
rect 239456 223196 255504 223224
rect 239456 223184 239462 223196
rect 255498 223184 255504 223196
rect 255556 223184 255562 223236
rect 326338 223184 326344 223236
rect 326396 223224 326402 223236
rect 369118 223224 369124 223236
rect 326396 223196 369124 223224
rect 326396 223184 326402 223196
rect 369118 223184 369124 223196
rect 369176 223184 369182 223236
rect 400122 223184 400128 223236
rect 400180 223224 400186 223236
rect 406470 223224 406476 223236
rect 400180 223196 406476 223224
rect 400180 223184 400186 223196
rect 406470 223184 406476 223196
rect 406528 223184 406534 223236
rect 406562 223184 406568 223236
rect 406620 223224 406626 223236
rect 536558 223224 536564 223236
rect 406620 223196 536564 223224
rect 406620 223184 406626 223196
rect 536558 223184 536564 223196
rect 536616 223184 536622 223236
rect 536650 223184 536656 223236
rect 536708 223224 536714 223236
rect 615034 223224 615040 223236
rect 536708 223196 615040 223224
rect 536708 223184 536714 223196
rect 615034 223184 615040 223196
rect 615092 223184 615098 223236
rect 140130 223116 140136 223168
rect 140188 223156 140194 223168
rect 230014 223156 230020 223168
rect 140188 223128 230020 223156
rect 140188 223116 140194 223128
rect 230014 223116 230020 223128
rect 230072 223116 230078 223168
rect 235902 223116 235908 223168
rect 235960 223156 235966 223168
rect 249978 223156 249984 223168
rect 235960 223128 249984 223156
rect 235960 223116 235966 223128
rect 249978 223116 249984 223128
rect 250036 223116 250042 223168
rect 325602 223116 325608 223168
rect 325660 223156 325666 223168
rect 364978 223156 364984 223168
rect 325660 223128 364984 223156
rect 325660 223116 325666 223128
rect 364978 223116 364984 223128
rect 365036 223116 365042 223168
rect 399386 223116 399392 223168
rect 399444 223156 399450 223168
rect 541618 223156 541624 223168
rect 399444 223128 541624 223156
rect 399444 223116 399450 223128
rect 541618 223116 541624 223128
rect 541676 223116 541682 223168
rect 135162 223048 135168 223100
rect 135220 223088 135226 223100
rect 227530 223088 227536 223100
rect 135220 223060 227536 223088
rect 135220 223048 135226 223060
rect 227530 223048 227536 223060
rect 227588 223048 227594 223100
rect 232590 223048 232596 223100
rect 232648 223088 232654 223100
rect 242710 223088 242716 223100
rect 232648 223060 242716 223088
rect 232648 223048 232654 223060
rect 242710 223048 242716 223060
rect 242768 223048 242774 223100
rect 242802 223048 242808 223100
rect 242860 223088 242866 223100
rect 258810 223088 258816 223100
rect 242860 223060 258816 223088
rect 242860 223048 242866 223060
rect 258810 223048 258816 223060
rect 258868 223048 258874 223100
rect 271414 223048 271420 223100
rect 271472 223088 271478 223100
rect 285674 223088 285680 223100
rect 271472 223060 285680 223088
rect 271472 223048 271478 223060
rect 285674 223048 285680 223060
rect 285732 223048 285738 223100
rect 328454 223048 328460 223100
rect 328512 223088 328518 223100
rect 371694 223088 371700 223100
rect 328512 223060 371700 223088
rect 328512 223048 328518 223060
rect 371694 223048 371700 223060
rect 371752 223048 371758 223100
rect 400766 223048 400772 223100
rect 400824 223088 400830 223100
rect 545114 223088 545120 223100
rect 400824 223060 545120 223088
rect 400824 223048 400830 223060
rect 545114 223048 545120 223060
rect 545172 223048 545178 223100
rect 545758 223048 545764 223100
rect 545816 223088 545822 223100
rect 616874 223088 616880 223100
rect 545816 223060 616880 223088
rect 545816 223048 545822 223060
rect 616874 223048 616880 223060
rect 616932 223048 616938 223100
rect 133414 222980 133420 223032
rect 133472 223020 133478 223032
rect 227162 223020 227168 223032
rect 133472 222992 227168 223020
rect 133472 222980 133478 222992
rect 227162 222980 227168 222992
rect 227220 222980 227226 223032
rect 231026 222980 231032 223032
rect 231084 223020 231090 223032
rect 248506 223020 248512 223032
rect 231084 222992 248512 223020
rect 231084 222980 231090 222992
rect 248506 222980 248512 222992
rect 248564 222980 248570 223032
rect 323762 222980 323768 223032
rect 323820 223020 323826 223032
rect 364334 223020 364340 223032
rect 323820 222992 364340 223020
rect 323820 222980 323826 222992
rect 364334 222980 364340 222992
rect 364392 222980 364398 223032
rect 372062 222980 372068 223032
rect 372120 223020 372126 223032
rect 397730 223020 397736 223032
rect 372120 222992 397736 223020
rect 372120 222980 372126 222992
rect 397730 222980 397736 222992
rect 397788 222980 397794 223032
rect 401778 222980 401784 223032
rect 401836 223020 401842 223032
rect 401836 222992 406424 223020
rect 401836 222980 401842 222992
rect 128354 222912 128360 222964
rect 128412 222952 128418 222964
rect 224678 222952 224684 222964
rect 128412 222924 224684 222952
rect 128412 222912 128418 222924
rect 224678 222912 224684 222924
rect 224736 222912 224742 222964
rect 236086 222912 236092 222964
rect 236144 222952 236150 222964
rect 255314 222952 255320 222964
rect 236144 222924 255320 222952
rect 236144 222912 236150 222924
rect 255314 222912 255320 222924
rect 255372 222912 255378 222964
rect 263778 222912 263784 222964
rect 263836 222952 263842 222964
rect 280982 222952 280988 222964
rect 263836 222924 280988 222952
rect 263836 222912 263842 222924
rect 280982 222912 280988 222924
rect 281040 222912 281046 222964
rect 327350 222912 327356 222964
rect 327408 222952 327414 222964
rect 370038 222952 370044 222964
rect 327408 222924 370044 222952
rect 327408 222912 327414 222924
rect 370038 222912 370044 222924
rect 370096 222912 370102 222964
rect 396534 222912 396540 222964
rect 396592 222952 396598 222964
rect 401962 222952 401968 222964
rect 396592 222924 401968 222952
rect 396592 222912 396598 222924
rect 401962 222912 401968 222924
rect 402020 222912 402026 222964
rect 406396 222952 406424 222992
rect 406470 222980 406476 223032
rect 406528 223020 406534 223032
rect 543550 223020 543556 223032
rect 406528 222992 543556 223020
rect 406528 222980 406534 222992
rect 543550 222980 543556 222992
rect 543608 222980 543614 223032
rect 617334 223020 617340 223032
rect 548352 222992 617340 223020
rect 546678 222952 546684 222964
rect 406396 222924 546684 222952
rect 546678 222912 546684 222924
rect 546736 222912 546742 222964
rect 548352 222896 548380 222992
rect 617334 222980 617340 222992
rect 617392 222980 617398 223032
rect 565998 222912 566004 222964
rect 566056 222952 566062 222964
rect 620554 222952 620560 222964
rect 566056 222924 620560 222952
rect 566056 222912 566062 222924
rect 620554 222912 620560 222924
rect 620612 222912 620618 222964
rect 126698 222844 126704 222896
rect 126756 222884 126762 222896
rect 224034 222884 224040 222896
rect 126756 222856 224040 222884
rect 126756 222844 126762 222856
rect 224034 222844 224040 222856
rect 224092 222844 224098 222896
rect 232682 222844 232688 222896
rect 232740 222884 232746 222896
rect 255774 222884 255780 222896
rect 232740 222856 255780 222884
rect 232740 222844 232746 222856
rect 255774 222844 255780 222856
rect 255832 222844 255838 222896
rect 257062 222844 257068 222896
rect 257120 222884 257126 222896
rect 278130 222884 278136 222896
rect 257120 222856 278136 222884
rect 257120 222844 257126 222856
rect 278130 222844 278136 222856
rect 278188 222844 278194 222896
rect 325234 222844 325240 222896
rect 325292 222884 325298 222896
rect 367462 222884 367468 222896
rect 325292 222856 367468 222884
rect 325292 222844 325298 222856
rect 367462 222844 367468 222856
rect 367520 222844 367526 222896
rect 368566 222844 368572 222896
rect 368624 222884 368630 222896
rect 398558 222884 398564 222896
rect 368624 222856 398564 222884
rect 368624 222844 368630 222856
rect 398558 222844 398564 222856
rect 398616 222844 398622 222896
rect 402238 222844 402244 222896
rect 402296 222884 402302 222896
rect 548334 222884 548340 222896
rect 402296 222856 548340 222884
rect 402296 222844 402302 222856
rect 548334 222844 548340 222856
rect 548392 222844 548398 222896
rect 549346 222844 549352 222896
rect 549404 222884 549410 222896
rect 551094 222884 551100 222896
rect 549404 222856 551100 222884
rect 549404 222844 549410 222856
rect 551094 222844 551100 222856
rect 551152 222884 551158 222896
rect 617794 222884 617800 222896
rect 551152 222856 617800 222884
rect 551152 222844 551158 222856
rect 617794 222844 617800 222856
rect 617852 222844 617858 222896
rect 66990 222776 66996 222828
rect 67048 222816 67054 222828
rect 114278 222816 114284 222828
rect 67048 222788 114284 222816
rect 67048 222776 67054 222788
rect 114278 222776 114284 222788
rect 114336 222776 114342 222828
rect 116578 222776 116584 222828
rect 116636 222816 116642 222828
rect 220078 222816 220084 222828
rect 116636 222788 220084 222816
rect 116636 222776 116642 222788
rect 220078 222776 220084 222788
rect 220136 222776 220142 222828
rect 224310 222776 224316 222828
rect 224368 222816 224374 222828
rect 248414 222816 248420 222828
rect 224368 222788 248420 222816
rect 224368 222776 224374 222788
rect 248414 222776 248420 222788
rect 248472 222776 248478 222828
rect 264606 222776 264612 222828
rect 264664 222816 264670 222828
rect 282822 222816 282828 222828
rect 264664 222788 282828 222816
rect 264664 222776 264670 222788
rect 282822 222776 282828 222788
rect 282880 222776 282886 222828
rect 326614 222776 326620 222828
rect 326672 222816 326678 222828
rect 370866 222816 370872 222828
rect 326672 222788 370872 222816
rect 326672 222776 326678 222788
rect 370866 222776 370872 222788
rect 370924 222776 370930 222828
rect 401870 222776 401876 222828
rect 401928 222816 401934 222828
rect 547506 222816 547512 222828
rect 401928 222788 547512 222816
rect 401928 222776 401934 222788
rect 547506 222776 547512 222788
rect 547564 222776 547570 222828
rect 553762 222776 553768 222828
rect 553820 222816 553826 222828
rect 553820 222788 554360 222816
rect 553820 222776 553826 222788
rect 554332 222760 554360 222788
rect 91370 222708 91376 222760
rect 91428 222748 91434 222760
rect 201586 222748 201592 222760
rect 91428 222720 201592 222748
rect 91428 222708 91434 222720
rect 201586 222708 201592 222720
rect 201644 222708 201650 222760
rect 214190 222708 214196 222760
rect 214248 222748 214254 222760
rect 245654 222748 245660 222760
rect 214248 222720 245660 222748
rect 214248 222708 214254 222720
rect 245654 222708 245660 222720
rect 245712 222708 245718 222760
rect 246114 222708 246120 222760
rect 246172 222748 246178 222760
rect 258718 222748 258724 222760
rect 246172 222720 258724 222748
rect 246172 222708 246178 222720
rect 258718 222708 258724 222720
rect 258776 222708 258782 222760
rect 262950 222708 262956 222760
rect 263008 222748 263014 222760
rect 281718 222748 281724 222760
rect 263008 222720 281724 222748
rect 263008 222708 263014 222720
rect 281718 222708 281724 222720
rect 281776 222708 281782 222760
rect 327718 222708 327724 222760
rect 327776 222748 327782 222760
rect 372614 222748 372620 222760
rect 327776 222720 372620 222748
rect 327776 222708 327782 222720
rect 372614 222708 372620 222720
rect 372672 222708 372678 222760
rect 373994 222708 374000 222760
rect 374052 222748 374058 222760
rect 391014 222748 391020 222760
rect 374052 222720 391020 222748
rect 374052 222708 374058 222720
rect 391014 222708 391020 222720
rect 391072 222708 391078 222760
rect 404722 222708 404728 222760
rect 404780 222748 404786 222760
rect 554222 222748 554228 222760
rect 404780 222720 554228 222748
rect 404780 222708 404786 222720
rect 554222 222708 554228 222720
rect 554280 222708 554286 222760
rect 554314 222708 554320 222760
rect 554372 222748 554378 222760
rect 618254 222748 618260 222760
rect 554372 222720 618260 222748
rect 554372 222708 554378 222720
rect 618254 222708 618260 222720
rect 618312 222708 618318 222760
rect 89714 222640 89720 222692
rect 89772 222680 89778 222692
rect 201678 222680 201684 222692
rect 89772 222652 201684 222680
rect 89772 222640 89778 222652
rect 201678 222640 201684 222652
rect 201736 222640 201742 222692
rect 222562 222640 222568 222692
rect 222620 222680 222626 222692
rect 258166 222680 258172 222692
rect 222620 222652 258172 222680
rect 222620 222640 222626 222652
rect 258166 222640 258172 222652
rect 258224 222640 258230 222692
rect 260466 222640 260472 222692
rect 260524 222680 260530 222692
rect 279602 222680 279608 222692
rect 260524 222652 279608 222680
rect 260524 222640 260530 222652
rect 279602 222640 279608 222652
rect 279660 222640 279666 222692
rect 329466 222640 329472 222692
rect 329524 222680 329530 222692
rect 377582 222680 377588 222692
rect 329524 222652 377588 222680
rect 329524 222640 329530 222652
rect 377582 222640 377588 222652
rect 377640 222640 377646 222692
rect 391750 222640 391756 222692
rect 391808 222680 391814 222692
rect 402974 222680 402980 222692
rect 391808 222652 402980 222680
rect 391808 222640 391814 222652
rect 402974 222640 402980 222652
rect 403032 222640 403038 222692
rect 406102 222640 406108 222692
rect 406160 222680 406166 222692
rect 556706 222680 556712 222692
rect 406160 222652 556712 222680
rect 406160 222640 406166 222652
rect 556706 222640 556712 222652
rect 556764 222640 556770 222692
rect 568574 222640 568580 222692
rect 568632 222680 568638 222692
rect 621014 222680 621020 222692
rect 568632 222652 621020 222680
rect 568632 222640 568638 222652
rect 621014 222640 621020 222652
rect 621072 222640 621078 222692
rect 82170 222572 82176 222624
rect 82228 222612 82234 222624
rect 198734 222612 198740 222624
rect 82228 222584 198740 222612
rect 82228 222572 82234 222584
rect 198734 222572 198740 222584
rect 198792 222572 198798 222624
rect 207474 222572 207480 222624
rect 207532 222612 207538 222624
rect 246206 222612 246212 222624
rect 207532 222584 246212 222612
rect 207532 222572 207538 222584
rect 246206 222572 246212 222584
rect 246264 222572 246270 222624
rect 259362 222572 259368 222624
rect 259420 222612 259426 222624
rect 280338 222612 280344 222624
rect 259420 222584 280344 222612
rect 259420 222572 259426 222584
rect 280338 222572 280344 222584
rect 280396 222572 280402 222624
rect 329834 222572 329840 222624
rect 329892 222612 329898 222624
rect 375374 222612 375380 222624
rect 329892 222584 375380 222612
rect 329892 222572 329898 222584
rect 375374 222572 375380 222584
rect 375432 222572 375438 222624
rect 405090 222572 405096 222624
rect 405148 222612 405154 222624
rect 555050 222612 555056 222624
rect 405148 222584 555056 222612
rect 405148 222572 405154 222584
rect 555050 222572 555056 222584
rect 555108 222572 555114 222624
rect 556062 222572 556068 222624
rect 556120 222612 556126 222624
rect 618714 222612 618720 222624
rect 556120 222584 618720 222612
rect 556120 222572 556126 222584
rect 618714 222572 618720 222584
rect 618772 222572 618778 222624
rect 85482 222504 85488 222556
rect 85540 222544 85546 222556
rect 205450 222544 205456 222556
rect 85540 222516 205456 222544
rect 85540 222504 85546 222516
rect 205450 222504 205456 222516
rect 205508 222504 205514 222556
rect 215846 222504 215852 222556
rect 215904 222544 215910 222556
rect 259178 222544 259184 222556
rect 215904 222516 259184 222544
rect 215904 222504 215910 222516
rect 259178 222504 259184 222516
rect 259236 222504 259242 222556
rect 261294 222504 261300 222556
rect 261352 222544 261358 222556
rect 281350 222544 281356 222556
rect 261352 222516 281356 222544
rect 261352 222504 261358 222516
rect 281350 222504 281356 222516
rect 281408 222504 281414 222556
rect 284938 222544 284944 222556
rect 281460 222516 284944 222544
rect 81250 222436 81256 222488
rect 81308 222476 81314 222488
rect 204714 222476 204720 222488
rect 81308 222448 204720 222476
rect 81308 222436 81314 222448
rect 204714 222436 204720 222448
rect 204772 222436 204778 222488
rect 209130 222436 209136 222488
rect 209188 222476 209194 222488
rect 258626 222476 258632 222488
rect 209188 222448 258632 222476
rect 209188 222436 209194 222448
rect 258626 222436 258632 222448
rect 258684 222436 258690 222488
rect 262122 222436 262128 222488
rect 262180 222476 262186 222488
rect 280706 222476 280712 222488
rect 262180 222448 280712 222476
rect 262180 222436 262186 222448
rect 280706 222436 280712 222448
rect 280764 222436 280770 222488
rect 75362 222368 75368 222420
rect 75420 222408 75426 222420
rect 201126 222408 201132 222420
rect 75420 222380 201132 222408
rect 75420 222368 75426 222380
rect 201126 222368 201132 222380
rect 201184 222368 201190 222420
rect 205818 222368 205824 222420
rect 205876 222408 205882 222420
rect 257522 222408 257528 222420
rect 205876 222380 257528 222408
rect 205876 222368 205882 222380
rect 257522 222368 257528 222380
rect 257580 222368 257586 222420
rect 272242 222368 272248 222420
rect 272300 222408 272306 222420
rect 281460 222408 281488 222516
rect 284938 222504 284944 222516
rect 284996 222504 285002 222556
rect 331582 222504 331588 222556
rect 331640 222544 331646 222556
rect 378410 222544 378416 222556
rect 331640 222516 378416 222544
rect 331640 222504 331646 222516
rect 378410 222504 378416 222516
rect 378468 222504 378474 222556
rect 378502 222504 378508 222556
rect 378560 222544 378566 222556
rect 392670 222544 392676 222556
rect 378560 222516 392676 222544
rect 378560 222504 378566 222516
rect 392670 222504 392676 222516
rect 392728 222504 392734 222556
rect 406378 222504 406384 222556
rect 406436 222544 406442 222556
rect 558178 222544 558184 222556
rect 406436 222516 558184 222544
rect 406436 222504 406442 222516
rect 558178 222504 558184 222516
rect 558236 222504 558242 222556
rect 559098 222504 559104 222556
rect 559156 222544 559162 222556
rect 619174 222544 619180 222556
rect 559156 222516 619180 222544
rect 559156 222504 559162 222516
rect 619174 222504 619180 222516
rect 619232 222504 619238 222556
rect 283098 222436 283104 222488
rect 283156 222476 283162 222488
rect 290274 222476 290280 222488
rect 283156 222448 290280 222476
rect 283156 222436 283162 222448
rect 290274 222436 290280 222448
rect 290332 222436 290338 222488
rect 338298 222436 338304 222488
rect 338356 222476 338362 222488
rect 343082 222476 343088 222488
rect 338356 222448 343088 222476
rect 338356 222436 338362 222448
rect 343082 222436 343088 222448
rect 343140 222436 343146 222488
rect 343542 222436 343548 222488
rect 343600 222476 343606 222488
rect 376754 222476 376760 222488
rect 343600 222448 376760 222476
rect 343600 222436 343606 222448
rect 376754 222436 376760 222448
rect 376812 222436 376818 222488
rect 377030 222436 377036 222488
rect 377088 222476 377094 222488
rect 399478 222476 399484 222488
rect 377088 222448 399484 222476
rect 377088 222436 377094 222448
rect 399478 222436 399484 222448
rect 399536 222436 399542 222488
rect 407942 222436 407948 222488
rect 408000 222476 408006 222488
rect 561766 222476 561772 222488
rect 408000 222448 561772 222476
rect 408000 222436 408006 222448
rect 561766 222436 561772 222448
rect 561824 222436 561830 222488
rect 563698 222436 563704 222488
rect 563756 222476 563762 222488
rect 620094 222476 620100 222488
rect 563756 222448 620100 222476
rect 563756 222436 563762 222448
rect 620094 222436 620100 222448
rect 620152 222436 620158 222488
rect 272300 222380 281488 222408
rect 272300 222368 272306 222380
rect 328086 222368 328092 222420
rect 328144 222408 328150 222420
rect 338022 222408 338028 222420
rect 328144 222380 338028 222408
rect 328144 222368 328150 222380
rect 338022 222368 338028 222380
rect 338080 222368 338086 222420
rect 338206 222368 338212 222420
rect 338264 222408 338270 222420
rect 374178 222408 374184 222420
rect 338264 222380 374184 222408
rect 338264 222368 338270 222380
rect 374178 222368 374184 222380
rect 374236 222368 374242 222420
rect 375282 222368 375288 222420
rect 375340 222408 375346 222420
rect 394694 222408 394700 222420
rect 375340 222380 394700 222408
rect 375340 222368 375346 222380
rect 394694 222368 394700 222380
rect 394752 222368 394758 222420
rect 407574 222368 407580 222420
rect 407632 222408 407638 222420
rect 561582 222408 561588 222420
rect 407632 222380 561588 222408
rect 407632 222368 407638 222380
rect 561582 222368 561588 222380
rect 561640 222408 561646 222420
rect 619634 222408 619640 222420
rect 561640 222380 619640 222408
rect 561640 222368 561646 222380
rect 619634 222368 619640 222380
rect 619692 222368 619698 222420
rect 68646 222300 68652 222352
rect 68704 222340 68710 222352
rect 198274 222340 198280 222352
rect 68704 222312 198280 222340
rect 68704 222300 68710 222312
rect 198274 222300 198280 222312
rect 198332 222300 198338 222352
rect 202414 222300 202420 222352
rect 202472 222340 202478 222352
rect 256050 222340 256056 222352
rect 202472 222312 256056 222340
rect 202472 222300 202478 222312
rect 256050 222300 256056 222312
rect 256108 222300 256114 222352
rect 269666 222300 269672 222352
rect 269724 222340 269730 222352
rect 284570 222340 284576 222352
rect 269724 222312 284576 222340
rect 269724 222300 269730 222312
rect 284570 222300 284576 222312
rect 284628 222300 284634 222352
rect 332686 222300 332692 222352
rect 332744 222340 332750 222352
rect 381814 222340 381820 222352
rect 332744 222312 381820 222340
rect 332744 222300 332750 222312
rect 381814 222300 381820 222312
rect 381872 222300 381878 222352
rect 390830 222300 390836 222352
rect 390888 222340 390894 222352
rect 390888 222312 401548 222340
rect 390888 222300 390894 222312
rect 53558 222232 53564 222284
rect 53616 222272 53622 222284
rect 183002 222272 183008 222284
rect 53616 222244 183008 222272
rect 53616 222232 53622 222244
rect 183002 222232 183008 222244
rect 183060 222232 183066 222284
rect 187234 222232 187240 222284
rect 187292 222272 187298 222284
rect 235902 222272 235908 222284
rect 187292 222244 235908 222272
rect 187292 222232 187298 222244
rect 235902 222232 235908 222244
rect 235960 222232 235966 222284
rect 254578 222232 254584 222284
rect 254636 222272 254642 222284
rect 278498 222272 278504 222284
rect 254636 222244 278504 222272
rect 254636 222232 254642 222244
rect 278498 222232 278504 222244
rect 278556 222232 278562 222284
rect 310974 222232 310980 222284
rect 311032 222272 311038 222284
rect 333974 222272 333980 222284
rect 311032 222244 333980 222272
rect 311032 222232 311038 222244
rect 333974 222232 333980 222244
rect 334032 222232 334038 222284
rect 337654 222232 337660 222284
rect 337712 222272 337718 222284
rect 346486 222272 346492 222284
rect 337712 222244 346492 222272
rect 337712 222232 337718 222244
rect 346486 222232 346492 222244
rect 346544 222232 346550 222284
rect 346578 222232 346584 222284
rect 346636 222272 346642 222284
rect 385126 222272 385132 222284
rect 346636 222244 385132 222272
rect 346636 222232 346642 222244
rect 385126 222232 385132 222244
rect 385184 222232 385190 222284
rect 391842 222232 391848 222284
rect 391900 222272 391906 222284
rect 401134 222272 401140 222284
rect 391900 222244 401140 222272
rect 391900 222232 391906 222244
rect 401134 222232 401140 222244
rect 401192 222232 401198 222284
rect 41690 222164 41696 222216
rect 41748 222204 41754 222216
rect 59538 222204 59544 222216
rect 41748 222176 59544 222204
rect 41748 222164 41754 222176
rect 59538 222164 59544 222176
rect 59596 222164 59602 222216
rect 61930 222164 61936 222216
rect 61988 222204 61994 222216
rect 195422 222204 195428 222216
rect 61988 222176 195428 222204
rect 61988 222164 61994 222176
rect 195422 222164 195428 222176
rect 195480 222164 195486 222216
rect 200758 222164 200764 222216
rect 200816 222204 200822 222216
rect 255682 222204 255688 222216
rect 200816 222176 255688 222204
rect 200816 222164 200822 222176
rect 255682 222164 255688 222176
rect 255740 222164 255746 222216
rect 258810 222164 258816 222216
rect 258868 222204 258874 222216
rect 279234 222204 279240 222216
rect 258868 222176 279240 222204
rect 258868 222164 258874 222176
rect 279234 222164 279240 222176
rect 279292 222164 279298 222216
rect 312354 222164 312360 222216
rect 312412 222204 312418 222216
rect 337194 222204 337200 222216
rect 312412 222176 337200 222204
rect 312412 222164 312418 222176
rect 337194 222164 337200 222176
rect 337252 222164 337258 222216
rect 340966 222164 340972 222216
rect 341024 222204 341030 222216
rect 349798 222204 349804 222216
rect 341024 222176 349804 222204
rect 341024 222164 341030 222176
rect 349798 222164 349804 222176
rect 349856 222164 349862 222216
rect 349890 222164 349896 222216
rect 349948 222204 349954 222216
rect 393590 222204 393596 222216
rect 349948 222176 393596 222204
rect 349948 222164 349954 222176
rect 393590 222164 393596 222176
rect 393648 222164 393654 222216
rect 162026 222096 162032 222148
rect 162084 222136 162090 222148
rect 238938 222136 238944 222148
rect 162084 222108 238944 222136
rect 162084 222096 162090 222108
rect 238938 222096 238944 222108
rect 238996 222096 239002 222148
rect 244458 222096 244464 222148
rect 244516 222136 244522 222148
rect 256602 222136 256608 222148
rect 244516 222108 256608 222136
rect 244516 222096 244522 222108
rect 256602 222096 256608 222108
rect 256660 222096 256666 222148
rect 273070 222096 273076 222148
rect 273128 222136 273134 222148
rect 286042 222136 286048 222148
rect 273128 222108 286048 222136
rect 273128 222096 273134 222108
rect 286042 222096 286048 222108
rect 286100 222096 286106 222148
rect 322750 222096 322756 222148
rect 322808 222136 322814 222148
rect 358262 222136 358268 222148
rect 322808 222108 358268 222136
rect 322808 222096 322814 222108
rect 358262 222096 358268 222108
rect 358320 222096 358326 222148
rect 381906 222096 381912 222148
rect 381964 222136 381970 222148
rect 401410 222136 401416 222148
rect 381964 222108 401416 222136
rect 381964 222096 381970 222108
rect 401410 222096 401416 222108
rect 401468 222096 401474 222148
rect 401520 222136 401548 222312
rect 408310 222300 408316 222352
rect 408368 222340 408374 222352
rect 562962 222340 562968 222352
rect 408368 222312 562968 222340
rect 408368 222300 408374 222312
rect 562962 222300 562968 222312
rect 563020 222340 563026 222352
rect 634538 222340 634544 222352
rect 563020 222312 634544 222340
rect 563020 222300 563026 222312
rect 634538 222300 634544 222312
rect 634596 222300 634602 222352
rect 410058 222232 410064 222284
rect 410116 222272 410122 222284
rect 566826 222272 566832 222284
rect 410116 222244 566832 222272
rect 410116 222232 410122 222244
rect 566826 222232 566832 222244
rect 566884 222232 566890 222284
rect 570230 222232 570236 222284
rect 570288 222272 570294 222284
rect 570874 222272 570880 222284
rect 570288 222244 570880 222272
rect 570288 222232 570294 222244
rect 570874 222232 570880 222244
rect 570932 222272 570938 222284
rect 635918 222272 635924 222284
rect 570932 222244 635924 222272
rect 570932 222232 570938 222244
rect 635918 222232 635924 222244
rect 635976 222232 635982 222284
rect 410426 222164 410432 222216
rect 410484 222204 410490 222216
rect 567654 222204 567660 222216
rect 410484 222176 567660 222204
rect 410484 222164 410490 222176
rect 567654 222164 567660 222176
rect 567712 222164 567718 222216
rect 521654 222136 521660 222148
rect 401520 222108 521660 222136
rect 521654 222096 521660 222108
rect 521712 222096 521718 222148
rect 536282 222096 536288 222148
rect 536340 222136 536346 222148
rect 541434 222136 541440 222148
rect 536340 222108 541440 222136
rect 536340 222096 536346 222108
rect 541434 222096 541440 222108
rect 541492 222096 541498 222148
rect 615494 222136 615500 222148
rect 542556 222108 615500 222136
rect 160370 222028 160376 222080
rect 160428 222068 160434 222080
rect 238294 222068 238300 222080
rect 160428 222040 238300 222068
rect 160428 222028 160434 222040
rect 238294 222028 238300 222040
rect 238352 222028 238358 222080
rect 274726 222028 274732 222080
rect 274784 222068 274790 222080
rect 287054 222068 287060 222080
rect 274784 222040 287060 222068
rect 274784 222028 274790 222040
rect 287054 222028 287060 222040
rect 287112 222028 287118 222080
rect 320910 222028 320916 222080
rect 320968 222068 320974 222080
rect 357342 222068 357348 222080
rect 320968 222040 357348 222068
rect 320968 222028 320974 222040
rect 357342 222028 357348 222040
rect 357400 222028 357406 222080
rect 393222 222028 393228 222080
rect 393280 222068 393286 222080
rect 526438 222068 526444 222080
rect 393280 222040 526444 222068
rect 393280 222028 393286 222040
rect 526438 222028 526444 222040
rect 526496 222028 526502 222080
rect 538858 222028 538864 222080
rect 538916 222068 538922 222080
rect 542556 222068 542584 222108
rect 615494 222096 615500 222108
rect 615552 222096 615558 222148
rect 538916 222040 542584 222068
rect 538916 222028 538922 222040
rect 552566 222028 552572 222080
rect 552624 222068 552630 222080
rect 553210 222068 553216 222080
rect 552624 222040 553216 222068
rect 552624 222028 552630 222040
rect 553210 222028 553216 222040
rect 553268 222068 553274 222080
rect 632698 222068 632704 222080
rect 553268 222040 632704 222068
rect 553268 222028 553274 222040
rect 632698 222028 632704 222040
rect 632756 222028 632762 222080
rect 90542 221960 90548 222012
rect 90600 222000 90606 222012
rect 160094 222000 160100 222012
rect 90600 221972 160100 222000
rect 90600 221960 90606 221972
rect 160094 221960 160100 221972
rect 160152 221960 160158 222012
rect 170490 221960 170496 222012
rect 170548 222000 170554 222012
rect 232590 222000 232596 222012
rect 170548 221972 232596 222000
rect 170548 221960 170554 221972
rect 232590 221960 232596 221972
rect 232648 221960 232654 222012
rect 241790 222000 241796 222012
rect 232792 221972 241796 222000
rect 168742 221892 168748 221944
rect 168800 221932 168806 221944
rect 232792 221932 232820 221972
rect 241790 221960 241796 221972
rect 241848 221960 241854 222012
rect 319806 221960 319812 222012
rect 319864 222000 319870 222012
rect 354030 222000 354036 222012
rect 319864 221972 354036 222000
rect 319864 221960 319870 221972
rect 354030 221960 354036 221972
rect 354088 221960 354094 222012
rect 388714 221960 388720 222012
rect 388772 222000 388778 222012
rect 516410 222000 516416 222012
rect 388772 221972 516416 222000
rect 388772 221960 388778 221972
rect 516410 221960 516416 221972
rect 516468 221960 516474 222012
rect 532694 221960 532700 222012
rect 532752 222000 532758 222012
rect 533430 222000 533436 222012
rect 532752 221972 533436 222000
rect 532752 221960 532758 221972
rect 533430 221960 533436 221972
rect 533488 222000 533494 222012
rect 614574 222000 614580 222012
rect 533488 221972 614580 222000
rect 533488 221960 533494 221972
rect 614574 221960 614580 221972
rect 614632 221960 614638 222012
rect 168800 221904 232820 221932
rect 168800 221892 168806 221904
rect 234338 221892 234344 221944
rect 234396 221932 234402 221944
rect 248598 221932 248604 221944
rect 234396 221904 248604 221932
rect 234396 221892 234402 221904
rect 248598 221892 248604 221904
rect 248656 221892 248662 221944
rect 273898 221892 273904 221944
rect 273956 221932 273962 221944
rect 285306 221932 285312 221944
rect 273956 221904 285312 221932
rect 273956 221892 273962 221904
rect 285306 221892 285312 221904
rect 285364 221892 285370 221944
rect 287054 221892 287060 221944
rect 287112 221932 287118 221944
rect 289262 221932 289268 221944
rect 287112 221904 289268 221932
rect 287112 221892 287118 221904
rect 289262 221892 289268 221904
rect 289320 221892 289326 221944
rect 318058 221892 318064 221944
rect 318116 221932 318122 221944
rect 350626 221932 350632 221944
rect 318116 221904 350632 221932
rect 318116 221892 318122 221904
rect 350626 221892 350632 221904
rect 350684 221892 350690 221944
rect 387610 221892 387616 221944
rect 387668 221932 387674 221944
rect 513834 221932 513840 221944
rect 387668 221904 513840 221932
rect 387668 221892 387674 221904
rect 513834 221892 513840 221904
rect 513892 221892 513898 221944
rect 530670 221892 530676 221944
rect 530728 221932 530734 221944
rect 614022 221932 614028 221944
rect 530728 221904 614028 221932
rect 530728 221892 530734 221904
rect 614022 221892 614028 221904
rect 614080 221892 614086 221944
rect 177206 221824 177212 221876
rect 177264 221864 177270 221876
rect 177264 221836 236040 221864
rect 177264 221824 177270 221836
rect 183922 221756 183928 221808
rect 183980 221796 183986 221808
rect 236012 221796 236040 221836
rect 281442 221824 281448 221876
rect 281500 221864 281506 221876
rect 289906 221864 289912 221876
rect 281500 221836 289912 221864
rect 281500 221824 281506 221836
rect 289906 221824 289912 221836
rect 289964 221824 289970 221876
rect 319898 221824 319904 221876
rect 319956 221864 319962 221876
rect 351454 221864 351460 221876
rect 319956 221836 351460 221864
rect 319956 221824 319962 221836
rect 351454 221824 351460 221836
rect 351512 221824 351518 221876
rect 386230 221824 386236 221876
rect 386288 221864 386294 221876
rect 510614 221864 510620 221876
rect 386288 221836 510620 221864
rect 386288 221824 386294 221836
rect 510614 221824 510620 221836
rect 510672 221824 510678 221876
rect 547506 221824 547512 221876
rect 547564 221864 547570 221876
rect 631778 221864 631784 221876
rect 547564 221836 631784 221864
rect 547564 221824 547570 221836
rect 631778 221824 631784 221836
rect 631836 221824 631842 221876
rect 245746 221796 245752 221808
rect 183980 221768 235948 221796
rect 236012 221768 245752 221796
rect 183980 221756 183986 221768
rect 182082 221688 182088 221740
rect 182140 221728 182146 221740
rect 233510 221728 233516 221740
rect 182140 221700 233516 221728
rect 182140 221688 182146 221700
rect 233510 221688 233516 221700
rect 233568 221688 233574 221740
rect 179690 221620 179696 221672
rect 179748 221660 179754 221672
rect 235626 221660 235632 221672
rect 179748 221632 235632 221660
rect 179748 221620 179754 221632
rect 235626 221620 235632 221632
rect 235684 221620 235690 221672
rect 235920 221660 235948 221768
rect 245746 221756 245752 221768
rect 245804 221756 245810 221808
rect 268010 221756 268016 221808
rect 268068 221796 268074 221808
rect 284202 221796 284208 221808
rect 268068 221768 284208 221796
rect 268068 221756 268074 221768
rect 284202 221756 284208 221768
rect 284260 221756 284266 221808
rect 321278 221756 321284 221808
rect 321336 221796 321342 221808
rect 354858 221796 354864 221808
rect 321336 221768 354864 221796
rect 321336 221756 321342 221768
rect 354858 221756 354864 221768
rect 354916 221756 354922 221808
rect 385494 221756 385500 221808
rect 385552 221796 385558 221808
rect 508774 221796 508780 221808
rect 385552 221768 508780 221796
rect 385552 221756 385558 221768
rect 508774 221756 508780 221768
rect 508832 221756 508838 221808
rect 528370 221756 528376 221808
rect 528428 221796 528434 221808
rect 613562 221796 613568 221808
rect 528428 221768 613568 221796
rect 528428 221756 528434 221768
rect 613562 221756 613568 221768
rect 613620 221756 613626 221808
rect 257890 221688 257896 221740
rect 257948 221728 257954 221740
rect 279970 221728 279976 221740
rect 257948 221700 279976 221728
rect 257948 221688 257954 221700
rect 279970 221688 279976 221700
rect 280028 221688 280034 221740
rect 284846 221688 284852 221740
rect 284904 221728 284910 221740
rect 291378 221728 291384 221740
rect 284904 221700 291384 221728
rect 284904 221688 284910 221700
rect 291378 221688 291384 221700
rect 291436 221688 291442 221740
rect 316678 221688 316684 221740
rect 316736 221728 316742 221740
rect 347314 221728 347320 221740
rect 316736 221700 347320 221728
rect 316736 221688 316742 221700
rect 347314 221688 347320 221700
rect 347372 221688 347378 221740
rect 347774 221688 347780 221740
rect 347832 221728 347838 221740
rect 380066 221728 380072 221740
rect 347832 221700 380072 221728
rect 347832 221688 347838 221700
rect 380066 221688 380072 221700
rect 380124 221688 380130 221740
rect 383378 221688 383384 221740
rect 383436 221728 383442 221740
rect 503714 221728 503720 221740
rect 383436 221700 503720 221728
rect 383436 221688 383442 221700
rect 503714 221688 503720 221700
rect 503772 221688 503778 221740
rect 542722 221688 542728 221740
rect 542780 221728 542786 221740
rect 630858 221728 630864 221740
rect 542780 221700 630864 221728
rect 542780 221688 542786 221700
rect 630858 221688 630864 221700
rect 630916 221688 630922 221740
rect 248322 221660 248328 221672
rect 235920 221632 248328 221660
rect 248322 221620 248328 221632
rect 248380 221620 248386 221672
rect 255406 221620 255412 221672
rect 255464 221660 255470 221672
rect 277854 221660 277860 221672
rect 255464 221632 277860 221660
rect 255464 221620 255470 221632
rect 277854 221620 277860 221632
rect 277912 221620 277918 221672
rect 286410 221660 286416 221672
rect 277964 221632 286416 221660
rect 194042 221552 194048 221604
rect 194100 221592 194106 221604
rect 196066 221592 196072 221604
rect 194100 221564 196072 221592
rect 194100 221552 194106 221564
rect 196066 221552 196072 221564
rect 196124 221552 196130 221604
rect 196158 221552 196164 221604
rect 196216 221592 196222 221604
rect 196216 221564 235948 221592
rect 196216 221552 196222 221564
rect 159542 221484 159548 221536
rect 159600 221524 159606 221536
rect 209682 221524 209688 221536
rect 159600 221496 209688 221524
rect 159600 221484 159606 221496
rect 209682 221484 209688 221496
rect 209740 221484 209746 221536
rect 213362 221484 213368 221536
rect 213420 221524 213426 221536
rect 235920 221524 235948 221564
rect 235994 221552 236000 221604
rect 236052 221592 236058 221604
rect 245378 221592 245384 221604
rect 236052 221564 245384 221592
rect 236052 221552 236058 221564
rect 245378 221552 245384 221564
rect 245436 221552 245442 221604
rect 275554 221552 275560 221604
rect 275612 221592 275618 221604
rect 277964 221592 277992 221632
rect 286410 221620 286416 221632
rect 286468 221620 286474 221672
rect 317046 221620 317052 221672
rect 317104 221660 317110 221672
rect 345014 221660 345020 221672
rect 317104 221632 345020 221660
rect 317104 221620 317110 221632
rect 345014 221620 345020 221632
rect 345072 221620 345078 221672
rect 345106 221620 345112 221672
rect 345164 221660 345170 221672
rect 373350 221660 373356 221672
rect 345164 221632 373356 221660
rect 345164 221620 345170 221632
rect 373350 221620 373356 221632
rect 373408 221620 373414 221672
rect 384022 221620 384028 221672
rect 384080 221660 384086 221672
rect 505738 221660 505744 221672
rect 384080 221632 505744 221660
rect 384080 221620 384086 221632
rect 505738 221620 505744 221632
rect 505796 221620 505802 221672
rect 538306 221620 538312 221672
rect 538364 221660 538370 221672
rect 540146 221660 540152 221672
rect 538364 221632 540152 221660
rect 538364 221620 538370 221632
rect 540146 221620 540152 221632
rect 540204 221660 540210 221672
rect 630398 221660 630404 221672
rect 540204 221632 630404 221660
rect 540204 221620 540210 221632
rect 630398 221620 630404 221632
rect 630456 221620 630462 221672
rect 275612 221564 277992 221592
rect 275612 221552 275618 221564
rect 278130 221552 278136 221604
rect 278188 221592 278194 221604
rect 288526 221592 288532 221604
rect 278188 221564 288532 221592
rect 278188 221552 278194 221564
rect 288526 221552 288532 221564
rect 288584 221552 288590 221604
rect 318426 221552 318432 221604
rect 318484 221592 318490 221604
rect 348142 221592 348148 221604
rect 318484 221564 348148 221592
rect 318484 221552 318490 221564
rect 348142 221552 348148 221564
rect 348200 221552 348206 221604
rect 381998 221552 382004 221604
rect 382056 221592 382062 221604
rect 389358 221592 389364 221604
rect 382056 221564 389364 221592
rect 382056 221552 382062 221564
rect 389358 221552 389364 221564
rect 389416 221552 389422 221604
rect 401410 221552 401416 221604
rect 401468 221592 401474 221604
rect 500402 221592 500408 221604
rect 401468 221564 500408 221592
rect 401468 221552 401474 221564
rect 500402 221552 500408 221564
rect 500460 221552 500466 221604
rect 502702 221552 502708 221604
rect 502760 221592 502766 221604
rect 503806 221592 503812 221604
rect 502760 221564 503812 221592
rect 502760 221552 502766 221564
rect 503806 221552 503812 221564
rect 503864 221552 503870 221604
rect 513374 221552 513380 221604
rect 513432 221592 513438 221604
rect 610802 221592 610808 221604
rect 513432 221564 610808 221592
rect 513432 221552 513438 221564
rect 610802 221552 610808 221564
rect 610860 221552 610866 221604
rect 250070 221524 250076 221536
rect 213420 221496 231716 221524
rect 235920 221496 250076 221524
rect 213420 221484 213426 221496
rect 149422 221416 149428 221468
rect 149480 221456 149486 221468
rect 188430 221456 188436 221468
rect 149480 221428 188436 221456
rect 149480 221416 149486 221428
rect 188430 221416 188436 221428
rect 188488 221416 188494 221468
rect 195698 221416 195704 221468
rect 195756 221456 195762 221468
rect 195756 221428 196020 221456
rect 195756 221416 195762 221428
rect 192294 221348 192300 221400
rect 192352 221388 192358 221400
rect 193030 221388 193036 221400
rect 192352 221360 193036 221388
rect 192352 221348 192358 221360
rect 193030 221348 193036 221360
rect 193088 221348 193094 221400
rect 193122 221348 193128 221400
rect 193180 221388 193186 221400
rect 195882 221388 195888 221400
rect 193180 221360 195888 221388
rect 193180 221348 193186 221360
rect 195882 221348 195888 221360
rect 195940 221348 195946 221400
rect 195992 221388 196020 221428
rect 196066 221416 196072 221468
rect 196124 221456 196130 221468
rect 231688 221456 231716 221496
rect 250070 221484 250076 221496
rect 250128 221484 250134 221536
rect 266354 221484 266360 221536
rect 266412 221524 266418 221536
rect 283190 221524 283196 221536
rect 266412 221496 283196 221524
rect 266412 221484 266418 221496
rect 283190 221484 283196 221496
rect 283248 221484 283254 221536
rect 286502 221484 286508 221536
rect 286560 221524 286566 221536
rect 291746 221524 291752 221536
rect 286560 221496 291752 221524
rect 286560 221484 286566 221496
rect 291746 221484 291752 221496
rect 291804 221484 291810 221536
rect 315206 221484 315212 221536
rect 315264 221524 315270 221536
rect 343910 221524 343916 221536
rect 315264 221496 343916 221524
rect 315264 221484 315270 221496
rect 343910 221484 343916 221496
rect 343968 221484 343974 221536
rect 345290 221484 345296 221536
rect 345348 221524 345354 221536
rect 366634 221524 366640 221536
rect 345348 221496 366640 221524
rect 345348 221484 345354 221496
rect 366634 221484 366640 221496
rect 366692 221484 366698 221536
rect 380526 221484 380532 221536
rect 380584 221524 380590 221536
rect 497366 221524 497372 221536
rect 380584 221496 497372 221524
rect 380584 221484 380590 221496
rect 497366 221484 497372 221496
rect 497424 221524 497430 221536
rect 499482 221524 499488 221536
rect 497424 221496 499488 221524
rect 497424 221484 497430 221496
rect 499482 221484 499488 221496
rect 499540 221484 499546 221536
rect 534902 221484 534908 221536
rect 534960 221524 534966 221536
rect 629478 221524 629484 221536
rect 534960 221496 629484 221524
rect 534960 221484 534966 221496
rect 629478 221484 629484 221496
rect 629536 221484 629542 221536
rect 237006 221456 237012 221468
rect 196124 221428 231624 221456
rect 231688 221428 237012 221456
rect 196124 221416 196130 221428
rect 195992 221360 231440 221388
rect 166258 221280 166264 221332
rect 166316 221320 166322 221332
rect 208946 221320 208952 221332
rect 166316 221292 208952 221320
rect 166316 221280 166322 221292
rect 208946 221280 208952 221292
rect 209004 221280 209010 221332
rect 220078 221280 220084 221332
rect 220136 221320 220142 221332
rect 231210 221320 231216 221332
rect 220136 221292 231216 221320
rect 220136 221280 220142 221292
rect 231210 221280 231216 221292
rect 231268 221280 231274 221332
rect 172974 221212 172980 221264
rect 173032 221252 173038 221264
rect 214926 221252 214932 221264
rect 173032 221224 214932 221252
rect 173032 221212 173038 221224
rect 214926 221212 214932 221224
rect 214984 221212 214990 221264
rect 178862 221144 178868 221196
rect 178920 221184 178926 221196
rect 181898 221184 181904 221196
rect 178920 221156 181904 221184
rect 178920 221144 178926 221156
rect 181898 221144 181904 221156
rect 181956 221144 181962 221196
rect 189810 221144 189816 221196
rect 189868 221184 189874 221196
rect 231302 221184 231308 221196
rect 189868 221156 231308 221184
rect 189868 221144 189874 221156
rect 231302 221144 231308 221156
rect 231360 221144 231366 221196
rect 231412 221184 231440 221360
rect 231596 221252 231624 221428
rect 237006 221416 237012 221428
rect 237064 221416 237070 221468
rect 249518 221416 249524 221468
rect 249576 221456 249582 221468
rect 258902 221456 258908 221468
rect 249576 221428 258908 221456
rect 249576 221416 249582 221428
rect 258902 221416 258908 221428
rect 258960 221416 258966 221468
rect 265526 221416 265532 221468
rect 265584 221456 265590 221468
rect 282086 221456 282092 221468
rect 265584 221428 282092 221456
rect 265584 221416 265590 221428
rect 282086 221416 282092 221428
rect 282144 221416 282150 221468
rect 283926 221416 283932 221468
rect 283984 221456 283990 221468
rect 283984 221428 284294 221456
rect 283984 221416 283990 221428
rect 236914 221348 236920 221400
rect 236972 221388 236978 221400
rect 241238 221388 241244 221400
rect 236972 221360 241244 221388
rect 236972 221348 236978 221360
rect 241238 221348 241244 221360
rect 241296 221348 241302 221400
rect 247862 221348 247868 221400
rect 247920 221388 247926 221400
rect 255958 221388 255964 221400
rect 247920 221360 255964 221388
rect 247920 221348 247926 221360
rect 255958 221348 255964 221360
rect 256016 221348 256022 221400
rect 256234 221348 256240 221400
rect 256292 221388 256298 221400
rect 259546 221388 259552 221400
rect 256292 221360 259552 221388
rect 256292 221348 256298 221360
rect 259546 221348 259552 221360
rect 259604 221348 259610 221400
rect 267182 221348 267188 221400
rect 267240 221388 267246 221400
rect 282454 221388 282460 221400
rect 267240 221360 282460 221388
rect 267240 221348 267246 221360
rect 282454 221348 282460 221360
rect 282512 221348 282518 221400
rect 233510 221280 233516 221332
rect 233568 221320 233574 221332
rect 239858 221320 239864 221332
rect 233568 221292 239864 221320
rect 233568 221280 233574 221292
rect 239858 221280 239864 221292
rect 239916 221280 239922 221332
rect 251082 221280 251088 221332
rect 251140 221320 251146 221332
rect 256510 221320 256516 221332
rect 251140 221292 256516 221320
rect 251140 221280 251146 221292
rect 256510 221280 256516 221292
rect 256568 221280 256574 221332
rect 270402 221280 270408 221332
rect 270460 221320 270466 221332
rect 283834 221320 283840 221332
rect 270460 221292 283840 221320
rect 270460 221280 270466 221292
rect 283834 221280 283840 221292
rect 283892 221280 283898 221332
rect 284266 221320 284294 221428
rect 288250 221416 288256 221468
rect 288308 221456 288314 221468
rect 292758 221456 292764 221468
rect 288308 221428 292764 221456
rect 288308 221416 288314 221428
rect 292758 221416 292764 221428
rect 292816 221416 292822 221468
rect 314562 221416 314568 221468
rect 314620 221456 314626 221468
rect 339678 221456 339684 221468
rect 314620 221428 339684 221456
rect 314620 221416 314626 221428
rect 339678 221416 339684 221428
rect 339736 221416 339742 221468
rect 380802 221416 380808 221468
rect 380860 221456 380866 221468
rect 497826 221456 497832 221468
rect 380860 221428 497832 221456
rect 380860 221416 380866 221428
rect 497826 221416 497832 221428
rect 497884 221416 497890 221468
rect 530118 221416 530124 221468
rect 530176 221456 530182 221468
rect 628466 221456 628472 221468
rect 530176 221428 628472 221456
rect 530176 221416 530182 221428
rect 628466 221416 628472 221428
rect 628524 221416 628530 221468
rect 289078 221348 289084 221400
rect 289136 221388 289142 221400
rect 292114 221388 292120 221400
rect 289136 221360 292120 221388
rect 289136 221348 289142 221360
rect 292114 221348 292120 221360
rect 292172 221348 292178 221400
rect 292390 221348 292396 221400
rect 292448 221388 292454 221400
rect 293494 221388 293500 221400
rect 292448 221360 293500 221388
rect 292448 221348 292454 221360
rect 293494 221348 293500 221360
rect 293552 221348 293558 221400
rect 314194 221348 314200 221400
rect 314252 221388 314258 221400
rect 338022 221388 338028 221400
rect 314252 221360 338028 221388
rect 314252 221348 314258 221360
rect 338022 221348 338028 221360
rect 338080 221348 338086 221400
rect 342898 221348 342904 221400
rect 342956 221388 342962 221400
rect 356514 221388 356520 221400
rect 342956 221360 356520 221388
rect 342956 221348 342962 221360
rect 356514 221348 356520 221360
rect 356572 221348 356578 221400
rect 379054 221348 379060 221400
rect 379112 221388 379118 221400
rect 494054 221388 494060 221400
rect 379112 221360 494060 221388
rect 379112 221348 379118 221360
rect 494054 221348 494060 221360
rect 494112 221348 494118 221400
rect 507946 221348 507952 221400
rect 508004 221388 508010 221400
rect 609882 221388 609888 221400
rect 508004 221360 609888 221388
rect 508004 221348 508010 221360
rect 609882 221348 609888 221360
rect 609940 221348 609946 221400
rect 289538 221320 289544 221332
rect 284266 221292 289544 221320
rect 289538 221280 289544 221292
rect 289596 221280 289602 221332
rect 291562 221280 291568 221332
rect 291620 221320 291626 221332
rect 294230 221320 294236 221332
rect 291620 221292 294236 221320
rect 291620 221280 291626 221292
rect 294230 221280 294236 221292
rect 294288 221280 294294 221332
rect 294966 221280 294972 221332
rect 295024 221320 295030 221332
rect 295610 221320 295616 221332
rect 295024 221292 295616 221320
rect 295024 221280 295030 221292
rect 295610 221280 295616 221292
rect 295668 221280 295674 221332
rect 313826 221280 313832 221332
rect 313884 221320 313890 221332
rect 340598 221320 340604 221332
rect 313884 221292 340604 221320
rect 313884 221280 313890 221292
rect 340598 221280 340604 221292
rect 340656 221280 340662 221332
rect 342070 221280 342076 221332
rect 342128 221320 342134 221332
rect 353294 221320 353300 221332
rect 342128 221292 353300 221320
rect 342128 221280 342134 221292
rect 353294 221280 353300 221292
rect 353352 221280 353358 221332
rect 377674 221280 377680 221332
rect 377732 221320 377738 221332
rect 490282 221320 490288 221332
rect 377732 221292 490288 221320
rect 377732 221280 377738 221292
rect 490282 221280 490288 221292
rect 490340 221280 490346 221332
rect 518986 221280 518992 221332
rect 519044 221320 519050 221332
rect 519998 221320 520004 221332
rect 519044 221292 520004 221320
rect 519044 221280 519050 221292
rect 519998 221280 520004 221292
rect 520056 221280 520062 221332
rect 525058 221280 525064 221332
rect 525116 221320 525122 221332
rect 627546 221320 627552 221332
rect 525116 221292 627552 221320
rect 525116 221280 525122 221292
rect 627546 221280 627552 221292
rect 627604 221280 627610 221332
rect 242986 221252 242992 221264
rect 231596 221224 242992 221252
rect 242986 221212 242992 221224
rect 243044 221212 243050 221264
rect 252922 221212 252928 221264
rect 252980 221252 252986 221264
rect 258350 221252 258356 221264
rect 252980 221224 258356 221252
rect 252980 221212 252986 221224
rect 258350 221212 258356 221224
rect 258408 221212 258414 221264
rect 268838 221212 268844 221264
rect 268896 221252 268902 221264
rect 283558 221252 283564 221264
rect 268896 221224 283564 221252
rect 268896 221212 268902 221224
rect 283558 221212 283564 221224
rect 283616 221212 283622 221264
rect 286686 221252 286692 221264
rect 283668 221224 286692 221252
rect 243078 221184 243084 221196
rect 231412 221156 243084 221184
rect 243078 221144 243084 221156
rect 243136 221144 243142 221196
rect 277302 221144 277308 221196
rect 277360 221184 277366 221196
rect 283668 221184 283696 221224
rect 286686 221212 286692 221224
rect 286744 221212 286750 221264
rect 289722 221212 289728 221264
rect 289780 221252 289786 221264
rect 293126 221252 293132 221264
rect 289780 221224 293132 221252
rect 289780 221212 289786 221224
rect 293126 221212 293132 221224
rect 293184 221212 293190 221264
rect 315574 221212 315580 221264
rect 315632 221252 315638 221264
rect 341426 221252 341432 221264
rect 315632 221224 341432 221252
rect 315632 221212 315638 221224
rect 341426 221212 341432 221224
rect 341484 221212 341490 221264
rect 371970 221212 371976 221264
rect 372028 221252 372034 221264
rect 476850 221252 476856 221264
rect 372028 221224 476856 221252
rect 372028 221212 372034 221224
rect 476850 221212 476856 221224
rect 476908 221212 476914 221264
rect 503162 221212 503168 221264
rect 503220 221252 503226 221264
rect 608962 221252 608968 221264
rect 503220 221224 608968 221252
rect 503220 221212 503226 221224
rect 608962 221212 608968 221224
rect 609020 221212 609026 221264
rect 277360 221156 283696 221184
rect 277360 221144 277366 221156
rect 283742 221144 283748 221196
rect 283800 221184 283806 221196
rect 287422 221184 287428 221196
rect 283800 221156 287428 221184
rect 283800 221144 283806 221156
rect 287422 221144 287428 221156
rect 287480 221144 287486 221196
rect 313090 221144 313096 221196
rect 313148 221184 313154 221196
rect 336734 221184 336740 221196
rect 313148 221156 336740 221184
rect 313148 221144 313154 221156
rect 336734 221144 336740 221156
rect 336792 221144 336798 221196
rect 337378 221144 337384 221196
rect 337436 221184 337442 221196
rect 349890 221184 349896 221196
rect 337436 221156 349896 221184
rect 337436 221144 337442 221156
rect 349890 221144 349896 221156
rect 349948 221144 349954 221196
rect 367278 221144 367284 221196
rect 367336 221184 367342 221196
rect 464246 221184 464252 221196
rect 367336 221156 464252 221184
rect 367336 221144 367342 221156
rect 464246 221144 464252 221156
rect 464304 221144 464310 221196
rect 519998 221144 520004 221196
rect 520056 221184 520062 221196
rect 626626 221184 626632 221196
rect 520056 221156 626632 221184
rect 520056 221144 520062 221156
rect 626626 221144 626632 221156
rect 626684 221144 626690 221196
rect 655698 221144 655704 221196
rect 655756 221184 655762 221196
rect 676030 221184 676036 221196
rect 655756 221156 676036 221184
rect 655756 221144 655762 221156
rect 676030 221144 676036 221156
rect 676088 221144 676094 221196
rect 183094 221076 183100 221128
rect 183152 221116 183158 221128
rect 216122 221116 216128 221128
rect 183152 221088 216128 221116
rect 183152 221076 183158 221088
rect 216122 221076 216128 221088
rect 216180 221076 216186 221128
rect 230106 221116 230112 221128
rect 226306 221088 230112 221116
rect 188982 221008 188988 221060
rect 189040 221048 189046 221060
rect 196158 221048 196164 221060
rect 189040 221020 196164 221048
rect 189040 221008 189046 221020
rect 196158 221008 196164 221020
rect 196216 221008 196222 221060
rect 199930 221008 199936 221060
rect 199988 221048 199994 221060
rect 226306 221048 226334 221088
rect 230106 221076 230112 221088
rect 230164 221076 230170 221128
rect 230198 221076 230204 221128
rect 230256 221116 230262 221128
rect 239766 221116 239772 221128
rect 230256 221088 239772 221116
rect 230256 221076 230262 221088
rect 239766 221076 239772 221088
rect 239824 221076 239830 221128
rect 282362 221076 282368 221128
rect 282420 221116 282426 221128
rect 287054 221116 287060 221128
rect 282420 221088 287060 221116
rect 282420 221076 282426 221088
rect 287054 221076 287060 221088
rect 287112 221076 287118 221128
rect 287330 221076 287336 221128
rect 287388 221116 287394 221128
rect 291010 221116 291016 221128
rect 287388 221088 291016 221116
rect 287388 221076 287394 221088
rect 291010 221076 291016 221088
rect 291068 221076 291074 221128
rect 330202 221076 330208 221128
rect 330260 221116 330266 221128
rect 343542 221116 343548 221128
rect 330260 221088 343548 221116
rect 330260 221076 330266 221088
rect 343542 221076 343548 221088
rect 343600 221076 343606 221128
rect 365714 221076 365720 221128
rect 365772 221116 365778 221128
rect 407022 221116 407028 221128
rect 365772 221088 407028 221116
rect 365772 221076 365778 221088
rect 407022 221076 407028 221088
rect 407080 221076 407086 221128
rect 517054 221076 517060 221128
rect 517112 221116 517118 221128
rect 517606 221116 517612 221128
rect 517112 221088 517612 221116
rect 517112 221076 517118 221088
rect 517606 221076 517612 221088
rect 517664 221116 517670 221128
rect 626166 221116 626172 221128
rect 517664 221088 626172 221116
rect 517664 221076 517670 221088
rect 626166 221076 626172 221088
rect 626224 221076 626230 221128
rect 199988 221020 226334 221048
rect 199988 221008 199994 221020
rect 226794 221008 226800 221060
rect 226852 221048 226858 221060
rect 239950 221048 239956 221060
rect 226852 221020 239956 221048
rect 226852 221008 226858 221020
rect 239950 221008 239956 221020
rect 240008 221008 240014 221060
rect 279786 221008 279792 221060
rect 279844 221048 279850 221060
rect 288894 221048 288900 221060
rect 279844 221020 288900 221048
rect 279844 221008 279850 221020
rect 288894 221008 288900 221020
rect 288952 221008 288958 221060
rect 342990 221008 342996 221060
rect 343048 221048 343054 221060
rect 359918 221048 359924 221060
rect 343048 221020 359924 221048
rect 343048 221008 343054 221020
rect 359918 221008 359924 221020
rect 359976 221008 359982 221060
rect 376846 221008 376852 221060
rect 376904 221048 376910 221060
rect 382642 221048 382648 221060
rect 376904 221020 382648 221048
rect 376904 221008 376910 221020
rect 382642 221008 382648 221020
rect 382700 221008 382706 221060
rect 389082 221008 389088 221060
rect 389140 221048 389146 221060
rect 396074 221048 396080 221060
rect 389140 221020 396080 221048
rect 389140 221008 389146 221020
rect 396074 221008 396080 221020
rect 396132 221008 396138 221060
rect 397638 221008 397644 221060
rect 397696 221048 397702 221060
rect 537386 221048 537392 221060
rect 397696 221020 537392 221048
rect 397696 221008 397702 221020
rect 537386 221008 537392 221020
rect 537444 221008 537450 221060
rect 558178 221008 558184 221060
rect 558236 221048 558242 221060
rect 633618 221048 633624 221060
rect 558236 221020 633624 221048
rect 558236 221008 558242 221020
rect 633618 221008 633624 221020
rect 633676 221008 633682 221060
rect 655514 221008 655520 221060
rect 655572 221048 655578 221060
rect 675846 221048 675852 221060
rect 655572 221020 675852 221048
rect 655572 221008 655578 221020
rect 675846 221008 675852 221020
rect 675904 221008 675910 221060
rect 206646 220940 206652 220992
rect 206704 220980 206710 220992
rect 236270 220980 236276 220992
rect 206704 220952 226334 220980
rect 206704 220940 206710 220952
rect 196526 220872 196532 220924
rect 196584 220912 196590 220924
rect 216582 220912 216588 220924
rect 196584 220884 216588 220912
rect 196584 220872 196590 220884
rect 216582 220872 216588 220884
rect 216640 220872 216646 220924
rect 164602 220804 164608 220856
rect 164660 220844 164666 220856
rect 166350 220844 166356 220856
rect 164660 220816 166356 220844
rect 164660 220804 164666 220816
rect 166350 220804 166356 220816
rect 166408 220804 166414 220856
rect 167914 220804 167920 220856
rect 167972 220844 167978 220856
rect 169110 220844 169116 220856
rect 167972 220816 169116 220844
rect 167972 220804 167978 220816
rect 169110 220804 169116 220816
rect 169168 220804 169174 220856
rect 174630 220804 174636 220856
rect 174688 220844 174694 220856
rect 176654 220844 176660 220856
rect 174688 220816 176660 220844
rect 174688 220804 174694 220816
rect 176654 220804 176660 220816
rect 176712 220804 176718 220856
rect 204070 220804 204076 220856
rect 204128 220844 204134 220856
rect 209222 220844 209228 220856
rect 204128 220816 209228 220844
rect 204128 220804 204134 220816
rect 209222 220804 209228 220816
rect 209280 220804 209286 220856
rect 226306 220844 226334 220952
rect 226812 220952 236276 220980
rect 226812 220844 226840 220952
rect 236270 220940 236276 220952
rect 236328 220940 236334 220992
rect 276474 220940 276480 220992
rect 276532 220980 276538 220992
rect 283742 220980 283748 220992
rect 276532 220952 283748 220980
rect 276532 220940 276538 220952
rect 283742 220940 283748 220952
rect 283800 220940 283806 220992
rect 285674 220940 285680 220992
rect 285732 220980 285738 220992
rect 290642 220980 290648 220992
rect 285732 220952 290648 220980
rect 285732 220940 285738 220952
rect 290642 220940 290648 220952
rect 290700 220940 290706 220992
rect 334158 220940 334164 220992
rect 334216 220980 334222 220992
rect 346578 220980 346584 220992
rect 334216 220952 346584 220980
rect 334216 220940 334222 220952
rect 346578 220940 346584 220952
rect 346636 220940 346642 220992
rect 512178 220940 512184 220992
rect 512236 220980 512242 220992
rect 625246 220980 625252 220992
rect 512236 220952 625252 220980
rect 512236 220940 512242 220952
rect 625246 220940 625252 220952
rect 625304 220940 625310 220992
rect 230106 220872 230112 220924
rect 230164 220912 230170 220924
rect 232038 220912 232044 220924
rect 230164 220884 232044 220912
rect 230164 220872 230170 220884
rect 232038 220872 232044 220884
rect 232096 220872 232102 220924
rect 280614 220872 280620 220924
rect 280672 220912 280678 220924
rect 288158 220912 288164 220924
rect 280672 220884 288164 220912
rect 280672 220872 280678 220884
rect 288158 220872 288164 220884
rect 288216 220872 288222 220924
rect 395430 220872 395436 220924
rect 395488 220912 395494 220924
rect 532694 220912 532700 220924
rect 395488 220884 532700 220912
rect 395488 220872 395494 220884
rect 532694 220872 532700 220884
rect 532752 220872 532758 220924
rect 541434 220872 541440 220924
rect 541492 220912 541498 220924
rect 615954 220912 615960 220924
rect 541492 220884 615960 220912
rect 541492 220872 541498 220884
rect 615954 220872 615960 220884
rect 616012 220872 616018 220924
rect 226306 220816 226840 220844
rect 231210 220804 231216 220856
rect 231268 220844 231274 220856
rect 236730 220844 236736 220856
rect 231268 220816 236736 220844
rect 231268 220804 231274 220816
rect 236730 220804 236736 220816
rect 236788 220804 236794 220856
rect 395062 220804 395068 220856
rect 395120 220844 395126 220856
rect 531498 220844 531504 220856
rect 395120 220816 531504 220844
rect 395120 220804 395126 220816
rect 531498 220804 531504 220816
rect 531556 220804 531562 220856
rect 543550 220804 543556 220856
rect 543608 220844 543614 220856
rect 616414 220844 616420 220856
rect 543608 220816 616420 220844
rect 543608 220804 543614 220816
rect 616414 220804 616420 220816
rect 616472 220804 616478 220856
rect 655422 220804 655428 220856
rect 655480 220844 655486 220856
rect 675938 220844 675944 220856
rect 655480 220816 675944 220844
rect 655480 220804 655486 220816
rect 675938 220804 675944 220816
rect 675996 220804 676002 220856
rect 42150 220736 42156 220788
rect 42208 220776 42214 220788
rect 56502 220776 56508 220788
rect 42208 220748 56508 220776
rect 42208 220736 42214 220748
rect 56502 220736 56508 220748
rect 56560 220736 56566 220788
rect 344830 220736 344836 220788
rect 344888 220776 344894 220788
rect 412910 220776 412916 220788
rect 344888 220748 412916 220776
rect 344888 220736 344894 220748
rect 412910 220736 412916 220748
rect 412968 220736 412974 220788
rect 349154 220668 349160 220720
rect 349212 220708 349218 220720
rect 423030 220708 423036 220720
rect 349212 220680 423036 220708
rect 349212 220668 349218 220680
rect 423030 220668 423036 220680
rect 423088 220668 423094 220720
rect 347682 220600 347688 220652
rect 347740 220640 347746 220652
rect 419718 220640 419724 220652
rect 347740 220612 419724 220640
rect 347740 220600 347746 220612
rect 419718 220600 419724 220612
rect 419776 220600 419782 220652
rect 350534 220532 350540 220584
rect 350592 220572 350598 220584
rect 426342 220572 426348 220584
rect 350592 220544 426348 220572
rect 350592 220532 350598 220544
rect 426342 220532 426348 220544
rect 426400 220532 426406 220584
rect 142706 220464 142712 220516
rect 142764 220504 142770 220516
rect 229646 220504 229652 220516
rect 142764 220476 229652 220504
rect 142764 220464 142770 220476
rect 229646 220464 229652 220476
rect 229704 220464 229710 220516
rect 352006 220464 352012 220516
rect 352064 220504 352070 220516
rect 429746 220504 429752 220516
rect 352064 220476 429752 220504
rect 352064 220464 352070 220476
rect 429746 220464 429752 220476
rect 429804 220464 429810 220516
rect 139302 220396 139308 220448
rect 139360 220436 139366 220448
rect 228266 220436 228272 220448
rect 139360 220408 228272 220436
rect 139360 220396 139366 220408
rect 228266 220396 228272 220408
rect 228324 220396 228330 220448
rect 353386 220396 353392 220448
rect 353444 220436 353450 220448
rect 433334 220436 433340 220448
rect 353444 220408 433340 220436
rect 353444 220396 353450 220408
rect 433334 220396 433340 220408
rect 433392 220396 433398 220448
rect 135990 220328 135996 220380
rect 136048 220368 136054 220380
rect 226610 220368 226616 220380
rect 136048 220340 226616 220368
rect 136048 220328 136054 220340
rect 226610 220328 226616 220340
rect 226668 220328 226674 220380
rect 357618 220328 357624 220380
rect 357676 220368 357682 220380
rect 440694 220368 440700 220380
rect 357676 220340 440700 220368
rect 357676 220328 357682 220340
rect 440694 220328 440700 220340
rect 440752 220328 440758 220380
rect 132402 220260 132408 220312
rect 132460 220300 132466 220312
rect 225414 220300 225420 220312
rect 132460 220272 225420 220300
rect 132460 220260 132466 220272
rect 225414 220260 225420 220272
rect 225472 220260 225478 220312
rect 355042 220260 355048 220312
rect 355100 220300 355106 220312
rect 436462 220300 436468 220312
rect 355100 220272 436468 220300
rect 355100 220260 355106 220272
rect 436462 220260 436468 220272
rect 436520 220260 436526 220312
rect 129274 220192 129280 220244
rect 129332 220232 129338 220244
rect 223942 220232 223948 220244
rect 129332 220204 223948 220232
rect 129332 220192 129338 220204
rect 223942 220192 223948 220204
rect 224000 220192 224006 220244
rect 360194 220192 360200 220244
rect 360252 220232 360258 220244
rect 447410 220232 447416 220244
rect 360252 220204 447416 220232
rect 360252 220192 360258 220204
rect 447410 220192 447416 220204
rect 447468 220192 447474 220244
rect 125870 220124 125876 220176
rect 125928 220164 125934 220176
rect 222286 220164 222292 220176
rect 125928 220136 222292 220164
rect 125928 220124 125934 220136
rect 222286 220124 222292 220136
rect 222344 220124 222350 220176
rect 367646 220124 367652 220176
rect 367704 220164 367710 220176
rect 466730 220164 466736 220176
rect 367704 220136 466736 220164
rect 367704 220124 367710 220136
rect 466730 220124 466736 220136
rect 466788 220124 466794 220176
rect 122466 220056 122472 220108
rect 122524 220096 122530 220108
rect 221090 220096 221096 220108
rect 122524 220068 221096 220096
rect 122524 220056 122530 220068
rect 221090 220056 221096 220068
rect 221148 220056 221154 220108
rect 370130 220056 370136 220108
rect 370188 220096 370194 220108
rect 470962 220096 470968 220108
rect 370188 220068 470968 220096
rect 370188 220056 370194 220068
rect 470962 220056 470968 220068
rect 471020 220056 471026 220108
rect 53742 219988 53748 220040
rect 53800 220028 53806 220040
rect 651282 220028 651288 220040
rect 53800 220000 651288 220028
rect 53800 219988 53806 220000
rect 651282 219988 651288 220000
rect 651340 219988 651346 220040
rect 53834 219920 53840 219972
rect 53892 219960 53898 219972
rect 655514 219960 655520 219972
rect 53892 219932 655520 219960
rect 53892 219920 53898 219932
rect 655514 219920 655520 219932
rect 655572 219920 655578 219972
rect 56594 219852 56600 219904
rect 56652 219892 56658 219904
rect 664346 219892 664352 219904
rect 56652 219864 664352 219892
rect 56652 219852 56658 219864
rect 664346 219852 664352 219864
rect 664404 219852 664410 219904
rect 56686 219784 56692 219836
rect 56744 219824 56750 219836
rect 663886 219824 663892 219836
rect 56744 219796 663892 219824
rect 56744 219784 56750 219796
rect 663886 219784 663892 219796
rect 663944 219784 663950 219836
rect 45738 219716 45744 219768
rect 45796 219756 45802 219768
rect 656894 219756 656900 219768
rect 45796 219728 656900 219756
rect 45796 219716 45802 219728
rect 656894 219716 656900 219728
rect 656952 219716 656958 219768
rect 50982 219648 50988 219700
rect 51040 219688 51046 219700
rect 662966 219688 662972 219700
rect 51040 219660 662972 219688
rect 51040 219648 51046 219660
rect 662966 219648 662972 219660
rect 663024 219648 663030 219700
rect 675570 219620 675576 219632
rect 675566 219592 675576 219620
rect 675570 219580 675576 219592
rect 675628 219620 675634 219632
rect 676030 219620 676036 219632
rect 675628 219592 676036 219620
rect 675628 219580 675634 219592
rect 676030 219580 676036 219592
rect 676088 219580 676094 219632
rect 675662 219552 675668 219564
rect 675660 219524 675668 219552
rect 675662 219512 675668 219524
rect 675720 219552 675726 219564
rect 675938 219552 675944 219564
rect 675720 219524 675944 219552
rect 675720 219512 675726 219524
rect 675938 219512 675944 219524
rect 675996 219512 676002 219564
rect 48590 219444 48596 219496
rect 48648 219484 48654 219496
rect 662506 219484 662512 219496
rect 48648 219456 662512 219484
rect 48648 219444 48654 219456
rect 662506 219444 662512 219456
rect 662564 219444 662570 219496
rect 346302 219308 346308 219360
rect 346360 219348 346366 219360
rect 416222 219348 416228 219360
rect 346360 219320 416228 219348
rect 346360 219308 346366 219320
rect 416222 219308 416228 219320
rect 416280 219308 416286 219360
rect 343450 219240 343456 219292
rect 343508 219280 343514 219292
rect 409506 219280 409512 219292
rect 343508 219252 409512 219280
rect 343508 219240 343514 219252
rect 409506 219240 409512 219252
rect 409564 219240 409570 219292
rect 525794 218424 525800 218476
rect 525852 218464 525858 218476
rect 613102 218464 613108 218476
rect 525852 218436 613108 218464
rect 525852 218424 525858 218436
rect 613102 218424 613108 218436
rect 613160 218424 613166 218476
rect 523402 218356 523408 218408
rect 523460 218396 523466 218408
rect 612642 218396 612648 218408
rect 523460 218368 612648 218396
rect 523460 218356 523466 218368
rect 612642 218356 612648 218368
rect 612700 218356 612706 218408
rect 520826 218288 520832 218340
rect 520884 218328 520890 218340
rect 612182 218328 612188 218340
rect 520884 218300 612188 218328
rect 520884 218288 520890 218300
rect 612182 218288 612188 218300
rect 612240 218288 612246 218340
rect 674466 218288 674472 218340
rect 674524 218328 674530 218340
rect 676030 218328 676036 218340
rect 674524 218300 676036 218328
rect 674524 218288 674530 218300
rect 676030 218288 676036 218300
rect 676088 218288 676094 218340
rect 518710 218220 518716 218272
rect 518768 218260 518774 218272
rect 611722 218260 611728 218272
rect 518768 218232 611728 218260
rect 518768 218220 518774 218232
rect 611722 218220 611728 218232
rect 611780 218220 611786 218272
rect 513466 218152 513472 218204
rect 513524 218192 513530 218204
rect 515766 218192 515772 218204
rect 513524 218164 515772 218192
rect 513524 218152 513530 218164
rect 515766 218152 515772 218164
rect 515824 218192 515830 218204
rect 611262 218192 611268 218204
rect 515824 218164 611268 218192
rect 515824 218152 515830 218164
rect 611262 218152 611268 218164
rect 611320 218152 611326 218204
rect 490282 218084 490288 218136
rect 490340 218124 490346 218136
rect 607122 218124 607128 218136
rect 490340 218096 607128 218124
rect 490340 218084 490346 218096
rect 607122 218084 607128 218096
rect 607180 218084 607186 218136
rect 487154 218016 487160 218068
rect 487212 218056 487218 218068
rect 606662 218056 606668 218068
rect 487212 218028 606668 218056
rect 487212 218016 487218 218028
rect 606662 218016 606668 218028
rect 606720 218016 606726 218068
rect 674742 218016 674748 218068
rect 674800 218056 674806 218068
rect 676030 218056 676036 218068
rect 674800 218028 676036 218056
rect 674800 218016 674806 218028
rect 676030 218016 676036 218028
rect 676088 218016 676094 218068
rect 8202 217880 8208 217932
rect 8260 217920 8266 217932
rect 8260 217892 33134 217920
rect 8260 217880 8266 217892
rect 33106 217580 33134 217892
rect 61838 217812 61844 217864
rect 61896 217852 61902 217864
rect 62942 217852 62948 217864
rect 61896 217824 62948 217852
rect 61896 217812 61902 217824
rect 62942 217812 62948 217824
rect 63000 217812 63006 217864
rect 418154 217812 418160 217864
rect 418212 217852 418218 217864
rect 418614 217852 418620 217864
rect 418212 217824 418620 217852
rect 418212 217812 418218 217824
rect 418614 217812 418620 217824
rect 418672 217812 418678 217864
rect 665726 217580 665732 217592
rect 33106 217552 665732 217580
rect 665726 217540 665732 217552
rect 665784 217540 665790 217592
rect 567976 217472 567982 217524
rect 568034 217512 568040 217524
rect 635458 217512 635464 217524
rect 568034 217484 635464 217512
rect 568034 217472 568040 217484
rect 635458 217472 635464 217484
rect 635516 217472 635522 217524
rect 560754 217404 560760 217456
rect 560812 217444 560818 217456
rect 634078 217444 634084 217456
rect 560812 217416 634084 217444
rect 560812 217404 560818 217416
rect 634078 217404 634084 217416
rect 634136 217404 634142 217456
rect 565722 217336 565728 217388
rect 565780 217376 565786 217388
rect 634998 217376 635004 217388
rect 565780 217348 635004 217376
rect 565780 217336 565786 217348
rect 634998 217336 635004 217348
rect 635056 217336 635062 217388
rect 555694 217268 555700 217320
rect 555752 217308 555758 217320
rect 633158 217308 633164 217320
rect 555752 217280 633164 217308
rect 555752 217268 555758 217280
rect 633158 217268 633164 217280
rect 633216 217268 633222 217320
rect 550634 217200 550640 217252
rect 550692 217240 550698 217252
rect 632238 217240 632244 217252
rect 550692 217212 632244 217240
rect 550692 217200 550698 217212
rect 632238 217200 632244 217212
rect 632296 217200 632302 217252
rect 511074 217132 511080 217184
rect 511132 217172 511138 217184
rect 523034 217172 523040 217184
rect 511132 217144 523040 217172
rect 511132 217132 511138 217144
rect 523034 217132 523040 217144
rect 523092 217132 523098 217184
rect 545390 217132 545396 217184
rect 545448 217172 545454 217184
rect 631318 217172 631324 217184
rect 545448 217144 631324 217172
rect 545448 217132 545454 217144
rect 631318 217132 631324 217144
rect 631376 217132 631382 217184
rect 489270 217064 489276 217116
rect 489328 217104 489334 217116
rect 500126 217104 500132 217116
rect 489328 217076 500132 217104
rect 489328 217064 489334 217076
rect 500126 217064 500132 217076
rect 500184 217064 500190 217116
rect 515306 217064 515312 217116
rect 515364 217104 515370 217116
rect 516042 217104 516048 217116
rect 515364 217076 516048 217104
rect 515364 217064 515370 217076
rect 516042 217064 516048 217076
rect 516100 217064 516106 217116
rect 532786 217064 532792 217116
rect 532844 217104 532850 217116
rect 628926 217104 628932 217116
rect 532844 217076 628932 217104
rect 532844 217064 532850 217076
rect 628926 217064 628932 217076
rect 628984 217064 628990 217116
rect 418522 216996 418528 217048
rect 418580 217036 418586 217048
rect 639690 217036 639696 217048
rect 418580 217008 639696 217036
rect 418580 216996 418586 217008
rect 639690 216996 639696 217008
rect 639748 216996 639754 217048
rect 418430 216928 418436 216980
rect 418488 216968 418494 216980
rect 640610 216968 640616 216980
rect 418488 216940 640616 216968
rect 418488 216928 418494 216940
rect 640610 216928 640616 216940
rect 640668 216928 640674 216980
rect 418614 216860 418620 216912
rect 418672 216900 418678 216912
rect 640150 216900 640156 216912
rect 418672 216872 640156 216900
rect 418672 216860 418678 216872
rect 640150 216860 640156 216872
rect 640208 216860 640214 216912
rect 417878 216792 417884 216844
rect 417936 216832 417942 216844
rect 641070 216832 641076 216844
rect 417936 216804 641076 216832
rect 417936 216792 417942 216804
rect 641070 216792 641076 216804
rect 641128 216792 641134 216844
rect 62022 216724 62028 216776
rect 62080 216764 62086 216776
rect 648522 216764 648528 216776
rect 62080 216736 648528 216764
rect 62080 216724 62086 216736
rect 648522 216724 648528 216736
rect 648580 216724 648586 216776
rect 41506 216656 41512 216708
rect 41564 216696 41570 216708
rect 59354 216696 59360 216708
rect 41564 216668 59360 216696
rect 41564 216656 41570 216668
rect 59354 216656 59360 216668
rect 59412 216656 59418 216708
rect 62942 216656 62948 216708
rect 63000 216696 63006 216708
rect 663426 216696 663432 216708
rect 63000 216668 663432 216696
rect 63000 216656 63006 216668
rect 663426 216656 663432 216668
rect 663484 216656 663490 216708
rect 674650 216656 674656 216708
rect 674708 216696 674714 216708
rect 676030 216696 676036 216708
rect 674708 216668 676036 216696
rect 674708 216656 674714 216668
rect 676030 216656 676036 216668
rect 676088 216656 676094 216708
rect 41414 216588 41420 216640
rect 41472 216628 41478 216640
rect 59262 216628 59268 216640
rect 41472 216600 59268 216628
rect 41472 216588 41478 216600
rect 59262 216588 59268 216600
rect 59320 216588 59326 216640
rect 499298 216520 499304 216572
rect 499356 216560 499362 216572
rect 499356 216532 500356 216560
rect 499356 216520 499362 216532
rect 492582 216452 492588 216504
rect 492640 216492 492646 216504
rect 492640 216464 500264 216492
rect 492640 216452 492646 216464
rect 484210 216384 484216 216436
rect 484268 216384 484274 216436
rect 486694 216384 486700 216436
rect 486752 216384 486758 216436
rect 490098 216384 490104 216436
rect 490156 216384 490162 216436
rect 496630 216384 496636 216436
rect 496688 216384 496694 216436
rect 500126 216384 500132 216436
rect 500184 216384 500190 216436
rect 484228 215540 484256 216384
rect 486712 215608 486740 216384
rect 490116 216356 490144 216384
rect 490116 216328 495204 216356
rect 495176 215676 495204 216328
rect 496648 215744 496676 216384
rect 500144 215812 500172 216384
rect 500236 215948 500264 216464
rect 500328 216288 500356 216532
rect 506106 216520 506112 216572
rect 506164 216560 506170 216572
rect 506164 216532 522988 216560
rect 506164 216520 506170 216532
rect 501046 216452 501052 216504
rect 501104 216492 501110 216504
rect 501104 216464 517560 216492
rect 501104 216452 501110 216464
rect 505002 216384 505008 216436
rect 505060 216424 505066 216436
rect 505060 216396 509832 216424
rect 505060 216384 505066 216396
rect 500328 216260 507854 216288
rect 507826 215948 507854 216260
rect 509804 216016 509832 216396
rect 509938 216404 509990 216410
rect 516042 216384 516048 216436
rect 516100 216384 516106 216436
rect 509938 216346 509990 216352
rect 509950 216084 509978 216346
rect 516060 216152 516088 216384
rect 517532 216220 517560 216464
rect 522850 216384 522856 216436
rect 522908 216384 522914 216436
rect 522868 216288 522896 216384
rect 522960 216356 522988 216532
rect 538030 216520 538036 216572
rect 538088 216560 538094 216572
rect 629938 216560 629944 216572
rect 538088 216532 629944 216560
rect 538088 216520 538094 216532
rect 629938 216520 629944 216532
rect 629996 216520 630002 216572
rect 666554 216520 666560 216572
rect 666612 216560 666618 216572
rect 666830 216560 666836 216572
rect 666612 216532 666836 216560
rect 666612 216520 666618 216532
rect 666830 216520 666836 216532
rect 666888 216520 666894 216572
rect 523034 216452 523040 216504
rect 523092 216492 523098 216504
rect 523092 216464 527174 216492
rect 523092 216452 523098 216464
rect 527146 216424 527174 216464
rect 527726 216452 527732 216504
rect 527784 216492 527790 216504
rect 628006 216492 628012 216504
rect 527784 216464 628012 216492
rect 527784 216452 527790 216464
rect 628006 216452 628012 216464
rect 628064 216452 628070 216504
rect 610342 216424 610348 216436
rect 527146 216396 610348 216424
rect 610342 216384 610348 216396
rect 610400 216384 610406 216436
rect 609422 216356 609428 216368
rect 522960 216328 609428 216356
rect 609422 216316 609428 216328
rect 609480 216316 609486 216368
rect 627086 216288 627092 216300
rect 522868 216260 627092 216288
rect 627086 216248 627092 216260
rect 627144 216248 627150 216300
rect 674282 216248 674288 216300
rect 674340 216288 674346 216300
rect 675938 216288 675944 216300
rect 674340 216260 675944 216288
rect 674340 216248 674346 216260
rect 675938 216248 675944 216260
rect 675996 216248 676002 216300
rect 608502 216220 608508 216232
rect 517532 216192 608508 216220
rect 608502 216180 608508 216192
rect 608560 216180 608566 216232
rect 625706 216152 625712 216164
rect 516060 216124 625712 216152
rect 625706 216112 625712 216124
rect 625764 216112 625770 216164
rect 624786 216084 624792 216096
rect 509950 216056 624792 216084
rect 624786 216044 624792 216056
rect 624844 216044 624850 216096
rect 623866 216016 623872 216028
rect 509804 215988 623872 216016
rect 623866 215976 623872 215988
rect 623924 215976 623930 216028
rect 622946 215948 622952 215960
rect 500236 215920 500448 215948
rect 507826 215920 622952 215948
rect 500420 215880 500448 215920
rect 622946 215908 622952 215920
rect 623004 215908 623010 215960
rect 622026 215880 622032 215892
rect 500420 215852 622032 215880
rect 622026 215840 622032 215852
rect 622084 215840 622090 215892
rect 674926 215840 674932 215892
rect 674984 215880 674990 215892
rect 675846 215880 675852 215892
rect 674984 215852 675852 215880
rect 674984 215840 674990 215852
rect 675846 215840 675852 215852
rect 675904 215840 675910 215892
rect 621474 215812 621480 215824
rect 500144 215784 621480 215812
rect 621474 215772 621480 215784
rect 621532 215772 621538 215824
rect 637390 215744 637396 215756
rect 496648 215716 637396 215744
rect 637390 215704 637396 215716
rect 637448 215704 637454 215756
rect 636378 215676 636384 215688
rect 495176 215648 636384 215676
rect 636378 215636 636384 215648
rect 636436 215636 636442 215688
rect 638310 215608 638316 215620
rect 486712 215580 638316 215608
rect 638310 215568 638316 215580
rect 638368 215568 638374 215620
rect 638770 215540 638776 215552
rect 484228 215512 638776 215540
rect 638770 215500 638776 215512
rect 638828 215500 638834 215552
rect 673546 215500 673552 215552
rect 673604 215540 673610 215552
rect 675754 215540 675760 215552
rect 673604 215512 675760 215540
rect 673604 215500 673610 215512
rect 675754 215500 675760 215512
rect 675812 215500 675818 215552
rect 48222 215432 48228 215484
rect 48280 215472 48286 215484
rect 666186 215472 666192 215484
rect 48280 215444 666192 215472
rect 48280 215432 48286 215444
rect 666186 215432 666192 215444
rect 666244 215432 666250 215484
rect 673730 215432 673736 215484
rect 673788 215472 673794 215484
rect 675846 215472 675852 215484
rect 673788 215444 675852 215472
rect 673788 215432 673794 215444
rect 675846 215432 675852 215444
rect 675904 215432 675910 215484
rect 31662 215364 31668 215416
rect 31720 215404 31726 215416
rect 665266 215404 665272 215416
rect 31720 215376 665272 215404
rect 31720 215364 31726 215376
rect 665266 215364 665272 215376
rect 665324 215364 665330 215416
rect 674558 215364 674564 215416
rect 674616 215404 674622 215416
rect 675938 215404 675944 215416
rect 674616 215376 675944 215404
rect 674616 215364 674622 215376
rect 675938 215364 675944 215376
rect 675996 215364 676002 215416
rect 582282 215296 582288 215348
rect 582340 215336 582346 215348
rect 600038 215336 600044 215348
rect 582340 215308 600044 215336
rect 582340 215296 582346 215308
rect 600038 215296 600044 215308
rect 600096 215296 600102 215348
rect 674834 215296 674840 215348
rect 674892 215336 674898 215348
rect 676030 215336 676036 215348
rect 674892 215308 676036 215336
rect 674892 215296 674898 215308
rect 676030 215296 676036 215308
rect 676088 215296 676094 215348
rect 673638 214616 673644 214668
rect 673696 214656 673702 214668
rect 676030 214656 676036 214668
rect 673696 214628 676036 214656
rect 673696 214616 673702 214628
rect 676030 214616 676036 214628
rect 676088 214616 676094 214668
rect 41506 213256 41512 213308
rect 41564 213296 41570 213308
rect 666922 213296 666928 213308
rect 41564 213268 666928 213296
rect 41564 213256 41570 213268
rect 666922 213256 666928 213268
rect 666980 213256 666986 213308
rect 582282 212576 582288 212628
rect 582340 212616 582346 212628
rect 599946 212616 599952 212628
rect 582340 212588 599952 212616
rect 582340 212576 582346 212588
rect 599946 212576 599952 212588
rect 600004 212576 600010 212628
rect 673454 212576 673460 212628
rect 673512 212616 673518 212628
rect 675938 212616 675944 212628
rect 673512 212588 675944 212616
rect 673512 212576 673518 212588
rect 675938 212576 675944 212588
rect 675996 212576 676002 212628
rect 580258 212508 580264 212560
rect 580316 212548 580322 212560
rect 599854 212548 599860 212560
rect 580316 212520 599860 212548
rect 580316 212508 580322 212520
rect 599854 212508 599860 212520
rect 599912 212508 599918 212560
rect 673822 212508 673828 212560
rect 673880 212548 673886 212560
rect 676030 212548 676036 212560
rect 673880 212520 676036 212548
rect 673880 212508 673886 212520
rect 676030 212508 676036 212520
rect 676088 212508 676094 212560
rect 672718 212032 672724 212084
rect 672776 212072 672782 212084
rect 676030 212072 676036 212084
rect 672776 212044 676036 212072
rect 672776 212032 672782 212044
rect 676030 212032 676036 212044
rect 676088 212032 676094 212084
rect 662782 210060 662788 210112
rect 662840 210100 662846 210112
rect 664438 210100 664444 210112
rect 662840 210072 664444 210100
rect 662840 210060 662846 210072
rect 664438 210060 664444 210072
rect 664496 210060 664502 210112
rect 582282 209856 582288 209908
rect 582340 209896 582346 209908
rect 601142 209896 601148 209908
rect 582340 209868 601148 209896
rect 582340 209856 582346 209868
rect 601142 209856 601148 209868
rect 601200 209856 601206 209908
rect 580074 209788 580080 209840
rect 580132 209828 580138 209840
rect 600774 209828 600780 209840
rect 580132 209800 600780 209828
rect 580132 209788 580138 209800
rect 600774 209788 600780 209800
rect 600832 209788 600838 209840
rect 641806 209788 641812 209840
rect 641864 209828 641870 209840
rect 642082 209828 642088 209840
rect 641864 209800 642088 209828
rect 641864 209788 641870 209800
rect 642082 209788 642088 209800
rect 642140 209788 642146 209840
rect 644658 209788 644664 209840
rect 644716 209828 644722 209840
rect 644934 209828 644940 209840
rect 644716 209800 644940 209828
rect 644716 209788 644722 209800
rect 644934 209788 644940 209800
rect 644992 209788 644998 209840
rect 647418 209788 647424 209840
rect 647476 209828 647482 209840
rect 647694 209828 647700 209840
rect 647476 209800 647700 209828
rect 647476 209788 647482 209800
rect 647694 209788 647700 209800
rect 647752 209788 647758 209840
rect 673454 207272 673460 207324
rect 673512 207272 673518 207324
rect 582282 207068 582288 207120
rect 582340 207108 582346 207120
rect 599670 207108 599676 207120
rect 582340 207080 599676 207108
rect 582340 207068 582346 207080
rect 599670 207068 599676 207080
rect 599728 207068 599734 207120
rect 673472 207052 673500 207272
rect 673546 207068 673552 207120
rect 673604 207108 673610 207120
rect 674926 207108 674932 207120
rect 673604 207080 674932 207108
rect 673604 207068 673610 207080
rect 674926 207068 674932 207080
rect 674984 207068 674990 207120
rect 581454 207000 581460 207052
rect 581512 207040 581518 207052
rect 601602 207040 601608 207052
rect 581512 207012 601608 207040
rect 581512 207000 581518 207012
rect 601602 207000 601608 207012
rect 601660 207000 601666 207052
rect 673454 207000 673460 207052
rect 673512 207000 673518 207052
rect 674926 206320 674932 206372
rect 674984 206360 674990 206372
rect 675386 206360 675392 206372
rect 674984 206332 675392 206360
rect 674984 206320 674990 206332
rect 675386 206320 675392 206332
rect 675444 206320 675450 206372
rect 675018 206252 675024 206304
rect 675076 206292 675082 206304
rect 675754 206292 675760 206304
rect 675076 206264 675760 206292
rect 675076 206252 675082 206264
rect 675754 206252 675760 206264
rect 675812 206252 675818 206304
rect 675202 206184 675208 206236
rect 675260 206224 675266 206236
rect 675478 206224 675484 206236
rect 675260 206196 675484 206224
rect 675260 206184 675266 206196
rect 675478 206184 675484 206196
rect 675536 206184 675542 206236
rect 675662 206184 675668 206236
rect 675720 206184 675726 206236
rect 674742 205572 674748 205624
rect 674800 205612 674806 205624
rect 675386 205612 675392 205624
rect 674800 205584 675392 205612
rect 674800 205572 674806 205584
rect 675386 205572 675392 205584
rect 675444 205572 675450 205624
rect 675680 205544 675708 206184
rect 674760 205516 675708 205544
rect 674760 205488 674788 205516
rect 674742 205436 674748 205488
rect 674800 205436 674806 205488
rect 38470 205028 38476 205080
rect 38528 205068 38534 205080
rect 43530 205068 43536 205080
rect 38528 205040 43536 205068
rect 38528 205028 38534 205040
rect 43530 205028 43536 205040
rect 43588 205028 43594 205080
rect 674834 204960 674840 205012
rect 674892 205000 674898 205012
rect 675386 205000 675392 205012
rect 674892 204972 675392 205000
rect 674892 204960 674898 204972
rect 675386 204960 675392 204972
rect 675444 204960 675450 205012
rect 38194 204416 38200 204468
rect 38252 204456 38258 204468
rect 43622 204456 43628 204468
rect 38252 204428 43628 204456
rect 38252 204416 38258 204428
rect 43622 204416 43628 204428
rect 43680 204416 43686 204468
rect 38102 204348 38108 204400
rect 38160 204388 38166 204400
rect 43346 204388 43352 204400
rect 38160 204360 43352 204388
rect 38160 204348 38166 204360
rect 43346 204348 43352 204360
rect 43404 204348 43410 204400
rect 674466 204348 674472 204400
rect 674524 204388 674530 204400
rect 675386 204388 675392 204400
rect 674524 204360 675392 204388
rect 674524 204348 674530 204360
rect 675386 204348 675392 204360
rect 675444 204348 675450 204400
rect 38562 204280 38568 204332
rect 38620 204320 38626 204332
rect 42242 204320 42248 204332
rect 38620 204292 42248 204320
rect 38620 204280 38626 204292
rect 42242 204280 42248 204292
rect 42300 204280 42306 204332
rect 582282 204280 582288 204332
rect 582340 204320 582346 204332
rect 599946 204320 599952 204332
rect 582340 204292 599952 204320
rect 582340 204280 582346 204292
rect 599946 204280 599952 204292
rect 600004 204280 600010 204332
rect 673362 204212 673368 204264
rect 673420 204252 673426 204264
rect 674466 204252 674472 204264
rect 673420 204224 674472 204252
rect 673420 204212 673426 204224
rect 674466 204212 674472 204224
rect 674524 204212 674530 204264
rect 674650 202716 674656 202768
rect 674708 202756 674714 202768
rect 675386 202756 675392 202768
rect 674708 202728 675392 202756
rect 674708 202716 674714 202728
rect 675386 202716 675392 202728
rect 675444 202716 675450 202768
rect 674558 201832 674564 201884
rect 674616 201872 674622 201884
rect 675386 201872 675392 201884
rect 674616 201844 675392 201872
rect 674616 201832 674622 201844
rect 675386 201832 675392 201844
rect 675444 201832 675450 201884
rect 581086 201560 581092 201612
rect 581144 201600 581150 201612
rect 599946 201600 599952 201612
rect 581144 201572 599952 201600
rect 581144 201560 581150 201572
rect 599946 201560 599952 201572
rect 600004 201560 600010 201612
rect 580718 201492 580724 201544
rect 580776 201532 580782 201544
rect 598934 201532 598940 201544
rect 580776 201504 598940 201532
rect 580776 201492 580782 201504
rect 598934 201492 598940 201504
rect 598992 201492 598998 201544
rect 673730 201492 673736 201544
rect 673788 201532 673794 201544
rect 675386 201532 675392 201544
rect 673788 201504 675392 201532
rect 673788 201492 673794 201504
rect 675386 201492 675392 201504
rect 675444 201492 675450 201544
rect 37918 201424 37924 201476
rect 37976 201464 37982 201476
rect 43714 201464 43720 201476
rect 37976 201436 43720 201464
rect 37976 201424 37982 201436
rect 43714 201424 43720 201436
rect 43772 201424 43778 201476
rect 38010 200880 38016 200932
rect 38068 200920 38074 200932
rect 43162 200920 43168 200932
rect 38068 200892 43168 200920
rect 38068 200880 38074 200892
rect 43162 200880 43168 200892
rect 43220 200880 43226 200932
rect 673822 200676 673828 200728
rect 673880 200716 673886 200728
rect 675386 200716 675392 200728
rect 673880 200688 675392 200716
rect 673880 200676 673886 200688
rect 675386 200676 675392 200688
rect 675444 200676 675450 200728
rect 581086 200064 581092 200116
rect 581144 200104 581150 200116
rect 599946 200104 599952 200116
rect 581144 200076 599952 200104
rect 581144 200064 581150 200076
rect 599946 200064 599952 200076
rect 600004 200064 600010 200116
rect 582282 198704 582288 198756
rect 582340 198744 582346 198756
rect 599946 198744 599952 198756
rect 582340 198716 599952 198744
rect 582340 198704 582346 198716
rect 599946 198704 599952 198716
rect 600004 198704 600010 198756
rect 674282 198364 674288 198416
rect 674340 198404 674346 198416
rect 675386 198404 675392 198416
rect 674340 198376 675392 198404
rect 674340 198364 674346 198376
rect 675386 198364 675392 198376
rect 675444 198364 675450 198416
rect 673454 197548 673460 197600
rect 673512 197588 673518 197600
rect 675478 197588 675484 197600
rect 673512 197560 675484 197588
rect 673512 197548 673518 197560
rect 675478 197548 675484 197560
rect 675536 197548 675542 197600
rect 582282 197344 582288 197396
rect 582340 197384 582346 197396
rect 599394 197384 599400 197396
rect 582340 197356 599400 197384
rect 582340 197344 582346 197356
rect 599394 197344 599400 197356
rect 599452 197344 599458 197396
rect 580718 197276 580724 197328
rect 580776 197316 580782 197328
rect 599946 197316 599952 197328
rect 580776 197288 599952 197316
rect 580776 197276 580782 197288
rect 599946 197276 599952 197288
rect 600004 197276 600010 197328
rect 673638 197140 673644 197192
rect 673696 197180 673702 197192
rect 675386 197180 675392 197192
rect 673696 197152 675392 197180
rect 673696 197140 673702 197152
rect 675386 197140 675392 197152
rect 675444 197140 675450 197192
rect 42242 196528 42248 196580
rect 42300 196568 42306 196580
rect 43162 196568 43168 196580
rect 42300 196540 43168 196568
rect 42300 196528 42306 196540
rect 43162 196528 43168 196540
rect 43220 196528 43226 196580
rect 675018 196528 675024 196580
rect 675076 196568 675082 196580
rect 675386 196568 675392 196580
rect 675076 196540 675392 196568
rect 675076 196528 675082 196540
rect 675386 196528 675392 196540
rect 675444 196528 675450 196580
rect 674742 196392 674748 196444
rect 674800 196432 674806 196444
rect 675018 196432 675024 196444
rect 674800 196404 675024 196432
rect 674800 196392 674806 196404
rect 675018 196392 675024 196404
rect 675076 196392 675082 196444
rect 674466 195304 674472 195356
rect 674524 195344 674530 195356
rect 675386 195344 675392 195356
rect 674524 195316 675392 195344
rect 674524 195304 674530 195316
rect 675386 195304 675392 195316
rect 675444 195304 675450 195356
rect 582190 194624 582196 194676
rect 582248 194664 582254 194676
rect 599946 194664 599952 194676
rect 582248 194636 599952 194664
rect 582248 194624 582254 194636
rect 599946 194624 599952 194636
rect 600004 194624 600010 194676
rect 582282 194556 582288 194608
rect 582340 194596 582346 194608
rect 599854 194596 599860 194608
rect 582340 194568 599860 194596
rect 582340 194556 582346 194568
rect 599854 194556 599860 194568
rect 599912 194556 599918 194608
rect 675294 193536 675300 193588
rect 675352 193536 675358 193588
rect 42058 193468 42064 193520
rect 42116 193508 42122 193520
rect 42702 193508 42708 193520
rect 42116 193480 42708 193508
rect 42116 193468 42122 193480
rect 42702 193468 42708 193480
rect 42760 193468 42766 193520
rect 675312 193384 675340 193536
rect 675294 193332 675300 193384
rect 675352 193332 675358 193384
rect 674926 192856 674932 192908
rect 674984 192896 674990 192908
rect 675202 192896 675208 192908
rect 674984 192868 675208 192896
rect 674984 192856 674990 192868
rect 675202 192856 675208 192868
rect 675260 192856 675266 192908
rect 582282 191836 582288 191888
rect 582340 191876 582346 191888
rect 599486 191876 599492 191888
rect 582340 191848 599492 191876
rect 582340 191836 582346 191848
rect 599486 191836 599492 191848
rect 599544 191836 599550 191888
rect 581270 191768 581276 191820
rect 581328 191808 581334 191820
rect 599946 191808 599952 191820
rect 581328 191780 599952 191808
rect 581328 191768 581334 191780
rect 599946 191768 599952 191780
rect 600004 191768 600010 191820
rect 42334 191632 42340 191684
rect 42392 191672 42398 191684
rect 43070 191672 43076 191684
rect 42392 191644 43076 191672
rect 42392 191632 42398 191644
rect 43070 191632 43076 191644
rect 43128 191632 43134 191684
rect 673546 191632 673552 191684
rect 673604 191672 673610 191684
rect 675386 191672 675392 191684
rect 673604 191644 675392 191672
rect 673604 191632 673610 191644
rect 675386 191632 675392 191644
rect 675444 191632 675450 191684
rect 42058 191428 42064 191480
rect 42116 191468 42122 191480
rect 43254 191468 43260 191480
rect 42116 191440 43260 191468
rect 42116 191428 42122 191440
rect 43254 191428 43260 191440
rect 43312 191428 43318 191480
rect 579706 190408 579712 190460
rect 579764 190448 579770 190460
rect 599946 190448 599952 190460
rect 579764 190420 599952 190448
rect 579764 190408 579770 190420
rect 599946 190408 599952 190420
rect 600004 190408 600010 190460
rect 42334 190340 42340 190392
rect 42392 190380 42398 190392
rect 43346 190380 43352 190392
rect 42392 190352 43352 190380
rect 42392 190340 42398 190352
rect 43346 190340 43352 190352
rect 43404 190340 43410 190392
rect 42242 189796 42248 189848
rect 42300 189836 42306 189848
rect 43438 189836 43444 189848
rect 42300 189808 43444 189836
rect 42300 189796 42306 189808
rect 43438 189796 43444 189808
rect 43496 189796 43502 189848
rect 42334 189728 42340 189780
rect 42392 189768 42398 189780
rect 43714 189768 43720 189780
rect 42392 189740 43720 189768
rect 42392 189728 42398 189740
rect 43714 189728 43720 189740
rect 43772 189728 43778 189780
rect 42426 189116 42432 189168
rect 42484 189156 42490 189168
rect 43622 189156 43628 189168
rect 42484 189128 43628 189156
rect 42484 189116 42490 189128
rect 43622 189116 43628 189128
rect 43680 189116 43686 189168
rect 582282 187620 582288 187672
rect 582340 187660 582346 187672
rect 601510 187660 601516 187672
rect 582340 187632 601516 187660
rect 582340 187620 582346 187632
rect 601510 187620 601516 187632
rect 601568 187620 601574 187672
rect 579890 187552 579896 187604
rect 579948 187592 579954 187604
rect 601602 187592 601608 187604
rect 579948 187564 601608 187592
rect 579948 187552 579954 187564
rect 601602 187552 601608 187564
rect 601660 187552 601666 187604
rect 42334 186668 42340 186720
rect 42392 186708 42398 186720
rect 43530 186708 43536 186720
rect 42392 186680 43536 186708
rect 42392 186668 42398 186680
rect 43530 186668 43536 186680
rect 43588 186668 43594 186720
rect 580258 184832 580264 184884
rect 580316 184872 580322 184884
rect 599946 184872 599952 184884
rect 580316 184844 599952 184872
rect 580316 184832 580322 184844
rect 599946 184832 599952 184844
rect 600004 184832 600010 184884
rect 580902 184764 580908 184816
rect 580960 184804 580966 184816
rect 599118 184804 599124 184816
rect 580960 184776 599124 184804
rect 580960 184764 580966 184776
rect 599118 184764 599124 184776
rect 599176 184764 599182 184816
rect 42150 182112 42156 182164
rect 42208 182152 42214 182164
rect 48498 182152 48504 182164
rect 42208 182124 48504 182152
rect 42208 182112 42214 182124
rect 48498 182112 48504 182124
rect 48556 182112 48562 182164
rect 580626 182112 580632 182164
rect 580684 182152 580690 182164
rect 600038 182152 600044 182164
rect 580684 182124 600044 182152
rect 580684 182112 580690 182124
rect 600038 182112 600044 182124
rect 600096 182112 600102 182164
rect 580534 182044 580540 182096
rect 580592 182084 580598 182096
rect 599854 182084 599860 182096
rect 580592 182056 599860 182084
rect 580592 182044 580598 182056
rect 599854 182044 599860 182056
rect 599912 182044 599918 182096
rect 580718 179324 580724 179376
rect 580776 179364 580782 179376
rect 598934 179364 598940 179376
rect 580776 179336 598940 179364
rect 580776 179324 580782 179336
rect 598934 179324 598940 179336
rect 598992 179324 598998 179376
rect 581086 179256 581092 179308
rect 581144 179296 581150 179308
rect 599946 179296 599952 179308
rect 581144 179268 599952 179296
rect 581144 179256 581150 179268
rect 599946 179256 599952 179268
rect 600004 179256 600010 179308
rect 666830 178032 666836 178084
rect 666888 178032 666894 178084
rect 666738 177828 666744 177880
rect 666796 177868 666802 177880
rect 666848 177868 666876 178032
rect 666796 177840 666876 177868
rect 666796 177828 666802 177840
rect 670326 177080 670332 177132
rect 670384 177120 670390 177132
rect 676030 177120 676036 177132
rect 670384 177092 676036 177120
rect 670384 177080 670390 177092
rect 676030 177080 676036 177092
rect 676088 177080 676094 177132
rect 670234 176944 670240 176996
rect 670292 176984 670298 176996
rect 675938 176984 675944 176996
rect 670292 176956 675944 176984
rect 670292 176944 670298 176956
rect 675938 176944 675944 176956
rect 675996 176944 676002 176996
rect 667014 176808 667020 176860
rect 667072 176848 667078 176860
rect 675846 176848 675852 176860
rect 667072 176820 675852 176848
rect 667072 176808 667078 176820
rect 675846 176808 675852 176820
rect 675904 176808 675910 176860
rect 581086 176672 581092 176724
rect 581144 176712 581150 176724
rect 599946 176712 599952 176724
rect 581144 176684 599952 176712
rect 581144 176672 581150 176684
rect 599946 176672 599952 176684
rect 600004 176672 600010 176724
rect 581454 176604 581460 176656
rect 581512 176644 581518 176656
rect 600038 176644 600044 176656
rect 581512 176616 600044 176644
rect 581512 176604 581518 176616
rect 600038 176604 600044 176616
rect 600096 176604 600102 176656
rect 675202 176604 675208 176656
rect 675260 176644 675266 176656
rect 676030 176644 676036 176656
rect 675260 176616 676036 176644
rect 675260 176604 675266 176616
rect 676030 176604 676036 176616
rect 676088 176604 676094 176656
rect 675018 176332 675024 176384
rect 675076 176372 675082 176384
rect 676030 176372 676036 176384
rect 675076 176344 676036 176372
rect 675076 176332 675082 176344
rect 676030 176332 676036 176344
rect 676088 176332 676094 176384
rect 673362 175992 673368 176044
rect 673420 176032 673426 176044
rect 675938 176032 675944 176044
rect 673420 176004 675944 176032
rect 673420 175992 673426 176004
rect 675938 175992 675944 176004
rect 675996 175992 676002 176044
rect 674742 175516 674748 175568
rect 674800 175556 674806 175568
rect 676030 175556 676036 175568
rect 674800 175528 676036 175556
rect 674800 175516 674806 175528
rect 676030 175516 676036 175528
rect 676088 175516 676094 175568
rect 581638 173884 581644 173936
rect 581696 173924 581702 173936
rect 599946 173924 599952 173936
rect 581696 173896 599952 173924
rect 581696 173884 581702 173896
rect 599946 173884 599952 173896
rect 600004 173884 600010 173936
rect 674742 173884 674748 173936
rect 674800 173924 674806 173936
rect 676030 173924 676036 173936
rect 674800 173896 676036 173924
rect 674800 173884 674806 173896
rect 676030 173884 676036 173896
rect 676088 173884 676094 173936
rect 579706 173816 579712 173868
rect 579764 173856 579770 173868
rect 599854 173856 599860 173868
rect 579764 173828 599860 173856
rect 579764 173816 579770 173828
rect 599854 173816 599860 173828
rect 599912 173816 599918 173868
rect 582282 173748 582288 173800
rect 582340 173788 582346 173800
rect 600130 173788 600136 173800
rect 582340 173760 600136 173788
rect 582340 173748 582346 173760
rect 600130 173748 600136 173760
rect 600188 173748 600194 173800
rect 673546 172864 673552 172916
rect 673604 172904 673610 172916
rect 676030 172904 676036 172916
rect 673604 172876 676036 172904
rect 673604 172864 673610 172876
rect 676030 172864 676036 172876
rect 676088 172864 676094 172916
rect 674282 172048 674288 172100
rect 674340 172088 674346 172100
rect 675938 172088 675944 172100
rect 674340 172060 675944 172088
rect 674340 172048 674346 172060
rect 675938 172048 675944 172060
rect 675996 172048 676002 172100
rect 674834 171232 674840 171284
rect 674892 171272 674898 171284
rect 676030 171272 676036 171284
rect 674892 171244 676036 171272
rect 674892 171232 674898 171244
rect 676030 171232 676036 171244
rect 676088 171232 676094 171284
rect 582098 171164 582104 171216
rect 582156 171204 582162 171216
rect 599946 171204 599952 171216
rect 582156 171176 599952 171204
rect 582156 171164 582162 171176
rect 599946 171164 599952 171176
rect 600004 171164 600010 171216
rect 674558 171164 674564 171216
rect 674616 171204 674622 171216
rect 675938 171204 675944 171216
rect 674616 171176 675944 171204
rect 674616 171164 674622 171176
rect 675938 171164 675944 171176
rect 675996 171164 676002 171216
rect 579890 171096 579896 171148
rect 579948 171136 579954 171148
rect 599486 171136 599492 171148
rect 579948 171108 599492 171136
rect 579948 171096 579954 171108
rect 599486 171096 599492 171108
rect 599544 171096 599550 171148
rect 674650 171096 674656 171148
rect 674708 171136 674714 171148
rect 676030 171136 676036 171148
rect 674708 171108 676036 171136
rect 674708 171096 674714 171108
rect 676030 171096 676036 171108
rect 676088 171096 676094 171148
rect 582006 171028 582012 171080
rect 582064 171068 582070 171080
rect 599762 171068 599768 171080
rect 582064 171040 599768 171068
rect 582064 171028 582070 171040
rect 599762 171028 599768 171040
rect 599820 171028 599826 171080
rect 580534 170960 580540 171012
rect 580592 171000 580598 171012
rect 599670 171000 599676 171012
rect 580592 170972 599676 171000
rect 580592 170960 580598 170972
rect 599670 170960 599676 170972
rect 599728 170960 599734 171012
rect 666646 170144 666652 170196
rect 666704 170144 666710 170196
rect 666664 169992 666692 170144
rect 673730 170008 673736 170060
rect 673788 170048 673794 170060
rect 675938 170048 675944 170060
rect 673788 170020 675944 170048
rect 673788 170008 673794 170020
rect 675938 170008 675944 170020
rect 675996 170008 676002 170060
rect 666646 169940 666652 169992
rect 666704 169940 666710 169992
rect 674926 169600 674932 169652
rect 674984 169640 674990 169652
rect 676030 169640 676036 169652
rect 674984 169612 676036 169640
rect 674984 169600 674990 169612
rect 676030 169600 676036 169612
rect 676088 169600 676094 169652
rect 673638 169192 673644 169244
rect 673696 169232 673702 169244
rect 675938 169232 675944 169244
rect 673696 169204 675944 169232
rect 673696 169192 673702 169204
rect 675938 169192 675944 169204
rect 675996 169192 676002 169244
rect 675018 168920 675024 168972
rect 675076 168960 675082 168972
rect 676030 168960 676036 168972
rect 675076 168932 676036 168960
rect 675076 168920 675082 168932
rect 676030 168920 676036 168932
rect 676088 168920 676094 168972
rect 674466 168580 674472 168632
rect 674524 168620 674530 168632
rect 675938 168620 675944 168632
rect 674524 168592 675944 168620
rect 674524 168580 674530 168592
rect 675938 168580 675944 168592
rect 675996 168580 676002 168632
rect 580442 168512 580448 168564
rect 580500 168552 580506 168564
rect 599946 168552 599952 168564
rect 580500 168524 599952 168552
rect 580500 168512 580506 168524
rect 599946 168512 599952 168524
rect 600004 168512 600010 168564
rect 673822 168512 673828 168564
rect 673880 168552 673886 168564
rect 676030 168552 676036 168564
rect 673880 168524 676036 168552
rect 673880 168512 673886 168524
rect 676030 168512 676036 168524
rect 676088 168512 676094 168564
rect 579798 168444 579804 168496
rect 579856 168484 579862 168496
rect 599854 168484 599860 168496
rect 579856 168456 599860 168484
rect 579856 168444 579862 168456
rect 599854 168444 599860 168456
rect 599912 168444 599918 168496
rect 580258 168376 580264 168428
rect 580316 168416 580322 168428
rect 599486 168416 599492 168428
rect 580316 168388 599492 168416
rect 580316 168376 580322 168388
rect 599486 168376 599492 168388
rect 599544 168376 599550 168428
rect 580166 168308 580172 168360
rect 580224 168348 580230 168360
rect 600406 168348 600412 168360
rect 580224 168320 600412 168348
rect 580224 168308 580230 168320
rect 600406 168308 600412 168320
rect 600464 168308 600470 168360
rect 671982 167016 671988 167068
rect 672040 167056 672046 167068
rect 676030 167056 676036 167068
rect 672040 167028 676036 167056
rect 672040 167016 672046 167028
rect 676030 167016 676036 167028
rect 676088 167016 676094 167068
rect 582282 165724 582288 165776
rect 582340 165764 582346 165776
rect 600038 165764 600044 165776
rect 582340 165736 600044 165764
rect 582340 165724 582346 165736
rect 600038 165724 600044 165736
rect 600096 165724 600102 165776
rect 582190 165656 582196 165708
rect 582248 165696 582254 165708
rect 599946 165696 599952 165708
rect 582248 165668 599952 165696
rect 582248 165656 582254 165668
rect 599946 165656 599952 165668
rect 600004 165656 600010 165708
rect 581270 165588 581276 165640
rect 581328 165628 581334 165640
rect 599486 165628 599492 165640
rect 581328 165600 599492 165628
rect 581328 165588 581334 165600
rect 599486 165588 599492 165600
rect 599544 165588 599550 165640
rect 581822 165520 581828 165572
rect 581880 165560 581886 165572
rect 601326 165560 601332 165572
rect 581880 165532 601332 165560
rect 581880 165520 581886 165532
rect 601326 165520 601332 165532
rect 601384 165520 601390 165572
rect 673454 164840 673460 164892
rect 673512 164880 673518 164892
rect 673730 164880 673736 164892
rect 673512 164852 673736 164880
rect 673512 164840 673518 164852
rect 673730 164840 673736 164852
rect 673788 164840 673794 164892
rect 673822 164568 673828 164620
rect 673880 164608 673886 164620
rect 674282 164608 674288 164620
rect 673880 164580 674288 164608
rect 673880 164568 673886 164580
rect 674282 164568 674288 164580
rect 674340 164568 674346 164620
rect 674282 164432 674288 164484
rect 674340 164472 674346 164484
rect 674466 164472 674472 164484
rect 674340 164444 674472 164472
rect 674340 164432 674346 164444
rect 674466 164432 674472 164444
rect 674524 164432 674530 164484
rect 675110 164432 675116 164484
rect 675168 164472 675174 164484
rect 675386 164472 675392 164484
rect 675168 164444 675392 164472
rect 675168 164432 675174 164444
rect 675386 164432 675392 164444
rect 675444 164432 675450 164484
rect 674466 164296 674472 164348
rect 674524 164336 674530 164348
rect 674650 164336 674656 164348
rect 674524 164308 674656 164336
rect 674524 164296 674530 164308
rect 674650 164296 674656 164308
rect 674708 164296 674714 164348
rect 674650 164160 674656 164212
rect 674708 164200 674714 164212
rect 674926 164200 674932 164212
rect 674708 164172 674932 164200
rect 674708 164160 674714 164172
rect 674926 164160 674932 164172
rect 674984 164160 674990 164212
rect 675018 163956 675024 164008
rect 675076 163996 675082 164008
rect 675662 163996 675668 164008
rect 675076 163968 675668 163996
rect 675076 163956 675082 163968
rect 675662 163956 675668 163968
rect 675720 163956 675726 164008
rect 580074 162936 580080 162988
rect 580132 162976 580138 162988
rect 600038 162976 600044 162988
rect 580132 162948 600044 162976
rect 580132 162936 580138 162948
rect 600038 162936 600044 162948
rect 600096 162936 600102 162988
rect 581178 162868 581184 162920
rect 581236 162908 581242 162920
rect 599946 162908 599952 162920
rect 581236 162880 599952 162908
rect 581236 162868 581242 162880
rect 599946 162868 599952 162880
rect 600004 162868 600010 162920
rect 675754 161168 675760 161220
rect 675812 161168 675818 161220
rect 666830 160964 666836 161016
rect 666888 161004 666894 161016
rect 675386 161004 675392 161016
rect 666888 160976 675392 161004
rect 666888 160964 666894 160976
rect 675386 160964 675392 160976
rect 675444 160964 675450 161016
rect 582098 160216 582104 160268
rect 582156 160256 582162 160268
rect 599946 160256 599952 160268
rect 582156 160228 599952 160256
rect 582156 160216 582162 160228
rect 599946 160216 599952 160228
rect 600004 160216 600010 160268
rect 581638 160148 581644 160200
rect 581696 160188 581702 160200
rect 599854 160188 599860 160200
rect 581696 160160 599860 160188
rect 581696 160148 581702 160160
rect 599854 160148 599860 160160
rect 599912 160148 599918 160200
rect 675018 160148 675024 160200
rect 675076 160188 675082 160200
rect 675294 160188 675300 160200
rect 675076 160160 675300 160188
rect 675076 160148 675082 160160
rect 675294 160148 675300 160160
rect 675352 160148 675358 160200
rect 581730 160080 581736 160132
rect 581788 160120 581794 160132
rect 600038 160120 600044 160132
rect 581788 160092 600044 160120
rect 581788 160080 581794 160092
rect 600038 160080 600044 160092
rect 600096 160080 600102 160132
rect 675018 160012 675024 160064
rect 675076 160052 675082 160064
rect 675772 160052 675800 161168
rect 675076 160024 675800 160052
rect 675076 160012 675082 160024
rect 674742 159332 674748 159384
rect 674800 159372 674806 159384
rect 675478 159372 675484 159384
rect 674800 159344 675484 159372
rect 674800 159332 674806 159344
rect 675478 159332 675484 159344
rect 675536 159332 675542 159384
rect 674650 158040 674656 158092
rect 674708 158080 674714 158092
rect 675294 158080 675300 158092
rect 674708 158052 675300 158080
rect 674708 158040 674714 158052
rect 675294 158040 675300 158052
rect 675352 158040 675358 158092
rect 674834 157700 674840 157752
rect 674892 157740 674898 157752
rect 675478 157740 675484 157752
rect 674892 157712 675484 157740
rect 674892 157700 674898 157712
rect 675478 157700 675484 157712
rect 675536 157700 675542 157752
rect 581086 157496 581092 157548
rect 581144 157536 581150 157548
rect 599854 157536 599860 157548
rect 581144 157508 599860 157536
rect 581144 157496 581150 157508
rect 599854 157496 599860 157508
rect 599912 157496 599918 157548
rect 580902 157428 580908 157480
rect 580960 157468 580966 157480
rect 599946 157468 599952 157480
rect 580960 157440 599952 157468
rect 580960 157428 580966 157440
rect 599946 157428 599952 157440
rect 600004 157428 600010 157480
rect 580626 157360 580632 157412
rect 580684 157400 580690 157412
rect 600038 157400 600044 157412
rect 580684 157372 600044 157400
rect 580684 157360 580690 157372
rect 600038 157360 600044 157372
rect 600096 157360 600102 157412
rect 674466 156884 674472 156936
rect 674524 156924 674530 156936
rect 675386 156924 675392 156936
rect 674524 156896 675392 156924
rect 674524 156884 674530 156896
rect 675386 156884 675392 156896
rect 675444 156884 675450 156936
rect 674926 155864 674932 155916
rect 674984 155904 674990 155916
rect 675478 155904 675484 155916
rect 674984 155876 675484 155904
rect 674984 155864 674990 155876
rect 675478 155864 675484 155876
rect 675536 155864 675542 155916
rect 674282 155796 674288 155848
rect 674340 155836 674346 155848
rect 675294 155836 675300 155848
rect 674340 155808 675300 155836
rect 674340 155796 674346 155808
rect 675294 155796 675300 155808
rect 675352 155796 675358 155848
rect 580718 154640 580724 154692
rect 580776 154680 580782 154692
rect 599946 154680 599952 154692
rect 580776 154652 599952 154680
rect 580776 154640 580782 154652
rect 599946 154640 599952 154652
rect 600004 154640 600010 154692
rect 580534 154572 580540 154624
rect 580592 154612 580598 154624
rect 599854 154612 599860 154624
rect 580592 154584 599860 154612
rect 580592 154572 580598 154584
rect 599854 154572 599860 154584
rect 599912 154572 599918 154624
rect 673822 153348 673828 153400
rect 673880 153388 673886 153400
rect 675386 153388 675392 153400
rect 673880 153360 675392 153388
rect 673880 153348 673886 153360
rect 675386 153348 675392 153360
rect 675444 153348 675450 153400
rect 673638 152192 673644 152244
rect 673696 152232 673702 152244
rect 675294 152232 675300 152244
rect 673696 152204 675300 152232
rect 673696 152192 673702 152204
rect 675294 152192 675300 152204
rect 675352 152192 675358 152244
rect 582282 151920 582288 151972
rect 582340 151960 582346 151972
rect 599854 151960 599860 151972
rect 582340 151932 599860 151960
rect 582340 151920 582346 151932
rect 599854 151920 599860 151932
rect 599912 151920 599918 151972
rect 581822 151852 581828 151904
rect 581880 151892 581886 151904
rect 599946 151892 599952 151904
rect 581880 151864 599952 151892
rect 581880 151852 581886 151864
rect 599946 151852 599952 151864
rect 600004 151852 600010 151904
rect 580810 151784 580816 151836
rect 580868 151824 580874 151836
rect 600038 151824 600044 151836
rect 580868 151796 600044 151824
rect 580868 151784 580874 151796
rect 600038 151784 600044 151796
rect 600096 151784 600102 151836
rect 673730 151512 673736 151564
rect 673788 151552 673794 151564
rect 675294 151552 675300 151564
rect 673788 151524 675300 151552
rect 673788 151512 673794 151524
rect 675294 151512 675300 151524
rect 675352 151512 675358 151564
rect 675110 150424 675116 150476
rect 675168 150464 675174 150476
rect 675294 150464 675300 150476
rect 675168 150436 675300 150464
rect 675168 150424 675174 150436
rect 675294 150424 675300 150436
rect 675352 150424 675358 150476
rect 673454 150356 673460 150408
rect 673512 150396 673518 150408
rect 675386 150396 675392 150408
rect 673512 150368 675392 150396
rect 673512 150356 673518 150368
rect 675386 150356 675392 150368
rect 675444 150356 675450 150408
rect 582006 149200 582012 149252
rect 582064 149240 582070 149252
rect 600038 149240 600044 149252
rect 582064 149212 600044 149240
rect 582064 149200 582070 149212
rect 600038 149200 600044 149212
rect 600096 149200 600102 149252
rect 581546 149132 581552 149184
rect 581604 149172 581610 149184
rect 599854 149172 599860 149184
rect 581604 149144 599860 149172
rect 581604 149132 581610 149144
rect 599854 149132 599860 149144
rect 599912 149132 599918 149184
rect 581362 149064 581368 149116
rect 581420 149104 581426 149116
rect 599946 149104 599952 149116
rect 581420 149076 599952 149104
rect 581420 149064 581426 149076
rect 599946 149064 599952 149076
rect 600004 149064 600010 149116
rect 673546 148520 673552 148572
rect 673604 148560 673610 148572
rect 675386 148560 675392 148572
rect 673604 148532 675392 148560
rect 673604 148520 673610 148532
rect 675386 148520 675392 148532
rect 675444 148520 675450 148572
rect 674558 146684 674564 146736
rect 674616 146724 674622 146736
rect 675386 146724 675392 146736
rect 674616 146696 675392 146724
rect 674616 146684 674622 146696
rect 675386 146684 675392 146696
rect 675444 146684 675450 146736
rect 582190 146344 582196 146396
rect 582248 146384 582254 146396
rect 599854 146384 599860 146396
rect 582248 146356 599860 146384
rect 582248 146344 582254 146356
rect 599854 146344 599860 146356
rect 599912 146344 599918 146396
rect 581454 146276 581460 146328
rect 581512 146316 581518 146328
rect 599946 146316 599952 146328
rect 581512 146288 599952 146316
rect 581512 146276 581518 146288
rect 599946 146276 599952 146288
rect 600004 146276 600010 146328
rect 581914 143692 581920 143744
rect 581972 143732 581978 143744
rect 599854 143732 599860 143744
rect 581972 143704 599860 143732
rect 581972 143692 581978 143704
rect 599854 143692 599860 143704
rect 599912 143692 599918 143744
rect 581730 143624 581736 143676
rect 581788 143664 581794 143676
rect 599946 143664 599952 143676
rect 581788 143636 599952 143664
rect 581788 143624 581794 143636
rect 599946 143624 599952 143636
rect 600004 143624 600010 143676
rect 581270 143556 581276 143608
rect 581328 143596 581334 143608
rect 600038 143596 600044 143608
rect 581328 143568 600044 143596
rect 581328 143556 581334 143568
rect 600038 143556 600044 143568
rect 600096 143556 600102 143608
rect 581638 140904 581644 140956
rect 581696 140944 581702 140956
rect 599946 140944 599952 140956
rect 581696 140916 599952 140944
rect 581696 140904 581702 140916
rect 599946 140904 599952 140916
rect 600004 140904 600010 140956
rect 580994 140836 581000 140888
rect 581052 140876 581058 140888
rect 600038 140876 600044 140888
rect 581052 140848 600044 140876
rect 581052 140836 581058 140848
rect 600038 140836 600044 140848
rect 600096 140836 600102 140888
rect 581178 140768 581184 140820
rect 581236 140808 581242 140820
rect 599854 140808 599860 140820
rect 581236 140780 599860 140808
rect 581236 140768 581242 140780
rect 599854 140768 599860 140780
rect 599912 140768 599918 140820
rect 581086 138116 581092 138168
rect 581144 138156 581150 138168
rect 599946 138156 599952 138168
rect 581144 138128 599952 138156
rect 581144 138116 581150 138128
rect 599946 138116 599952 138128
rect 600004 138116 600010 138168
rect 579706 138048 579712 138100
rect 579764 138088 579770 138100
rect 600038 138088 600044 138100
rect 579764 138060 600044 138088
rect 579764 138048 579770 138060
rect 600038 138048 600044 138060
rect 600096 138048 600102 138100
rect 579890 137980 579896 138032
rect 579948 138020 579954 138032
rect 599854 138020 599860 138032
rect 579948 137992 599860 138020
rect 579948 137980 579954 137992
rect 599854 137980 599860 137992
rect 599912 137980 599918 138032
rect 580074 135328 580080 135380
rect 580132 135368 580138 135380
rect 599854 135368 599860 135380
rect 580132 135340 599860 135368
rect 580132 135328 580138 135340
rect 599854 135328 599860 135340
rect 599912 135328 599918 135380
rect 580166 135260 580172 135312
rect 580224 135300 580230 135312
rect 599946 135300 599952 135312
rect 580224 135272 599952 135300
rect 580224 135260 580230 135272
rect 599946 135260 599952 135272
rect 600004 135260 600010 135312
rect 670142 132880 670148 132932
rect 670200 132920 670206 132932
rect 676214 132920 676220 132932
rect 670200 132892 676220 132920
rect 670200 132880 670206 132892
rect 676214 132880 676220 132892
rect 676272 132880 676278 132932
rect 670050 132744 670056 132796
rect 670108 132784 670114 132796
rect 676122 132784 676128 132796
rect 670108 132756 676128 132784
rect 670108 132744 670114 132756
rect 676122 132744 676128 132756
rect 676180 132744 676186 132796
rect 580902 132608 580908 132660
rect 580960 132648 580966 132660
rect 599946 132648 599952 132660
rect 580960 132620 599952 132648
rect 580960 132608 580966 132620
rect 599946 132608 599952 132620
rect 600004 132608 600010 132660
rect 669958 132608 669964 132660
rect 670016 132648 670022 132660
rect 676030 132648 676036 132660
rect 670016 132620 676036 132648
rect 670016 132608 670022 132620
rect 676030 132608 676036 132620
rect 676088 132608 676094 132660
rect 580258 132540 580264 132592
rect 580316 132580 580322 132592
rect 599854 132580 599860 132592
rect 580316 132552 599860 132580
rect 580316 132540 580322 132552
rect 599854 132540 599860 132552
rect 599912 132540 599918 132592
rect 579982 132472 579988 132524
rect 580040 132512 580046 132524
rect 600038 132512 600044 132524
rect 580040 132484 600044 132512
rect 580040 132472 580046 132484
rect 600038 132472 600044 132484
rect 600096 132472 600102 132524
rect 675202 132404 675208 132456
rect 675260 132444 675266 132456
rect 676030 132444 676036 132456
rect 675260 132416 676036 132444
rect 675260 132404 675266 132416
rect 676030 132404 676036 132416
rect 676088 132404 676094 132456
rect 672166 131656 672172 131708
rect 672224 131696 672230 131708
rect 673270 131696 673276 131708
rect 672224 131668 673276 131696
rect 672224 131656 672230 131668
rect 673270 131656 673276 131668
rect 673328 131696 673334 131708
rect 676030 131696 676036 131708
rect 673328 131668 676036 131696
rect 673328 131656 673334 131668
rect 676030 131656 676036 131668
rect 676088 131656 676094 131708
rect 673362 131452 673368 131504
rect 673420 131492 673426 131504
rect 676214 131492 676220 131504
rect 673420 131464 676220 131492
rect 673420 131452 673426 131464
rect 676214 131452 676220 131464
rect 676272 131452 676278 131504
rect 672258 130840 672264 130892
rect 672316 130880 672322 130892
rect 676030 130880 676036 130892
rect 672316 130852 676036 130880
rect 672316 130840 672322 130852
rect 676030 130840 676036 130852
rect 676088 130840 676094 130892
rect 671890 130024 671896 130076
rect 671948 130064 671954 130076
rect 672074 130064 672080 130076
rect 671948 130036 672080 130064
rect 671948 130024 671954 130036
rect 672074 130024 672080 130036
rect 672132 130064 672138 130076
rect 676030 130064 676036 130076
rect 672132 130036 676036 130064
rect 672132 130024 672138 130036
rect 676030 130024 676036 130036
rect 676088 130024 676094 130076
rect 580350 129888 580356 129940
rect 580408 129928 580414 129940
rect 600038 129928 600044 129940
rect 580408 129900 600044 129928
rect 580408 129888 580414 129900
rect 600038 129888 600044 129900
rect 600096 129888 600102 129940
rect 580626 129820 580632 129872
rect 580684 129860 580690 129872
rect 599854 129860 599860 129872
rect 580684 129832 599860 129860
rect 580684 129820 580690 129832
rect 599854 129820 599860 129832
rect 599912 129820 599918 129872
rect 580442 129752 580448 129804
rect 580500 129792 580506 129804
rect 599946 129792 599952 129804
rect 580500 129764 599952 129792
rect 580500 129752 580506 129764
rect 599946 129752 599952 129764
rect 600004 129752 600010 129804
rect 672350 129412 672356 129464
rect 672408 129452 672414 129464
rect 673086 129452 673092 129464
rect 672408 129424 673092 129452
rect 672408 129412 672414 129424
rect 673086 129412 673092 129424
rect 673144 129452 673150 129464
rect 676214 129452 676220 129464
rect 673144 129424 676220 129452
rect 673144 129412 673150 129424
rect 676214 129412 676220 129424
rect 676272 129412 676278 129464
rect 674742 127712 674748 127764
rect 674800 127752 674806 127764
rect 676030 127752 676036 127764
rect 674800 127724 676036 127752
rect 674800 127712 674806 127724
rect 676030 127712 676036 127724
rect 676088 127712 676094 127764
rect 673546 127304 673552 127356
rect 673604 127344 673610 127356
rect 675938 127344 675944 127356
rect 673604 127316 675944 127344
rect 673604 127304 673610 127316
rect 675938 127304 675944 127316
rect 675996 127304 676002 127356
rect 580718 127032 580724 127084
rect 580776 127072 580782 127084
rect 599854 127072 599860 127084
rect 580776 127044 599860 127072
rect 580776 127032 580782 127044
rect 599854 127032 599860 127044
rect 599912 127032 599918 127084
rect 673822 127032 673828 127084
rect 673880 127072 673886 127084
rect 675938 127072 675944 127084
rect 673880 127044 675944 127072
rect 673880 127032 673886 127044
rect 675938 127032 675944 127044
rect 675996 127032 676002 127084
rect 580534 126964 580540 127016
rect 580592 127004 580598 127016
rect 599946 127004 599952 127016
rect 580592 126976 599952 127004
rect 580592 126964 580598 126976
rect 599946 126964 599952 126976
rect 600004 126964 600010 127016
rect 674834 126964 674840 127016
rect 674892 127004 674898 127016
rect 676030 127004 676036 127016
rect 674892 126976 676036 127004
rect 674892 126964 674898 126976
rect 676030 126964 676036 126976
rect 676088 126964 676094 127016
rect 674650 126488 674656 126540
rect 674708 126528 674714 126540
rect 676030 126528 676036 126540
rect 674708 126500 676036 126528
rect 674708 126488 674714 126500
rect 676030 126488 676036 126500
rect 676088 126488 676094 126540
rect 673638 124856 673644 124908
rect 673696 124896 673702 124908
rect 675938 124896 675944 124908
rect 673696 124868 675944 124896
rect 673696 124856 673702 124868
rect 675938 124856 675944 124868
rect 675996 124856 676002 124908
rect 673730 124448 673736 124500
rect 673788 124488 673794 124500
rect 675938 124488 675944 124500
rect 673788 124460 675944 124488
rect 673788 124448 673794 124460
rect 675938 124448 675944 124460
rect 675996 124448 676002 124500
rect 582282 124312 582288 124364
rect 582340 124352 582346 124364
rect 599854 124352 599860 124364
rect 582340 124324 599860 124352
rect 582340 124312 582346 124324
rect 599854 124312 599860 124324
rect 599912 124312 599918 124364
rect 581822 124244 581828 124296
rect 581880 124284 581886 124296
rect 599762 124284 599768 124296
rect 581880 124256 599768 124284
rect 581880 124244 581886 124256
rect 599762 124244 599768 124256
rect 599820 124244 599826 124296
rect 674926 124244 674932 124296
rect 674984 124284 674990 124296
rect 675938 124284 675944 124296
rect 674984 124256 675944 124284
rect 674984 124244 674990 124256
rect 675938 124244 675944 124256
rect 675996 124244 676002 124296
rect 580810 124176 580816 124228
rect 580868 124216 580874 124228
rect 599946 124216 599952 124228
rect 580868 124188 599952 124216
rect 580868 124176 580874 124188
rect 599946 124176 599952 124188
rect 600004 124176 600010 124228
rect 675018 124176 675024 124228
rect 675076 124216 675082 124228
rect 676030 124216 676036 124228
rect 675076 124188 676036 124216
rect 675076 124176 675082 124188
rect 676030 124176 676036 124188
rect 676088 124176 676094 124228
rect 582190 121592 582196 121644
rect 582248 121632 582254 121644
rect 599946 121632 599952 121644
rect 582248 121604 599952 121632
rect 582248 121592 582254 121604
rect 599946 121592 599952 121604
rect 600004 121592 600010 121644
rect 672442 121592 672448 121644
rect 672500 121632 672506 121644
rect 676214 121632 676220 121644
rect 672500 121604 676220 121632
rect 672500 121592 672506 121604
rect 676214 121592 676220 121604
rect 676272 121592 676278 121644
rect 582006 121524 582012 121576
rect 582064 121564 582070 121576
rect 599854 121564 599860 121576
rect 582064 121536 599860 121564
rect 582064 121524 582070 121536
rect 599854 121524 599860 121536
rect 599912 121524 599918 121576
rect 674282 121524 674288 121576
rect 674340 121564 674346 121576
rect 675938 121564 675944 121576
rect 674340 121536 675944 121564
rect 674340 121524 674346 121536
rect 675938 121524 675944 121536
rect 675996 121524 676002 121576
rect 582098 121456 582104 121508
rect 582156 121496 582162 121508
rect 600038 121496 600044 121508
rect 582156 121468 600044 121496
rect 582156 121456 582162 121468
rect 600038 121456 600044 121468
rect 600096 121456 600102 121508
rect 674466 121456 674472 121508
rect 674524 121496 674530 121508
rect 676030 121496 676036 121508
rect 674524 121468 676036 121496
rect 674524 121456 674530 121468
rect 676030 121456 676036 121468
rect 676088 121456 676094 121508
rect 674926 121388 674932 121440
rect 674984 121388 674990 121440
rect 674742 121320 674748 121372
rect 674800 121320 674806 121372
rect 674760 121168 674788 121320
rect 674944 121168 674972 121388
rect 674742 121116 674748 121168
rect 674800 121116 674806 121168
rect 674926 121116 674932 121168
rect 674984 121116 674990 121168
rect 583662 118804 583668 118856
rect 583720 118844 583726 118856
rect 599946 118844 599952 118856
rect 583720 118816 599952 118844
rect 583720 118804 583726 118816
rect 599946 118804 599952 118816
rect 600004 118804 600010 118856
rect 581914 118736 581920 118788
rect 581972 118776 581978 118788
rect 600038 118776 600044 118788
rect 581972 118748 600044 118776
rect 581972 118736 581978 118748
rect 600038 118736 600044 118748
rect 600096 118736 600102 118788
rect 581454 118668 581460 118720
rect 581512 118708 581518 118720
rect 599854 118708 599860 118720
rect 581512 118680 599860 118708
rect 581512 118668 581518 118680
rect 599854 118668 599860 118680
rect 599912 118668 599918 118720
rect 581730 116016 581736 116068
rect 581788 116056 581794 116068
rect 599946 116056 599952 116068
rect 581788 116028 599952 116056
rect 581788 116016 581794 116028
rect 599946 116016 599952 116028
rect 600004 116016 600010 116068
rect 581270 115948 581276 116000
rect 581328 115988 581334 116000
rect 600038 115988 600044 116000
rect 581328 115960 600044 115988
rect 581328 115948 581334 115960
rect 600038 115948 600044 115960
rect 600096 115948 600102 116000
rect 666738 115880 666744 115932
rect 666796 115920 666802 115932
rect 675386 115920 675392 115932
rect 666796 115892 675392 115920
rect 666796 115880 666802 115892
rect 675386 115880 675392 115892
rect 675444 115880 675450 115932
rect 675018 114996 675024 115048
rect 675076 115036 675082 115048
rect 675294 115036 675300 115048
rect 675076 115008 675300 115036
rect 675076 114996 675082 115008
rect 675294 114996 675300 115008
rect 675352 114996 675358 115048
rect 674742 114316 674748 114368
rect 674800 114356 674806 114368
rect 675294 114356 675300 114368
rect 674800 114328 675300 114356
rect 674800 114316 674806 114328
rect 675294 114316 675300 114328
rect 675352 114316 675358 114368
rect 674834 113704 674840 113756
rect 674892 113744 674898 113756
rect 675294 113744 675300 113756
rect 674892 113716 675300 113744
rect 674892 113704 674898 113716
rect 675294 113704 675300 113716
rect 675352 113704 675358 113756
rect 581638 113228 581644 113280
rect 581696 113268 581702 113280
rect 599946 113268 599952 113280
rect 581696 113240 599952 113268
rect 581696 113228 581702 113240
rect 599946 113228 599952 113240
rect 600004 113228 600010 113280
rect 581362 113160 581368 113212
rect 581420 113200 581426 113212
rect 599854 113200 599860 113212
rect 581420 113172 599860 113200
rect 581420 113160 581426 113172
rect 599854 113160 599860 113172
rect 599912 113160 599918 113212
rect 581546 110508 581552 110560
rect 581604 110548 581610 110560
rect 599854 110548 599860 110560
rect 581604 110520 599860 110548
rect 581604 110508 581610 110520
rect 599854 110508 599860 110520
rect 599912 110508 599918 110560
rect 580994 110440 581000 110492
rect 581052 110480 581058 110492
rect 599946 110480 599952 110492
rect 581052 110452 599952 110480
rect 581052 110440 581058 110452
rect 599946 110440 599952 110452
rect 600004 110440 600010 110492
rect 673730 110032 673736 110084
rect 673788 110072 673794 110084
rect 675110 110072 675116 110084
rect 673788 110044 675116 110072
rect 673788 110032 673794 110044
rect 675110 110032 675116 110044
rect 675168 110032 675174 110084
rect 673822 108196 673828 108248
rect 673880 108236 673886 108248
rect 675386 108236 675392 108248
rect 673880 108208 675392 108236
rect 673880 108196 673886 108208
rect 675386 108196 675392 108208
rect 675444 108196 675450 108248
rect 581178 107652 581184 107704
rect 581236 107692 581242 107704
rect 599302 107692 599308 107704
rect 581236 107664 599308 107692
rect 581236 107652 581242 107664
rect 599302 107652 599308 107664
rect 599360 107652 599366 107704
rect 674466 107516 674472 107568
rect 674524 107556 674530 107568
rect 675386 107556 675392 107568
rect 674524 107528 675392 107556
rect 674524 107516 674530 107528
rect 675386 107516 675392 107528
rect 675444 107516 675450 107568
rect 674282 106360 674288 106412
rect 674340 106400 674346 106412
rect 675386 106400 675392 106412
rect 674340 106372 675392 106400
rect 674340 106360 674346 106372
rect 675386 106360 675392 106372
rect 675444 106360 675450 106412
rect 673638 106292 673644 106344
rect 673696 106332 673702 106344
rect 675110 106332 675116 106344
rect 673696 106304 675116 106332
rect 673696 106292 673702 106304
rect 675110 106292 675116 106304
rect 675168 106292 675174 106344
rect 581086 104864 581092 104916
rect 581144 104904 581150 104916
rect 599946 104904 599952 104916
rect 581144 104876 599952 104904
rect 581144 104864 581150 104876
rect 599946 104864 599952 104876
rect 600004 104864 600010 104916
rect 673546 104524 673552 104576
rect 673604 104564 673610 104576
rect 675110 104564 675116 104576
rect 673604 104536 675116 104564
rect 673604 104524 673610 104536
rect 675110 104524 675116 104536
rect 675168 104524 675174 104576
rect 657722 99764 657728 99816
rect 657780 99804 657786 99816
rect 660896 99804 660902 99816
rect 657780 99776 660902 99804
rect 657780 99764 657786 99776
rect 660896 99764 660902 99776
rect 660954 99764 660960 99816
rect 580902 99356 580908 99408
rect 580960 99396 580966 99408
rect 599946 99396 599952 99408
rect 580960 99368 599952 99396
rect 580960 99356 580966 99368
rect 599946 99356 599952 99368
rect 600004 99356 600010 99408
rect 633066 96568 633072 96620
rect 633124 96608 633130 96620
rect 635274 96608 635280 96620
rect 633124 96580 635280 96608
rect 633124 96568 633130 96580
rect 635274 96568 635280 96580
rect 635332 96568 635338 96620
rect 636286 96568 636292 96620
rect 636344 96608 636350 96620
rect 640978 96608 640984 96620
rect 636344 96580 640984 96608
rect 636344 96568 636350 96580
rect 640978 96568 640984 96580
rect 641036 96568 641042 96620
rect 655974 96568 655980 96620
rect 656032 96608 656038 96620
rect 659562 96608 659568 96620
rect 656032 96580 659568 96608
rect 656032 96568 656038 96580
rect 659562 96568 659568 96580
rect 659620 96568 659626 96620
rect 661862 96568 661868 96620
rect 661920 96608 661926 96620
rect 663058 96608 663064 96620
rect 661920 96580 663064 96608
rect 661920 96568 661926 96580
rect 663058 96568 663064 96580
rect 663116 96568 663122 96620
rect 633802 96500 633808 96552
rect 633860 96540 633866 96552
rect 636378 96540 636384 96552
rect 633860 96512 636384 96540
rect 633860 96500 633866 96512
rect 636378 96500 636384 96512
rect 636436 96500 636442 96552
rect 637022 96500 637028 96552
rect 637080 96540 637086 96552
rect 642358 96540 642364 96552
rect 637080 96512 642364 96540
rect 637080 96500 637086 96512
rect 642358 96500 642364 96512
rect 642416 96500 642422 96552
rect 654686 96500 654692 96552
rect 654744 96540 654750 96552
rect 658274 96540 658280 96552
rect 654744 96512 658280 96540
rect 654744 96500 654750 96512
rect 658274 96500 658280 96512
rect 658332 96500 658338 96552
rect 659102 96500 659108 96552
rect 659160 96540 659166 96552
rect 662506 96540 662512 96552
rect 659160 96512 662512 96540
rect 659160 96500 659166 96512
rect 662506 96500 662512 96512
rect 662564 96500 662570 96552
rect 634446 96432 634452 96484
rect 634504 96472 634510 96484
rect 637574 96472 637580 96484
rect 634504 96444 637580 96472
rect 634504 96432 634510 96444
rect 637574 96432 637580 96444
rect 637632 96432 637638 96484
rect 635734 96364 635740 96416
rect 635792 96404 635798 96416
rect 639874 96404 639880 96416
rect 635792 96376 639880 96404
rect 635792 96364 635798 96376
rect 639874 96364 639880 96376
rect 639932 96364 639938 96416
rect 647510 96296 647516 96348
rect 647568 96336 647574 96348
rect 653950 96336 653956 96348
rect 647568 96308 653956 96336
rect 647568 96296 647574 96308
rect 653950 96296 653956 96308
rect 654008 96296 654014 96348
rect 631134 96024 631140 96076
rect 631192 96064 631198 96076
rect 632100 96064 632106 96076
rect 631192 96036 632106 96064
rect 631192 96024 631198 96036
rect 632100 96024 632106 96036
rect 632158 96024 632164 96076
rect 632422 96024 632428 96076
rect 632480 96064 632486 96076
rect 634400 96064 634406 96076
rect 632480 96036 634406 96064
rect 632480 96024 632486 96036
rect 634400 96024 634406 96036
rect 634458 96024 634464 96076
rect 635090 96024 635096 96076
rect 635148 96064 635154 96076
rect 639000 96064 639006 96076
rect 635148 96036 639006 96064
rect 635148 96024 635154 96036
rect 639000 96024 639006 96036
rect 639058 96024 639064 96076
rect 631778 95888 631784 95940
rect 631836 95928 631842 95940
rect 632974 95928 632980 95940
rect 631836 95900 632980 95928
rect 631836 95888 631842 95900
rect 632974 95888 632980 95900
rect 633032 95888 633038 95940
rect 640058 95888 640064 95940
rect 640116 95928 640122 95940
rect 646038 95928 646044 95940
rect 640116 95900 646044 95928
rect 640116 95888 640122 95900
rect 646038 95888 646044 95900
rect 646096 95888 646102 95940
rect 638862 95820 638868 95872
rect 638920 95860 638926 95872
rect 645854 95860 645860 95872
rect 638920 95832 645860 95860
rect 638920 95820 638926 95832
rect 645854 95820 645860 95832
rect 645912 95820 645918 95872
rect 646130 95820 646136 95872
rect 646188 95860 646194 95872
rect 663518 95860 663524 95872
rect 646188 95832 663524 95860
rect 646188 95820 646194 95832
rect 663518 95820 663524 95832
rect 663576 95820 663582 95872
rect 614758 95752 614764 95804
rect 614816 95792 614822 95804
rect 614816 95764 632054 95792
rect 614816 95752 614822 95764
rect 616138 95684 616144 95736
rect 616196 95724 616202 95736
rect 622486 95724 622492 95736
rect 616196 95696 622492 95724
rect 616196 95684 616202 95696
rect 622486 95684 622492 95696
rect 622544 95684 622550 95736
rect 621290 95616 621296 95668
rect 621348 95656 621354 95668
rect 623314 95656 623320 95668
rect 621348 95628 623320 95656
rect 621348 95616 621354 95628
rect 623314 95616 623320 95628
rect 623372 95616 623378 95668
rect 604454 95548 604460 95600
rect 604512 95588 604518 95600
rect 606386 95588 606392 95600
rect 604512 95560 606392 95588
rect 604512 95548 604518 95560
rect 606386 95548 606392 95560
rect 606444 95548 606450 95600
rect 607490 95548 607496 95600
rect 607548 95588 607554 95600
rect 608962 95588 608968 95600
rect 607548 95560 608968 95588
rect 607548 95548 607554 95560
rect 608962 95548 608968 95560
rect 609020 95548 609026 95600
rect 610250 95548 610256 95600
rect 610308 95588 610314 95600
rect 611538 95588 611544 95600
rect 610308 95560 611544 95588
rect 610308 95548 610314 95560
rect 611538 95548 611544 95560
rect 611596 95548 611602 95600
rect 618254 95548 618260 95600
rect 618312 95588 618318 95600
rect 620094 95588 620100 95600
rect 618312 95560 620100 95588
rect 618312 95548 618318 95560
rect 620094 95548 620100 95560
rect 620152 95548 620158 95600
rect 621474 95548 621480 95600
rect 621532 95588 621538 95600
rect 622670 95588 622676 95600
rect 621532 95560 622676 95588
rect 621532 95548 621538 95560
rect 622670 95548 622676 95560
rect 622728 95548 622734 95600
rect 621198 95480 621204 95532
rect 621256 95520 621262 95532
rect 622026 95520 622032 95532
rect 621256 95492 622032 95520
rect 621256 95480 621262 95492
rect 622026 95480 622032 95492
rect 622084 95480 622090 95532
rect 620002 95412 620008 95464
rect 620060 95452 620066 95464
rect 623406 95452 623412 95464
rect 620060 95424 623412 95452
rect 620060 95412 620066 95424
rect 623406 95412 623412 95424
rect 623464 95412 623470 95464
rect 591942 95344 591948 95396
rect 592000 95384 592006 95396
rect 610342 95384 610348 95396
rect 592000 95356 610348 95384
rect 592000 95344 592006 95356
rect 610342 95344 610348 95356
rect 610400 95344 610406 95396
rect 617426 95344 617432 95396
rect 617484 95384 617490 95396
rect 622118 95384 622124 95396
rect 617484 95356 622124 95384
rect 617484 95344 617490 95356
rect 622118 95344 622124 95356
rect 622176 95344 622182 95396
rect 589182 95276 589188 95328
rect 589240 95316 589246 95328
rect 612182 95316 612188 95328
rect 589240 95288 612188 95316
rect 589240 95276 589246 95288
rect 612182 95276 612188 95288
rect 612240 95276 612246 95328
rect 575658 95208 575664 95260
rect 575716 95248 575722 95260
rect 607674 95248 607680 95260
rect 575716 95220 607680 95248
rect 575716 95208 575722 95220
rect 607674 95208 607680 95220
rect 607732 95208 607738 95260
rect 632026 95180 632054 95764
rect 639598 95752 639604 95804
rect 639656 95792 639662 95804
rect 639656 95764 646084 95792
rect 639656 95752 639662 95764
rect 637482 95684 637488 95736
rect 637540 95724 637546 95736
rect 640518 95724 640524 95736
rect 637540 95696 640524 95724
rect 637540 95684 637546 95696
rect 640518 95684 640524 95696
rect 640576 95684 640582 95736
rect 640886 95684 640892 95736
rect 640944 95724 640950 95736
rect 645946 95724 645952 95736
rect 640944 95696 645952 95724
rect 640944 95684 640950 95696
rect 645946 95684 645952 95696
rect 646004 95684 646010 95736
rect 641622 95616 641628 95668
rect 641680 95656 641686 95668
rect 642818 95656 642824 95668
rect 641680 95628 642824 95656
rect 641680 95616 641686 95628
rect 642818 95616 642824 95628
rect 642876 95616 642882 95668
rect 638310 95548 638316 95600
rect 638368 95548 638374 95600
rect 642266 95548 642272 95600
rect 642324 95588 642330 95600
rect 642910 95588 642916 95600
rect 642324 95560 642916 95588
rect 642324 95548 642330 95560
rect 642910 95548 642916 95560
rect 642968 95548 642974 95600
rect 638328 95520 638356 95548
rect 642726 95520 642732 95532
rect 638328 95492 642732 95520
rect 642726 95480 642732 95492
rect 642784 95480 642790 95532
rect 646056 95464 646084 95764
rect 652018 95752 652024 95804
rect 652076 95792 652082 95804
rect 661954 95792 661960 95804
rect 652076 95764 661960 95792
rect 652076 95752 652082 95764
rect 661954 95752 661960 95764
rect 662012 95752 662018 95804
rect 652662 95616 652668 95668
rect 652720 95656 652726 95668
rect 663886 95656 663892 95668
rect 652720 95628 663892 95656
rect 652720 95616 652726 95628
rect 663886 95616 663892 95628
rect 663944 95616 663950 95668
rect 651834 95548 651840 95600
rect 651892 95588 651898 95600
rect 653398 95588 653404 95600
rect 651892 95560 653404 95588
rect 651892 95548 651898 95560
rect 653398 95548 653404 95560
rect 653456 95548 653462 95600
rect 656986 95548 656992 95600
rect 657044 95588 657050 95600
rect 659194 95588 659200 95600
rect 657044 95560 659200 95588
rect 657044 95548 657050 95560
rect 659194 95548 659200 95560
rect 659252 95548 659258 95600
rect 660574 95480 660580 95532
rect 660632 95520 660638 95532
rect 661402 95520 661408 95532
rect 660632 95492 661408 95520
rect 660632 95480 660638 95492
rect 661402 95480 661408 95492
rect 661460 95480 661466 95532
rect 646038 95412 646044 95464
rect 646096 95412 646102 95464
rect 646774 95412 646780 95464
rect 646832 95452 646838 95464
rect 646832 95424 651374 95452
rect 646832 95412 646838 95424
rect 648614 95344 648620 95396
rect 648672 95384 648678 95396
rect 650730 95384 650736 95396
rect 648672 95356 650736 95384
rect 648672 95344 648678 95356
rect 650730 95344 650736 95356
rect 650788 95344 650794 95396
rect 651346 95384 651374 95424
rect 663426 95384 663432 95396
rect 651346 95356 663432 95384
rect 663426 95344 663432 95356
rect 663484 95344 663490 95396
rect 657078 95208 657084 95260
rect 657136 95248 657142 95260
rect 657906 95248 657912 95260
rect 657136 95220 657912 95248
rect 657136 95208 657142 95220
rect 657906 95208 657912 95220
rect 657964 95208 657970 95260
rect 665174 95180 665180 95192
rect 632026 95152 665180 95180
rect 665174 95140 665180 95152
rect 665232 95140 665238 95192
rect 619358 95072 619364 95124
rect 619416 95112 619422 95124
rect 623498 95112 623504 95124
rect 619416 95084 623504 95112
rect 619416 95072 619422 95084
rect 623498 95072 623504 95084
rect 623556 95072 623562 95124
rect 643462 95072 643468 95124
rect 643520 95112 643526 95124
rect 644842 95112 644848 95124
rect 643520 95084 644848 95112
rect 643520 95072 643526 95084
rect 644842 95072 644848 95084
rect 644900 95072 644906 95124
rect 648798 94936 648804 94988
rect 648856 94976 648862 94988
rect 650086 94976 650092 94988
rect 648856 94948 650092 94976
rect 648856 94936 648862 94948
rect 650086 94936 650092 94948
rect 650144 94936 650150 94988
rect 616782 94868 616788 94920
rect 616840 94908 616846 94920
rect 623222 94908 623228 94920
rect 616840 94880 623228 94908
rect 616840 94868 616846 94880
rect 623222 94868 623228 94880
rect 623280 94868 623286 94920
rect 648890 94800 648896 94852
rect 648948 94840 648954 94852
rect 649442 94840 649448 94852
rect 648948 94812 649448 94840
rect 648948 94800 648954 94812
rect 649442 94800 649448 94812
rect 649500 94800 649506 94852
rect 618714 94732 618720 94784
rect 618772 94772 618778 94784
rect 623314 94772 623320 94784
rect 618772 94744 623320 94772
rect 618772 94732 618778 94744
rect 623314 94732 623320 94744
rect 623372 94732 623378 94784
rect 646590 94732 646596 94784
rect 646648 94772 646654 94784
rect 648154 94772 648160 94784
rect 646648 94744 648160 94772
rect 646648 94732 646654 94744
rect 648154 94732 648160 94744
rect 648212 94732 648218 94784
rect 653306 94732 653312 94784
rect 653364 94772 653370 94784
rect 663794 94772 663800 94784
rect 653364 94744 663800 94772
rect 653364 94732 653370 94744
rect 663794 94732 663800 94744
rect 663852 94732 663858 94784
rect 656618 94664 656624 94716
rect 656676 94704 656682 94716
rect 663702 94704 663708 94716
rect 656676 94676 663708 94704
rect 656676 94664 656682 94676
rect 663702 94664 663708 94676
rect 663760 94664 663766 94716
rect 657262 94596 657268 94648
rect 657320 94636 657326 94648
rect 663610 94636 663616 94648
rect 657320 94608 663616 94636
rect 657320 94596 657326 94608
rect 663610 94596 663616 94608
rect 663668 94596 663674 94648
rect 656894 94528 656900 94580
rect 656952 94568 656958 94580
rect 658550 94568 658556 94580
rect 656952 94540 658556 94568
rect 656952 94528 656958 94540
rect 658550 94528 658556 94540
rect 658608 94528 658614 94580
rect 648062 94460 648068 94512
rect 648120 94500 648126 94512
rect 659838 94500 659844 94512
rect 648120 94472 659844 94500
rect 648120 94460 648126 94472
rect 659838 94460 659844 94472
rect 659896 94460 659902 94512
rect 660390 94460 660396 94512
rect 660448 94460 660454 94512
rect 643554 94188 643560 94240
rect 643612 94228 643618 94240
rect 660408 94228 660436 94460
rect 643612 94200 660436 94228
rect 643612 94188 643618 94200
rect 618070 94120 618076 94172
rect 618128 94160 618134 94172
rect 623130 94160 623136 94172
rect 618128 94132 623136 94160
rect 618128 94120 618134 94132
rect 623130 94120 623136 94132
rect 623188 94120 623194 94172
rect 644198 94052 644204 94104
rect 644256 94092 644262 94104
rect 654042 94092 654048 94104
rect 644256 94064 654048 94092
rect 644256 94052 644262 94064
rect 654042 94052 654048 94064
rect 654100 94052 654106 94104
rect 649350 93984 649356 94036
rect 649408 94024 649414 94036
rect 656894 94024 656900 94036
rect 649408 93996 656900 94024
rect 649408 93984 649414 93996
rect 656894 93984 656900 93996
rect 656952 93984 656958 94036
rect 607214 93848 607220 93900
rect 607272 93888 607278 93900
rect 612918 93888 612924 93900
rect 607272 93860 612924 93888
rect 607272 93848 607278 93860
rect 612918 93848 612924 93860
rect 612976 93848 612982 93900
rect 644750 93848 644756 93900
rect 644808 93888 644814 93900
rect 653122 93888 653128 93900
rect 644808 93860 653128 93888
rect 644808 93848 644814 93860
rect 653122 93848 653128 93860
rect 653180 93848 653186 93900
rect 613010 93644 613016 93696
rect 613068 93684 613074 93696
rect 614850 93684 614856 93696
rect 613068 93656 614856 93684
rect 613068 93644 613074 93656
rect 614850 93644 614856 93656
rect 614908 93644 614914 93696
rect 663242 91060 663248 91112
rect 663300 91100 663306 91112
rect 663886 91100 663892 91112
rect 663300 91072 663892 91100
rect 663300 91060 663306 91072
rect 663886 91060 663892 91072
rect 663944 91060 663950 91112
rect 657078 88816 657084 88868
rect 657136 88856 657142 88868
rect 657998 88856 658004 88868
rect 657136 88828 658004 88856
rect 657136 88816 657142 88828
rect 657998 88816 658004 88828
rect 658056 88816 658062 88868
rect 659470 88748 659476 88800
rect 659528 88788 659534 88800
rect 663150 88788 663156 88800
rect 659528 88760 663156 88788
rect 659528 88748 659534 88760
rect 663150 88748 663156 88760
rect 663208 88748 663214 88800
rect 648614 85484 648620 85536
rect 648672 85524 648678 85536
rect 657170 85524 657176 85536
rect 648672 85496 657176 85524
rect 648672 85484 648678 85496
rect 657170 85484 657176 85496
rect 657228 85484 657234 85536
rect 651834 85416 651840 85468
rect 651892 85456 651898 85468
rect 658826 85456 658832 85468
rect 651892 85428 658832 85456
rect 651892 85416 651898 85428
rect 658826 85416 658832 85428
rect 658884 85416 658890 85468
rect 648890 85348 648896 85400
rect 648948 85388 648954 85400
rect 660666 85388 660672 85400
rect 648948 85360 660672 85388
rect 648948 85348 648954 85360
rect 660666 85348 660672 85360
rect 660724 85348 660730 85400
rect 648798 85280 648804 85332
rect 648856 85320 648862 85332
rect 657722 85320 657728 85332
rect 648856 85292 657728 85320
rect 648856 85280 648862 85292
rect 657722 85280 657728 85292
rect 657780 85280 657786 85332
rect 643462 85212 643468 85264
rect 643520 85252 643526 85264
rect 660114 85252 660120 85264
rect 643520 85224 660120 85252
rect 643520 85212 643526 85224
rect 660114 85212 660120 85224
rect 660172 85212 660178 85264
rect 646590 85144 646596 85196
rect 646648 85184 646654 85196
rect 661402 85184 661408 85196
rect 646648 85156 661408 85184
rect 646648 85144 646654 85156
rect 661402 85144 661408 85156
rect 661460 85144 661466 85196
rect 583754 84600 583760 84652
rect 583812 84640 583818 84652
rect 600314 84640 600320 84652
rect 583812 84612 600320 84640
rect 583812 84600 583818 84612
rect 600314 84600 600320 84612
rect 600372 84600 600378 84652
rect 582190 84532 582196 84584
rect 582248 84572 582254 84584
rect 600406 84572 600412 84584
rect 582248 84544 600412 84572
rect 582248 84532 582254 84544
rect 600406 84532 600412 84544
rect 600464 84532 600470 84584
rect 582282 84464 582288 84516
rect 582340 84504 582346 84516
rect 600682 84504 600688 84516
rect 582340 84476 600688 84504
rect 582340 84464 582346 84476
rect 600682 84464 600688 84476
rect 600740 84464 600746 84516
rect 581822 84396 581828 84448
rect 581880 84436 581886 84448
rect 600498 84436 600504 84448
rect 581880 84408 600504 84436
rect 581880 84396 581886 84408
rect 600498 84396 600504 84408
rect 600556 84396 600562 84448
rect 582006 84328 582012 84380
rect 582064 84368 582070 84380
rect 600774 84368 600780 84380
rect 582064 84340 600780 84368
rect 582064 84328 582070 84340
rect 600774 84328 600780 84340
rect 600832 84328 600838 84380
rect 582098 84260 582104 84312
rect 582156 84300 582162 84312
rect 600866 84300 600872 84312
rect 582156 84272 600872 84300
rect 582156 84260 582162 84272
rect 600866 84260 600872 84272
rect 600924 84260 600930 84312
rect 580718 84192 580724 84244
rect 580776 84232 580782 84244
rect 600222 84232 600228 84244
rect 580776 84204 600228 84232
rect 580776 84192 580782 84204
rect 600222 84192 600228 84204
rect 600280 84192 600286 84244
rect 580810 84124 580816 84176
rect 580868 84164 580874 84176
rect 600590 84164 600596 84176
rect 580868 84136 600596 84164
rect 580868 84124 580874 84136
rect 600590 84124 600596 84136
rect 600648 84124 600654 84176
rect 596910 83104 596916 83156
rect 596968 83144 596974 83156
rect 607214 83144 607220 83156
rect 596968 83116 607220 83144
rect 596968 83104 596974 83116
rect 607214 83104 607220 83116
rect 607272 83104 607278 83156
rect 597462 82832 597468 82884
rect 597520 82872 597526 82884
rect 604454 82872 604460 82884
rect 597520 82844 604460 82872
rect 597520 82832 597526 82844
rect 604454 82832 604460 82844
rect 604512 82832 604518 82884
rect 579614 82628 579620 82680
rect 579672 82668 579678 82680
rect 583662 82668 583668 82680
rect 579672 82640 583668 82668
rect 579672 82628 579678 82640
rect 583662 82628 583668 82640
rect 583720 82628 583726 82680
rect 600222 80112 600228 80164
rect 600280 80152 600286 80164
rect 612826 80152 612832 80164
rect 600280 80124 612832 80152
rect 600280 80112 600286 80124
rect 612826 80112 612832 80124
rect 612884 80112 612890 80164
rect 575842 78616 575848 78668
rect 575900 78656 575906 78668
rect 596910 78656 596916 78668
rect 575900 78628 596916 78656
rect 575900 78616 575906 78628
rect 596910 78616 596916 78628
rect 596968 78616 596974 78668
rect 575750 74944 575756 74996
rect 575808 74984 575814 74996
rect 589182 74984 589188 74996
rect 575808 74956 589188 74984
rect 575808 74944 575814 74956
rect 589182 74944 589188 74956
rect 589240 74944 589246 74996
rect 583662 73108 583668 73160
rect 583720 73148 583726 73160
rect 610158 73148 610164 73160
rect 583720 73120 610164 73148
rect 583720 73108 583726 73120
rect 610158 73108 610164 73120
rect 610216 73108 610222 73160
rect 586422 72632 586428 72684
rect 586480 72672 586486 72684
rect 591942 72672 591948 72684
rect 586480 72644 591948 72672
rect 586480 72632 586486 72644
rect 591942 72632 591948 72644
rect 592000 72632 592006 72684
rect 594702 66240 594708 66292
rect 594760 66280 594766 66292
rect 600222 66280 600228 66292
rect 594760 66252 600228 66280
rect 594760 66240 594766 66252
rect 600222 66240 600228 66252
rect 600280 66240 600286 66292
rect 602982 66240 602988 66292
rect 603040 66280 603046 66292
rect 610342 66280 610348 66292
rect 603040 66252 610348 66280
rect 603040 66240 603046 66252
rect 610342 66240 610348 66252
rect 610400 66240 610406 66292
rect 579614 66172 579620 66224
rect 579672 66212 579678 66224
rect 583754 66212 583760 66224
rect 579672 66184 583760 66212
rect 579672 66172 579678 66184
rect 583754 66172 583760 66184
rect 583812 66172 583818 66224
rect 587894 62296 587900 62348
rect 587952 62336 587958 62348
rect 597462 62336 597468 62348
rect 587952 62308 597468 62336
rect 587952 62296 587958 62308
rect 597462 62296 597468 62308
rect 597520 62296 597526 62348
rect 581638 53184 581644 53236
rect 581696 53224 581702 53236
rect 587894 53224 587900 53236
rect 581696 53196 587900 53224
rect 581696 53184 581702 53196
rect 587894 53184 587900 53196
rect 587952 53184 587958 53236
rect 145374 52436 145380 52488
rect 145432 52476 145438 52488
rect 198642 52476 198648 52488
rect 145432 52448 198648 52476
rect 145432 52436 145438 52448
rect 198642 52436 198648 52448
rect 198700 52436 198706 52488
rect 346854 52368 346860 52420
rect 346912 52408 346918 52420
rect 642910 52408 642916 52420
rect 346912 52380 642916 52408
rect 346912 52368 346918 52380
rect 642910 52368 642916 52380
rect 642968 52368 642974 52420
rect 52086 51076 52092 51128
rect 52144 51116 52150 51128
rect 213822 51116 213828 51128
rect 52144 51088 213828 51116
rect 52144 51076 52150 51088
rect 213822 51076 213828 51088
rect 213880 51116 213886 51128
rect 346486 51116 346492 51128
rect 213880 51088 346492 51116
rect 213880 51076 213886 51088
rect 346486 51076 346492 51088
rect 346544 51076 346550 51128
rect 198642 51008 198648 51060
rect 198700 51048 198706 51060
rect 207014 51048 207020 51060
rect 198700 51020 207020 51048
rect 198700 51008 198706 51020
rect 207014 51008 207020 51020
rect 207072 51048 207078 51060
rect 631870 51048 631876 51060
rect 207072 51020 631876 51048
rect 207072 51008 207078 51020
rect 631870 51008 631876 51020
rect 631928 51008 631934 51060
rect 478138 48424 478144 48476
rect 478196 48464 478202 48476
rect 526162 48464 526168 48476
rect 478196 48436 526168 48464
rect 478196 48424 478202 48436
rect 526162 48424 526168 48436
rect 526220 48424 526226 48476
rect 412634 48356 412640 48408
rect 412692 48396 412698 48408
rect 506382 48396 506388 48408
rect 412692 48368 506388 48396
rect 412692 48356 412698 48368
rect 506382 48356 506388 48368
rect 506440 48356 506446 48408
rect 571794 48356 571800 48408
rect 571852 48396 571858 48408
rect 581638 48396 581644 48408
rect 571852 48368 581644 48396
rect 571852 48356 571858 48368
rect 581638 48356 581644 48368
rect 581696 48356 581702 48408
rect 150342 48288 150348 48340
rect 150400 48328 150406 48340
rect 218054 48328 218060 48340
rect 150400 48300 218060 48328
rect 150400 48288 150406 48300
rect 218054 48288 218060 48300
rect 218112 48288 218118 48340
rect 281442 48288 281448 48340
rect 281500 48328 281506 48340
rect 502242 48328 502248 48340
rect 281500 48300 502248 48328
rect 281500 48288 281506 48300
rect 502242 48288 502248 48300
rect 502300 48288 502306 48340
rect 549254 48288 549260 48340
rect 549312 48328 549318 48340
rect 594702 48328 594708 48340
rect 549312 48300 594708 48328
rect 549312 48288 549318 48300
rect 594702 48288 594708 48300
rect 594760 48288 594766 48340
rect 568574 47200 568580 47252
rect 568632 47240 568638 47252
rect 575750 47240 575756 47252
rect 568632 47212 575756 47240
rect 568632 47200 568638 47212
rect 575750 47200 575756 47212
rect 575808 47200 575814 47252
rect 52270 47064 52276 47116
rect 52328 47104 52334 47116
rect 150342 47104 150348 47116
rect 52328 47076 150348 47104
rect 52328 47064 52334 47076
rect 150342 47064 150348 47076
rect 150400 47064 150406 47116
rect 577958 47064 577964 47116
rect 578016 47104 578022 47116
rect 583662 47104 583668 47116
rect 578016 47076 583668 47104
rect 578016 47064 578022 47076
rect 583662 47064 583668 47076
rect 583720 47064 583726 47116
rect 218054 46860 218060 46912
rect 218112 46900 218118 46912
rect 642634 46900 642640 46912
rect 218112 46872 642640 46900
rect 218112 46860 218118 46872
rect 642634 46860 642640 46872
rect 642692 46860 642698 46912
rect 460658 45976 460664 46028
rect 460716 46016 460722 46028
rect 610250 46016 610256 46028
rect 460716 45988 610256 46016
rect 460716 45976 460722 45988
rect 610250 45976 610256 45988
rect 610308 45976 610314 46028
rect 367094 45908 367100 45960
rect 367152 45948 367158 45960
rect 607306 45948 607312 45960
rect 367152 45920 607312 45948
rect 367152 45908 367158 45920
rect 607306 45908 607312 45920
rect 607364 45908 607370 45960
rect 311894 45840 311900 45892
rect 311952 45880 311958 45892
rect 607582 45880 607588 45892
rect 311952 45852 607588 45880
rect 311952 45840 311958 45852
rect 607582 45840 607588 45852
rect 607640 45840 607646 45892
rect 230934 45772 230940 45824
rect 230992 45812 230998 45824
rect 613010 45812 613016 45824
rect 230992 45784 613016 45812
rect 230992 45772 230998 45784
rect 613010 45772 613016 45784
rect 613068 45772 613074 45824
rect 85114 45704 85120 45756
rect 85172 45744 85178 45756
rect 475562 45744 475568 45756
rect 85172 45716 475568 45744
rect 85172 45704 85178 45716
rect 475562 45704 475568 45716
rect 475620 45704 475626 45756
rect 230382 45636 230388 45688
rect 230440 45676 230446 45688
rect 621382 45676 621388 45688
rect 230440 45648 621388 45676
rect 230440 45636 230446 45648
rect 621382 45636 621388 45648
rect 621440 45636 621446 45688
rect 233142 45568 233148 45620
rect 233200 45608 233206 45620
rect 642818 45608 642824 45620
rect 233200 45580 642824 45608
rect 233200 45568 233206 45580
rect 642818 45568 642824 45580
rect 642876 45568 642882 45620
rect 212442 45500 212448 45552
rect 212500 45540 212506 45552
rect 639322 45540 639328 45552
rect 212500 45512 639328 45540
rect 212500 45500 212506 45512
rect 639322 45500 639328 45512
rect 639380 45500 639386 45552
rect 194410 44072 194416 44124
rect 194468 44112 194474 44124
rect 661126 44112 661132 44124
rect 194468 44084 661132 44112
rect 194468 44072 194474 44084
rect 661126 44072 661132 44084
rect 661184 44072 661190 44124
rect 365162 43868 365168 43920
rect 365220 43908 365226 43920
rect 367094 43908 367100 43920
rect 365220 43880 367100 43908
rect 365220 43868 365226 43880
rect 367094 43868 367100 43880
rect 367152 43868 367158 43920
rect 310422 43800 310428 43852
rect 310480 43840 310486 43852
rect 311894 43840 311900 43852
rect 310480 43812 311900 43840
rect 310480 43800 310486 43812
rect 311894 43800 311900 43812
rect 311952 43800 311958 43852
rect 230474 43460 230480 43512
rect 230532 43500 230538 43512
rect 618254 43500 618260 43512
rect 230532 43472 618260 43500
rect 230532 43460 230538 43472
rect 618254 43460 618260 43472
rect 618312 43460 618318 43512
rect 230658 43392 230664 43444
rect 230716 43432 230722 43444
rect 621474 43432 621480 43444
rect 230716 43404 621480 43432
rect 230716 43392 230722 43404
rect 621474 43392 621480 43404
rect 621532 43392 621538 43444
rect 230842 43324 230848 43376
rect 230900 43364 230906 43376
rect 621198 43364 621204 43376
rect 230900 43336 621204 43364
rect 230900 43324 230906 43336
rect 621198 43324 621204 43336
rect 621256 43324 621262 43376
rect 230566 43256 230572 43308
rect 230624 43296 230630 43308
rect 621106 43296 621112 43308
rect 230624 43268 621112 43296
rect 230624 43256 230630 43268
rect 621106 43256 621112 43268
rect 621164 43256 621170 43308
rect 230750 43188 230756 43240
rect 230808 43228 230814 43240
rect 621290 43228 621296 43240
rect 230808 43200 621296 43228
rect 230808 43188 230814 43200
rect 621290 43188 621296 43200
rect 621348 43188 621354 43240
rect 226242 43120 226248 43172
rect 226300 43160 226306 43172
rect 622486 43160 622492 43172
rect 226300 43132 622492 43160
rect 226300 43120 226306 43132
rect 622486 43120 622492 43132
rect 622544 43120 622550 43172
rect 223482 43052 223488 43104
rect 223540 43092 223546 43104
rect 622302 43092 622308 43104
rect 223540 43064 622308 43092
rect 223540 43052 223546 43064
rect 622302 43052 622308 43064
rect 622360 43052 622366 43104
rect 52178 42712 52184 42764
rect 52236 42752 52242 42764
rect 215294 42752 215300 42764
rect 52236 42724 215300 42752
rect 52236 42712 52242 42724
rect 215294 42712 215300 42724
rect 215352 42712 215358 42764
rect 529658 42712 529664 42764
rect 529716 42752 529722 42764
rect 542998 42752 543004 42764
rect 529716 42724 543004 42752
rect 529716 42712 529722 42724
rect 542998 42712 543004 42724
rect 543056 42712 543062 42764
rect 475470 42616 475476 42628
rect 474490 42588 475476 42616
rect 475470 42576 475476 42588
rect 475528 42576 475534 42628
rect 513926 41964 513932 42016
rect 513984 42004 513990 42016
rect 520366 42004 520372 42016
rect 513984 41976 520372 42004
rect 513984 41964 513990 41976
rect 520366 41964 520372 41976
rect 520424 41964 520430 42016
rect 405826 41896 405832 41948
rect 405884 41936 405890 41948
rect 426342 41936 426348 41948
rect 405884 41908 426348 41936
rect 405884 41896 405890 41908
rect 426342 41896 426348 41908
rect 426400 41896 426406 41948
rect 514018 41896 514024 41948
rect 514076 41936 514082 41948
rect 514846 41936 514852 41948
rect 514076 41908 514852 41936
rect 514076 41896 514082 41908
rect 514846 41896 514852 41908
rect 514904 41896 514910 41948
rect 426342 41420 426348 41472
rect 426400 41460 426406 41472
rect 607490 41460 607496 41472
rect 426400 41432 607496 41460
rect 426400 41420 426406 41432
rect 607490 41420 607496 41432
rect 607548 41420 607554 41472
rect 506382 41352 506388 41404
rect 506440 41392 506446 41404
rect 513282 41392 513288 41404
rect 506440 41364 513288 41392
rect 506440 41352 506446 41364
rect 513282 41352 513288 41364
rect 513340 41352 513346 41404
rect 530394 41352 530400 41404
rect 530452 41392 530458 41404
rect 602982 41392 602988 41404
rect 530452 41364 602988 41392
rect 530452 41352 530458 41364
rect 602982 41352 602988 41364
rect 603040 41352 603046 41404
rect 530302 41284 530308 41336
rect 530360 41324 530366 41336
rect 571794 41324 571800 41336
rect 530360 41296 571800 41324
rect 530360 41284 530366 41296
rect 571794 41284 571800 41296
rect 571852 41284 571858 41336
rect 475562 38564 475568 38616
rect 475620 38604 475626 38616
rect 514018 38604 514024 38616
rect 475620 38576 514024 38604
rect 475620 38564 475626 38576
rect 514018 38564 514024 38576
rect 514076 38564 514082 38616
rect 502334 38496 502340 38548
rect 502392 38536 502398 38548
rect 513926 38536 513932 38548
rect 502392 38508 513932 38536
rect 502392 38496 502398 38508
rect 513926 38496 513932 38508
rect 513984 38496 513990 38548
rect 213178 24760 213184 24812
rect 213236 24800 213242 24812
rect 213822 24800 213828 24812
rect 213236 24772 213828 24800
rect 213236 24760 213242 24772
rect 213822 24760 213828 24772
rect 213880 24760 213886 24812
rect 224586 22992 224592 23044
rect 224644 23032 224650 23044
rect 226242 23032 226248 23044
rect 224644 23004 226248 23032
rect 224644 22992 224650 23004
rect 226242 22992 226248 23004
rect 226300 22992 226306 23044
rect 221734 22516 221740 22568
rect 221792 22556 221798 22568
rect 223482 22556 223488 22568
rect 221792 22528 223488 22556
rect 221792 22516 221798 22528
rect 223482 22516 223488 22528
rect 223540 22516 223546 22568
rect 229370 6468 229376 6520
rect 229428 6508 229434 6520
rect 233142 6508 233148 6520
rect 229428 6480 233148 6508
rect 229428 6468 229434 6480
rect 233142 6468 233148 6480
rect 233200 6468 233206 6520
<< via1 >>
rect 483572 1004640 483624 1004692
rect 655520 896996 655572 897048
rect 676036 896996 676088 897048
rect 673368 894616 673420 894668
rect 675852 894616 675904 894668
rect 655428 894480 655480 894532
rect 676036 894480 676088 894532
rect 670516 894412 670568 894464
rect 676128 894412 676180 894464
rect 655704 894344 655756 894396
rect 675944 894344 675996 894396
rect 670608 893800 670660 893852
rect 676036 893800 676088 893852
rect 670424 892984 670476 893036
rect 676036 892984 676088 893036
rect 674288 891488 674340 891540
rect 676036 891488 676088 891540
rect 674748 890672 674800 890724
rect 676036 890672 676088 890724
rect 674564 888768 674616 888820
rect 675944 888768 675996 888820
rect 675024 888700 675076 888752
rect 676036 888700 676088 888752
rect 673828 887816 673880 887868
rect 676036 887816 676088 887868
rect 673736 886048 673788 886100
rect 675944 886048 675996 886100
rect 674472 885980 674524 886032
rect 676036 885980 676088 886032
rect 655612 883260 655664 883312
rect 675392 883260 675444 883312
rect 671988 883192 672040 883244
rect 679532 883192 679584 883244
rect 675300 883124 675352 883176
rect 678980 883124 679032 883176
rect 675760 883056 675812 883108
rect 679348 883056 679400 883108
rect 674840 882988 674892 883040
rect 679624 882988 679676 883040
rect 674932 880404 674984 880456
rect 679072 880404 679124 880456
rect 675208 880336 675260 880388
rect 679164 880336 679216 880388
rect 675116 880268 675168 880320
rect 679256 880268 679308 880320
rect 674656 880200 674708 880252
rect 679440 880200 679492 880252
rect 675760 878364 675812 878416
rect 675760 877752 675812 877804
rect 674840 877276 674892 877328
rect 675300 877276 675352 877328
rect 674656 873740 674708 873792
rect 675116 873740 675168 873792
rect 673736 873604 673788 873656
rect 674656 873604 674708 873656
rect 675024 872720 675076 872772
rect 675024 872516 675076 872568
rect 674748 872448 674800 872500
rect 675208 872448 675260 872500
rect 673828 872312 673880 872364
rect 674748 872312 674800 872364
rect 655796 872176 655848 872228
rect 675116 872176 675168 872228
rect 674472 869932 674524 869984
rect 675208 869932 675260 869984
rect 674748 869388 674800 869440
rect 675208 869388 675260 869440
rect 674656 868708 674708 868760
rect 675208 868708 675260 868760
rect 674564 867552 674616 867604
rect 675116 867552 675168 867604
rect 674288 865716 674340 865768
rect 675208 865716 675260 865768
rect 656808 863812 656860 863864
rect 675116 863812 675168 863864
rect 41788 817640 41840 817692
rect 50988 817640 51040 817692
rect 41788 817232 41840 817284
rect 48320 817232 48372 817284
rect 41788 808256 41840 808308
rect 43536 808256 43588 808308
rect 42340 805944 42392 805996
rect 62120 805944 62172 805996
rect 41880 805876 41932 805928
rect 43352 805876 43404 805928
rect 41972 804244 42024 804296
rect 43260 804244 43312 804296
rect 42340 800436 42392 800488
rect 58256 800436 58308 800488
rect 42248 799280 42300 799332
rect 42708 799280 42760 799332
rect 42340 796832 42392 796884
rect 42616 796832 42668 796884
rect 42248 794996 42300 795048
rect 42892 794996 42944 795048
rect 42708 794860 42760 794912
rect 42892 794860 42944 794912
rect 42156 794248 42208 794300
rect 43260 794248 43312 794300
rect 42156 793772 42208 793824
rect 43536 793772 43588 793824
rect 42248 792616 42300 792668
rect 43076 792616 43128 792668
rect 655520 792140 655572 792192
rect 675392 792140 675444 792192
rect 42156 790644 42208 790696
rect 43352 790644 43404 790696
rect 42156 790100 42208 790152
rect 43904 790100 43956 790152
rect 42340 789352 42392 789404
rect 58072 789352 58124 789404
rect 42432 789284 42484 789336
rect 58532 789284 58584 789336
rect 42156 789216 42208 789268
rect 43812 789216 43864 789268
rect 42156 788808 42208 788860
rect 42892 788808 42944 788860
rect 42156 786972 42208 787024
rect 43444 786972 43496 787024
rect 48320 786564 48372 786616
rect 58440 786564 58492 786616
rect 50988 786496 51040 786548
rect 58532 786496 58584 786548
rect 42064 786224 42116 786276
rect 43720 786224 43772 786276
rect 673736 784728 673788 784780
rect 675116 784728 675168 784780
rect 656532 783844 656584 783896
rect 674656 783844 674708 783896
rect 673644 780920 673696 780972
rect 675208 780920 675260 780972
rect 674564 780104 674616 780156
rect 675484 780104 675536 780156
rect 675024 780036 675076 780088
rect 675024 779696 675076 779748
rect 674656 779560 674708 779612
rect 675116 779560 675168 779612
rect 674288 779084 674340 779136
rect 675208 779084 675260 779136
rect 673828 778608 673880 778660
rect 675208 778608 675260 778660
rect 674472 777316 674524 777368
rect 675392 777316 675444 777368
rect 654968 775480 655020 775532
rect 675116 775480 675168 775532
rect 41512 774732 41564 774784
rect 53748 774732 53800 774784
rect 41512 773848 41564 773900
rect 50988 773848 51040 773900
rect 41512 773440 41564 773492
rect 45468 773440 45520 773492
rect 675024 773372 675076 773424
rect 675668 773372 675720 773424
rect 674748 773304 674800 773356
rect 675760 773304 675812 773356
rect 674840 769632 674892 769684
rect 675300 769632 675352 769684
rect 42432 767388 42484 767440
rect 48228 767388 48280 767440
rect 38292 764464 38344 764516
rect 42248 764464 42300 764516
rect 41604 762832 41656 762884
rect 48320 762832 48372 762884
rect 38200 761676 38252 761728
rect 42156 761676 42208 761728
rect 41512 759296 41564 759348
rect 43536 759296 43588 759348
rect 42708 759092 42760 759144
rect 43352 759092 43404 759144
rect 38568 758956 38620 759008
rect 42708 758956 42760 759008
rect 43904 757732 43956 757784
rect 44180 757732 44232 757784
rect 43628 757596 43680 757648
rect 43904 757596 43956 757648
rect 42432 757460 42484 757512
rect 43628 757460 43680 757512
rect 42156 756984 42208 757036
rect 44272 756984 44324 757036
rect 42248 756236 42300 756288
rect 59268 756236 59320 756288
rect 42156 754876 42208 754928
rect 42340 754876 42392 754928
rect 42340 754264 42392 754316
rect 43076 754264 43128 754316
rect 43168 754196 43220 754248
rect 43168 753924 43220 753976
rect 42156 753312 42208 753364
rect 43260 753312 43312 753364
rect 42156 753040 42208 753092
rect 43168 753040 43220 753092
rect 42248 751748 42300 751800
rect 42708 751748 42760 751800
rect 42248 751204 42300 751256
rect 43352 751204 43404 751256
rect 42156 751068 42208 751120
rect 43076 751068 43128 751120
rect 43352 751068 43404 751120
rect 44088 751068 44140 751120
rect 42064 750592 42116 750644
rect 43536 750592 43588 750644
rect 42248 749368 42300 749420
rect 43812 749368 43864 749420
rect 655980 747940 656032 747992
rect 675392 747940 675444 747992
rect 43260 747872 43312 747924
rect 58440 747872 58492 747924
rect 42156 747464 42208 747516
rect 43536 747464 43588 747516
rect 42248 746240 42300 746292
rect 43996 746240 44048 746292
rect 42432 745220 42484 745272
rect 58440 745220 58492 745272
rect 45468 745152 45520 745204
rect 58532 745152 58584 745204
rect 42340 745084 42392 745136
rect 43352 745084 43404 745136
rect 673552 744132 673604 744184
rect 675760 744132 675812 744184
rect 42340 743248 42392 743300
rect 43904 743248 43956 743300
rect 42156 743044 42208 743096
rect 44088 743044 44140 743096
rect 50988 742364 51040 742416
rect 58440 742364 58492 742416
rect 53748 742296 53800 742348
rect 57980 742296 58032 742348
rect 674564 737264 674616 737316
rect 675208 737264 675260 737316
rect 655152 736992 655204 737044
rect 675208 736992 675260 737044
rect 656072 736924 656124 736976
rect 674840 736924 674892 736976
rect 674656 735632 674708 735684
rect 675392 735632 675444 735684
rect 674748 734748 674800 734800
rect 675392 734748 675444 734800
rect 673828 734136 673880 734188
rect 675392 734136 675444 734188
rect 673552 733864 673604 733916
rect 675392 733864 675444 733916
rect 675300 733796 675352 733848
rect 675300 733456 675352 733508
rect 673460 732300 673512 732352
rect 675392 732300 675444 732352
rect 674840 732028 674892 732080
rect 675392 732028 675444 732080
rect 41512 731076 41564 731128
rect 43628 731076 43680 731128
rect 674748 730464 674800 730516
rect 675392 730464 675444 730516
rect 674656 728764 674708 728816
rect 674656 728628 674708 728680
rect 675392 728628 675444 728680
rect 674564 728084 674616 728136
rect 676128 728084 676180 728136
rect 675208 728016 675260 728068
rect 678980 728016 679032 728068
rect 674564 727948 674616 728000
rect 673276 727880 673328 727932
rect 675208 727880 675260 727932
rect 674840 727812 674892 727864
rect 675116 727812 675168 727864
rect 673552 718836 673604 718888
rect 675576 718836 675628 718888
rect 673460 718700 673512 718752
rect 674656 718700 674708 718752
rect 41512 717612 41564 717664
rect 53748 717612 53800 717664
rect 41420 717476 41472 717528
rect 43536 717476 43588 717528
rect 670516 715368 670568 715420
rect 676036 715368 676088 715420
rect 655796 715232 655848 715284
rect 675944 715232 675996 715284
rect 655612 715096 655664 715148
rect 675760 715096 675812 715148
rect 655428 714960 655480 715012
rect 675852 714960 675904 715012
rect 675208 714892 675260 714944
rect 675760 714892 675812 714944
rect 42432 714824 42484 714876
rect 59360 714824 59412 714876
rect 670516 714824 670568 714876
rect 676036 714824 676088 714876
rect 673368 714484 673420 714536
rect 676036 714484 676088 714536
rect 43168 714144 43220 714196
rect 44364 714144 44416 714196
rect 673276 714008 673328 714060
rect 676036 714008 676088 714060
rect 41788 713804 41840 713856
rect 41788 713532 41840 713584
rect 669872 713396 669924 713448
rect 670424 713396 670476 713448
rect 676036 712512 676088 712564
rect 670608 712376 670660 712428
rect 669872 712308 669924 712360
rect 675944 712308 675996 712360
rect 43812 712240 43864 712292
rect 44272 712240 44324 712292
rect 670332 712240 670384 712292
rect 676036 712240 676088 712292
rect 670424 712172 670476 712224
rect 675852 712172 675904 712224
rect 43812 712104 43864 712156
rect 59268 712104 59320 712156
rect 675024 712104 675076 712156
rect 675944 712104 675996 712156
rect 42156 711696 42208 711748
rect 43352 711696 43404 711748
rect 673736 711492 673788 711544
rect 676036 711492 676088 711544
rect 42156 710880 42208 710932
rect 42432 710880 42484 710932
rect 42340 710268 42392 710320
rect 42708 710268 42760 710320
rect 42708 710132 42760 710184
rect 43260 710132 43312 710184
rect 43444 709860 43496 709912
rect 43904 709860 43956 709912
rect 43352 709792 43404 709844
rect 43996 709792 44048 709844
rect 43996 709588 44048 709640
rect 44272 709588 44324 709640
rect 44088 709520 44140 709572
rect 44364 709520 44416 709572
rect 43812 709384 43864 709436
rect 42248 709316 42300 709368
rect 674472 708840 674524 708892
rect 676036 708840 676088 708892
rect 42156 708568 42208 708620
rect 43628 708568 43680 708620
rect 674288 708228 674340 708280
rect 676036 708228 676088 708280
rect 673644 707820 673696 707872
rect 676036 707820 676088 707872
rect 42432 706732 42484 706784
rect 43444 706732 43496 706784
rect 42248 706188 42300 706240
rect 43536 706188 43588 706240
rect 42340 705916 42392 705968
rect 43260 705916 43312 705968
rect 672080 705100 672132 705152
rect 676036 705100 676088 705152
rect 42064 704216 42116 704268
rect 42708 704216 42760 704268
rect 42432 703808 42484 703860
rect 58532 703808 58584 703860
rect 655980 703808 656032 703860
rect 675392 703808 675444 703860
rect 42340 702448 42392 702500
rect 43352 702448 43404 702500
rect 42340 701904 42392 701956
rect 43812 701904 43864 701956
rect 42248 701768 42300 701820
rect 44088 701768 44140 701820
rect 42340 699388 42392 699440
rect 43996 699388 44048 699440
rect 654232 692860 654284 692912
rect 675208 692860 675260 692912
rect 673736 690140 673788 690192
rect 675300 690140 675352 690192
rect 654140 690004 654192 690056
rect 675300 690004 675352 690056
rect 673644 689120 673696 689172
rect 675484 689120 675536 689172
rect 675208 688712 675260 688764
rect 675484 688712 675536 688764
rect 673368 688576 673420 688628
rect 675392 688576 675444 688628
rect 41512 688304 41564 688356
rect 53840 688304 53892 688356
rect 673552 687828 673604 687880
rect 675116 687828 675168 687880
rect 41788 687624 41840 687676
rect 50988 687624 51040 687676
rect 674472 687284 674524 687336
rect 675392 687284 675444 687336
rect 41788 687216 41840 687268
rect 45744 687216 45796 687268
rect 675116 684224 675168 684276
rect 675208 684224 675260 684276
rect 675024 684020 675076 684072
rect 674288 683884 674340 683936
rect 675024 683884 675076 683936
rect 675208 683884 675260 683936
rect 675116 683612 675168 683664
rect 675392 683612 675444 683664
rect 673736 680348 673788 680400
rect 674288 680348 674340 680400
rect 675300 678920 675352 678972
rect 679072 678920 679124 678972
rect 41788 678580 41840 678632
rect 44088 678580 44140 678632
rect 41788 676608 41840 676660
rect 43168 676608 43220 676660
rect 5540 675724 5592 675776
rect 30564 675724 30616 675776
rect 5448 674772 5500 674824
rect 43352 674772 43404 674824
rect 43076 672528 43128 672580
rect 43536 672528 43588 672580
rect 41880 672392 41932 672444
rect 43076 672392 43128 672444
rect 43444 672120 43496 672172
rect 43996 672120 44048 672172
rect 43260 671984 43312 672036
rect 43444 671984 43496 672036
rect 42340 671780 42392 671832
rect 43168 671780 43220 671832
rect 655888 670896 655940 670948
rect 676220 670896 676272 670948
rect 43536 670828 43588 670880
rect 43996 670828 44048 670880
rect 42340 670760 42392 670812
rect 60648 670760 60700 670812
rect 655704 670760 655756 670812
rect 676036 670760 676088 670812
rect 42432 670692 42484 670744
rect 43536 670692 43588 670744
rect 43720 670624 43772 670676
rect 44272 670624 44324 670676
rect 41788 670556 41840 670608
rect 41788 670352 41840 670404
rect 673276 669332 673328 669384
rect 676036 669332 676088 669384
rect 669596 669264 669648 669316
rect 670516 669264 670568 669316
rect 669596 668176 669648 668228
rect 676128 668176 676180 668228
rect 670424 668108 670476 668160
rect 676220 668108 676272 668160
rect 655520 668040 655572 668092
rect 678980 668040 679032 668092
rect 670608 667972 670660 668024
rect 676312 667972 676364 668024
rect 42248 667836 42300 667888
rect 43168 667836 43220 667888
rect 675208 667836 675260 667888
rect 676036 667836 676088 667888
rect 42156 667700 42208 667752
rect 42340 667700 42392 667752
rect 43168 667700 43220 667752
rect 44180 667700 44232 667752
rect 42156 666680 42208 666732
rect 43628 666680 43680 666732
rect 674564 665932 674616 665984
rect 676036 665932 676088 665984
rect 670240 665252 670292 665304
rect 676220 665252 676272 665304
rect 42156 665184 42208 665236
rect 43260 665184 43312 665236
rect 670332 665184 670384 665236
rect 678980 665184 679032 665236
rect 675024 665116 675076 665168
rect 676036 665116 676088 665168
rect 674748 665048 674800 665100
rect 676128 665048 676180 665100
rect 42156 664640 42208 664692
rect 43536 664640 43588 664692
rect 43628 664504 43680 664556
rect 44272 664504 44324 664556
rect 674656 664300 674708 664352
rect 676036 664300 676088 664352
rect 42156 664164 42208 664216
rect 43168 664164 43220 664216
rect 42156 663348 42208 663400
rect 43076 663348 43128 663400
rect 673828 663076 673880 663128
rect 676036 663076 676088 663128
rect 42156 661036 42208 661088
rect 43352 661036 43404 661088
rect 42156 660492 42208 660544
rect 43260 660492 43312 660544
rect 42432 659676 42484 659728
rect 58440 659676 58492 659728
rect 672172 659676 672224 659728
rect 678980 659676 679032 659728
rect 42248 659608 42300 659660
rect 58532 659608 58584 659660
rect 45744 659540 45796 659592
rect 58624 659540 58676 659592
rect 42248 659472 42300 659524
rect 43628 659472 43680 659524
rect 42156 659200 42208 659252
rect 44088 659200 44140 659252
rect 42156 657364 42208 657416
rect 43536 657364 43588 657416
rect 655704 656888 655756 656940
rect 675392 656888 675444 656940
rect 50988 656820 51040 656872
rect 58440 656820 58492 656872
rect 53840 656752 53892 656804
rect 58992 656752 59044 656804
rect 42156 656004 42208 656056
rect 43904 656004 43956 656056
rect 673736 649544 673788 649596
rect 675392 649544 675444 649596
rect 674656 648932 674708 648984
rect 675116 648932 675168 648984
rect 674564 648864 674616 648916
rect 675300 648864 675352 648916
rect 654416 648592 654468 648644
rect 675116 648592 675168 648644
rect 673460 647708 673512 647760
rect 675392 647708 675444 647760
rect 656440 645872 656492 645924
rect 675208 645872 675260 645924
rect 674748 645192 674800 645244
rect 675392 645192 675444 645244
rect 41512 645056 41564 645108
rect 53840 645056 53892 645108
rect 41788 644988 41840 645040
rect 56508 644988 56560 645040
rect 673828 644580 673880 644632
rect 675392 644580 675444 644632
rect 673276 644240 673328 644292
rect 673736 644240 673788 644292
rect 673736 644104 673788 644156
rect 675392 644104 675444 644156
rect 41788 644036 41840 644088
rect 50988 644036 51040 644088
rect 675484 643560 675536 643612
rect 675116 643492 675168 643544
rect 675392 643492 675444 643544
rect 675208 643356 675260 643408
rect 674656 642200 674708 642252
rect 675116 642200 675168 642252
rect 674656 642064 674708 642116
rect 675392 642064 675444 642116
rect 675116 640772 675168 640824
rect 675300 640704 675352 640756
rect 675024 640228 675076 640280
rect 675392 640228 675444 640280
rect 675208 638664 675260 638716
rect 675208 638460 675260 638512
rect 675116 638392 675168 638444
rect 675484 638392 675536 638444
rect 674564 638188 674616 638240
rect 675760 638188 675812 638240
rect 673736 638052 673788 638104
rect 674564 638052 674616 638104
rect 673276 637916 673328 637968
rect 673736 637916 673788 637968
rect 674748 637780 674800 637832
rect 675208 637780 675260 637832
rect 675668 637508 675720 637560
rect 679072 637508 679124 637560
rect 673828 637236 673880 637288
rect 674656 637236 674708 637288
rect 673460 637100 673512 637152
rect 673828 637100 673880 637152
rect 41512 633224 41564 633276
rect 48412 633224 48464 633276
rect 20628 632612 20680 632664
rect 30196 632612 30248 632664
rect 42432 630912 42484 630964
rect 43720 630912 43772 630964
rect 43168 630844 43220 630896
rect 43812 630844 43864 630896
rect 20628 630776 20680 630828
rect 43720 630776 43772 630828
rect 24768 630708 24820 630760
rect 43168 630708 43220 630760
rect 43076 629348 43128 629400
rect 43996 629348 44048 629400
rect 38476 629212 38528 629264
rect 43076 629212 43128 629264
rect 43352 626832 43404 626884
rect 43628 626832 43680 626884
rect 42708 626696 42760 626748
rect 43352 626696 43404 626748
rect 42708 626560 42760 626612
rect 58532 626560 58584 626612
rect 42156 625268 42208 625320
rect 42340 625268 42392 625320
rect 42340 624452 42392 624504
rect 42708 624452 42760 624504
rect 655796 624112 655848 624164
rect 678980 624112 679032 624164
rect 670608 624044 670660 624096
rect 676220 624044 676272 624096
rect 655612 623976 655664 624028
rect 676312 623976 676364 624028
rect 670516 623908 670568 623960
rect 676128 623908 676180 623960
rect 655428 623840 655480 623892
rect 676036 623840 676088 623892
rect 673276 623772 673328 623824
rect 675944 623772 675996 623824
rect 674932 623704 674984 623756
rect 676036 623704 676088 623756
rect 42156 623432 42208 623484
rect 43260 623432 43312 623484
rect 42248 622412 42300 622464
rect 42708 622412 42760 622464
rect 42340 622208 42392 622260
rect 43076 622208 43128 622260
rect 42340 621664 42392 621716
rect 43444 621664 43496 621716
rect 670608 621120 670660 621172
rect 676128 621120 676180 621172
rect 670424 621052 670476 621104
rect 676220 621052 676272 621104
rect 670240 620984 670292 621036
rect 676312 620984 676364 621036
rect 674288 620916 674340 620968
rect 676036 620916 676088 620968
rect 42064 620780 42116 620832
rect 43628 620780 43680 620832
rect 42064 620168 42116 620220
rect 43076 620168 43128 620220
rect 673552 620100 673604 620152
rect 676036 620100 676088 620152
rect 42432 619148 42484 619200
rect 43168 619148 43220 619200
rect 42708 618196 42760 618248
rect 58164 618196 58216 618248
rect 674472 618196 674524 618248
rect 676036 618196 676088 618248
rect 673644 618060 673696 618112
rect 676036 618060 676088 618112
rect 42064 617312 42116 617364
rect 43352 617312 43404 617364
rect 673368 616700 673420 616752
rect 676220 616700 676272 616752
rect 42340 616020 42392 616072
rect 44088 616020 44140 616072
rect 42248 615952 42300 616004
rect 43720 615952 43772 616004
rect 42156 615816 42208 615868
rect 43812 615816 43864 615868
rect 42432 615476 42484 615528
rect 58532 615476 58584 615528
rect 50988 615408 51040 615460
rect 58164 615408 58216 615460
rect 672264 614592 672316 614644
rect 679072 614592 679124 614644
rect 42156 614184 42208 614236
rect 43996 614184 44048 614236
rect 655428 612824 655480 612876
rect 675668 612824 675720 612876
rect 56508 612688 56560 612740
rect 57980 612688 58032 612740
rect 53840 612076 53892 612128
rect 57980 612076 58032 612128
rect 674288 608948 674340 609000
rect 675576 608948 675628 609000
rect 674472 605072 674524 605124
rect 675208 605072 675260 605124
rect 673644 603440 673696 603492
rect 675484 603440 675536 603492
rect 656808 601740 656860 601792
rect 675208 601740 675260 601792
rect 41788 601672 41840 601724
rect 56508 601672 56560 601724
rect 655612 601672 655664 601724
rect 675300 601672 675352 601724
rect 673552 600380 673604 600432
rect 674472 600380 674524 600432
rect 674472 600244 674524 600296
rect 675484 600244 675536 600296
rect 674288 599904 674340 599956
rect 674656 599904 674708 599956
rect 674288 599768 674340 599820
rect 675484 599768 675536 599820
rect 674932 598952 674984 599004
rect 675392 598952 675444 599004
rect 675208 598884 675260 598936
rect 675300 598816 675352 598868
rect 675392 598680 675444 598732
rect 675300 598612 675352 598664
rect 673460 598544 673512 598596
rect 675484 598544 675536 598596
rect 673552 597252 673604 597304
rect 675208 597252 675260 597304
rect 673552 597116 673604 597168
rect 675392 597116 675444 597168
rect 674656 595416 674708 595468
rect 675208 595416 675260 595468
rect 674656 595280 674708 595332
rect 675392 595280 675444 595332
rect 675300 593512 675352 593564
rect 675208 593172 675260 593224
rect 675576 593172 675628 593224
rect 43076 592968 43128 593020
rect 43352 592968 43404 593020
rect 43352 592832 43404 592884
rect 44088 592832 44140 592884
rect 678980 592752 679032 592804
rect 674932 589364 674984 589416
rect 675300 589364 675352 589416
rect 41512 589228 41564 589280
rect 53840 589228 53892 589280
rect 674472 589228 674524 589280
rect 674932 589228 674984 589280
rect 38568 587800 38620 587852
rect 42340 587800 42392 587852
rect 43076 585148 43128 585200
rect 58532 585148 58584 585200
rect 42432 584196 42484 584248
rect 44272 584196 44324 584248
rect 43352 583856 43404 583908
rect 673460 583720 673512 583772
rect 674472 583720 674524 583772
rect 674656 583720 674708 583772
rect 675208 583720 675260 583772
rect 43536 583652 43588 583704
rect 673552 583584 673604 583636
rect 674656 583584 674708 583636
rect 42248 582564 42300 582616
rect 59360 582564 59412 582616
rect 42156 582088 42208 582140
rect 43260 582088 43312 582140
rect 43260 581952 43312 582004
rect 43536 581952 43588 582004
rect 42156 581476 42208 581528
rect 43076 581476 43128 581528
rect 43444 580388 43496 580440
rect 43996 580388 44048 580440
rect 42248 580320 42300 580372
rect 44088 580320 44140 580372
rect 42248 580116 42300 580168
rect 44088 580116 44140 580168
rect 656164 580048 656216 580100
rect 676220 580048 676272 580100
rect 655980 579912 656032 579964
rect 676128 579912 676180 579964
rect 655520 579776 655572 579828
rect 676312 579776 676364 579828
rect 670516 579640 670568 579692
rect 676220 579640 676272 579692
rect 673276 579028 673328 579080
rect 676036 579028 676088 579080
rect 42248 578960 42300 579012
rect 43628 578960 43680 579012
rect 42156 578756 42208 578808
rect 43168 578756 43220 578808
rect 42156 578416 42208 578468
rect 43812 578416 43864 578468
rect 43904 578416 43956 578468
rect 673368 578416 673420 578468
rect 676220 578416 676272 578468
rect 43904 578212 43956 578264
rect 42248 577124 42300 577176
rect 44088 577124 44140 577176
rect 42156 576920 42208 576972
rect 43076 576920 43128 576972
rect 670424 576920 670476 576972
rect 676220 576920 676272 576972
rect 670608 576852 670660 576904
rect 676128 576852 676180 576904
rect 675024 576784 675076 576836
rect 676036 576784 676088 576836
rect 673736 576716 673788 576768
rect 675944 576716 675996 576768
rect 675116 576036 675168 576088
rect 676036 576036 676088 576088
rect 42340 575968 42392 576020
rect 43536 575968 43588 576020
rect 42432 574064 42484 574116
rect 60648 574064 60700 574116
rect 42156 573792 42208 573844
rect 43352 573792 43404 573844
rect 674748 573656 674800 573708
rect 676036 573656 676088 573708
rect 42340 572840 42392 572892
rect 43444 572840 43496 572892
rect 674564 572772 674616 572824
rect 676036 572772 676088 572824
rect 673828 572364 673880 572416
rect 676036 572364 676088 572416
rect 42248 571956 42300 572008
rect 44088 571956 44140 572008
rect 42340 571616 42392 571668
rect 43720 571616 43772 571668
rect 56508 571276 56560 571328
rect 58716 571276 58768 571328
rect 42064 570936 42116 570988
rect 43260 570936 43312 570988
rect 673460 568760 673512 568812
rect 675392 568760 675444 568812
rect 655980 568624 656032 568676
rect 675392 568624 675444 568676
rect 672356 568556 672408 568608
rect 678980 568556 679032 568608
rect 673828 564408 673880 564460
rect 675300 564408 675352 564460
rect 675024 559512 675076 559564
rect 675484 559512 675536 559564
rect 41512 558764 41564 558816
rect 56508 558764 56560 558816
rect 41512 558628 41564 558680
rect 53932 558628 53984 558680
rect 674288 558220 674340 558272
rect 675392 558220 675444 558272
rect 674564 558016 674616 558068
rect 675300 558016 675352 558068
rect 41512 557540 41564 557592
rect 50988 557540 51040 557592
rect 654232 557540 654284 557592
rect 675116 557540 675168 557592
rect 674748 555228 674800 555280
rect 675392 555228 675444 555280
rect 654140 554752 654192 554804
rect 675300 554752 675352 554804
rect 673092 554684 673144 554736
rect 673460 554684 673512 554736
rect 673460 554548 673512 554600
rect 675392 554548 675444 554600
rect 673736 553800 673788 553852
rect 675576 553800 675628 553852
rect 675484 553732 675536 553784
rect 675116 553460 675168 553512
rect 675392 553460 675444 553512
rect 675116 553324 675168 553376
rect 673184 552168 673236 552220
rect 673828 552168 673880 552220
rect 673828 552032 673880 552084
rect 674564 552032 674616 552084
rect 674564 551896 674616 551948
rect 675392 551896 675444 551948
rect 673276 548972 673328 549024
rect 673460 548972 673512 549024
rect 673460 548836 673512 548888
rect 675300 548836 675352 548888
rect 41512 548632 41564 548684
rect 43628 548632 43680 548684
rect 41512 548428 41564 548480
rect 43260 548428 43312 548480
rect 673092 547952 673144 548004
rect 675392 547952 675444 548004
rect 673184 547612 673236 547664
rect 677600 547612 677652 547664
rect 41512 546864 41564 546916
rect 45744 546864 45796 546916
rect 41604 546388 41656 546440
rect 43720 546388 43772 546440
rect 41420 546320 41472 546372
rect 43444 546320 43496 546372
rect 673828 545232 673880 545284
rect 675576 545232 675628 545284
rect 673828 545096 673880 545148
rect 674288 545096 674340 545148
rect 674748 545096 674800 545148
rect 675024 545096 675076 545148
rect 674840 544756 674892 544808
rect 675116 544756 675168 544808
rect 673736 544552 673788 544604
rect 674288 544552 674340 544604
rect 673276 544416 673328 544468
rect 673736 544416 673788 544468
rect 675392 543668 675444 543720
rect 679440 543668 679492 543720
rect 674840 542104 674892 542156
rect 675300 542104 675352 542156
rect 41788 541016 41840 541068
rect 42248 541016 42300 541068
rect 43076 541016 43128 541068
rect 59268 541016 59320 541068
rect 59452 540948 59504 541000
rect 41788 540744 41840 540796
rect 42064 538908 42116 538960
rect 43352 538908 43404 538960
rect 42248 538092 42300 538144
rect 43076 538092 43128 538144
rect 42064 537072 42116 537124
rect 43168 537072 43220 537124
rect 655888 535712 655940 535764
rect 676036 535712 676088 535764
rect 42156 535576 42208 535628
rect 43260 535576 43312 535628
rect 655704 535576 655756 535628
rect 676220 535576 676272 535628
rect 42064 535032 42116 535084
rect 43720 535032 43772 535084
rect 42156 534420 42208 534472
rect 43628 534420 43680 534472
rect 673368 534080 673420 534132
rect 676036 534080 676088 534132
rect 42156 533944 42208 533996
rect 43352 533944 43404 533996
rect 655796 532856 655848 532908
rect 678980 532856 679032 532908
rect 674932 532788 674984 532840
rect 675208 532720 675260 532772
rect 676220 532720 676272 532772
rect 678980 532720 679032 532772
rect 42156 531428 42208 531480
rect 43444 531428 43496 531480
rect 42156 530680 42208 530732
rect 42340 530680 42392 530732
rect 43260 529932 43312 529984
rect 58532 529932 58584 529984
rect 50988 529864 51040 529916
rect 58348 529864 58400 529916
rect 674656 529864 674708 529916
rect 676036 529864 676088 529916
rect 673644 529796 673696 529848
rect 675760 529796 675812 529848
rect 42156 529456 42208 529508
rect 43076 529456 43128 529508
rect 42156 527756 42208 527808
rect 42432 527756 42484 527808
rect 56508 527076 56560 527128
rect 60648 527076 60700 527128
rect 674472 527076 674524 527128
rect 676036 527076 676088 527128
rect 53932 527008 53984 527060
rect 59360 527008 59412 527060
rect 42156 526396 42208 526448
rect 43168 526396 43220 526448
rect 42156 525716 42208 525768
rect 43260 525716 43312 525768
rect 672448 524424 672500 524476
rect 678980 524424 679032 524476
rect 674748 493348 674800 493400
rect 675852 493348 675904 493400
rect 673460 492532 673512 492584
rect 675484 492532 675536 492584
rect 675392 492328 675444 492380
rect 676036 492328 676088 492380
rect 655612 491648 655664 491700
rect 676036 491648 676088 491700
rect 655520 491512 655572 491564
rect 676036 491512 676088 491564
rect 655428 491376 655480 491428
rect 675944 491376 675996 491428
rect 676220 491240 676272 491292
rect 677416 491240 677468 491292
rect 676220 488520 676272 488572
rect 677488 488520 677540 488572
rect 674840 485732 674892 485784
rect 676036 485732 676088 485784
rect 674564 485664 674616 485716
rect 675944 485664 675996 485716
rect 673828 485596 673880 485648
rect 675852 485596 675904 485648
rect 675024 485460 675076 485512
rect 676036 485460 676088 485512
rect 673552 483420 673604 483472
rect 676036 483420 676088 483472
rect 674288 482944 674340 482996
rect 676036 482944 676088 482996
rect 673736 482876 673788 482928
rect 675944 482876 675996 482928
rect 672540 480700 672592 480752
rect 676036 480700 676088 480752
rect 676128 475396 676180 475448
rect 679166 475396 679218 475448
rect 676036 475208 676088 475260
rect 679624 475208 679676 475260
rect 675944 475016 675996 475068
rect 679440 475016 679492 475068
rect 41788 430856 41840 430908
rect 56508 430856 56560 430908
rect 41788 419432 41840 419484
rect 45928 419432 45980 419484
rect 41972 416644 42024 416696
rect 43168 416644 43220 416696
rect 41880 416576 41932 416628
rect 43076 416576 43128 416628
rect 42340 411204 42392 411256
rect 43076 411204 43128 411256
rect 43076 410796 43128 410848
rect 43812 410796 43864 410848
rect 43812 409844 43864 409896
rect 43996 409844 44048 409896
rect 43996 409708 44048 409760
rect 44180 409708 44232 409760
rect 42248 409504 42300 409556
rect 42340 409300 42392 409352
rect 42064 408008 42116 408060
rect 43260 408008 43312 408060
rect 42156 407872 42208 407924
rect 42340 407872 42392 407924
rect 42156 407600 42208 407652
rect 43168 407600 43220 407652
rect 42064 406784 42116 406836
rect 43352 406784 43404 406836
rect 42156 406172 42208 406224
rect 43628 406172 43680 406224
rect 42248 405628 42300 405680
rect 58164 405628 58216 405680
rect 42248 405492 42300 405544
rect 43076 405492 43128 405544
rect 42432 405152 42484 405204
rect 42708 405152 42760 405204
rect 42156 403860 42208 403912
rect 43996 403860 44048 403912
rect 42156 403316 42208 403368
rect 44088 403316 44140 403368
rect 655704 403112 655756 403164
rect 676220 403112 676272 403164
rect 655520 403044 655572 403096
rect 676312 403044 676364 403096
rect 655428 402976 655480 403028
rect 675852 402976 675904 403028
rect 42340 402908 42392 402960
rect 58164 402908 58216 402960
rect 42340 402772 42392 402824
rect 43536 402772 43588 402824
rect 42340 400596 42392 400648
rect 43444 400596 43496 400648
rect 42340 399644 42392 399696
rect 43812 399644 43864 399696
rect 56508 399644 56560 399696
rect 58164 399644 58216 399696
rect 674472 398216 674524 398268
rect 676036 398216 676088 398268
rect 674564 397604 674616 397656
rect 675944 397604 675996 397656
rect 673736 397536 673788 397588
rect 676128 397536 676180 397588
rect 674656 397468 674708 397520
rect 676036 397468 676088 397520
rect 674288 396992 674340 397044
rect 676036 396992 676088 397044
rect 673460 395360 673512 395412
rect 675852 395360 675904 395412
rect 674840 394952 674892 395004
rect 675944 394952 675996 395004
rect 673552 394884 673604 394936
rect 675852 394884 675904 394936
rect 675024 394816 675076 394868
rect 676128 394816 676180 394868
rect 675116 394748 675168 394800
rect 675944 394748 675996 394800
rect 675208 394680 675260 394732
rect 676036 394680 676088 394732
rect 42156 394612 42208 394664
rect 58900 394612 58952 394664
rect 673644 394136 673696 394188
rect 676036 394136 676088 394188
rect 672816 392028 672868 392080
rect 678980 392028 679032 392080
rect 673828 391960 673880 392012
rect 676036 391960 676088 392012
rect 41512 387812 41564 387864
rect 53932 387812 53984 387864
rect 41788 387744 41840 387796
rect 56508 387744 56560 387796
rect 41512 386656 41564 386708
rect 50988 386656 51040 386708
rect 675760 386588 675812 386640
rect 673368 385976 673420 386028
rect 674564 385976 674616 386028
rect 675392 385976 675444 386028
rect 675760 385976 675812 386028
rect 674564 385840 674616 385892
rect 675208 385568 675260 385620
rect 675392 385568 675444 385620
rect 673736 384956 673788 385008
rect 675208 384956 675260 385008
rect 674472 384752 674524 384804
rect 675392 384752 675444 384804
rect 673368 384684 673420 384736
rect 673644 384684 673696 384736
rect 674656 383120 674708 383172
rect 675392 383120 675444 383172
rect 675024 382440 675076 382492
rect 675392 382440 675444 382492
rect 674840 381896 674892 381948
rect 675392 381896 675444 381948
rect 675116 381284 675168 381336
rect 675392 381284 675444 381336
rect 674288 381148 674340 381200
rect 675116 381148 675168 381200
rect 43444 379448 43496 379500
rect 43352 379176 43404 379228
rect 43536 379312 43588 379364
rect 44088 379312 44140 379364
rect 673644 378768 673696 378820
rect 675392 378768 675444 378820
rect 673736 378156 673788 378208
rect 675484 378156 675536 378208
rect 673552 377408 673604 377460
rect 675392 377408 675444 377460
rect 673828 376932 673880 376984
rect 675484 376932 675536 376984
rect 41788 376184 41840 376236
rect 46020 376184 46072 376236
rect 673460 375708 673512 375760
rect 675392 375708 675444 375760
rect 38200 375300 38252 375352
rect 42248 375300 42300 375352
rect 41420 375232 41472 375284
rect 43260 375232 43312 375284
rect 42340 374212 42392 374264
rect 42708 374212 42760 374264
rect 675024 373464 675076 373516
rect 675300 373464 675352 373516
rect 41604 372784 41656 372836
rect 43996 372784 44048 372836
rect 654508 372512 654560 372564
rect 674564 372512 674616 372564
rect 41512 371424 41564 371476
rect 42708 371424 42760 371476
rect 43720 371288 43772 371340
rect 43812 371084 43864 371136
rect 41972 370200 42024 370252
rect 42248 369316 42300 369368
rect 42156 368092 42208 368144
rect 42340 368092 42392 368144
rect 42156 366256 42208 366308
rect 43168 366256 43220 366308
rect 42340 366120 42392 366172
rect 43168 366120 43220 366172
rect 42340 365032 42392 365084
rect 42156 364760 42208 364812
rect 42708 364760 42760 364812
rect 42708 364624 42760 364676
rect 42248 364080 42300 364132
rect 43444 364080 43496 364132
rect 43444 363944 43496 363996
rect 43904 363944 43956 363996
rect 42156 363808 42208 363860
rect 43260 363808 43312 363860
rect 43168 363740 43220 363792
rect 43996 363740 44048 363792
rect 42156 363128 42208 363180
rect 43536 363128 43588 363180
rect 42432 361904 42484 361956
rect 43076 361904 43128 361956
rect 42340 361564 42392 361616
rect 58348 361496 58400 361548
rect 42708 361292 42760 361344
rect 58164 361292 58216 361344
rect 42064 360612 42116 360664
rect 43904 360612 43956 360664
rect 42340 360272 42392 360324
rect 43444 360272 43496 360324
rect 42156 359932 42208 359984
rect 43996 359932 44048 359984
rect 50988 358708 51040 358760
rect 58532 358708 58584 358760
rect 42432 358300 42484 358352
rect 43352 358300 43404 358352
rect 673092 357008 673144 357060
rect 675668 357008 675720 357060
rect 42432 356464 42484 356516
rect 43628 356464 43680 356516
rect 655520 356464 655572 356516
rect 675944 356464 675996 356516
rect 42340 356396 42392 356448
rect 43812 356396 43864 356448
rect 655428 356328 655480 356380
rect 676036 356328 676088 356380
rect 655612 356192 655664 356244
rect 675852 356192 675904 356244
rect 673368 356124 673420 356176
rect 676036 356124 676088 356176
rect 56508 355988 56560 356040
rect 58072 355988 58124 356040
rect 53932 355920 53984 355972
rect 59360 355920 59412 355972
rect 673184 355376 673236 355428
rect 676036 355376 676088 355428
rect 673276 354560 673328 354612
rect 676036 354560 676088 354612
rect 674656 353472 674708 353524
rect 676036 353472 676088 353524
rect 675116 353268 675168 353320
rect 676036 353268 676088 353320
rect 674840 351432 674892 351484
rect 676036 351432 676088 351484
rect 673736 351024 673788 351076
rect 675944 351024 675996 351076
rect 673552 350820 673604 350872
rect 675852 350820 675904 350872
rect 673460 350684 673512 350736
rect 675852 350684 675904 350736
rect 674564 350616 674616 350668
rect 675944 350616 675996 350668
rect 675208 350548 675260 350600
rect 676036 350548 676088 350600
rect 42156 350480 42208 350532
rect 58624 350480 58676 350532
rect 674288 349800 674340 349852
rect 676036 349800 676088 349852
rect 673644 347896 673696 347948
rect 675852 347896 675904 347948
rect 674472 347828 674524 347880
rect 675944 347828 675996 347880
rect 675024 347760 675076 347812
rect 676036 347760 676088 347812
rect 672908 347216 672960 347268
rect 676036 347216 676088 347268
rect 41512 344224 41564 344276
rect 46572 344224 46624 344276
rect 41512 343816 41564 343868
rect 46388 343816 46440 343868
rect 41512 343408 41564 343460
rect 46480 343408 46532 343460
rect 41512 342864 41564 342916
rect 44088 342864 44140 342916
rect 673828 341776 673880 341828
rect 674288 341776 674340 341828
rect 674288 341640 674340 341692
rect 674472 341640 674524 341692
rect 674564 341368 674616 341420
rect 675392 341368 675444 341420
rect 675116 340824 675168 340876
rect 675024 340756 675076 340808
rect 675484 340756 675536 340808
rect 675024 340620 675076 340672
rect 675392 340620 675444 340672
rect 675116 340416 675168 340468
rect 674656 339532 674708 339584
rect 675484 339532 675536 339584
rect 674840 337900 674892 337952
rect 675484 337900 675536 337952
rect 674472 336676 674524 336728
rect 675208 336676 675260 336728
rect 674288 335452 674340 335504
rect 675116 335452 675168 335504
rect 673736 335384 673788 335436
rect 675208 335384 675260 335436
rect 655980 335316 656032 335368
rect 675024 335316 675076 335368
rect 41604 332800 41656 332852
rect 46204 332800 46256 332852
rect 673828 332392 673880 332444
rect 675116 332392 675168 332444
rect 673644 331712 673696 331764
rect 675116 331712 675168 331764
rect 41420 331168 41472 331220
rect 43536 331168 43588 331220
rect 673460 331100 673512 331152
rect 675116 331100 675168 331152
rect 41512 330080 41564 330132
rect 43076 330080 43128 330132
rect 33048 329944 33100 329996
rect 42248 329944 42300 329996
rect 674564 328720 674616 328772
rect 675392 328720 675444 328772
rect 41788 326952 41840 327004
rect 673552 326884 673604 326936
rect 675392 326884 675444 326936
rect 41788 326748 41840 326800
rect 42248 323144 42300 323196
rect 42248 322940 42300 322992
rect 42248 321988 42300 322040
rect 43720 321988 43772 322040
rect 42248 321784 42300 321836
rect 43260 321784 43312 321836
rect 42156 321580 42208 321632
rect 43444 321580 43496 321632
rect 42248 320560 42300 320612
rect 43168 320560 43220 320612
rect 42156 320424 42208 320476
rect 43628 320424 43680 320476
rect 42432 318724 42484 318776
rect 42708 318724 42760 318776
rect 43720 318724 43772 318776
rect 58440 318724 58492 318776
rect 42340 317364 42392 317416
rect 58164 317364 58216 317416
rect 42432 316888 42484 316940
rect 43076 316888 43128 316940
rect 42340 316820 42392 316872
rect 43536 316820 43588 316872
rect 46480 314576 46532 314628
rect 58532 314576 58584 314628
rect 46572 314508 46624 314560
rect 58164 314508 58216 314560
rect 673092 312400 673144 312452
rect 676036 312400 676088 312452
rect 655428 312128 655480 312180
rect 676220 312128 676272 312180
rect 655704 311992 655756 312044
rect 676312 311992 676364 312044
rect 655520 311924 655572 311976
rect 676128 311924 676180 311976
rect 671620 311856 671672 311908
rect 676220 311856 676272 311908
rect 46388 311788 46440 311840
rect 58532 311788 58584 311840
rect 673368 311652 673420 311704
rect 676036 311652 676088 311704
rect 673368 311040 673420 311092
rect 676220 311040 676272 311092
rect 673184 310632 673236 310684
rect 676220 310632 676272 310684
rect 671712 310224 671764 310276
rect 676220 310224 676272 310276
rect 673276 309816 673328 309868
rect 676220 309816 676272 309868
rect 671804 309408 671856 309460
rect 676220 309408 676272 309460
rect 674656 309136 674708 309188
rect 676036 309136 676088 309188
rect 673460 308048 673512 308100
rect 676036 308048 676088 308100
rect 674472 306824 674524 306876
rect 676036 306824 676088 306876
rect 674564 306416 674616 306468
rect 676036 306416 676088 306468
rect 673552 306348 673604 306400
rect 676128 306348 676180 306400
rect 42064 306280 42116 306332
rect 58348 306280 58400 306332
rect 675208 306008 675260 306060
rect 676036 306008 676088 306060
rect 673644 305056 673696 305108
rect 676128 305056 676180 305108
rect 675024 304784 675076 304836
rect 676036 304784 676088 304836
rect 673828 304308 673880 304360
rect 676128 304308 676180 304360
rect 674840 304172 674892 304224
rect 676036 304172 676088 304224
rect 674288 303900 674340 303952
rect 676128 303900 676180 303952
rect 673736 303696 673788 303748
rect 676036 303696 676088 303748
rect 41880 301384 41932 301436
rect 54024 301384 54076 301436
rect 41788 301316 41840 301368
rect 57888 301316 57940 301368
rect 41788 301180 41840 301232
rect 43352 301180 43404 301232
rect 673000 300840 673052 300892
rect 678980 300840 679032 300892
rect 675116 298256 675168 298308
rect 675392 298256 675444 298308
rect 655060 298120 655112 298172
rect 675392 298120 675444 298172
rect 674656 295400 674708 295452
rect 675300 295400 675352 295452
rect 42340 295332 42392 295384
rect 58532 295332 58584 295384
rect 674564 295196 674616 295248
rect 675392 295196 675444 295248
rect 674472 294108 674524 294160
rect 675300 294108 675352 294160
rect 674564 293904 674616 293956
rect 675116 293904 675168 293956
rect 43352 292544 43404 292596
rect 58348 292544 58400 292596
rect 41788 291864 41840 291916
rect 43444 291864 43496 291916
rect 674840 291252 674892 291304
rect 675116 291048 675168 291100
rect 674288 290436 674340 290488
rect 675116 290436 675168 290488
rect 41788 289824 41840 289876
rect 42708 289824 42760 289876
rect 54024 289756 54076 289808
rect 58532 289756 58584 289808
rect 654140 289076 654192 289128
rect 667020 289076 667072 289128
rect 30012 288804 30064 288856
rect 673552 288600 673604 288652
rect 675392 288600 675444 288652
rect 42248 288396 42300 288448
rect 673828 287376 673880 287428
rect 675116 287376 675168 287428
rect 656808 287240 656860 287292
rect 666836 287240 666888 287292
rect 56508 287104 56560 287156
rect 57980 287104 58032 287156
rect 46112 287036 46164 287088
rect 58532 287036 58584 287088
rect 654140 287036 654192 287088
rect 670240 287036 670292 287088
rect 673460 286764 673512 286816
rect 675116 286764 675168 286816
rect 673644 286696 673696 286748
rect 675208 286696 675260 286748
rect 673460 286628 673512 286680
rect 674564 286628 674616 286680
rect 673736 286560 673788 286612
rect 675392 286560 675444 286612
rect 43076 285608 43128 285660
rect 43720 285608 43772 285660
rect 42432 285472 42484 285524
rect 43076 285472 43128 285524
rect 53932 285132 53984 285184
rect 57980 285132 58032 285184
rect 655244 284928 655296 284980
rect 670332 284928 670384 284980
rect 654508 284656 654560 284708
rect 666744 284656 666796 284708
rect 51080 284316 51132 284368
rect 58532 284316 58584 284368
rect 43996 284248 44048 284300
rect 44272 284248 44324 284300
rect 41880 283772 41932 283824
rect 41880 283568 41932 283620
rect 654232 283160 654284 283212
rect 669964 283160 670016 283212
rect 673460 282820 673512 282872
rect 675116 282820 675168 282872
rect 42156 281732 42208 281784
rect 43628 281732 43680 281784
rect 43628 281596 43680 281648
rect 44272 281596 44324 281648
rect 48504 281528 48556 281580
rect 57980 281528 58032 281580
rect 655244 281528 655296 281580
rect 670056 281528 670108 281580
rect 42156 281052 42208 281104
rect 42340 281052 42392 281104
rect 42340 280440 42392 280492
rect 43444 280440 43496 280492
rect 654140 280372 654192 280424
rect 670148 280372 670200 280424
rect 42156 279828 42208 279880
rect 43168 279828 43220 279880
rect 42156 279216 42208 279268
rect 43352 279216 43404 279268
rect 654876 278740 654928 278792
rect 666652 278740 666704 278792
rect 42064 278604 42116 278656
rect 42708 278604 42760 278656
rect 42708 278468 42760 278520
rect 43904 278468 43956 278520
rect 671620 278332 671672 278384
rect 678980 278332 679032 278384
rect 671712 278264 671764 278316
rect 679072 278264 679124 278316
rect 671804 278060 671856 278112
rect 679164 278060 679216 278112
rect 48320 277584 48372 277636
rect 648620 277584 648672 277636
rect 48412 277516 48464 277568
rect 654140 277516 654192 277568
rect 48228 277380 48280 277432
rect 666560 277380 666612 277432
rect 42340 276768 42392 276820
rect 43812 276768 43864 276820
rect 42248 276700 42300 276752
rect 43076 276700 43128 276752
rect 42064 276564 42116 276616
rect 43536 276564 43588 276616
rect 387248 276020 387300 276072
rect 405096 276020 405148 276072
rect 347780 275952 347832 276004
rect 478328 275952 478380 276004
rect 350172 275884 350224 275936
rect 485504 275884 485556 275936
rect 353208 275816 353260 275868
rect 492588 275816 492640 275868
rect 355784 275748 355836 275800
rect 499672 275748 499724 275800
rect 358544 275680 358596 275732
rect 506756 275680 506808 275732
rect 361488 275612 361540 275664
rect 513840 275612 513892 275664
rect 42432 275544 42484 275596
rect 42708 275544 42760 275596
rect 363972 275544 364024 275596
rect 520924 275544 520976 275596
rect 366456 275476 366508 275528
rect 528008 275476 528060 275528
rect 369124 275408 369176 275460
rect 535092 275408 535144 275460
rect 371792 275340 371844 275392
rect 542176 275340 542228 275392
rect 375288 275272 375340 275324
rect 550456 275272 550508 275324
rect 377956 275204 378008 275256
rect 557540 275204 557592 275256
rect 380348 275136 380400 275188
rect 564624 275136 564676 275188
rect 382924 275068 382976 275120
rect 571708 275068 571760 275120
rect 385592 275000 385644 275052
rect 578884 275000 578936 275052
rect 401600 274932 401652 274984
rect 585968 274932 586020 274984
rect 320272 274864 320324 274916
rect 387248 274864 387300 274916
rect 405372 274864 405424 274916
rect 627276 274864 627328 274916
rect 319904 274728 319956 274780
rect 401692 274796 401744 274848
rect 593052 274796 593104 274848
rect 403900 274728 403952 274780
rect 404268 274728 404320 274780
rect 628472 274728 628524 274780
rect 321008 274660 321060 274712
rect 407488 274660 407540 274712
rect 409236 274660 409288 274712
rect 322756 274592 322808 274644
rect 410984 274592 411036 274644
rect 429108 274660 429160 274712
rect 634360 274660 634412 274712
rect 641444 274592 641496 274644
rect 343732 274524 343784 274576
rect 467748 274524 467800 274576
rect 345112 274456 345164 274508
rect 471244 274456 471296 274508
rect 342536 274388 342588 274440
rect 464160 274388 464212 274440
rect 339776 274320 339828 274372
rect 457076 274320 457128 274372
rect 42156 274252 42208 274304
rect 44088 274252 44140 274304
rect 337108 274252 337160 274304
rect 449992 274252 450044 274304
rect 335728 274184 335780 274236
rect 446496 274184 446548 274236
rect 334348 274116 334400 274168
rect 442908 274116 442960 274168
rect 333428 274048 333480 274100
rect 439320 274048 439372 274100
rect 331680 273980 331732 274032
rect 435824 273980 435876 274032
rect 330760 273912 330812 273964
rect 432236 273912 432288 273964
rect 329012 273844 329064 273896
rect 428740 273844 428792 273896
rect 327724 273776 327776 273828
rect 425152 273776 425204 273828
rect 325516 273708 325568 273760
rect 418068 273708 418120 273760
rect 326344 273640 326396 273692
rect 421656 273640 421708 273692
rect 323676 273572 323728 273624
rect 414572 273572 414624 273624
rect 42064 273504 42116 273556
rect 43628 273504 43680 273556
rect 388260 273504 388312 273556
rect 401600 273504 401652 273556
rect 406568 273436 406620 273488
rect 429108 273504 429160 273556
rect 391020 273232 391072 273284
rect 401692 273232 401744 273284
rect 154488 273164 154540 273216
rect 225328 273164 225380 273216
rect 263232 273164 263284 273216
rect 266728 273164 266780 273216
rect 291200 273164 291252 273216
rect 328276 273164 328328 273216
rect 345480 273164 345532 273216
rect 472440 273164 472492 273216
rect 472532 273164 472584 273216
rect 610716 273164 610768 273216
rect 156880 273096 156932 273148
rect 208308 273096 208360 273148
rect 260932 273096 260984 273148
rect 265808 273096 265860 273148
rect 292120 273096 292172 273148
rect 330576 273096 330628 273148
rect 356244 273096 356296 273148
rect 500868 273096 500920 273148
rect 149796 273028 149848 273080
rect 224408 273028 224460 273080
rect 243176 273028 243228 273080
rect 259184 273028 259236 273080
rect 259736 273028 259788 273080
rect 265348 273028 265400 273080
rect 293868 273028 293920 273080
rect 335360 273028 335412 273080
rect 342812 273028 342864 273080
rect 465356 273028 465408 273080
rect 467748 273028 467800 273080
rect 617800 273028 617852 273080
rect 143908 272960 143960 273012
rect 221280 272960 221332 273012
rect 241980 272960 242032 273012
rect 258724 272960 258776 273012
rect 296076 272960 296128 273012
rect 341248 272960 341300 273012
rect 347872 272960 347924 273012
rect 351920 272960 351972 273012
rect 361580 272960 361632 273012
rect 515036 272960 515088 273012
rect 148600 272892 148652 272944
rect 223212 272892 223264 272944
rect 236092 272892 236144 272944
rect 256424 272892 256476 272944
rect 294880 272892 294932 272944
rect 337752 272892 337804 272944
rect 350080 272892 350132 272944
rect 484308 272892 484360 272944
rect 485044 272892 485096 272944
rect 635556 272892 635608 272944
rect 145104 272824 145156 272876
rect 222200 272824 222252 272876
rect 234896 272824 234948 272876
rect 256056 272824 256108 272876
rect 301412 272824 301464 272876
rect 355416 272824 355468 272876
rect 372804 272824 372856 272876
rect 381452 272824 381504 272876
rect 383660 272824 383712 272876
rect 388536 272824 388588 272876
rect 390468 272824 390520 272876
rect 526812 272824 526864 272876
rect 146208 272756 146260 272808
rect 223028 272756 223080 272808
rect 238484 272756 238536 272808
rect 257436 272756 257488 272808
rect 301872 272756 301924 272808
rect 356612 272756 356664 272808
rect 363880 272756 363932 272808
rect 519728 272756 519780 272808
rect 139124 272688 139176 272740
rect 220360 272688 220412 272740
rect 239588 272688 239640 272740
rect 257804 272688 257856 272740
rect 295248 272688 295300 272740
rect 338856 272688 338908 272740
rect 339408 272688 339460 272740
rect 455880 272688 455932 272740
rect 455972 272688 456024 272740
rect 624976 272688 625028 272740
rect 137928 272620 137980 272672
rect 219440 272620 219492 272672
rect 232504 272620 232556 272672
rect 255136 272620 255188 272672
rect 304080 272620 304132 272672
rect 362500 272620 362552 272672
rect 375380 272620 375432 272672
rect 551652 272620 551704 272672
rect 136824 272552 136876 272604
rect 218612 272552 218664 272604
rect 237288 272552 237340 272604
rect 257252 272552 257304 272604
rect 304540 272552 304592 272604
rect 363696 272552 363748 272604
rect 378048 272552 378100 272604
rect 558736 272552 558788 272604
rect 130844 272484 130896 272536
rect 216864 272484 216916 272536
rect 233700 272484 233752 272536
rect 255596 272484 255648 272536
rect 288164 272484 288216 272536
rect 319996 272484 320048 272536
rect 320088 272484 320140 272536
rect 377864 272484 377916 272536
rect 132040 272416 132092 272468
rect 217692 272416 217744 272468
rect 227812 272416 227864 272468
rect 253388 272416 253440 272468
rect 293408 272416 293460 272468
rect 334164 272416 334216 272468
rect 334256 272416 334308 272468
rect 391572 272484 391624 272536
rect 572904 272484 572956 272536
rect 441712 272416 441764 272468
rect 441804 272416 441856 272468
rect 632060 272416 632112 272468
rect 129648 272348 129700 272400
rect 215668 272348 215720 272400
rect 231308 272348 231360 272400
rect 254676 272348 254728 272400
rect 307208 272348 307260 272400
rect 370780 272348 370832 272400
rect 372068 272348 372120 272400
rect 390468 272348 390520 272400
rect 391204 272348 391256 272400
rect 579988 272348 580040 272400
rect 124956 272280 125008 272332
rect 215024 272280 215076 272332
rect 229008 272280 229060 272332
rect 253756 272280 253808 272332
rect 287612 272280 287664 272332
rect 318800 272280 318852 272332
rect 318892 272280 318944 272332
rect 384948 272280 385000 272332
rect 390008 272280 390060 272332
rect 123760 272212 123812 272264
rect 214196 272212 214248 272264
rect 230204 272212 230256 272264
rect 254216 272212 254268 272264
rect 288900 272212 288952 272264
rect 321192 272212 321244 272264
rect 325332 272212 325384 272264
rect 390928 272212 390980 272264
rect 391112 272280 391164 272332
rect 587072 272280 587124 272332
rect 590660 272212 590712 272264
rect 104900 272144 104952 272196
rect 206284 272144 206336 272196
rect 226616 272144 226668 272196
rect 252928 272144 252980 272196
rect 286692 272144 286744 272196
rect 315212 272144 315264 272196
rect 315304 272144 315356 272196
rect 392124 272144 392176 272196
rect 394056 272144 394108 272196
rect 601332 272144 601384 272196
rect 97816 272076 97868 272128
rect 203892 272076 203944 272128
rect 205364 272076 205416 272128
rect 244924 272076 244976 272128
rect 91836 272008 91888 272060
rect 195980 272008 196032 272060
rect 201776 272008 201828 272060
rect 240140 272008 240192 272060
rect 89536 271940 89588 271992
rect 200764 271940 200816 271992
rect 208308 271940 208360 271992
rect 227076 271940 227128 271992
rect 240784 271940 240836 271992
rect 258264 272076 258316 272128
rect 292580 272076 292632 272128
rect 331772 272076 331824 272128
rect 331864 272076 331916 272128
rect 434628 272076 434680 272128
rect 435732 272076 435784 272128
rect 642640 272076 642692 272128
rect 82452 271872 82504 271924
rect 198556 271872 198608 271924
rect 245568 271872 245620 271924
rect 260012 272008 260064 272060
rect 287152 272008 287204 272060
rect 317604 272008 317656 272060
rect 317880 272008 317932 272060
rect 399208 272008 399260 272060
rect 399576 272008 399628 272060
rect 611912 272008 611964 272060
rect 262128 271940 262180 271992
rect 266268 271940 266320 271992
rect 286968 271940 287020 271992
rect 316408 271940 316460 271992
rect 318800 271940 318852 271992
rect 401508 271940 401560 271992
rect 407396 271940 407448 271992
rect 65892 271804 65944 271856
rect 176844 271804 176896 271856
rect 194692 271804 194744 271856
rect 240876 271804 240928 271856
rect 244372 271804 244424 271856
rect 259552 271872 259604 271924
rect 289544 271872 289596 271924
rect 322388 271872 322440 271924
rect 246764 271804 246816 271856
rect 260472 271804 260524 271856
rect 264428 271804 264480 271856
rect 267188 271804 267240 271856
rect 289636 271804 289688 271856
rect 155684 271736 155736 271788
rect 225880 271736 225932 271788
rect 249064 271736 249116 271788
rect 261392 271736 261444 271788
rect 291660 271736 291712 271788
rect 313372 271736 313424 271788
rect 161572 271668 161624 271720
rect 227996 271668 228048 271720
rect 251456 271668 251508 271720
rect 262220 271668 262272 271720
rect 285404 271668 285456 271720
rect 312912 271668 312964 271720
rect 163964 271600 164016 271652
rect 229744 271600 229796 271652
rect 253848 271600 253900 271652
rect 263140 271600 263192 271652
rect 290740 271600 290792 271652
rect 313280 271600 313332 271652
rect 313556 271804 313608 271856
rect 320548 271804 320600 271856
rect 406292 271872 406344 271924
rect 411444 271872 411496 271924
rect 413652 271940 413704 271992
rect 622584 271940 622636 271992
rect 323216 271804 323268 271856
rect 413376 271804 413428 271856
rect 636752 271872 636804 271924
rect 647424 271804 647476 271856
rect 329472 271736 329524 271788
rect 353576 271736 353628 271788
rect 493692 271736 493744 271788
rect 498660 271736 498712 271788
rect 603632 271736 603684 271788
rect 313556 271668 313608 271720
rect 349528 271668 349580 271720
rect 350908 271668 350960 271720
rect 486608 271668 486660 271720
rect 323492 271600 323544 271652
rect 348240 271600 348292 271652
rect 479524 271600 479576 271652
rect 162768 271532 162820 271584
rect 228824 271532 228876 271584
rect 257344 271532 257396 271584
rect 264520 271532 264572 271584
rect 289820 271532 289872 271584
rect 324688 271532 324740 271584
rect 347596 271532 347648 271584
rect 477224 271532 477276 271584
rect 171048 271464 171100 271516
rect 232412 271464 232464 271516
rect 258540 271464 258592 271516
rect 264888 271464 264940 271516
rect 266820 271464 266872 271516
rect 268016 271464 268068 271516
rect 290280 271464 290332 271516
rect 134432 271396 134484 271448
rect 195796 271396 195848 271448
rect 197084 271396 197136 271448
rect 241796 271396 241848 271448
rect 254952 271396 255004 271448
rect 263600 271396 263652 271448
rect 285864 271396 285916 271448
rect 168748 271328 168800 271380
rect 230664 271328 230716 271380
rect 252652 271328 252704 271380
rect 262864 271328 262916 271380
rect 284208 271328 284260 271380
rect 309324 271328 309376 271380
rect 169852 271260 169904 271312
rect 231492 271260 231544 271312
rect 250260 271260 250312 271312
rect 261852 271260 261904 271312
rect 313280 271464 313332 271516
rect 327080 271464 327132 271516
rect 314660 271396 314712 271448
rect 344836 271464 344888 271516
rect 344928 271464 344980 271516
rect 470140 271464 470192 271516
rect 342168 271396 342220 271448
rect 462964 271396 463016 271448
rect 325884 271328 325936 271380
rect 340144 271328 340196 271380
rect 458272 271328 458324 271380
rect 314108 271260 314160 271312
rect 336464 271260 336516 271312
rect 448796 271260 448848 271312
rect 176844 271192 176896 271244
rect 192116 271192 192168 271244
rect 178132 271124 178184 271176
rect 197360 271192 197412 271244
rect 233332 271192 233384 271244
rect 337476 271192 337528 271244
rect 451188 271192 451240 271244
rect 231860 271124 231912 271176
rect 334808 271124 334860 271176
rect 444104 271124 444156 271176
rect 175832 271056 175884 271108
rect 197176 271056 197228 271108
rect 197268 271056 197320 271108
rect 234160 271056 234212 271108
rect 247868 271056 247920 271108
rect 260932 271056 260984 271108
rect 332140 271056 332192 271108
rect 437020 271056 437072 271108
rect 182916 270988 182968 271040
rect 236000 270988 236052 271040
rect 332416 270988 332468 271040
rect 429936 270988 429988 271040
rect 187608 270920 187660 270972
rect 238208 270920 238260 270972
rect 328644 270920 328696 270972
rect 427544 270920 427596 270972
rect 186412 270852 186464 270904
rect 237288 270852 237340 270904
rect 325976 270852 326028 270904
rect 420460 270852 420512 270904
rect 142712 270784 142764 270836
rect 146208 270784 146260 270836
rect 188804 270784 188856 270836
rect 239128 270784 239180 270836
rect 324136 270784 324188 270836
rect 415768 270784 415820 270836
rect 176936 270716 176988 270768
rect 197268 270716 197320 270768
rect 133236 270512 133288 270564
rect 191196 270512 191248 270564
rect 234620 270716 234672 270768
rect 327172 270716 327224 270768
rect 383844 270716 383896 270768
rect 386236 270716 386288 270768
rect 391204 270716 391256 270768
rect 402060 270716 402112 270768
rect 413652 270716 413704 270768
rect 199568 270648 199620 270700
rect 242624 270648 242676 270700
rect 256148 270648 256200 270700
rect 264060 270648 264112 270700
rect 320180 270648 320232 270700
rect 374368 270648 374420 270700
rect 383476 270648 383528 270700
rect 391572 270648 391624 270700
rect 198280 270580 198332 270632
rect 242256 270580 242308 270632
rect 327540 270580 327592 270632
rect 376760 270580 376812 270632
rect 388996 270580 389048 270632
rect 391112 270580 391164 270632
rect 312544 270512 312596 270564
rect 342444 270512 342496 270564
rect 147404 270444 147456 270496
rect 208124 270444 208176 270496
rect 141516 270376 141568 270428
rect 220820 270444 220872 270496
rect 225420 270444 225472 270496
rect 252468 270444 252520 270496
rect 265624 270444 265676 270496
rect 267556 270444 267608 270496
rect 269396 270444 269448 270496
rect 270316 270444 270368 270496
rect 271144 270444 271196 270496
rect 275100 270444 275152 270496
rect 276940 270444 276992 270496
rect 290464 270444 290516 270496
rect 295616 270444 295668 270496
rect 340052 270444 340104 270496
rect 140320 270308 140372 270360
rect 219992 270376 220044 270428
rect 224224 270376 224276 270428
rect 252008 270376 252060 270428
rect 269856 270376 269908 270428
rect 271512 270376 271564 270428
rect 271604 270376 271656 270428
rect 276204 270376 276256 270428
rect 277492 270376 277544 270428
rect 207848 270240 207900 270292
rect 207940 270240 207992 270292
rect 215484 270240 215536 270292
rect 135628 270172 135680 270224
rect 219072 270308 219124 270360
rect 221924 270308 221976 270360
rect 251088 270308 251140 270360
rect 272064 270308 272116 270360
rect 277400 270308 277452 270360
rect 277860 270308 277912 270360
rect 296996 270376 297048 270428
rect 343640 270376 343692 270428
rect 218336 270240 218388 270292
rect 249800 270240 249852 270292
rect 220728 270172 220780 270224
rect 250720 270172 250772 270224
rect 270684 270172 270736 270224
rect 273904 270172 273956 270224
rect 278688 270172 278740 270224
rect 291568 270308 291620 270360
rect 298284 270308 298336 270360
rect 347136 270512 347188 270564
rect 346032 270444 346084 270496
rect 473636 270444 473688 270496
rect 346860 270376 346912 270428
rect 476028 270376 476080 270428
rect 348608 270308 348660 270360
rect 480720 270308 480772 270360
rect 297916 270240 297968 270292
rect 345940 270240 345992 270292
rect 349528 270240 349580 270292
rect 483112 270240 483164 270292
rect 126152 270104 126204 270156
rect 213460 270104 213512 270156
rect 213644 270104 213696 270156
rect 248052 270104 248104 270156
rect 272984 270104 273036 270156
rect 279792 270104 279844 270156
rect 292764 270172 292816 270224
rect 300124 270172 300176 270224
rect 347872 270172 347924 270224
rect 351276 270172 351328 270224
rect 487804 270172 487856 270224
rect 295156 270104 295208 270156
rect 298744 270104 298796 270156
rect 348332 270104 348384 270156
rect 359372 270104 359424 270156
rect 509056 270104 509108 270156
rect 127348 270036 127400 270088
rect 207940 270036 207992 270088
rect 208124 270036 208176 270088
rect 222660 270036 222712 270088
rect 223120 270036 223172 270088
rect 251548 270036 251600 270088
rect 273720 270036 273772 270088
rect 280988 270036 281040 270088
rect 281080 270036 281132 270088
rect 293960 270036 294012 270088
rect 300584 270036 300636 270088
rect 353116 270036 353168 270088
rect 360200 270036 360252 270088
rect 511448 270036 511500 270088
rect 121460 269968 121512 270020
rect 213736 269968 213788 270020
rect 215944 269968 215996 270020
rect 248880 269968 248932 270020
rect 272524 269968 272576 270020
rect 278596 269968 278648 270020
rect 279148 269968 279200 270020
rect 296352 269968 296404 270020
rect 303252 269968 303304 270020
rect 359924 269968 359976 270020
rect 364708 269968 364760 270020
rect 523316 269968 523368 270020
rect 119068 269900 119120 269952
rect 211896 269900 211948 269952
rect 217140 269900 217192 269952
rect 249340 269900 249392 269952
rect 279608 269900 279660 269952
rect 297548 269900 297600 269952
rect 302792 269900 302844 269952
rect 359004 269900 359056 269952
rect 367376 269900 367428 269952
rect 530400 269900 530452 269952
rect 114376 269832 114428 269884
rect 211068 269832 211120 269884
rect 212448 269832 212500 269884
rect 247592 269832 247644 269884
rect 280068 269832 280120 269884
rect 298468 269832 298520 269884
rect 305460 269832 305512 269884
rect 366088 269832 366140 269884
rect 368204 269832 368256 269884
rect 532700 269832 532752 269884
rect 113180 269764 113232 269816
rect 210148 269764 210200 269816
rect 214840 269764 214892 269816
rect 248420 269764 248472 269816
rect 280528 269764 280580 269816
rect 299848 269764 299900 269816
rect 306748 269764 306800 269816
rect 369584 269764 369636 269816
rect 372712 269764 372764 269816
rect 544568 269764 544620 269816
rect 109592 269696 109644 269748
rect 208860 269696 208912 269748
rect 211252 269696 211304 269748
rect 247132 269696 247184 269748
rect 278320 269696 278372 269748
rect 281080 269696 281132 269748
rect 108396 269628 108448 269680
rect 207940 269628 207992 269680
rect 208032 269628 208084 269680
rect 245752 269628 245804 269680
rect 274732 269628 274784 269680
rect 284484 269696 284536 269748
rect 305920 269696 305972 269748
rect 367284 269696 367336 269748
rect 374000 269696 374052 269748
rect 548064 269696 548116 269748
rect 281816 269628 281868 269680
rect 303436 269628 303488 269680
rect 308220 269628 308272 269680
rect 373172 269628 373224 269680
rect 379336 269628 379388 269680
rect 562324 269628 562376 269680
rect 102508 269560 102560 269612
rect 206192 269560 206244 269612
rect 210056 269560 210108 269612
rect 246672 269560 246724 269612
rect 281448 269560 281500 269612
rect 302240 269560 302292 269612
rect 310796 269560 310848 269612
rect 380256 269560 380308 269612
rect 384672 269560 384724 269612
rect 576492 269560 576544 269612
rect 94228 269492 94280 269544
rect 202604 269492 202656 269544
rect 209136 269492 209188 269544
rect 246212 269492 246264 269544
rect 280988 269492 281040 269544
rect 301044 269492 301096 269544
rect 313464 269492 313516 269544
rect 386972 269492 387024 269544
rect 387340 269492 387392 269544
rect 583576 269492 583628 269544
rect 95424 269424 95476 269476
rect 203524 269424 203576 269476
rect 206560 269424 206612 269476
rect 245292 269424 245344 269476
rect 282736 269424 282788 269476
rect 305828 269424 305880 269476
rect 316132 269424 316184 269476
rect 42432 269356 42484 269408
rect 43260 269356 43312 269408
rect 87144 269356 87196 269408
rect 200396 269356 200448 269408
rect 202972 269356 203024 269408
rect 244004 269356 244056 269408
rect 282276 269356 282328 269408
rect 304632 269356 304684 269408
rect 316592 269356 316644 269408
rect 392768 269424 392820 269476
rect 597744 269424 597796 269476
rect 75368 269288 75420 269340
rect 195428 269288 195480 269340
rect 204168 269288 204220 269340
rect 244464 269288 244516 269340
rect 283656 269288 283708 269340
rect 308128 269288 308180 269340
rect 317512 269288 317564 269340
rect 387432 269288 387484 269340
rect 394424 269356 394476 269408
rect 396724 269356 396776 269408
rect 608416 269356 608468 269408
rect 395620 269288 395672 269340
rect 399392 269288 399444 269340
rect 615500 269288 615552 269340
rect 72976 269220 73028 269272
rect 195060 269220 195112 269272
rect 200580 269220 200632 269272
rect 243084 269220 243136 269272
rect 283196 269220 283248 269272
rect 307024 269220 307076 269272
rect 319260 269220 319312 269272
rect 195888 269152 195940 269204
rect 241336 269152 241388 269204
rect 284944 269152 284996 269204
rect 311716 269152 311768 269204
rect 321928 269152 321980 269204
rect 397184 269152 397236 269204
rect 400772 269220 400824 269272
rect 618996 269220 619048 269272
rect 402704 269152 402756 269204
rect 408776 269152 408828 269204
rect 640340 269152 640392 269204
rect 67088 269084 67140 269136
rect 192760 269084 192812 269136
rect 193496 269084 193548 269136
rect 240416 269084 240468 269136
rect 270316 269084 270368 269136
rect 272708 269084 272760 269136
rect 284484 269084 284536 269136
rect 310520 269084 310572 269136
rect 322848 269084 322900 269136
rect 401600 269084 401652 269136
rect 403900 269084 403952 269136
rect 405372 269084 405424 269136
rect 411904 269084 411956 269136
rect 648712 269084 648764 269136
rect 153384 269016 153436 269068
rect 225788 269016 225840 269068
rect 234620 269016 234672 269068
rect 239588 269016 239640 269068
rect 294328 269016 294380 269068
rect 336556 269016 336608 269068
rect 343272 269016 343324 269068
rect 466552 269016 466604 269068
rect 152188 268948 152240 269000
rect 224868 268948 224920 269000
rect 292948 268948 293000 269000
rect 332968 268948 333020 269000
rect 344192 268948 344244 269000
rect 468944 268948 468996 269000
rect 165160 268880 165212 268932
rect 229284 268880 229336 268932
rect 297456 268880 297508 268932
rect 314660 268880 314712 268932
rect 341524 268880 341576 268932
rect 461860 268880 461912 268932
rect 160468 268812 160520 268864
rect 228456 268812 228508 268864
rect 340604 268812 340656 268864
rect 459468 268812 459520 268864
rect 167552 268744 167604 268796
rect 231124 268744 231176 268796
rect 296536 268744 296588 268796
rect 312544 268744 312596 268796
rect 338856 268744 338908 268796
rect 454684 268744 454736 268796
rect 166356 268676 166408 268728
rect 230204 268676 230256 268728
rect 273812 268676 273864 268728
rect 282184 268676 282236 268728
rect 309876 268676 309928 268728
rect 320088 268676 320140 268728
rect 337936 268676 337988 268728
rect 452384 268676 452436 268728
rect 172244 268608 172296 268660
rect 231952 268608 232004 268660
rect 274272 268608 274324 268660
rect 283380 268608 283432 268660
rect 299204 268608 299256 268660
rect 313556 268608 313608 268660
rect 336188 268608 336240 268660
rect 447600 268608 447652 268660
rect 173440 268540 173492 268592
rect 232872 268540 232924 268592
rect 312544 268540 312596 268592
rect 318892 268540 318944 268592
rect 335268 268540 335320 268592
rect 445300 268540 445352 268592
rect 174636 268472 174688 268524
rect 233792 268472 233844 268524
rect 240140 268472 240192 268524
rect 243544 268472 243596 268524
rect 331312 268472 331364 268524
rect 331864 268472 331916 268524
rect 333520 268472 333572 268524
rect 440516 268472 440568 268524
rect 179328 268404 179380 268456
rect 234620 268404 234672 268456
rect 332600 268404 332652 268456
rect 438216 268404 438268 268456
rect 181720 268336 181772 268388
rect 236460 268336 236512 268388
rect 330852 268336 330904 268388
rect 433432 268336 433484 268388
rect 180524 268268 180576 268320
rect 235540 268268 235592 268320
rect 275192 268268 275244 268320
rect 285680 268268 285732 268320
rect 329932 268268 329984 268320
rect 431132 268268 431184 268320
rect 184112 268200 184164 268252
rect 236920 268200 236972 268252
rect 275652 268200 275704 268252
rect 286876 268200 286928 268252
rect 309416 268200 309468 268252
rect 327540 268200 327592 268252
rect 328184 268200 328236 268252
rect 426348 268200 426400 268252
rect 185216 268132 185268 268184
rect 237748 268132 237800 268184
rect 312084 268132 312136 268184
rect 327172 268132 327224 268184
rect 327264 268132 327316 268184
rect 423956 268132 424008 268184
rect 190000 268064 190052 268116
rect 238668 268064 238720 268116
rect 313924 268064 313976 268116
rect 192392 267996 192444 268048
rect 239956 267996 240008 268048
rect 314844 267996 314896 268048
rect 325332 267996 325384 268048
rect 329472 267996 329524 268048
rect 332416 267996 332468 268048
rect 332692 268064 332744 268116
rect 383660 267996 383712 268048
rect 387432 267996 387484 268048
rect 398012 267996 398064 268048
rect 401600 268064 401652 268116
rect 412180 268064 412232 268116
rect 656164 268064 656216 268116
rect 676220 268064 676272 268116
rect 416872 267996 416924 268048
rect 195796 267928 195848 267980
rect 218152 267928 218204 267980
rect 219532 267928 219584 267980
rect 250260 267928 250312 267980
rect 276480 267928 276532 267980
rect 289268 267928 289320 267980
rect 311256 267928 311308 267980
rect 74172 267860 74224 267912
rect 195888 267860 195940 267912
rect 207848 267860 207900 267912
rect 217324 267860 217376 267912
rect 231860 267860 231912 267912
rect 235080 267860 235132 267912
rect 276296 267860 276348 267912
rect 288072 267860 288124 267912
rect 324596 267860 324648 267912
rect 332692 267860 332744 267912
rect 371332 267928 371384 267980
rect 372528 267928 372580 267980
rect 397184 267928 397236 267980
rect 409788 267928 409840 267980
rect 655980 267928 656032 267980
rect 676036 267928 676088 267980
rect 372804 267860 372856 267912
rect 308588 267792 308640 267844
rect 320180 267792 320232 267844
rect 213460 267724 213512 267776
rect 214656 267724 214708 267776
rect 398104 267724 398156 267776
rect 399576 267724 399628 267776
rect 655796 267724 655848 267776
rect 676128 267724 676180 267776
rect 367744 267656 367796 267708
rect 531596 267656 531648 267708
rect 370504 267588 370556 267640
rect 538680 267588 538732 267640
rect 373172 267520 373224 267572
rect 545764 267520 545816 267572
rect 373540 267452 373592 267504
rect 546960 267452 547012 267504
rect 374460 267384 374512 267436
rect 549260 267384 549312 267436
rect 376208 267316 376260 267368
rect 554044 267316 554096 267368
rect 375840 267248 375892 267300
rect 552848 267248 552900 267300
rect 377128 267180 377180 267232
rect 556344 267180 556396 267232
rect 299664 267112 299716 267164
rect 350724 267112 350776 267164
rect 378508 267112 378560 267164
rect 559932 267112 559984 267164
rect 300952 267044 301004 267096
rect 354220 267044 354272 267096
rect 378876 267044 378928 267096
rect 561128 267044 561180 267096
rect 302332 266976 302384 267028
rect 357808 266976 357860 267028
rect 379796 266976 379848 267028
rect 563428 266976 563480 267028
rect 303712 266908 303764 266960
rect 361396 266908 361448 266960
rect 381636 266908 381688 266960
rect 568212 266908 568264 266960
rect 305000 266840 305052 266892
rect 364892 266840 364944 266892
rect 381176 266840 381228 266892
rect 567016 266840 567068 266892
rect 306380 266772 306432 266824
rect 368480 266772 368532 266824
rect 382464 266772 382516 266824
rect 570604 266772 570656 266824
rect 307668 266704 307720 266756
rect 371976 266704 372028 266756
rect 384304 266704 384356 266756
rect 575296 266704 575348 266756
rect 309048 266636 309100 266688
rect 375564 266636 375616 266688
rect 383844 266636 383896 266688
rect 574100 266636 574152 266688
rect 673368 266636 673420 266688
rect 676036 266636 676088 266688
rect 310336 266568 310388 266620
rect 379060 266568 379112 266620
rect 385132 266568 385184 266620
rect 577688 266568 577740 266620
rect 311716 266500 311768 266552
rect 382648 266500 382700 266552
rect 386512 266500 386564 266552
rect 581184 266500 581236 266552
rect 313004 266432 313056 266484
rect 386144 266432 386196 266484
rect 387800 266432 387852 266484
rect 584772 266432 584824 266484
rect 116676 266364 116728 266416
rect 211528 266364 211580 266416
rect 389180 266364 389232 266416
rect 588268 266364 588320 266416
rect 68192 266296 68244 266348
rect 193220 266296 193272 266348
rect 315672 266296 315724 266348
rect 392216 266296 392268 266348
rect 392308 266296 392360 266348
rect 596548 266296 596600 266348
rect 365076 266228 365128 266280
rect 524512 266228 524564 266280
rect 362408 266160 362460 266212
rect 517336 266160 517388 266212
rect 359740 266092 359792 266144
rect 510252 266092 510304 266144
rect 357072 266024 357124 266076
rect 503168 266024 503220 266076
rect 354404 265956 354456 266008
rect 496084 265956 496136 266008
rect 351736 265888 351788 265940
rect 489000 265888 489052 265940
rect 349068 265820 349120 265872
rect 481916 265820 481968 265872
rect 346400 265752 346452 265804
rect 474832 265752 474884 265804
rect 341064 265684 341116 265736
rect 460664 265684 460716 265736
rect 338396 265616 338448 265668
rect 453580 265616 453632 265668
rect 317052 265548 317104 265600
rect 394700 265548 394752 265600
rect 394976 265548 395028 265600
rect 498660 265548 498712 265600
rect 675208 265548 675260 265600
rect 676036 265548 676088 265600
rect 326804 265480 326856 265532
rect 422852 265480 422904 265532
rect 325608 265412 325660 265464
rect 419264 265412 419316 265464
rect 321468 265344 321520 265396
rect 314384 265276 314436 265328
rect 389732 265276 389784 265328
rect 394700 265344 394752 265396
rect 396816 265344 396868 265396
rect 408592 265344 408644 265396
rect 409604 265344 409656 265396
rect 435732 265344 435784 265396
rect 400312 265276 400364 265328
rect 467748 265276 467800 265328
rect 318340 265208 318392 265260
rect 400220 265208 400272 265260
rect 42156 264732 42208 264784
rect 59452 264732 59504 264784
rect 673828 263032 673880 263084
rect 676036 263032 676088 263084
rect 673460 262488 673512 262540
rect 676128 262488 676180 262540
rect 673552 262284 673604 262336
rect 676128 262284 676180 262336
rect 674472 262216 674524 262268
rect 676036 262216 676088 262268
rect 674932 261808 674984 261860
rect 676036 261808 676088 261860
rect 673644 260176 673696 260228
rect 675668 260176 675720 260228
rect 673736 259700 673788 259752
rect 675668 259700 675720 259752
rect 674748 259632 674800 259684
rect 676128 259632 676180 259684
rect 674656 259564 674708 259616
rect 675944 259564 675996 259616
rect 674840 259496 674892 259548
rect 676128 259496 676180 259548
rect 675024 259428 675076 259480
rect 676036 259428 676088 259480
rect 674288 258952 674340 259004
rect 676036 258952 676088 259004
rect 41788 258068 41840 258120
rect 53932 258068 53984 258120
rect 41512 257932 41564 257984
rect 51080 257932 51132 257984
rect 41512 257524 41564 257576
rect 46112 257524 46164 257576
rect 672632 256776 672684 256828
rect 678980 256776 679032 256828
rect 52276 256708 52328 256760
rect 184940 256708 184992 256760
rect 674564 256708 674616 256760
rect 676036 256708 676088 256760
rect 673552 252696 673604 252748
rect 673552 252492 673604 252544
rect 673736 252288 673788 252340
rect 674288 252288 674340 252340
rect 674288 252152 674340 252204
rect 674564 252152 674616 252204
rect 674656 251880 674708 251932
rect 674840 251880 674892 251932
rect 675668 251336 675720 251388
rect 675760 251336 675812 251388
rect 416780 251200 416832 251252
rect 567108 251200 567160 251252
rect 674748 251200 674800 251252
rect 675300 251200 675352 251252
rect 675300 250928 675352 250980
rect 675760 250724 675812 250776
rect 675024 250180 675076 250232
rect 675484 250180 675536 250232
rect 675024 249772 675076 249824
rect 675300 249772 675352 249824
rect 674472 249636 674524 249688
rect 675300 249636 675352 249688
rect 673828 249568 673880 249620
rect 675392 249568 675444 249620
rect 673368 249500 673420 249552
rect 674472 249500 674524 249552
rect 416780 248412 416832 248464
rect 564348 248412 564400 248464
rect 41420 247664 41472 247716
rect 45652 247664 45704 247716
rect 674840 247256 674892 247308
rect 675392 247256 675444 247308
rect 674932 246984 674984 247036
rect 675208 246984 675260 247036
rect 41512 246916 41564 246968
rect 43352 246916 43404 246968
rect 674564 246508 674616 246560
rect 675392 246508 675444 246560
rect 674656 246032 674708 246084
rect 675392 246032 675444 246084
rect 20720 245828 20772 245880
rect 30104 245828 30156 245880
rect 52184 245760 52236 245812
rect 184940 245760 184992 245812
rect 41512 245692 41564 245744
rect 56692 245692 56744 245744
rect 41420 245624 41472 245676
rect 56600 245624 56652 245676
rect 416780 245624 416832 245676
rect 564532 245624 564584 245676
rect 43260 245556 43312 245608
rect 655612 245556 655664 245608
rect 675300 245556 675352 245608
rect 43444 245488 43496 245540
rect 38108 245420 38160 245472
rect 43260 245420 43312 245472
rect 674288 245420 674340 245472
rect 675300 245420 675352 245472
rect 38200 245352 38252 245404
rect 43076 245352 43128 245404
rect 43720 244808 43772 244860
rect 43904 244808 43956 244860
rect 43444 244672 43496 244724
rect 43720 244672 43772 244724
rect 42340 244536 42392 244588
rect 43444 244536 43496 244588
rect 20720 244332 20772 244384
rect 42248 244332 42300 244384
rect 673552 243584 673604 243636
rect 675392 243584 675444 243636
rect 673736 242904 673788 242956
rect 675392 242904 675444 242956
rect 673644 242156 673696 242208
rect 675392 242156 675444 242208
rect 673460 241068 673512 241120
rect 675300 241068 675352 241120
rect 674472 239912 674524 239964
rect 675300 239912 675352 239964
rect 42248 239708 42300 239760
rect 42708 239708 42760 239760
rect 42156 238484 42208 238536
rect 43812 238484 43864 238536
rect 42248 236036 42300 236088
rect 43076 236036 43128 236088
rect 42156 235356 42208 235408
rect 43352 235356 43404 235408
rect 42156 234608 42208 234660
rect 43168 234608 43220 234660
rect 42248 233520 42300 233572
rect 43260 233520 43312 233572
rect 42156 233316 42208 233368
rect 43536 233316 43588 233368
rect 52092 230796 52144 230848
rect 184940 237396 184992 237448
rect 674932 235560 674984 235612
rect 675760 235560 675812 235612
rect 674748 235492 674800 235544
rect 675668 235492 675720 235544
rect 345940 231140 345992 231192
rect 414020 231140 414072 231192
rect 355876 231072 355928 231124
rect 437296 231072 437348 231124
rect 347320 231004 347372 231056
rect 417148 231004 417200 231056
rect 356244 230936 356296 230988
rect 439780 230936 439832 230988
rect 348792 230868 348844 230920
rect 420460 230868 420512 230920
rect 351644 230800 351696 230852
rect 427176 230800 427228 230852
rect 354496 230732 354548 230784
rect 433892 230732 433944 230784
rect 45928 230664 45980 230716
rect 656900 230664 656952 230716
rect 46204 230596 46256 230648
rect 659752 230596 659804 230648
rect 42248 230528 42300 230580
rect 43720 230528 43772 230580
rect 46020 230528 46072 230580
rect 659660 230528 659712 230580
rect 45652 230460 45704 230512
rect 662788 230460 662840 230512
rect 42156 230324 42208 230376
rect 43996 230324 44048 230376
rect 359096 230324 359148 230376
rect 446588 230324 446640 230376
rect 357716 230256 357768 230308
rect 443184 230256 443236 230308
rect 363052 230188 363104 230240
rect 454132 230188 454184 230240
rect 361948 230120 362000 230172
rect 453304 230120 453356 230172
rect 360568 230052 360620 230104
rect 449900 230052 449952 230104
rect 364800 229984 364852 230036
rect 460020 229984 460072 230036
rect 363420 229916 363472 229968
rect 456616 229916 456668 229968
rect 42156 229848 42208 229900
rect 43904 229848 43956 229900
rect 364064 229848 364116 229900
rect 455788 229848 455840 229900
rect 366916 229780 366968 229832
rect 462504 229780 462556 229832
rect 366272 229712 366324 229764
rect 463700 229712 463752 229764
rect 372620 229644 372672 229696
rect 476028 229644 476080 229696
rect 370504 229576 370556 229628
rect 473452 229576 473504 229628
rect 369124 229508 369176 229560
rect 470140 229508 470192 229560
rect 371240 229440 371292 229492
rect 472624 229440 472676 229492
rect 373356 229372 373408 229424
rect 480352 229372 480404 229424
rect 374828 229304 374880 229356
rect 483020 229304 483072 229356
rect 376208 229236 376260 229288
rect 487160 229236 487212 229288
rect 393688 229168 393740 229220
rect 528376 229168 528428 229220
rect 396908 229100 396960 229152
rect 536656 229100 536708 229152
rect 158720 229032 158772 229084
rect 237564 229032 237616 229084
rect 246212 229032 246264 229084
rect 258540 229032 258592 229084
rect 296352 229032 296404 229084
rect 298468 229032 298520 229084
rect 298836 229032 298888 229084
rect 302700 229032 302752 229084
rect 304172 229032 304224 229084
rect 314660 229032 314712 229084
rect 339132 229032 339184 229084
rect 377036 229032 377088 229084
rect 152832 228964 152884 229016
rect 233976 228964 234028 229016
rect 243544 228964 243596 229016
rect 272432 228964 272484 229016
rect 293224 228964 293276 229016
rect 294604 228964 294656 229016
rect 297456 228964 297508 229016
rect 299388 228964 299440 229016
rect 303528 228964 303580 229016
rect 315304 228964 315356 229016
rect 318800 228964 318852 229016
rect 340972 228964 341024 229016
rect 342352 228964 342404 229016
rect 380900 228964 380952 229016
rect 388352 228964 388404 229016
rect 397368 229032 397420 229084
rect 401508 229032 401560 229084
rect 458180 229032 458232 229084
rect 392124 228964 392176 229016
rect 467012 228964 467064 229016
rect 156972 228896 157024 228948
rect 237196 228896 237248 228948
rect 241244 228896 241296 228948
rect 269580 228896 269632 228948
rect 296720 228896 296772 228948
rect 300216 228896 300268 228948
rect 304540 228896 304592 228948
rect 316132 228896 316184 228948
rect 336280 228896 336332 228948
rect 378508 228896 378560 228948
rect 389732 228896 389784 228948
rect 464436 228896 464488 228948
rect 150256 228828 150308 228880
rect 234344 228828 234396 228880
rect 239772 228828 239824 228880
rect 266728 228828 266780 228880
rect 308496 228828 308548 228880
rect 324596 228828 324648 228880
rect 340880 228828 340932 228880
rect 383752 228828 383804 228880
rect 387248 228828 387300 228880
rect 401508 228828 401560 228880
rect 151728 228760 151780 228812
rect 234712 228760 234764 228812
rect 239956 228760 240008 228812
rect 265348 228760 265400 228812
rect 305644 228760 305696 228812
rect 317880 228760 317932 228812
rect 340604 228760 340656 228812
rect 391756 228760 391808 228812
rect 394056 228760 394108 228812
rect 469956 228828 470008 228880
rect 403348 228760 403400 228812
rect 416780 228760 416832 228812
rect 416872 228760 416924 228812
rect 477500 228760 477552 228812
rect 146024 228692 146076 228744
rect 231124 228692 231176 228744
rect 241980 228692 242032 228744
rect 272156 228692 272208 228744
rect 306656 228692 306708 228744
rect 323860 228692 323912 228744
rect 337752 228692 337804 228744
rect 389088 228692 389140 228744
rect 396172 228692 396224 228744
rect 473268 228692 473320 228744
rect 138480 228624 138532 228676
rect 229008 228624 229060 228676
rect 245292 228624 245344 228676
rect 273536 228624 273588 228676
rect 304908 228624 304960 228676
rect 318708 228624 318760 228676
rect 323492 228624 323544 228676
rect 362408 228624 362460 228676
rect 376576 228624 376628 228676
rect 460940 228624 460992 228676
rect 143448 228556 143500 228608
rect 231492 228556 231544 228608
rect 239864 228556 239916 228608
rect 268200 228556 268252 228608
rect 307392 228556 307444 228608
rect 322940 228556 322992 228608
rect 336648 228556 336700 228608
rect 375288 228556 375340 228608
rect 377956 228556 378008 228608
rect 474740 228556 474792 228608
rect 145196 228488 145248 228540
rect 231860 228488 231912 228540
rect 240140 228488 240192 228540
rect 271052 228488 271104 228540
rect 308864 228488 308916 228540
rect 326252 228488 326304 228540
rect 335176 228488 335228 228540
rect 374000 228488 374052 228540
rect 375472 228488 375524 228540
rect 480260 228488 480312 228540
rect 136824 228420 136876 228472
rect 228640 228420 228692 228472
rect 238576 228420 238628 228472
rect 270684 228420 270736 228472
rect 307760 228420 307812 228472
rect 325700 228420 325752 228472
rect 332048 228420 332100 228472
rect 376852 228420 376904 228472
rect 379428 228420 379480 228472
rect 494520 228420 494572 228472
rect 131764 228352 131816 228404
rect 226156 228352 226208 228404
rect 235264 228352 235316 228404
rect 269304 228352 269356 228404
rect 302792 228352 302844 228404
rect 311164 228352 311216 228404
rect 317420 228352 317472 228404
rect 125048 228284 125100 228336
rect 223304 228284 223356 228336
rect 229284 228284 229336 228336
rect 267464 228284 267516 228336
rect 308128 228284 308180 228336
rect 327080 228284 327132 228336
rect 130108 228216 130160 228268
rect 225788 228216 225840 228268
rect 227628 228216 227680 228268
rect 267096 228216 267148 228268
rect 300952 228216 301004 228268
rect 310244 228216 310296 228268
rect 123392 228148 123444 228200
rect 222936 228148 222988 228200
rect 231676 228148 231728 228200
rect 267832 228148 267884 228200
rect 307024 228148 307076 228200
rect 321192 228148 321244 228200
rect 329196 228352 329248 228404
rect 375932 228352 375984 228404
rect 382280 228352 382332 228404
rect 501236 228352 501288 228404
rect 334900 228284 334952 228336
rect 382004 228284 382056 228336
rect 384396 228284 384448 228336
rect 506296 228284 506348 228336
rect 330576 228216 330628 228268
rect 379244 228216 379296 228268
rect 386512 228216 386564 228268
rect 511356 228216 511408 228268
rect 337660 228148 337712 228200
rect 339500 228148 339552 228200
rect 391848 228148 391900 228200
rect 400496 228148 400548 228200
rect 416872 228148 416924 228200
rect 416964 228148 417016 228200
rect 550272 228148 550324 228200
rect 114928 228080 114980 228132
rect 218980 228080 219032 228132
rect 223488 228080 223540 228132
rect 263876 228080 263928 228132
rect 309508 228080 309560 228132
rect 330484 228080 330536 228132
rect 333428 228080 333480 228132
rect 385960 228080 386012 228132
rect 403624 228080 403676 228132
rect 552020 228080 552072 228132
rect 108212 228012 108264 228064
rect 216128 228012 216180 228064
rect 216680 228012 216732 228064
rect 261024 228012 261076 228064
rect 311716 228012 311768 228064
rect 332968 228012 333020 228064
rect 337016 228012 337068 228064
rect 391940 228012 391992 228064
rect 402980 228012 403032 228064
rect 416964 228012 417016 228064
rect 417056 228012 417108 228064
rect 549260 228012 549312 228064
rect 72056 227944 72108 227996
rect 199752 227944 199804 227996
rect 203248 227944 203300 227996
rect 255320 227944 255372 227996
rect 255964 227944 256016 227996
rect 275652 227944 275704 227996
rect 311348 227944 311400 227996
rect 331312 227944 331364 227996
rect 341248 227944 341300 227996
rect 396540 227944 396592 227996
rect 406844 227944 406896 227996
rect 559288 227944 559340 227996
rect 78772 227876 78824 227928
rect 193772 227876 193824 227928
rect 69480 227808 69532 227860
rect 200120 227876 200172 227928
rect 209596 227876 209648 227928
rect 258172 227876 258224 227928
rect 258356 227876 258408 227928
rect 277492 227876 277544 227928
rect 301688 227876 301740 227928
rect 309416 227876 309468 227928
rect 310612 227876 310664 227928
rect 332140 227876 332192 227928
rect 338396 227876 338448 227928
rect 392952 227876 393004 227928
rect 409052 227876 409104 227928
rect 564440 227876 564492 227928
rect 198740 227808 198792 227860
rect 203984 227808 204036 227860
rect 65340 227740 65392 227792
rect 196900 227740 196952 227792
rect 198924 227740 198976 227792
rect 254676 227808 254728 227860
rect 259552 227808 259604 227860
rect 278872 227808 278924 227860
rect 312084 227808 312136 227860
rect 335544 227808 335596 227860
rect 341616 227808 341668 227860
rect 403624 227808 403676 227860
rect 409328 227808 409380 227860
rect 565452 227808 565504 227860
rect 52736 227672 52788 227724
rect 192944 227672 192996 227724
rect 197360 227672 197412 227724
rect 254308 227740 254360 227792
rect 256516 227740 256568 227792
rect 277124 227740 277176 227792
rect 312728 227740 312780 227792
rect 334716 227740 334768 227792
rect 341984 227740 342036 227792
rect 402980 227740 403032 227792
rect 407212 227740 407264 227792
rect 560392 227740 560444 227792
rect 204260 227672 204312 227724
rect 251824 227672 251876 227724
rect 253756 227672 253808 227724
rect 276756 227672 276808 227724
rect 315948 227672 316000 227724
rect 338304 227672 338356 227724
rect 344468 227672 344520 227724
rect 410340 227672 410392 227724
rect 411536 227672 411588 227724
rect 570236 227672 570288 227724
rect 156144 227604 156196 227656
rect 235356 227604 235408 227656
rect 248696 227604 248748 227656
rect 275008 227604 275060 227656
rect 306012 227604 306064 227656
rect 319536 227604 319588 227656
rect 322020 227604 322072 227656
rect 359096 227604 359148 227656
rect 385132 227604 385184 227656
rect 453856 227604 453908 227656
rect 162768 227536 162820 227588
rect 238208 227536 238260 227588
rect 250352 227536 250404 227588
rect 275284 227536 275336 227588
rect 320272 227536 320324 227588
rect 342076 227536 342128 227588
rect 343732 227536 343784 227588
rect 378140 227536 378192 227588
rect 383016 227536 383068 227588
rect 452568 227536 452620 227588
rect 165436 227468 165488 227520
rect 240416 227468 240468 227520
rect 252008 227468 252060 227520
rect 276388 227468 276440 227520
rect 305276 227468 305328 227520
rect 320364 227468 320416 227520
rect 320640 227468 320692 227520
rect 356060 227468 356112 227520
rect 374460 227468 374512 227520
rect 435732 227468 435784 227520
rect 163688 227400 163740 227452
rect 240048 227400 240100 227452
rect 258724 227400 258776 227452
rect 274272 227400 274324 227452
rect 303804 227400 303856 227452
rect 317420 227400 317472 227452
rect 321652 227400 321704 227452
rect 342904 227400 342956 227452
rect 371608 227400 371660 227452
rect 433156 227400 433208 227452
rect 42064 227332 42116 227384
rect 43444 227332 43496 227384
rect 167092 227332 167144 227384
rect 241428 227332 241480 227384
rect 253572 227332 253624 227384
rect 272800 227332 272852 227384
rect 303160 227332 303212 227384
rect 312820 227332 312872 227384
rect 323124 227332 323176 227384
rect 342996 227332 343048 227384
rect 365904 227332 365956 227384
rect 425428 227332 425480 227384
rect 173624 227264 173676 227316
rect 244280 227264 244332 227316
rect 253204 227264 253256 227316
rect 271420 227264 271472 227316
rect 295248 227264 295300 227316
rect 296812 227264 296864 227316
rect 298744 227264 298796 227316
rect 301044 227264 301096 227316
rect 302424 227264 302476 227316
rect 313648 227264 313700 227316
rect 325976 227264 326028 227316
rect 345296 227264 345348 227316
rect 350172 227264 350224 227316
rect 408500 227264 408552 227316
rect 169576 227196 169628 227248
rect 241060 227196 241112 227248
rect 248512 227196 248564 227248
rect 268568 227196 268620 227248
rect 302056 227196 302108 227248
rect 311992 227196 312044 227248
rect 368756 227196 368808 227248
rect 430396 227196 430448 227248
rect 172152 227128 172204 227180
rect 243268 227128 243320 227180
rect 256608 227128 256660 227180
rect 258724 227128 258776 227180
rect 181904 227060 181956 227112
rect 246120 227060 246172 227112
rect 247040 227060 247092 227112
rect 273904 227128 273956 227180
rect 309232 227128 309284 227180
rect 328828 227128 328880 227180
rect 331680 227128 331732 227180
rect 347780 227128 347832 227180
rect 353024 227128 353076 227180
rect 413192 227128 413244 227180
rect 258908 227060 258960 227112
rect 276020 227060 276072 227112
rect 306380 227060 306432 227112
rect 322020 227060 322072 227112
rect 358728 227060 358780 227112
rect 415308 227060 415360 227112
rect 176384 226992 176436 227044
rect 243912 226992 243964 227044
rect 255504 226992 255556 227044
rect 271788 226992 271840 227044
rect 338028 226992 338080 227044
rect 372068 226992 372120 227044
rect 372988 226992 373040 227044
rect 433248 226992 433300 227044
rect 180524 226924 180576 226976
rect 247132 226924 247184 226976
rect 190368 226856 190420 226908
rect 251456 226924 251508 226976
rect 258724 226924 258776 226976
rect 274640 226924 274692 226976
rect 298100 226924 298152 226976
rect 301964 226924 302016 226976
rect 310520 226924 310572 226976
rect 329656 226924 329708 226976
rect 364432 226924 364484 226976
rect 422300 226924 422352 226976
rect 248604 226856 248656 226908
rect 269948 226856 270000 226908
rect 290740 226856 290792 226908
rect 292396 226856 292448 226908
rect 300676 226856 300728 226908
rect 308588 226856 308640 226908
rect 361580 226856 361632 226908
rect 416872 226856 416924 226908
rect 42156 226788 42208 226840
rect 43628 226788 43680 226840
rect 189264 226788 189316 226840
rect 248972 226788 249024 226840
rect 186412 226720 186464 226772
rect 248236 226720 248288 226772
rect 248420 226720 248472 226772
rect 265716 226788 265768 226840
rect 299572 226788 299624 226840
rect 306932 226788 306984 226840
rect 359832 226788 359884 226840
rect 404544 226788 404596 226840
rect 409696 226788 409748 226840
rect 447140 226788 447192 226840
rect 255780 226720 255832 226772
rect 268936 226720 268988 226772
rect 299204 226720 299256 226772
rect 305276 226720 305328 226772
rect 368388 226720 368440 226772
rect 408776 226720 408828 226772
rect 195888 226652 195940 226704
rect 251088 226652 251140 226704
rect 258816 226652 258868 226704
rect 273168 226652 273220 226704
rect 297824 226652 297876 226704
rect 301872 226652 301924 226704
rect 301964 226652 302016 226704
rect 303620 226652 303672 226704
rect 329104 226652 329156 226704
rect 345112 226652 345164 226704
rect 365536 226652 365588 226704
rect 405832 226652 405884 226704
rect 408684 226652 408736 226704
rect 444380 226652 444432 226704
rect 193036 226584 193088 226636
rect 204260 226584 204312 226636
rect 236276 226584 236328 226636
rect 256792 226584 256844 226636
rect 300308 226584 300360 226636
rect 306380 226584 306432 226636
rect 395804 226584 395856 226636
rect 438768 226584 438820 226636
rect 193772 226516 193824 226568
rect 202604 226516 202656 226568
rect 301320 226516 301372 226568
rect 307760 226516 307812 226568
rect 402612 226516 402664 226568
rect 417056 226516 417108 226568
rect 255320 226448 255372 226500
rect 270316 226448 270368 226500
rect 374092 226448 374144 226500
rect 405740 226448 405792 226500
rect 201592 226380 201644 226432
rect 209044 226380 209096 226432
rect 233516 226380 233568 226432
rect 247500 226380 247552 226432
rect 404360 226380 404412 226432
rect 441620 226516 441672 226568
rect 183008 226312 183060 226364
rect 192300 226312 192352 226364
rect 258172 226312 258224 226364
rect 264612 226312 264664 226364
rect 299940 226312 299992 226364
rect 304356 226312 304408 226364
rect 309876 226312 309928 226364
rect 327908 226312 327960 226364
rect 144368 226244 144420 226296
rect 230756 226244 230808 226296
rect 349436 226244 349488 226296
rect 425060 226244 425112 226296
rect 430396 226244 430448 226296
rect 467564 226244 467616 226296
rect 147772 226176 147824 226228
rect 232228 226176 232280 226228
rect 352656 226176 352708 226228
rect 428924 226176 428976 226228
rect 433156 226176 433208 226228
rect 474280 226176 474332 226228
rect 141056 226108 141108 226160
rect 229376 226108 229428 226160
rect 353760 226108 353812 226160
rect 434812 226108 434864 226160
rect 137652 226040 137704 226092
rect 227904 226040 227956 226092
rect 352288 226040 352340 226092
rect 431408 226040 431460 226092
rect 433248 226040 433300 226092
rect 477776 226040 477828 226092
rect 134248 225972 134300 226024
rect 226524 225972 226576 226024
rect 356980 225972 357032 226024
rect 439044 225972 439096 226024
rect 130936 225904 130988 225956
rect 225052 225904 225104 225956
rect 243084 225904 243136 225956
rect 252928 225904 252980 225956
rect 355508 225904 355560 225956
rect 435640 225904 435692 225956
rect 435732 225904 435784 225956
rect 480996 225972 481048 226024
rect 127532 225836 127584 225888
rect 223672 225836 223724 225888
rect 242992 225836 243044 225888
rect 252836 225836 252888 225888
rect 356612 225836 356664 225888
rect 429108 225836 429160 225888
rect 119160 225768 119212 225820
rect 219716 225768 219768 225820
rect 231308 225768 231360 225820
rect 249616 225768 249668 225820
rect 359464 225768 359516 225820
rect 448244 225836 448296 225888
rect 474740 225836 474792 225888
rect 491300 225836 491352 225888
rect 124128 225700 124180 225752
rect 222200 225700 222252 225752
rect 232044 225700 232096 225752
rect 253940 225700 253992 225752
rect 362316 225700 362368 225752
rect 114100 225632 114152 225684
rect 217968 225632 218020 225684
rect 110696 225564 110748 225616
rect 216496 225564 216548 225616
rect 216588 225564 216640 225616
rect 252468 225632 252520 225684
rect 360844 225632 360896 225684
rect 451556 225700 451608 225752
rect 452568 225768 452620 225820
rect 503168 225768 503220 225820
rect 454960 225700 455012 225752
rect 460940 225700 460992 225752
rect 487804 225700 487856 225752
rect 228456 225564 228508 225616
rect 266452 225564 266504 225616
rect 362684 225564 362736 225616
rect 440332 225564 440384 225616
rect 105728 225496 105780 225548
rect 214012 225496 214064 225548
rect 218428 225496 218480 225548
rect 262128 225496 262180 225548
rect 365168 225496 365220 225548
rect 461676 225632 461728 225684
rect 467012 225632 467064 225684
rect 523960 225632 524012 225684
rect 440516 225564 440568 225616
rect 452660 225564 452712 225616
rect 453856 225564 453908 225616
rect 507952 225564 508004 225616
rect 107384 225428 107436 225480
rect 215116 225428 215168 225480
rect 221740 225428 221792 225480
rect 263600 225428 263652 225480
rect 363696 225428 363748 225480
rect 458456 225496 458508 225548
rect 464436 225496 464488 225548
rect 518900 225496 518952 225548
rect 458180 225428 458232 225480
rect 513380 225428 513432 225480
rect 100668 225360 100720 225412
rect 192760 225360 192812 225412
rect 97264 225292 97316 225344
rect 207020 225360 207072 225412
rect 225144 225360 225196 225412
rect 264980 225360 265032 225412
rect 355140 225360 355192 225412
rect 438124 225360 438176 225412
rect 438768 225360 438820 225412
rect 532700 225360 532752 225412
rect 95608 225224 95660 225276
rect 209688 225292 209740 225344
rect 215024 225292 215076 225344
rect 260748 225292 260800 225344
rect 366548 225292 366600 225344
rect 465080 225292 465132 225344
rect 469956 225292 470008 225344
rect 529020 225292 529072 225344
rect 211712 225224 211764 225276
rect 259276 225224 259328 225276
rect 343088 225224 343140 225276
rect 365720 225224 365772 225276
rect 368020 225224 368072 225276
rect 468392 225224 468444 225276
rect 473268 225224 473320 225276
rect 533988 225224 534040 225276
rect 88892 225156 88944 225208
rect 192668 225156 192720 225208
rect 192760 225156 192812 225208
rect 197452 225156 197504 225208
rect 208308 225156 208360 225208
rect 257896 225156 257948 225208
rect 313464 225156 313516 225208
rect 338856 225156 338908 225208
rect 339868 225156 339920 225208
rect 368572 225156 368624 225208
rect 369768 225156 369820 225208
rect 469220 225156 469272 225208
rect 477500 225156 477552 225208
rect 544108 225156 544160 225208
rect 92204 225088 92256 225140
rect 208032 225088 208084 225140
rect 209228 225088 209280 225140
rect 257160 225088 257212 225140
rect 314936 225088 314988 225140
rect 342536 225088 342588 225140
rect 358360 225088 358412 225140
rect 73712 225020 73764 225072
rect 200856 225020 200908 225072
rect 201408 225020 201460 225072
rect 255044 225020 255096 225072
rect 317788 225020 317840 225072
rect 348976 225020 349028 225072
rect 357992 225020 358044 225072
rect 441620 225088 441672 225140
rect 554320 225088 554372 225140
rect 60280 224952 60332 225004
rect 195152 224952 195204 225004
rect 195244 224952 195296 225004
rect 252192 224952 252244 225004
rect 319168 224952 319220 225004
rect 352380 224952 352432 225004
rect 361212 224952 361264 225004
rect 434628 224952 434680 225004
rect 442356 225020 442408 225072
rect 444380 225020 444432 225072
rect 563704 225020 563756 225072
rect 55128 224884 55180 224936
rect 192576 224884 192628 224936
rect 192668 224884 192720 224936
rect 206836 224884 206888 224936
rect 206928 224884 206980 224936
rect 250720 224884 250772 224936
rect 316316 224884 316368 224936
rect 345664 224884 345716 224936
rect 346584 224884 346636 224936
rect 416688 224884 416740 224936
rect 416780 224884 416832 224936
rect 444840 224952 444892 225004
rect 447140 224952 447192 225004
rect 566004 224952 566056 225004
rect 549352 224884 549404 224936
rect 114284 224816 114336 224868
rect 198004 224816 198056 224868
rect 198188 224816 198240 224868
rect 253296 224816 253348 224868
rect 350908 224816 350960 224868
rect 428004 224816 428056 224868
rect 434628 224816 434680 224868
rect 449072 224816 449124 224868
rect 154488 224748 154540 224800
rect 235080 224748 235132 224800
rect 354128 224748 354180 224800
rect 425244 224748 425296 224800
rect 151084 224680 151136 224732
rect 233608 224680 233660 224732
rect 351276 224680 351328 224732
rect 425520 224748 425572 224800
rect 429108 224748 429160 224800
rect 441620 224748 441672 224800
rect 425428 224680 425480 224732
rect 460940 224680 460992 224732
rect 161204 224612 161256 224664
rect 237932 224612 237984 224664
rect 349804 224612 349856 224664
rect 401508 224612 401560 224664
rect 416688 224612 416740 224664
rect 417976 224612 418028 224664
rect 422300 224612 422352 224664
rect 457444 224612 457496 224664
rect 157800 224544 157852 224596
rect 236460 224544 236512 224596
rect 342720 224544 342772 224596
rect 405648 224544 405700 224596
rect 405740 224544 405792 224596
rect 479340 224544 479392 224596
rect 169116 224476 169168 224528
rect 240784 224476 240836 224528
rect 348056 224476 348108 224528
rect 421288 224476 421340 224528
rect 425244 224476 425296 224528
rect 432236 224476 432288 224528
rect 166356 224408 166408 224460
rect 239312 224408 239364 224460
rect 346952 224408 347004 224460
rect 415400 224408 415452 224460
rect 416872 224408 416924 224460
rect 450728 224408 450780 224460
rect 171048 224340 171100 224392
rect 242164 224340 242216 224392
rect 348424 224340 348476 224392
rect 418804 224340 418856 224392
rect 176660 224272 176712 224324
rect 243636 224272 243688 224324
rect 345204 224272 345256 224324
rect 414572 224272 414624 224324
rect 415308 224272 415360 224324
rect 444380 224272 444432 224324
rect 181352 224204 181404 224256
rect 246488 224204 246540 224256
rect 345572 224204 345624 224256
rect 412088 224204 412140 224256
rect 413192 224204 413244 224256
rect 430580 224204 430632 224256
rect 178040 224136 178092 224188
rect 245016 224136 245068 224188
rect 344100 224136 344152 224188
rect 408684 224136 408736 224188
rect 408776 224136 408828 224188
rect 465908 224136 465960 224188
rect 184756 224068 184808 224120
rect 247868 224068 247920 224120
rect 340236 224068 340288 224120
rect 400404 224068 400456 224120
rect 405832 224068 405884 224120
rect 459192 224068 459244 224120
rect 146300 224000 146352 224052
rect 197452 224000 197504 224052
rect 212264 224000 212316 224052
rect 216128 224000 216180 224052
rect 246764 224000 246816 224052
rect 383752 224000 383804 224052
rect 404452 224000 404504 224052
rect 404544 224000 404596 224052
rect 445668 224000 445720 224052
rect 188160 223932 188212 223984
rect 249340 223932 249392 223984
rect 378140 223932 378192 223984
rect 204904 223864 204956 223916
rect 256424 223864 256476 223916
rect 380900 223864 380952 223916
rect 401508 223932 401560 223984
rect 422300 223932 422352 223984
rect 188436 223796 188488 223848
rect 232504 223796 232556 223848
rect 407856 223796 407908 223848
rect 411260 223796 411312 223848
rect 191472 223728 191524 223780
rect 206928 223728 206980 223780
rect 208952 223728 209004 223780
rect 239680 223728 239732 223780
rect 185584 223592 185636 223644
rect 189264 223592 189316 223644
rect 209688 223660 209740 223712
rect 236828 223660 236880 223712
rect 209412 223592 209464 223644
rect 214932 223592 214984 223644
rect 242532 223592 242584 223644
rect 408500 223592 408552 223644
rect 423864 223592 423916 223644
rect 480260 223592 480312 223644
rect 484400 223592 484452 223644
rect 155316 223524 155368 223576
rect 236092 223524 236144 223576
rect 278688 223524 278740 223576
rect 287796 223524 287848 223576
rect 324504 223524 324556 223576
rect 363236 223524 363288 223576
rect 392952 223524 393004 223576
rect 395252 223524 395304 223576
rect 402980 223524 403032 223576
rect 406200 223524 406252 223576
rect 503812 223524 503864 223576
rect 623412 223524 623464 223576
rect 93768 223456 93820 223508
rect 146300 223456 146352 223508
rect 153660 223456 153712 223508
rect 235724 223456 235776 223508
rect 241152 223456 241204 223508
rect 253572 223456 253624 223508
rect 322388 223456 322440 223508
rect 360752 223456 360804 223508
rect 494060 223456 494112 223508
rect 607588 223456 607640 223508
rect 146944 223388 146996 223440
rect 232872 223388 232924 223440
rect 324136 223388 324188 223440
rect 361764 223388 361816 223440
rect 397276 223388 397328 223440
rect 406568 223388 406620 223440
rect 499488 223388 499540 223440
rect 608048 223388 608100 223440
rect 148600 223320 148652 223372
rect 233240 223320 233292 223372
rect 237748 223320 237800 223372
rect 253204 223320 253256 223372
rect 324872 223320 324924 223372
rect 365812 223320 365864 223372
rect 398288 223320 398340 223372
rect 539048 223320 539100 223372
rect 87144 223252 87196 223304
rect 172428 223252 172480 223304
rect 175464 223252 175516 223304
rect 244648 223252 244700 223304
rect 326988 223252 327040 223304
rect 368296 223252 368348 223304
rect 399024 223252 399076 223304
rect 536288 223252 536340 223304
rect 536380 223252 536432 223304
rect 141884 223184 141936 223236
rect 230388 223184 230440 223236
rect 239404 223184 239456 223236
rect 255504 223184 255556 223236
rect 326344 223184 326396 223236
rect 369124 223184 369176 223236
rect 400128 223184 400180 223236
rect 406476 223184 406528 223236
rect 406568 223184 406620 223236
rect 536564 223184 536616 223236
rect 536656 223184 536708 223236
rect 615040 223184 615092 223236
rect 140136 223116 140188 223168
rect 230020 223116 230072 223168
rect 235908 223116 235960 223168
rect 249984 223116 250036 223168
rect 325608 223116 325660 223168
rect 364984 223116 365036 223168
rect 399392 223116 399444 223168
rect 541624 223116 541676 223168
rect 135168 223048 135220 223100
rect 227536 223048 227588 223100
rect 232596 223048 232648 223100
rect 242716 223048 242768 223100
rect 242808 223048 242860 223100
rect 258816 223048 258868 223100
rect 271420 223048 271472 223100
rect 285680 223048 285732 223100
rect 328460 223048 328512 223100
rect 371700 223048 371752 223100
rect 400772 223048 400824 223100
rect 545120 223048 545172 223100
rect 545764 223048 545816 223100
rect 616880 223048 616932 223100
rect 133420 222980 133472 223032
rect 227168 222980 227220 223032
rect 231032 222980 231084 223032
rect 248512 222980 248564 223032
rect 323768 222980 323820 223032
rect 364340 222980 364392 223032
rect 372068 222980 372120 223032
rect 397736 222980 397788 223032
rect 401784 222980 401836 223032
rect 128360 222912 128412 222964
rect 224684 222912 224736 222964
rect 236092 222912 236144 222964
rect 255320 222912 255372 222964
rect 263784 222912 263836 222964
rect 280988 222912 281040 222964
rect 327356 222912 327408 222964
rect 370044 222912 370096 222964
rect 396540 222912 396592 222964
rect 401968 222912 402020 222964
rect 406476 222980 406528 223032
rect 543556 222980 543608 223032
rect 546684 222912 546736 222964
rect 617340 222980 617392 223032
rect 566004 222912 566056 222964
rect 620560 222912 620612 222964
rect 126704 222844 126756 222896
rect 224040 222844 224092 222896
rect 232688 222844 232740 222896
rect 255780 222844 255832 222896
rect 257068 222844 257120 222896
rect 278136 222844 278188 222896
rect 325240 222844 325292 222896
rect 367468 222844 367520 222896
rect 368572 222844 368624 222896
rect 398564 222844 398616 222896
rect 402244 222844 402296 222896
rect 548340 222844 548392 222896
rect 549352 222844 549404 222896
rect 551100 222844 551152 222896
rect 617800 222844 617852 222896
rect 66996 222776 67048 222828
rect 114284 222776 114336 222828
rect 116584 222776 116636 222828
rect 220084 222776 220136 222828
rect 224316 222776 224368 222828
rect 248420 222776 248472 222828
rect 264612 222776 264664 222828
rect 282828 222776 282880 222828
rect 326620 222776 326672 222828
rect 370872 222776 370924 222828
rect 401876 222776 401928 222828
rect 547512 222776 547564 222828
rect 553768 222776 553820 222828
rect 91376 222708 91428 222760
rect 201592 222708 201644 222760
rect 214196 222708 214248 222760
rect 245660 222708 245712 222760
rect 246120 222708 246172 222760
rect 258724 222708 258776 222760
rect 262956 222708 263008 222760
rect 281724 222708 281776 222760
rect 327724 222708 327776 222760
rect 372620 222708 372672 222760
rect 374000 222708 374052 222760
rect 391020 222708 391072 222760
rect 404728 222708 404780 222760
rect 554228 222708 554280 222760
rect 554320 222708 554372 222760
rect 618260 222708 618312 222760
rect 89720 222640 89772 222692
rect 201684 222640 201736 222692
rect 222568 222640 222620 222692
rect 258172 222640 258224 222692
rect 260472 222640 260524 222692
rect 279608 222640 279660 222692
rect 329472 222640 329524 222692
rect 377588 222640 377640 222692
rect 391756 222640 391808 222692
rect 402980 222640 403032 222692
rect 406108 222640 406160 222692
rect 556712 222640 556764 222692
rect 568580 222640 568632 222692
rect 621020 222640 621072 222692
rect 82176 222572 82228 222624
rect 198740 222572 198792 222624
rect 207480 222572 207532 222624
rect 246212 222572 246264 222624
rect 259368 222572 259420 222624
rect 280344 222572 280396 222624
rect 329840 222572 329892 222624
rect 375380 222572 375432 222624
rect 405096 222572 405148 222624
rect 555056 222572 555108 222624
rect 556068 222572 556120 222624
rect 618720 222572 618772 222624
rect 85488 222504 85540 222556
rect 205456 222504 205508 222556
rect 215852 222504 215904 222556
rect 259184 222504 259236 222556
rect 261300 222504 261352 222556
rect 281356 222504 281408 222556
rect 81256 222436 81308 222488
rect 204720 222436 204772 222488
rect 209136 222436 209188 222488
rect 258632 222436 258684 222488
rect 262128 222436 262180 222488
rect 280712 222436 280764 222488
rect 75368 222368 75420 222420
rect 201132 222368 201184 222420
rect 205824 222368 205876 222420
rect 257528 222368 257580 222420
rect 272248 222368 272300 222420
rect 284944 222504 284996 222556
rect 331588 222504 331640 222556
rect 378416 222504 378468 222556
rect 378508 222504 378560 222556
rect 392676 222504 392728 222556
rect 406384 222504 406436 222556
rect 558184 222504 558236 222556
rect 559104 222504 559156 222556
rect 619180 222504 619232 222556
rect 283104 222436 283156 222488
rect 290280 222436 290332 222488
rect 338304 222436 338356 222488
rect 343088 222436 343140 222488
rect 343548 222436 343600 222488
rect 376760 222436 376812 222488
rect 377036 222436 377088 222488
rect 399484 222436 399536 222488
rect 407948 222436 408000 222488
rect 561772 222436 561824 222488
rect 563704 222436 563756 222488
rect 620100 222436 620152 222488
rect 328092 222368 328144 222420
rect 338028 222368 338080 222420
rect 338212 222368 338264 222420
rect 374184 222368 374236 222420
rect 375288 222368 375340 222420
rect 394700 222368 394752 222420
rect 407580 222368 407632 222420
rect 561588 222368 561640 222420
rect 619640 222368 619692 222420
rect 68652 222300 68704 222352
rect 198280 222300 198332 222352
rect 202420 222300 202472 222352
rect 256056 222300 256108 222352
rect 269672 222300 269724 222352
rect 284576 222300 284628 222352
rect 332692 222300 332744 222352
rect 381820 222300 381872 222352
rect 390836 222300 390888 222352
rect 53564 222232 53616 222284
rect 183008 222232 183060 222284
rect 187240 222232 187292 222284
rect 235908 222232 235960 222284
rect 254584 222232 254636 222284
rect 278504 222232 278556 222284
rect 310980 222232 311032 222284
rect 333980 222232 334032 222284
rect 337660 222232 337712 222284
rect 346492 222232 346544 222284
rect 346584 222232 346636 222284
rect 385132 222232 385184 222284
rect 391848 222232 391900 222284
rect 401140 222232 401192 222284
rect 41696 222164 41748 222216
rect 59544 222164 59596 222216
rect 61936 222164 61988 222216
rect 195428 222164 195480 222216
rect 200764 222164 200816 222216
rect 255688 222164 255740 222216
rect 258816 222164 258868 222216
rect 279240 222164 279292 222216
rect 312360 222164 312412 222216
rect 337200 222164 337252 222216
rect 340972 222164 341024 222216
rect 349804 222164 349856 222216
rect 349896 222164 349948 222216
rect 393596 222164 393648 222216
rect 162032 222096 162084 222148
rect 238944 222096 238996 222148
rect 244464 222096 244516 222148
rect 256608 222096 256660 222148
rect 273076 222096 273128 222148
rect 286048 222096 286100 222148
rect 322756 222096 322808 222148
rect 358268 222096 358320 222148
rect 381912 222096 381964 222148
rect 401416 222096 401468 222148
rect 408316 222300 408368 222352
rect 562968 222300 563020 222352
rect 634544 222300 634596 222352
rect 410064 222232 410116 222284
rect 566832 222232 566884 222284
rect 570236 222232 570288 222284
rect 570880 222232 570932 222284
rect 635924 222232 635976 222284
rect 410432 222164 410484 222216
rect 567660 222164 567712 222216
rect 521660 222096 521712 222148
rect 536288 222096 536340 222148
rect 541440 222096 541492 222148
rect 160376 222028 160428 222080
rect 238300 222028 238352 222080
rect 274732 222028 274784 222080
rect 287060 222028 287112 222080
rect 320916 222028 320968 222080
rect 357348 222028 357400 222080
rect 393228 222028 393280 222080
rect 526444 222028 526496 222080
rect 538864 222028 538916 222080
rect 615500 222096 615552 222148
rect 552572 222028 552624 222080
rect 553216 222028 553268 222080
rect 632704 222028 632756 222080
rect 90548 221960 90600 222012
rect 160100 221960 160152 222012
rect 170496 221960 170548 222012
rect 232596 221960 232648 222012
rect 168748 221892 168800 221944
rect 241796 221960 241848 222012
rect 319812 221960 319864 222012
rect 354036 221960 354088 222012
rect 388720 221960 388772 222012
rect 516416 221960 516468 222012
rect 532700 221960 532752 222012
rect 533436 221960 533488 222012
rect 614580 221960 614632 222012
rect 234344 221892 234396 221944
rect 248604 221892 248656 221944
rect 273904 221892 273956 221944
rect 285312 221892 285364 221944
rect 287060 221892 287112 221944
rect 289268 221892 289320 221944
rect 318064 221892 318116 221944
rect 350632 221892 350684 221944
rect 387616 221892 387668 221944
rect 513840 221892 513892 221944
rect 530676 221892 530728 221944
rect 614028 221892 614080 221944
rect 177212 221824 177264 221876
rect 183928 221756 183980 221808
rect 281448 221824 281500 221876
rect 289912 221824 289964 221876
rect 319904 221824 319956 221876
rect 351460 221824 351512 221876
rect 386236 221824 386288 221876
rect 510620 221824 510672 221876
rect 547512 221824 547564 221876
rect 631784 221824 631836 221876
rect 182088 221688 182140 221740
rect 233516 221688 233568 221740
rect 179696 221620 179748 221672
rect 235632 221620 235684 221672
rect 245752 221756 245804 221808
rect 268016 221756 268068 221808
rect 284208 221756 284260 221808
rect 321284 221756 321336 221808
rect 354864 221756 354916 221808
rect 385500 221756 385552 221808
rect 508780 221756 508832 221808
rect 528376 221756 528428 221808
rect 613568 221756 613620 221808
rect 257896 221688 257948 221740
rect 279976 221688 280028 221740
rect 284852 221688 284904 221740
rect 291384 221688 291436 221740
rect 316684 221688 316736 221740
rect 347320 221688 347372 221740
rect 347780 221688 347832 221740
rect 380072 221688 380124 221740
rect 383384 221688 383436 221740
rect 503720 221688 503772 221740
rect 542728 221688 542780 221740
rect 630864 221688 630916 221740
rect 248328 221620 248380 221672
rect 255412 221620 255464 221672
rect 277860 221620 277912 221672
rect 194048 221552 194100 221604
rect 196072 221552 196124 221604
rect 196164 221552 196216 221604
rect 159548 221484 159600 221536
rect 209688 221484 209740 221536
rect 213368 221484 213420 221536
rect 236000 221552 236052 221604
rect 245384 221552 245436 221604
rect 275560 221552 275612 221604
rect 286416 221620 286468 221672
rect 317052 221620 317104 221672
rect 345020 221620 345072 221672
rect 345112 221620 345164 221672
rect 373356 221620 373408 221672
rect 384028 221620 384080 221672
rect 505744 221620 505796 221672
rect 538312 221620 538364 221672
rect 540152 221620 540204 221672
rect 630404 221620 630456 221672
rect 278136 221552 278188 221604
rect 288532 221552 288584 221604
rect 318432 221552 318484 221604
rect 348148 221552 348200 221604
rect 382004 221552 382056 221604
rect 389364 221552 389416 221604
rect 401416 221552 401468 221604
rect 500408 221552 500460 221604
rect 502708 221552 502760 221604
rect 503812 221552 503864 221604
rect 513380 221552 513432 221604
rect 610808 221552 610860 221604
rect 149428 221416 149480 221468
rect 188436 221416 188488 221468
rect 195704 221416 195756 221468
rect 192300 221348 192352 221400
rect 193036 221348 193088 221400
rect 193128 221348 193180 221400
rect 195888 221348 195940 221400
rect 196072 221416 196124 221468
rect 250076 221484 250128 221536
rect 266360 221484 266412 221536
rect 283196 221484 283248 221536
rect 286508 221484 286560 221536
rect 291752 221484 291804 221536
rect 315212 221484 315264 221536
rect 343916 221484 343968 221536
rect 345296 221484 345348 221536
rect 366640 221484 366692 221536
rect 380532 221484 380584 221536
rect 497372 221484 497424 221536
rect 499488 221484 499540 221536
rect 534908 221484 534960 221536
rect 629484 221484 629536 221536
rect 166264 221280 166316 221332
rect 208952 221280 209004 221332
rect 220084 221280 220136 221332
rect 231216 221280 231268 221332
rect 172980 221212 173032 221264
rect 214932 221212 214984 221264
rect 178868 221144 178920 221196
rect 181904 221144 181956 221196
rect 189816 221144 189868 221196
rect 231308 221144 231360 221196
rect 237012 221416 237064 221468
rect 249524 221416 249576 221468
rect 258908 221416 258960 221468
rect 265532 221416 265584 221468
rect 282092 221416 282144 221468
rect 283932 221416 283984 221468
rect 236920 221348 236972 221400
rect 241244 221348 241296 221400
rect 247868 221348 247920 221400
rect 255964 221348 256016 221400
rect 256240 221348 256292 221400
rect 259552 221348 259604 221400
rect 267188 221348 267240 221400
rect 282460 221348 282512 221400
rect 233516 221280 233568 221332
rect 239864 221280 239916 221332
rect 251088 221280 251140 221332
rect 256516 221280 256568 221332
rect 270408 221280 270460 221332
rect 283840 221280 283892 221332
rect 288256 221416 288308 221468
rect 292764 221416 292816 221468
rect 314568 221416 314620 221468
rect 339684 221416 339736 221468
rect 380808 221416 380860 221468
rect 497832 221416 497884 221468
rect 530124 221416 530176 221468
rect 628472 221416 628524 221468
rect 289084 221348 289136 221400
rect 292120 221348 292172 221400
rect 292396 221348 292448 221400
rect 293500 221348 293552 221400
rect 314200 221348 314252 221400
rect 338028 221348 338080 221400
rect 342904 221348 342956 221400
rect 356520 221348 356572 221400
rect 379060 221348 379112 221400
rect 494060 221348 494112 221400
rect 507952 221348 508004 221400
rect 609888 221348 609940 221400
rect 289544 221280 289596 221332
rect 291568 221280 291620 221332
rect 294236 221280 294288 221332
rect 294972 221280 295024 221332
rect 295616 221280 295668 221332
rect 313832 221280 313884 221332
rect 340604 221280 340656 221332
rect 342076 221280 342128 221332
rect 353300 221280 353352 221332
rect 377680 221280 377732 221332
rect 490288 221280 490340 221332
rect 518992 221280 519044 221332
rect 520004 221280 520056 221332
rect 525064 221280 525116 221332
rect 627552 221280 627604 221332
rect 242992 221212 243044 221264
rect 252928 221212 252980 221264
rect 258356 221212 258408 221264
rect 268844 221212 268896 221264
rect 283564 221212 283616 221264
rect 243084 221144 243136 221196
rect 277308 221144 277360 221196
rect 286692 221212 286744 221264
rect 289728 221212 289780 221264
rect 293132 221212 293184 221264
rect 315580 221212 315632 221264
rect 341432 221212 341484 221264
rect 371976 221212 372028 221264
rect 476856 221212 476908 221264
rect 503168 221212 503220 221264
rect 608968 221212 609020 221264
rect 283748 221144 283800 221196
rect 287428 221144 287480 221196
rect 313096 221144 313148 221196
rect 336740 221144 336792 221196
rect 337384 221144 337436 221196
rect 349896 221144 349948 221196
rect 367284 221144 367336 221196
rect 464252 221144 464304 221196
rect 520004 221144 520056 221196
rect 626632 221144 626684 221196
rect 655704 221144 655756 221196
rect 676036 221144 676088 221196
rect 183100 221076 183152 221128
rect 216128 221076 216180 221128
rect 188988 221008 189040 221060
rect 196164 221008 196216 221060
rect 199936 221008 199988 221060
rect 230112 221076 230164 221128
rect 230204 221076 230256 221128
rect 239772 221076 239824 221128
rect 282368 221076 282420 221128
rect 287060 221076 287112 221128
rect 287336 221076 287388 221128
rect 291016 221076 291068 221128
rect 330208 221076 330260 221128
rect 343548 221076 343600 221128
rect 365720 221076 365772 221128
rect 407028 221076 407080 221128
rect 517060 221076 517112 221128
rect 517612 221076 517664 221128
rect 626172 221076 626224 221128
rect 226800 221008 226852 221060
rect 239956 221008 240008 221060
rect 279792 221008 279844 221060
rect 288900 221008 288952 221060
rect 342996 221008 343048 221060
rect 359924 221008 359976 221060
rect 376852 221008 376904 221060
rect 382648 221008 382700 221060
rect 389088 221008 389140 221060
rect 396080 221008 396132 221060
rect 397644 221008 397696 221060
rect 537392 221008 537444 221060
rect 558184 221008 558236 221060
rect 633624 221008 633676 221060
rect 655520 221008 655572 221060
rect 675852 221008 675904 221060
rect 206652 220940 206704 220992
rect 196532 220872 196584 220924
rect 216588 220872 216640 220924
rect 164608 220804 164660 220856
rect 166356 220804 166408 220856
rect 167920 220804 167972 220856
rect 169116 220804 169168 220856
rect 174636 220804 174688 220856
rect 176660 220804 176712 220856
rect 204076 220804 204128 220856
rect 209228 220804 209280 220856
rect 236276 220940 236328 220992
rect 276480 220940 276532 220992
rect 283748 220940 283800 220992
rect 285680 220940 285732 220992
rect 290648 220940 290700 220992
rect 334164 220940 334216 220992
rect 346584 220940 346636 220992
rect 512184 220940 512236 220992
rect 625252 220940 625304 220992
rect 230112 220872 230164 220924
rect 232044 220872 232096 220924
rect 280620 220872 280672 220924
rect 288164 220872 288216 220924
rect 395436 220872 395488 220924
rect 532700 220872 532752 220924
rect 541440 220872 541492 220924
rect 615960 220872 616012 220924
rect 231216 220804 231268 220856
rect 236736 220804 236788 220856
rect 395068 220804 395120 220856
rect 531504 220804 531556 220856
rect 543556 220804 543608 220856
rect 616420 220804 616472 220856
rect 655428 220804 655480 220856
rect 675944 220804 675996 220856
rect 42156 220736 42208 220788
rect 56508 220736 56560 220788
rect 344836 220736 344888 220788
rect 412916 220736 412968 220788
rect 349160 220668 349212 220720
rect 423036 220668 423088 220720
rect 347688 220600 347740 220652
rect 419724 220600 419776 220652
rect 350540 220532 350592 220584
rect 426348 220532 426400 220584
rect 142712 220464 142764 220516
rect 229652 220464 229704 220516
rect 352012 220464 352064 220516
rect 429752 220464 429804 220516
rect 139308 220396 139360 220448
rect 228272 220396 228324 220448
rect 353392 220396 353444 220448
rect 433340 220396 433392 220448
rect 135996 220328 136048 220380
rect 226616 220328 226668 220380
rect 357624 220328 357676 220380
rect 440700 220328 440752 220380
rect 132408 220260 132460 220312
rect 225420 220260 225472 220312
rect 355048 220260 355100 220312
rect 436468 220260 436520 220312
rect 129280 220192 129332 220244
rect 223948 220192 224000 220244
rect 360200 220192 360252 220244
rect 447416 220192 447468 220244
rect 125876 220124 125928 220176
rect 222292 220124 222344 220176
rect 367652 220124 367704 220176
rect 466736 220124 466788 220176
rect 122472 220056 122524 220108
rect 221096 220056 221148 220108
rect 370136 220056 370188 220108
rect 470968 220056 471020 220108
rect 53748 219988 53800 220040
rect 651288 219988 651340 220040
rect 53840 219920 53892 219972
rect 655520 219920 655572 219972
rect 56600 219852 56652 219904
rect 664352 219852 664404 219904
rect 56692 219784 56744 219836
rect 663892 219784 663944 219836
rect 45744 219716 45796 219768
rect 656900 219716 656952 219768
rect 50988 219648 51040 219700
rect 662972 219648 663024 219700
rect 675576 219580 675628 219632
rect 676036 219580 676088 219632
rect 675668 219512 675720 219564
rect 675944 219512 675996 219564
rect 48596 219444 48648 219496
rect 662512 219444 662564 219496
rect 346308 219308 346360 219360
rect 416228 219308 416280 219360
rect 343456 219240 343508 219292
rect 409512 219240 409564 219292
rect 525800 218424 525852 218476
rect 613108 218424 613160 218476
rect 523408 218356 523460 218408
rect 612648 218356 612700 218408
rect 520832 218288 520884 218340
rect 612188 218288 612240 218340
rect 674472 218288 674524 218340
rect 676036 218288 676088 218340
rect 518716 218220 518768 218272
rect 611728 218220 611780 218272
rect 513472 218152 513524 218204
rect 515772 218152 515824 218204
rect 611268 218152 611320 218204
rect 490288 218084 490340 218136
rect 607128 218084 607180 218136
rect 487160 218016 487212 218068
rect 606668 218016 606720 218068
rect 674748 218016 674800 218068
rect 676036 218016 676088 218068
rect 8208 217880 8260 217932
rect 61844 217812 61896 217864
rect 62948 217812 63000 217864
rect 418160 217812 418212 217864
rect 418620 217812 418672 217864
rect 665732 217540 665784 217592
rect 567982 217472 568034 217524
rect 635464 217472 635516 217524
rect 560760 217404 560812 217456
rect 634084 217404 634136 217456
rect 565728 217336 565780 217388
rect 635004 217336 635056 217388
rect 555700 217268 555752 217320
rect 633164 217268 633216 217320
rect 550640 217200 550692 217252
rect 632244 217200 632296 217252
rect 511080 217132 511132 217184
rect 523040 217132 523092 217184
rect 545396 217132 545448 217184
rect 631324 217132 631376 217184
rect 489276 217064 489328 217116
rect 500132 217064 500184 217116
rect 515312 217064 515364 217116
rect 516048 217064 516100 217116
rect 532792 217064 532844 217116
rect 628932 217064 628984 217116
rect 418528 216996 418580 217048
rect 639696 216996 639748 217048
rect 418436 216928 418488 216980
rect 640616 216928 640668 216980
rect 418620 216860 418672 216912
rect 640156 216860 640208 216912
rect 417884 216792 417936 216844
rect 641076 216792 641128 216844
rect 62028 216724 62080 216776
rect 648528 216724 648580 216776
rect 41512 216656 41564 216708
rect 59360 216656 59412 216708
rect 62948 216656 63000 216708
rect 663432 216656 663484 216708
rect 674656 216656 674708 216708
rect 676036 216656 676088 216708
rect 41420 216588 41472 216640
rect 59268 216588 59320 216640
rect 499304 216520 499356 216572
rect 492588 216452 492640 216504
rect 484216 216384 484268 216436
rect 486700 216384 486752 216436
rect 490104 216384 490156 216436
rect 496636 216384 496688 216436
rect 500132 216384 500184 216436
rect 506112 216520 506164 216572
rect 501052 216452 501104 216504
rect 505008 216384 505060 216436
rect 509938 216352 509990 216404
rect 516048 216384 516100 216436
rect 522856 216384 522908 216436
rect 538036 216520 538088 216572
rect 629944 216520 629996 216572
rect 666560 216520 666612 216572
rect 666836 216520 666888 216572
rect 523040 216452 523092 216504
rect 527732 216452 527784 216504
rect 628012 216452 628064 216504
rect 610348 216384 610400 216436
rect 609428 216316 609480 216368
rect 627092 216248 627144 216300
rect 674288 216248 674340 216300
rect 675944 216248 675996 216300
rect 608508 216180 608560 216232
rect 625712 216112 625764 216164
rect 624792 216044 624844 216096
rect 623872 215976 623924 216028
rect 622952 215908 623004 215960
rect 622032 215840 622084 215892
rect 674932 215840 674984 215892
rect 675852 215840 675904 215892
rect 621480 215772 621532 215824
rect 637396 215704 637448 215756
rect 636384 215636 636436 215688
rect 638316 215568 638368 215620
rect 638776 215500 638828 215552
rect 673552 215500 673604 215552
rect 675760 215500 675812 215552
rect 48228 215432 48280 215484
rect 666192 215432 666244 215484
rect 673736 215432 673788 215484
rect 675852 215432 675904 215484
rect 31668 215364 31720 215416
rect 665272 215364 665324 215416
rect 674564 215364 674616 215416
rect 675944 215364 675996 215416
rect 582288 215296 582340 215348
rect 600044 215296 600096 215348
rect 674840 215296 674892 215348
rect 676036 215296 676088 215348
rect 673644 214616 673696 214668
rect 676036 214616 676088 214668
rect 41512 213256 41564 213308
rect 666928 213256 666980 213308
rect 582288 212576 582340 212628
rect 599952 212576 600004 212628
rect 673460 212576 673512 212628
rect 675944 212576 675996 212628
rect 580264 212508 580316 212560
rect 599860 212508 599912 212560
rect 673828 212508 673880 212560
rect 676036 212508 676088 212560
rect 672724 212032 672776 212084
rect 676036 212032 676088 212084
rect 662788 210060 662840 210112
rect 664444 210060 664496 210112
rect 582288 209856 582340 209908
rect 601148 209856 601200 209908
rect 580080 209788 580132 209840
rect 600780 209788 600832 209840
rect 641812 209788 641864 209840
rect 642088 209788 642140 209840
rect 644664 209788 644716 209840
rect 644940 209788 644992 209840
rect 647424 209788 647476 209840
rect 647700 209788 647752 209840
rect 673460 207272 673512 207324
rect 582288 207068 582340 207120
rect 599676 207068 599728 207120
rect 673552 207068 673604 207120
rect 674932 207068 674984 207120
rect 581460 207000 581512 207052
rect 601608 207000 601660 207052
rect 673460 207000 673512 207052
rect 674932 206320 674984 206372
rect 675392 206320 675444 206372
rect 675024 206252 675076 206304
rect 675760 206252 675812 206304
rect 675208 206184 675260 206236
rect 675484 206184 675536 206236
rect 675668 206184 675720 206236
rect 674748 205572 674800 205624
rect 675392 205572 675444 205624
rect 674748 205436 674800 205488
rect 38476 205028 38528 205080
rect 43536 205028 43588 205080
rect 674840 204960 674892 205012
rect 675392 204960 675444 205012
rect 38200 204416 38252 204468
rect 43628 204416 43680 204468
rect 38108 204348 38160 204400
rect 43352 204348 43404 204400
rect 674472 204348 674524 204400
rect 675392 204348 675444 204400
rect 38568 204280 38620 204332
rect 42248 204280 42300 204332
rect 582288 204280 582340 204332
rect 599952 204280 600004 204332
rect 673368 204212 673420 204264
rect 674472 204212 674524 204264
rect 674656 202716 674708 202768
rect 675392 202716 675444 202768
rect 674564 201832 674616 201884
rect 675392 201832 675444 201884
rect 581092 201560 581144 201612
rect 599952 201560 600004 201612
rect 580724 201492 580776 201544
rect 598940 201492 598992 201544
rect 673736 201492 673788 201544
rect 675392 201492 675444 201544
rect 37924 201424 37976 201476
rect 43720 201424 43772 201476
rect 38016 200880 38068 200932
rect 43168 200880 43220 200932
rect 673828 200676 673880 200728
rect 675392 200676 675444 200728
rect 581092 200064 581144 200116
rect 599952 200064 600004 200116
rect 582288 198704 582340 198756
rect 599952 198704 600004 198756
rect 674288 198364 674340 198416
rect 675392 198364 675444 198416
rect 673460 197548 673512 197600
rect 675484 197548 675536 197600
rect 582288 197344 582340 197396
rect 599400 197344 599452 197396
rect 580724 197276 580776 197328
rect 599952 197276 600004 197328
rect 673644 197140 673696 197192
rect 675392 197140 675444 197192
rect 42248 196528 42300 196580
rect 43168 196528 43220 196580
rect 675024 196528 675076 196580
rect 675392 196528 675444 196580
rect 674748 196392 674800 196444
rect 675024 196392 675076 196444
rect 674472 195304 674524 195356
rect 675392 195304 675444 195356
rect 582196 194624 582248 194676
rect 599952 194624 600004 194676
rect 582288 194556 582340 194608
rect 599860 194556 599912 194608
rect 675300 193536 675352 193588
rect 42064 193468 42116 193520
rect 42708 193468 42760 193520
rect 675300 193332 675352 193384
rect 674932 192856 674984 192908
rect 675208 192856 675260 192908
rect 582288 191836 582340 191888
rect 599492 191836 599544 191888
rect 581276 191768 581328 191820
rect 599952 191768 600004 191820
rect 42340 191632 42392 191684
rect 43076 191632 43128 191684
rect 673552 191632 673604 191684
rect 675392 191632 675444 191684
rect 42064 191428 42116 191480
rect 43260 191428 43312 191480
rect 579712 190408 579764 190460
rect 599952 190408 600004 190460
rect 42340 190340 42392 190392
rect 43352 190340 43404 190392
rect 42248 189796 42300 189848
rect 43444 189796 43496 189848
rect 42340 189728 42392 189780
rect 43720 189728 43772 189780
rect 42432 189116 42484 189168
rect 43628 189116 43680 189168
rect 582288 187620 582340 187672
rect 601516 187620 601568 187672
rect 579896 187552 579948 187604
rect 601608 187552 601660 187604
rect 42340 186668 42392 186720
rect 43536 186668 43588 186720
rect 580264 184832 580316 184884
rect 599952 184832 600004 184884
rect 580908 184764 580960 184816
rect 599124 184764 599176 184816
rect 42156 182112 42208 182164
rect 48504 182112 48556 182164
rect 580632 182112 580684 182164
rect 600044 182112 600096 182164
rect 580540 182044 580592 182096
rect 599860 182044 599912 182096
rect 580724 179324 580776 179376
rect 598940 179324 598992 179376
rect 581092 179256 581144 179308
rect 599952 179256 600004 179308
rect 666836 178032 666888 178084
rect 666744 177828 666796 177880
rect 670332 177080 670384 177132
rect 676036 177080 676088 177132
rect 670240 176944 670292 176996
rect 675944 176944 675996 176996
rect 667020 176808 667072 176860
rect 675852 176808 675904 176860
rect 581092 176672 581144 176724
rect 599952 176672 600004 176724
rect 581460 176604 581512 176656
rect 600044 176604 600096 176656
rect 675208 176604 675260 176656
rect 676036 176604 676088 176656
rect 675024 176332 675076 176384
rect 676036 176332 676088 176384
rect 673368 175992 673420 176044
rect 675944 175992 675996 176044
rect 674748 175516 674800 175568
rect 676036 175516 676088 175568
rect 581644 173884 581696 173936
rect 599952 173884 600004 173936
rect 674748 173884 674800 173936
rect 676036 173884 676088 173936
rect 579712 173816 579764 173868
rect 599860 173816 599912 173868
rect 582288 173748 582340 173800
rect 600136 173748 600188 173800
rect 673552 172864 673604 172916
rect 676036 172864 676088 172916
rect 674288 172048 674340 172100
rect 675944 172048 675996 172100
rect 674840 171232 674892 171284
rect 676036 171232 676088 171284
rect 582104 171164 582156 171216
rect 599952 171164 600004 171216
rect 674564 171164 674616 171216
rect 675944 171164 675996 171216
rect 579896 171096 579948 171148
rect 599492 171096 599544 171148
rect 674656 171096 674708 171148
rect 676036 171096 676088 171148
rect 582012 171028 582064 171080
rect 599768 171028 599820 171080
rect 580540 170960 580592 171012
rect 599676 170960 599728 171012
rect 666652 170144 666704 170196
rect 673736 170008 673788 170060
rect 675944 170008 675996 170060
rect 666652 169940 666704 169992
rect 674932 169600 674984 169652
rect 676036 169600 676088 169652
rect 673644 169192 673696 169244
rect 675944 169192 675996 169244
rect 675024 168920 675076 168972
rect 676036 168920 676088 168972
rect 674472 168580 674524 168632
rect 675944 168580 675996 168632
rect 580448 168512 580500 168564
rect 599952 168512 600004 168564
rect 673828 168512 673880 168564
rect 676036 168512 676088 168564
rect 579804 168444 579856 168496
rect 599860 168444 599912 168496
rect 580264 168376 580316 168428
rect 599492 168376 599544 168428
rect 580172 168308 580224 168360
rect 600412 168308 600464 168360
rect 671988 167016 672040 167068
rect 676036 167016 676088 167068
rect 582288 165724 582340 165776
rect 600044 165724 600096 165776
rect 582196 165656 582248 165708
rect 599952 165656 600004 165708
rect 581276 165588 581328 165640
rect 599492 165588 599544 165640
rect 581828 165520 581880 165572
rect 601332 165520 601384 165572
rect 673460 164840 673512 164892
rect 673736 164840 673788 164892
rect 673828 164568 673880 164620
rect 674288 164568 674340 164620
rect 674288 164432 674340 164484
rect 674472 164432 674524 164484
rect 675116 164432 675168 164484
rect 675392 164432 675444 164484
rect 674472 164296 674524 164348
rect 674656 164296 674708 164348
rect 674656 164160 674708 164212
rect 674932 164160 674984 164212
rect 675024 163956 675076 164008
rect 675668 163956 675720 164008
rect 580080 162936 580132 162988
rect 600044 162936 600096 162988
rect 581184 162868 581236 162920
rect 599952 162868 600004 162920
rect 675760 161168 675812 161220
rect 666836 160964 666888 161016
rect 675392 160964 675444 161016
rect 582104 160216 582156 160268
rect 599952 160216 600004 160268
rect 581644 160148 581696 160200
rect 599860 160148 599912 160200
rect 675024 160148 675076 160200
rect 675300 160148 675352 160200
rect 581736 160080 581788 160132
rect 600044 160080 600096 160132
rect 675024 160012 675076 160064
rect 674748 159332 674800 159384
rect 675484 159332 675536 159384
rect 674656 158040 674708 158092
rect 675300 158040 675352 158092
rect 674840 157700 674892 157752
rect 675484 157700 675536 157752
rect 581092 157496 581144 157548
rect 599860 157496 599912 157548
rect 580908 157428 580960 157480
rect 599952 157428 600004 157480
rect 580632 157360 580684 157412
rect 600044 157360 600096 157412
rect 674472 156884 674524 156936
rect 675392 156884 675444 156936
rect 674932 155864 674984 155916
rect 675484 155864 675536 155916
rect 674288 155796 674340 155848
rect 675300 155796 675352 155848
rect 580724 154640 580776 154692
rect 599952 154640 600004 154692
rect 580540 154572 580592 154624
rect 599860 154572 599912 154624
rect 673828 153348 673880 153400
rect 675392 153348 675444 153400
rect 673644 152192 673696 152244
rect 675300 152192 675352 152244
rect 582288 151920 582340 151972
rect 599860 151920 599912 151972
rect 581828 151852 581880 151904
rect 599952 151852 600004 151904
rect 580816 151784 580868 151836
rect 600044 151784 600096 151836
rect 673736 151512 673788 151564
rect 675300 151512 675352 151564
rect 675116 150424 675168 150476
rect 675300 150424 675352 150476
rect 673460 150356 673512 150408
rect 675392 150356 675444 150408
rect 582012 149200 582064 149252
rect 600044 149200 600096 149252
rect 581552 149132 581604 149184
rect 599860 149132 599912 149184
rect 581368 149064 581420 149116
rect 599952 149064 600004 149116
rect 673552 148520 673604 148572
rect 675392 148520 675444 148572
rect 674564 146684 674616 146736
rect 675392 146684 675444 146736
rect 582196 146344 582248 146396
rect 599860 146344 599912 146396
rect 581460 146276 581512 146328
rect 599952 146276 600004 146328
rect 581920 143692 581972 143744
rect 599860 143692 599912 143744
rect 581736 143624 581788 143676
rect 599952 143624 600004 143676
rect 581276 143556 581328 143608
rect 600044 143556 600096 143608
rect 581644 140904 581696 140956
rect 599952 140904 600004 140956
rect 581000 140836 581052 140888
rect 600044 140836 600096 140888
rect 581184 140768 581236 140820
rect 599860 140768 599912 140820
rect 581092 138116 581144 138168
rect 599952 138116 600004 138168
rect 579712 138048 579764 138100
rect 600044 138048 600096 138100
rect 579896 137980 579948 138032
rect 599860 137980 599912 138032
rect 580080 135328 580132 135380
rect 599860 135328 599912 135380
rect 580172 135260 580224 135312
rect 599952 135260 600004 135312
rect 670148 132880 670200 132932
rect 676220 132880 676272 132932
rect 670056 132744 670108 132796
rect 676128 132744 676180 132796
rect 580908 132608 580960 132660
rect 599952 132608 600004 132660
rect 669964 132608 670016 132660
rect 676036 132608 676088 132660
rect 580264 132540 580316 132592
rect 599860 132540 599912 132592
rect 579988 132472 580040 132524
rect 600044 132472 600096 132524
rect 675208 132404 675260 132456
rect 676036 132404 676088 132456
rect 672172 131656 672224 131708
rect 673276 131656 673328 131708
rect 676036 131656 676088 131708
rect 673368 131452 673420 131504
rect 676220 131452 676272 131504
rect 672264 130840 672316 130892
rect 676036 130840 676088 130892
rect 671896 130024 671948 130076
rect 672080 130024 672132 130076
rect 676036 130024 676088 130076
rect 580356 129888 580408 129940
rect 600044 129888 600096 129940
rect 580632 129820 580684 129872
rect 599860 129820 599912 129872
rect 580448 129752 580500 129804
rect 599952 129752 600004 129804
rect 672356 129412 672408 129464
rect 673092 129412 673144 129464
rect 676220 129412 676272 129464
rect 674748 127712 674800 127764
rect 676036 127712 676088 127764
rect 673552 127304 673604 127356
rect 675944 127304 675996 127356
rect 580724 127032 580776 127084
rect 599860 127032 599912 127084
rect 673828 127032 673880 127084
rect 675944 127032 675996 127084
rect 580540 126964 580592 127016
rect 599952 126964 600004 127016
rect 674840 126964 674892 127016
rect 676036 126964 676088 127016
rect 674656 126488 674708 126540
rect 676036 126488 676088 126540
rect 673644 124856 673696 124908
rect 675944 124856 675996 124908
rect 673736 124448 673788 124500
rect 675944 124448 675996 124500
rect 582288 124312 582340 124364
rect 599860 124312 599912 124364
rect 581828 124244 581880 124296
rect 599768 124244 599820 124296
rect 674932 124244 674984 124296
rect 675944 124244 675996 124296
rect 580816 124176 580868 124228
rect 599952 124176 600004 124228
rect 675024 124176 675076 124228
rect 676036 124176 676088 124228
rect 582196 121592 582248 121644
rect 599952 121592 600004 121644
rect 672448 121592 672500 121644
rect 676220 121592 676272 121644
rect 582012 121524 582064 121576
rect 599860 121524 599912 121576
rect 674288 121524 674340 121576
rect 675944 121524 675996 121576
rect 582104 121456 582156 121508
rect 600044 121456 600096 121508
rect 674472 121456 674524 121508
rect 676036 121456 676088 121508
rect 674932 121388 674984 121440
rect 674748 121320 674800 121372
rect 674748 121116 674800 121168
rect 674932 121116 674984 121168
rect 583668 118804 583720 118856
rect 599952 118804 600004 118856
rect 581920 118736 581972 118788
rect 600044 118736 600096 118788
rect 581460 118668 581512 118720
rect 599860 118668 599912 118720
rect 581736 116016 581788 116068
rect 599952 116016 600004 116068
rect 581276 115948 581328 116000
rect 600044 115948 600096 116000
rect 666744 115880 666796 115932
rect 675392 115880 675444 115932
rect 675024 114996 675076 115048
rect 675300 114996 675352 115048
rect 674748 114316 674800 114368
rect 675300 114316 675352 114368
rect 674840 113704 674892 113756
rect 675300 113704 675352 113756
rect 581644 113228 581696 113280
rect 599952 113228 600004 113280
rect 581368 113160 581420 113212
rect 599860 113160 599912 113212
rect 581552 110508 581604 110560
rect 599860 110508 599912 110560
rect 581000 110440 581052 110492
rect 599952 110440 600004 110492
rect 673736 110032 673788 110084
rect 675116 110032 675168 110084
rect 673828 108196 673880 108248
rect 675392 108196 675444 108248
rect 581184 107652 581236 107704
rect 599308 107652 599360 107704
rect 674472 107516 674524 107568
rect 675392 107516 675444 107568
rect 674288 106360 674340 106412
rect 675392 106360 675444 106412
rect 673644 106292 673696 106344
rect 675116 106292 675168 106344
rect 581092 104864 581144 104916
rect 599952 104864 600004 104916
rect 673552 104524 673604 104576
rect 675116 104524 675168 104576
rect 657728 99764 657780 99816
rect 660902 99764 660954 99816
rect 580908 99356 580960 99408
rect 599952 99356 600004 99408
rect 633072 96568 633124 96620
rect 635280 96568 635332 96620
rect 636292 96568 636344 96620
rect 640984 96568 641036 96620
rect 655980 96568 656032 96620
rect 659568 96568 659620 96620
rect 661868 96568 661920 96620
rect 663064 96568 663116 96620
rect 633808 96500 633860 96552
rect 636384 96500 636436 96552
rect 637028 96500 637080 96552
rect 642364 96500 642416 96552
rect 654692 96500 654744 96552
rect 658280 96500 658332 96552
rect 659108 96500 659160 96552
rect 662512 96500 662564 96552
rect 634452 96432 634504 96484
rect 637580 96432 637632 96484
rect 635740 96364 635792 96416
rect 639880 96364 639932 96416
rect 647516 96296 647568 96348
rect 653956 96296 654008 96348
rect 631140 96024 631192 96076
rect 632106 96024 632158 96076
rect 632428 96024 632480 96076
rect 634406 96024 634458 96076
rect 635096 96024 635148 96076
rect 639006 96024 639058 96076
rect 631784 95888 631836 95940
rect 632980 95888 633032 95940
rect 640064 95888 640116 95940
rect 646044 95888 646096 95940
rect 638868 95820 638920 95872
rect 645860 95820 645912 95872
rect 646136 95820 646188 95872
rect 663524 95820 663576 95872
rect 614764 95752 614816 95804
rect 616144 95684 616196 95736
rect 622492 95684 622544 95736
rect 621296 95616 621348 95668
rect 623320 95616 623372 95668
rect 604460 95548 604512 95600
rect 606392 95548 606444 95600
rect 607496 95548 607548 95600
rect 608968 95548 609020 95600
rect 610256 95548 610308 95600
rect 611544 95548 611596 95600
rect 618260 95548 618312 95600
rect 620100 95548 620152 95600
rect 621480 95548 621532 95600
rect 622676 95548 622728 95600
rect 621204 95480 621256 95532
rect 622032 95480 622084 95532
rect 620008 95412 620060 95464
rect 623412 95412 623464 95464
rect 591948 95344 592000 95396
rect 610348 95344 610400 95396
rect 617432 95344 617484 95396
rect 622124 95344 622176 95396
rect 589188 95276 589240 95328
rect 612188 95276 612240 95328
rect 575664 95208 575716 95260
rect 607680 95208 607732 95260
rect 639604 95752 639656 95804
rect 637488 95684 637540 95736
rect 640524 95684 640576 95736
rect 640892 95684 640944 95736
rect 645952 95684 646004 95736
rect 641628 95616 641680 95668
rect 642824 95616 642876 95668
rect 638316 95548 638368 95600
rect 642272 95548 642324 95600
rect 642916 95548 642968 95600
rect 642732 95480 642784 95532
rect 652024 95752 652076 95804
rect 661960 95752 662012 95804
rect 652668 95616 652720 95668
rect 663892 95616 663944 95668
rect 651840 95548 651892 95600
rect 653404 95548 653456 95600
rect 656992 95548 657044 95600
rect 659200 95548 659252 95600
rect 660580 95480 660632 95532
rect 661408 95480 661460 95532
rect 646044 95412 646096 95464
rect 646780 95412 646832 95464
rect 648620 95344 648672 95396
rect 650736 95344 650788 95396
rect 663432 95344 663484 95396
rect 657084 95208 657136 95260
rect 657912 95208 657964 95260
rect 665180 95140 665232 95192
rect 619364 95072 619416 95124
rect 623504 95072 623556 95124
rect 643468 95072 643520 95124
rect 644848 95072 644900 95124
rect 648804 94936 648856 94988
rect 650092 94936 650144 94988
rect 616788 94868 616840 94920
rect 623228 94868 623280 94920
rect 648896 94800 648948 94852
rect 649448 94800 649500 94852
rect 618720 94732 618772 94784
rect 623320 94732 623372 94784
rect 646596 94732 646648 94784
rect 648160 94732 648212 94784
rect 653312 94732 653364 94784
rect 663800 94732 663852 94784
rect 656624 94664 656676 94716
rect 663708 94664 663760 94716
rect 657268 94596 657320 94648
rect 663616 94596 663668 94648
rect 656900 94528 656952 94580
rect 658556 94528 658608 94580
rect 648068 94460 648120 94512
rect 659844 94460 659896 94512
rect 660396 94460 660448 94512
rect 643560 94188 643612 94240
rect 618076 94120 618128 94172
rect 623136 94120 623188 94172
rect 644204 94052 644256 94104
rect 654048 94052 654100 94104
rect 649356 93984 649408 94036
rect 656900 93984 656952 94036
rect 607220 93848 607272 93900
rect 612924 93848 612976 93900
rect 644756 93848 644808 93900
rect 653128 93848 653180 93900
rect 613016 93644 613068 93696
rect 614856 93644 614908 93696
rect 663248 91060 663300 91112
rect 663892 91060 663944 91112
rect 657084 88816 657136 88868
rect 658004 88816 658056 88868
rect 659476 88748 659528 88800
rect 663156 88748 663208 88800
rect 648620 85484 648672 85536
rect 657176 85484 657228 85536
rect 651840 85416 651892 85468
rect 658832 85416 658884 85468
rect 648896 85348 648948 85400
rect 660672 85348 660724 85400
rect 648804 85280 648856 85332
rect 657728 85280 657780 85332
rect 643468 85212 643520 85264
rect 660120 85212 660172 85264
rect 646596 85144 646648 85196
rect 661408 85144 661460 85196
rect 583760 84600 583812 84652
rect 600320 84600 600372 84652
rect 582196 84532 582248 84584
rect 600412 84532 600464 84584
rect 582288 84464 582340 84516
rect 600688 84464 600740 84516
rect 581828 84396 581880 84448
rect 600504 84396 600556 84448
rect 582012 84328 582064 84380
rect 600780 84328 600832 84380
rect 582104 84260 582156 84312
rect 600872 84260 600924 84312
rect 580724 84192 580776 84244
rect 600228 84192 600280 84244
rect 580816 84124 580868 84176
rect 600596 84124 600648 84176
rect 596916 83104 596968 83156
rect 607220 83104 607272 83156
rect 597468 82832 597520 82884
rect 604460 82832 604512 82884
rect 579620 82628 579672 82680
rect 583668 82628 583720 82680
rect 600228 80112 600280 80164
rect 612832 80112 612884 80164
rect 575848 78616 575900 78668
rect 596916 78616 596968 78668
rect 575756 74944 575808 74996
rect 589188 74944 589240 74996
rect 583668 73108 583720 73160
rect 610164 73108 610216 73160
rect 586428 72632 586480 72684
rect 591948 72632 592000 72684
rect 594708 66240 594760 66292
rect 600228 66240 600280 66292
rect 602988 66240 603040 66292
rect 610348 66240 610400 66292
rect 579620 66172 579672 66224
rect 583760 66172 583812 66224
rect 587900 62296 587952 62348
rect 597468 62296 597520 62348
rect 581644 53184 581696 53236
rect 587900 53184 587952 53236
rect 145380 52436 145432 52488
rect 198648 52436 198700 52488
rect 346860 52368 346912 52420
rect 642916 52368 642968 52420
rect 52092 51076 52144 51128
rect 213828 51076 213880 51128
rect 346492 51076 346544 51128
rect 198648 51008 198700 51060
rect 207020 51008 207072 51060
rect 631876 51008 631928 51060
rect 478144 48424 478196 48476
rect 526168 48424 526220 48476
rect 412640 48356 412692 48408
rect 506388 48356 506440 48408
rect 571800 48356 571852 48408
rect 581644 48356 581696 48408
rect 150348 48288 150400 48340
rect 218060 48288 218112 48340
rect 281448 48288 281500 48340
rect 502248 48288 502300 48340
rect 549260 48288 549312 48340
rect 594708 48288 594760 48340
rect 568580 47200 568632 47252
rect 575756 47200 575808 47252
rect 52276 47064 52328 47116
rect 150348 47064 150400 47116
rect 577964 47064 578016 47116
rect 583668 47064 583720 47116
rect 218060 46860 218112 46912
rect 642640 46860 642692 46912
rect 460664 45976 460716 46028
rect 610256 45976 610308 46028
rect 367100 45908 367152 45960
rect 607312 45908 607364 45960
rect 311900 45840 311952 45892
rect 607588 45840 607640 45892
rect 230940 45772 230992 45824
rect 613016 45772 613068 45824
rect 85120 45704 85172 45756
rect 475568 45704 475620 45756
rect 230388 45636 230440 45688
rect 621388 45636 621440 45688
rect 233148 45568 233200 45620
rect 642824 45568 642876 45620
rect 212448 45500 212500 45552
rect 639328 45500 639380 45552
rect 194416 44072 194468 44124
rect 661132 44072 661184 44124
rect 365168 43868 365220 43920
rect 367100 43868 367152 43920
rect 310428 43800 310480 43852
rect 311900 43800 311952 43852
rect 230480 43460 230532 43512
rect 618260 43460 618312 43512
rect 230664 43392 230716 43444
rect 621480 43392 621532 43444
rect 230848 43324 230900 43376
rect 621204 43324 621256 43376
rect 230572 43256 230624 43308
rect 621112 43256 621164 43308
rect 230756 43188 230808 43240
rect 621296 43188 621348 43240
rect 226248 43120 226300 43172
rect 622492 43120 622544 43172
rect 223488 43052 223540 43104
rect 622308 43052 622360 43104
rect 52184 42712 52236 42764
rect 215300 42712 215352 42764
rect 529664 42712 529716 42764
rect 543004 42712 543056 42764
rect 475476 42576 475528 42628
rect 513932 41964 513984 42016
rect 520372 41964 520424 42016
rect 405832 41896 405884 41948
rect 426348 41896 426400 41948
rect 514024 41896 514076 41948
rect 514852 41896 514904 41948
rect 426348 41420 426400 41472
rect 607496 41420 607548 41472
rect 506388 41352 506440 41404
rect 513288 41352 513340 41404
rect 530400 41352 530452 41404
rect 602988 41352 603040 41404
rect 530308 41284 530360 41336
rect 571800 41284 571852 41336
rect 475568 38564 475620 38616
rect 514024 38564 514076 38616
rect 502340 38496 502392 38548
rect 513932 38496 513984 38548
rect 213184 24760 213236 24812
rect 213828 24760 213880 24812
rect 224592 22992 224644 23044
rect 226248 22992 226300 23044
rect 221740 22516 221792 22568
rect 223488 22516 223540 22568
rect 229376 6468 229428 6520
rect 233148 6468 233200 6520
<< metal2 >>
rect 483570 1004728 483626 1004737
rect 483570 1004663 483572 1004672
rect 483624 1004663 483626 1004672
rect 483572 1004634 483624 1004640
rect 703694 897668 703722 897804
rect 704154 897668 704182 897804
rect 704614 897668 704642 897804
rect 705074 897668 705102 897804
rect 705534 897668 705562 897804
rect 705994 897668 706022 897804
rect 706454 897668 706482 897804
rect 706914 897668 706942 897804
rect 707374 897668 707402 897804
rect 707834 897668 707862 897804
rect 708294 897668 708322 897804
rect 708754 897668 708782 897804
rect 709214 897668 709242 897804
rect 676034 897152 676090 897161
rect 676034 897087 676090 897096
rect 676048 897054 676076 897087
rect 655520 897048 655572 897054
rect 655520 896990 655572 896996
rect 676036 897048 676088 897054
rect 676036 896990 676088 896996
rect 655428 894532 655480 894538
rect 655428 894474 655480 894480
rect 655440 866561 655468 894474
rect 655532 867649 655560 896990
rect 675942 896744 675998 896753
rect 675942 896679 675998 896688
rect 675850 894704 675906 894713
rect 673368 894668 673420 894674
rect 675850 894639 675852 894648
rect 673368 894610 673420 894616
rect 675904 894639 675906 894648
rect 675852 894610 675904 894616
rect 670516 894464 670568 894470
rect 670516 894406 670568 894412
rect 655704 894396 655756 894402
rect 655704 894338 655756 894344
rect 655612 883312 655664 883318
rect 655612 883254 655664 883260
rect 655518 867640 655574 867649
rect 655518 867575 655574 867584
rect 655426 866552 655482 866561
rect 655426 866487 655482 866496
rect 655624 865337 655652 883254
rect 655716 868873 655744 894338
rect 670424 893036 670476 893042
rect 670424 892978 670476 892984
rect 655796 872228 655848 872234
rect 655796 872170 655848 872176
rect 655702 868864 655758 868873
rect 655702 868799 655758 868808
rect 655610 865328 655666 865337
rect 655610 865263 655666 865272
rect 655808 863841 655836 872170
rect 656808 863864 656860 863870
rect 655794 863832 655850 863841
rect 656808 863806 656860 863812
rect 655794 863767 655850 863776
rect 656820 862617 656848 863806
rect 656806 862608 656862 862617
rect 656806 862543 656862 862552
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 41786 817728 41842 817737
rect 41786 817663 41788 817672
rect 41840 817663 41842 817672
rect 50988 817692 51040 817698
rect 41788 817634 41840 817640
rect 50988 817634 51040 817640
rect 41786 817320 41842 817329
rect 41786 817255 41788 817264
rect 41840 817255 41842 817264
rect 48320 817284 48372 817290
rect 41788 817226 41840 817232
rect 48320 817226 48372 817232
rect 41786 816912 41842 816921
rect 41786 816847 41842 816856
rect 41800 814609 41828 816847
rect 44610 816140 44638 816142
rect 44594 816130 44654 816140
rect 44594 816060 44654 816070
rect 43626 815280 43682 815289
rect 43626 815215 43682 815224
rect 41786 814600 41842 814609
rect 41786 814535 41842 814544
rect 43442 813240 43498 813249
rect 43442 813175 43498 813184
rect 42706 812832 42762 812841
rect 42706 812767 42762 812776
rect 42246 811200 42302 811209
rect 42246 811135 42302 811144
rect 41970 809160 42026 809169
rect 41970 809095 42026 809104
rect 41878 808752 41934 808761
rect 41878 808687 41934 808696
rect 41786 808344 41842 808353
rect 41786 808279 41788 808288
rect 41840 808279 41842 808288
rect 41788 808250 41840 808256
rect 41786 807528 41842 807537
rect 41786 807463 41842 807472
rect 41800 806313 41828 807463
rect 41786 806304 41842 806313
rect 41786 806239 41842 806248
rect 41892 805934 41920 808687
rect 41880 805928 41932 805934
rect 41880 805870 41932 805876
rect 41984 804302 42012 809095
rect 41972 804296 42024 804302
rect 41972 804238 42024 804244
rect 42260 799459 42288 811135
rect 42614 809568 42670 809577
rect 42614 809503 42670 809512
rect 42338 806304 42394 806313
rect 42338 806239 42394 806248
rect 42352 806002 42380 806239
rect 42340 805996 42392 806002
rect 42340 805938 42392 805944
rect 42340 800488 42392 800494
rect 42340 800430 42392 800436
rect 42182 799431 42288 799459
rect 42248 799332 42300 799338
rect 42248 799274 42300 799280
rect 42260 797619 42288 799274
rect 42182 797591 42288 797619
rect 42352 796974 42380 800430
rect 42182 796946 42380 796974
rect 42628 796890 42656 809503
rect 42720 799338 42748 812767
rect 43074 812424 43130 812433
rect 43074 812359 43130 812368
rect 42798 812016 42854 812025
rect 42798 811951 42854 811960
rect 42708 799332 42760 799338
rect 42708 799274 42760 799280
rect 42812 799218 42840 811951
rect 42890 811608 42946 811617
rect 42890 811543 42946 811552
rect 42720 799190 42840 799218
rect 42340 796884 42392 796890
rect 42340 796826 42392 796832
rect 42616 796884 42668 796890
rect 42616 796826 42668 796832
rect 42352 795779 42380 796826
rect 42182 795751 42380 795779
rect 42182 795110 42380 795138
rect 42248 795048 42300 795054
rect 41878 795016 41934 795025
rect 42248 794990 42300 794996
rect 41878 794951 41934 794960
rect 41892 794580 41920 794951
rect 42156 794300 42208 794306
rect 42156 794242 42208 794248
rect 42168 793900 42196 794242
rect 42156 793824 42208 793830
rect 42156 793766 42208 793772
rect 42168 793288 42196 793766
rect 42260 792758 42288 794990
rect 42182 792730 42288 792758
rect 42248 792668 42300 792674
rect 42248 792610 42300 792616
rect 42156 790696 42208 790702
rect 42156 790638 42208 790644
rect 42168 790228 42196 790638
rect 42156 790152 42208 790158
rect 42156 790094 42208 790100
rect 42168 789616 42196 790094
rect 42156 789268 42208 789274
rect 42156 789210 42208 789216
rect 42168 788936 42196 789210
rect 42156 788860 42208 788866
rect 42156 788802 42208 788808
rect 42168 788392 42196 788802
rect 42156 787024 42208 787030
rect 42156 786966 42208 786972
rect 42168 786556 42196 786966
rect 42064 786276 42116 786282
rect 42064 786218 42116 786224
rect 42076 785944 42104 786218
rect 42260 785278 42288 792610
rect 42352 791874 42380 795110
rect 42720 794918 42748 799190
rect 42904 795054 42932 811543
rect 42892 795048 42944 795054
rect 42892 794990 42944 794996
rect 42708 794912 42760 794918
rect 42708 794854 42760 794860
rect 42892 794912 42944 794918
rect 42892 794854 42944 794860
rect 42352 791846 42472 791874
rect 42340 789404 42392 789410
rect 42340 789346 42392 789352
rect 42182 785250 42288 785278
rect 42352 784734 42380 789346
rect 42444 789342 42472 791846
rect 42432 789336 42484 789342
rect 42432 789278 42484 789284
rect 42904 788866 42932 794854
rect 43088 792674 43116 812359
rect 43352 805928 43404 805934
rect 43352 805870 43404 805876
rect 43260 804296 43312 804302
rect 43260 804238 43312 804244
rect 43272 794306 43300 804238
rect 43260 794300 43312 794306
rect 43260 794242 43312 794248
rect 43076 792668 43128 792674
rect 43076 792610 43128 792616
rect 43364 790702 43392 805870
rect 43352 790696 43404 790702
rect 43352 790638 43404 790644
rect 42892 788860 42944 788866
rect 42892 788802 42944 788808
rect 43456 787030 43484 813175
rect 43536 808308 43588 808314
rect 43536 808250 43588 808256
rect 43548 793830 43576 808250
rect 43536 793824 43588 793830
rect 43536 793766 43588 793772
rect 43444 787024 43496 787030
rect 43444 786966 43496 786972
rect 42182 784706 42380 784734
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 41512 774784 41564 774790
rect 41510 774752 41512 774761
rect 41564 774752 41566 774761
rect 41510 774687 41566 774696
rect 41510 773936 41566 773945
rect 41510 773871 41512 773880
rect 41564 773871 41566 773880
rect 41512 773842 41564 773848
rect 41510 773528 41566 773537
rect 41510 773463 41512 773472
rect 41564 773463 41566 773472
rect 41512 773434 41564 773440
rect 43640 772449 43668 815215
rect 43718 810792 43774 810801
rect 43718 810727 43774 810736
rect 43732 786282 43760 810727
rect 43810 810384 43866 810393
rect 43810 810319 43866 810328
rect 43824 789274 43852 810319
rect 43902 809976 43958 809985
rect 43902 809911 43958 809920
rect 43916 790158 43944 809911
rect 43904 790152 43956 790158
rect 43904 790094 43956 790100
rect 43812 789268 43864 789274
rect 43812 789210 43864 789216
rect 43720 786276 43772 786282
rect 43720 786218 43772 786224
rect 44610 773324 44638 816060
rect 44702 814478 44730 814482
rect 44686 814468 44746 814478
rect 44686 814398 44746 814408
rect 44594 773314 44654 773324
rect 44594 773244 44654 773254
rect 44610 773236 44638 773244
rect 44594 772930 44654 772940
rect 44594 772860 44654 772870
rect 43626 772440 43682 772449
rect 43626 772375 43682 772384
rect 43718 772032 43774 772041
rect 43718 771967 43774 771976
rect 42338 769584 42394 769593
rect 42338 769519 42394 769528
rect 38290 767816 38346 767825
rect 38290 767751 38346 767760
rect 38198 767408 38254 767417
rect 38198 767343 38254 767352
rect 38212 761734 38240 767343
rect 38304 764522 38332 767751
rect 41510 764960 41566 764969
rect 41510 764895 41566 764904
rect 38566 764552 38622 764561
rect 38292 764516 38344 764522
rect 38566 764487 38622 764496
rect 38292 764458 38344 764464
rect 38200 761728 38252 761734
rect 38200 761670 38252 761676
rect 38580 759014 38608 764487
rect 41524 759354 41552 764895
rect 42248 764516 42300 764522
rect 42248 764458 42300 764464
rect 41602 764144 41658 764153
rect 41602 764079 41658 764088
rect 41616 762929 41644 764079
rect 41602 762920 41658 762929
rect 41602 762855 41604 762864
rect 41656 762855 41658 762864
rect 41604 762826 41656 762832
rect 42156 761728 42208 761734
rect 42156 761670 42208 761676
rect 41512 759348 41564 759354
rect 41512 759290 41564 759296
rect 38568 759008 38620 759014
rect 38568 758950 38620 758956
rect 42168 757042 42196 761670
rect 42156 757036 42208 757042
rect 42156 756978 42208 756984
rect 42260 756786 42288 764458
rect 42168 756758 42288 756786
rect 42168 756228 42196 756758
rect 42248 756288 42300 756294
rect 42248 756230 42300 756236
rect 42156 754928 42208 754934
rect 42156 754870 42208 754876
rect 42168 754392 42196 754870
rect 42168 753370 42196 753780
rect 42156 753364 42208 753370
rect 42156 753306 42208 753312
rect 42156 753092 42208 753098
rect 42156 753034 42208 753040
rect 42168 752556 42196 753034
rect 42168 751890 42196 751944
rect 42260 751890 42288 756230
rect 42352 754934 42380 769519
rect 43626 769176 43682 769185
rect 43626 769111 43682 769120
rect 43074 768768 43130 768777
rect 43074 768703 43130 768712
rect 42706 768360 42762 768369
rect 42706 768295 42762 768304
rect 42432 767440 42484 767446
rect 42484 767388 42605 767394
rect 42432 767382 42605 767388
rect 42444 767366 42605 767382
rect 42430 765504 42486 765513
rect 42430 765439 42486 765448
rect 42444 757518 42472 765439
rect 42720 759150 42748 768295
rect 42708 759144 42760 759150
rect 42708 759086 42760 759092
rect 42708 759008 42760 759014
rect 42708 758950 42760 758956
rect 42432 757512 42484 757518
rect 42432 757454 42484 757460
rect 42340 754928 42392 754934
rect 42340 754870 42392 754876
rect 42340 754316 42392 754322
rect 42340 754258 42392 754264
rect 42168 751862 42288 751890
rect 42248 751800 42300 751806
rect 42248 751742 42300 751748
rect 42260 751383 42288 751742
rect 42182 751355 42288 751383
rect 42248 751256 42300 751262
rect 42248 751198 42300 751204
rect 42156 751120 42208 751126
rect 42156 751062 42208 751068
rect 42168 750720 42196 751062
rect 42064 750644 42116 750650
rect 42064 750586 42116 750592
rect 42076 750108 42104 750586
rect 42260 749543 42288 751198
rect 42182 749515 42288 749543
rect 42248 749420 42300 749426
rect 42248 749362 42300 749368
rect 42156 747516 42208 747522
rect 42156 747458 42208 747464
rect 42168 747048 42196 747458
rect 42260 746415 42288 749362
rect 42182 746387 42288 746415
rect 42248 746292 42300 746298
rect 42248 746234 42300 746240
rect 42260 745770 42288 746234
rect 42182 745742 42288 745770
rect 42352 745226 42380 754258
rect 42720 751806 42748 758950
rect 43088 754322 43116 768703
rect 43166 766320 43222 766329
rect 43166 766255 43222 766264
rect 43076 754316 43128 754322
rect 43076 754258 43128 754264
rect 43180 754254 43208 766255
rect 43258 765912 43314 765921
rect 43258 765847 43314 765856
rect 43168 754248 43220 754254
rect 43168 754190 43220 754196
rect 43272 754066 43300 765847
rect 43536 759348 43588 759354
rect 43536 759290 43588 759296
rect 43352 759144 43404 759150
rect 43352 759086 43404 759092
rect 43088 754038 43300 754066
rect 42708 751800 42760 751806
rect 42708 751742 42760 751748
rect 43088 751126 43116 754038
rect 43168 753976 43220 753982
rect 43168 753918 43220 753924
rect 43180 753098 43208 753918
rect 43260 753364 43312 753370
rect 43260 753306 43312 753312
rect 43168 753092 43220 753098
rect 43168 753034 43220 753040
rect 43076 751120 43128 751126
rect 43076 751062 43128 751068
rect 43272 747930 43300 753306
rect 43364 751262 43392 759086
rect 43352 751256 43404 751262
rect 43352 751198 43404 751204
rect 43352 751120 43404 751126
rect 43352 751062 43404 751068
rect 43260 747924 43312 747930
rect 43260 747866 43312 747872
rect 42182 745198 42380 745226
rect 42432 745272 42484 745278
rect 42432 745214 42484 745220
rect 42340 745136 42392 745142
rect 42340 745078 42392 745084
rect 42352 743390 42380 745078
rect 42182 743362 42380 743390
rect 42340 743300 42392 743306
rect 42340 743242 42392 743248
rect 42156 743096 42208 743102
rect 42156 743038 42208 743044
rect 42168 742696 42196 743038
rect 42352 742098 42380 743242
rect 42182 742070 42380 742098
rect 42444 741554 42472 745214
rect 43364 745142 43392 751062
rect 43548 750650 43576 759290
rect 43640 757654 43668 769111
rect 43628 757648 43680 757654
rect 43628 757590 43680 757596
rect 43628 757512 43680 757518
rect 43628 757454 43680 757460
rect 43536 750644 43588 750650
rect 43536 750586 43588 750592
rect 43640 750530 43668 757454
rect 43548 750502 43668 750530
rect 43548 747522 43576 750502
rect 43732 747974 43760 771967
rect 44086 769992 44142 770001
rect 44086 769927 44142 769936
rect 43902 767136 43958 767145
rect 43902 767071 43958 767080
rect 43810 766728 43866 766737
rect 43810 766663 43866 766672
rect 43824 749426 43852 766663
rect 43916 757790 43944 767071
rect 43904 757784 43956 757790
rect 43904 757726 43956 757732
rect 43904 757648 43956 757654
rect 43904 757590 43956 757596
rect 43812 749420 43864 749426
rect 43812 749362 43864 749368
rect 43640 747946 43760 747974
rect 43536 747516 43588 747522
rect 43536 747458 43588 747464
rect 43352 745136 43404 745142
rect 43352 745078 43404 745084
rect 42182 741526 42472 741554
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 43640 731134 43668 747946
rect 43916 743306 43944 757590
rect 44100 751126 44128 769927
rect 44180 757784 44232 757790
rect 44180 757726 44232 757732
rect 44088 751120 44140 751126
rect 44088 751062 44140 751068
rect 44192 750938 44220 757726
rect 44272 757036 44324 757042
rect 44272 756978 44324 756984
rect 44008 750910 44220 750938
rect 44008 746298 44036 750910
rect 44284 750802 44312 756978
rect 44100 750774 44312 750802
rect 43996 746292 44048 746298
rect 43996 746234 44048 746240
rect 43904 743300 43956 743306
rect 43904 743242 43956 743248
rect 44100 743102 44128 750774
rect 44088 743096 44140 743102
rect 44088 743038 44140 743044
rect 41512 731128 41564 731134
rect 41512 731070 41564 731076
rect 43628 731128 43680 731134
rect 43628 731070 43680 731076
rect 44306 731096 44362 731105
rect 41524 729473 41552 731070
rect 44306 731031 44362 731040
rect 44148 730697 44176 730712
rect 44128 730688 44184 730697
rect 44128 730623 44184 730632
rect 43902 730280 43958 730289
rect 43902 730215 43958 730224
rect 41510 729464 41566 729473
rect 41510 729399 41566 729408
rect 43916 728929 43944 730215
rect 44148 729065 44176 730623
rect 44320 729201 44348 731031
rect 44610 730124 44638 772860
rect 44702 771688 44730 814398
rect 44794 813685 44822 813694
rect 44778 813676 44838 813685
rect 44778 813607 44838 813616
rect 44686 771678 44746 771688
rect 44686 771608 44746 771618
rect 44702 771590 44730 771608
rect 44702 771278 44730 771294
rect 44686 771268 44746 771278
rect 44686 771198 44746 771208
rect 44594 730114 44654 730124
rect 44594 730044 44654 730054
rect 44610 730036 44638 730044
rect 44594 729730 44654 729740
rect 44594 729660 44654 729670
rect 44306 729192 44362 729201
rect 44306 729127 44362 729136
rect 44138 729056 44194 729065
rect 44138 728991 44194 729000
rect 43718 728920 43774 728929
rect 43718 728855 43774 728864
rect 43902 728920 43958 728929
rect 43902 728855 43958 728864
rect 43166 726880 43222 726889
rect 43166 726815 43222 726824
rect 41786 724840 41842 724849
rect 41786 724775 41842 724784
rect 41418 723344 41474 723353
rect 41418 723279 41474 723288
rect 41432 717534 41460 723279
rect 41510 720896 41566 720905
rect 41510 720831 41566 720840
rect 41524 719681 41552 720831
rect 41510 719672 41566 719681
rect 41510 719607 41566 719616
rect 41524 717670 41552 719607
rect 41512 717664 41564 717670
rect 41512 717606 41564 717612
rect 41420 717528 41472 717534
rect 41420 717470 41472 717476
rect 41800 713862 41828 724775
rect 42246 723208 42302 723217
rect 42246 723143 42302 723152
rect 41788 713856 41840 713862
rect 41788 713798 41840 713804
rect 41788 713584 41840 713590
rect 41788 713526 41840 713532
rect 41800 713048 41828 713526
rect 42156 711748 42208 711754
rect 42156 711690 42208 711696
rect 42168 711212 42196 711690
rect 42156 710932 42208 710938
rect 42156 710874 42208 710880
rect 42168 710561 42196 710874
rect 42260 709866 42288 723143
rect 42706 722800 42762 722809
rect 42706 722735 42762 722744
rect 42338 721984 42394 721993
rect 42338 721919 42394 721928
rect 42352 710410 42380 721919
rect 42432 714876 42484 714882
rect 42432 714818 42484 714824
rect 42444 710938 42472 714818
rect 42432 710932 42484 710938
rect 42432 710874 42484 710880
rect 42352 710382 42472 710410
rect 42340 710320 42392 710326
rect 42340 710262 42392 710268
rect 42076 709838 42288 709866
rect 42076 709376 42104 709838
rect 42248 709368 42300 709374
rect 42248 709310 42300 709316
rect 42260 709050 42288 709310
rect 42168 709022 42288 709050
rect 42168 708696 42196 709022
rect 42156 708620 42208 708626
rect 42156 708562 42208 708568
rect 42168 708152 42196 708562
rect 42352 707554 42380 710262
rect 42182 707526 42380 707554
rect 42168 706982 42288 707010
rect 42168 706860 42196 706982
rect 42260 706874 42288 706982
rect 42444 706874 42472 710382
rect 42720 710326 42748 722735
rect 43180 714202 43208 726815
rect 43350 726472 43406 726481
rect 43350 726407 43406 726416
rect 43258 722392 43314 722401
rect 43258 722327 43314 722336
rect 43168 714196 43220 714202
rect 43168 714138 43220 714144
rect 42708 710320 42760 710326
rect 42708 710262 42760 710268
rect 43272 710190 43300 722327
rect 43364 711754 43392 726407
rect 43442 724024 43498 724033
rect 43442 723959 43498 723968
rect 43352 711748 43404 711754
rect 43352 711690 43404 711696
rect 42708 710184 42760 710190
rect 42708 710126 42760 710132
rect 43260 710184 43312 710190
rect 43260 710126 43312 710132
rect 42260 706846 42472 706874
rect 42432 706784 42484 706790
rect 42432 706726 42484 706732
rect 42444 706330 42472 706726
rect 42182 706302 42472 706330
rect 42248 706240 42300 706246
rect 42248 706182 42300 706188
rect 42064 704268 42116 704274
rect 42064 704210 42116 704216
rect 42076 703868 42104 704210
rect 42260 703202 42288 706182
rect 42340 705968 42392 705974
rect 42340 705910 42392 705916
rect 42182 703174 42288 703202
rect 42352 702590 42380 705910
rect 42720 704274 42748 710126
rect 43456 710002 43484 723959
rect 43626 721576 43682 721585
rect 43626 721511 43682 721520
rect 43536 717528 43588 717534
rect 43536 717470 43588 717476
rect 43272 709974 43484 710002
rect 43272 705974 43300 709974
rect 43444 709912 43496 709918
rect 43444 709854 43496 709860
rect 43352 709844 43404 709850
rect 43352 709786 43404 709792
rect 43260 705968 43312 705974
rect 43260 705910 43312 705916
rect 42708 704268 42760 704274
rect 42708 704210 42760 704216
rect 42432 703860 42484 703866
rect 42432 703802 42484 703808
rect 42168 702522 42196 702576
rect 42260 702562 42380 702590
rect 42260 702522 42288 702562
rect 42168 702494 42288 702522
rect 42340 702500 42392 702506
rect 42340 702442 42392 702448
rect 42352 702046 42380 702442
rect 42168 701978 42196 702032
rect 42260 702018 42380 702046
rect 42260 701978 42288 702018
rect 42168 701950 42288 701978
rect 42340 701956 42392 701962
rect 42340 701898 42392 701904
rect 42248 701820 42300 701826
rect 42248 701762 42300 701768
rect 42260 700179 42288 701762
rect 42182 700151 42288 700179
rect 42352 699530 42380 701898
rect 42182 699502 42380 699530
rect 42340 699440 42392 699446
rect 42340 699382 42392 699388
rect 42352 698918 42380 699382
rect 42168 698850 42196 698904
rect 42260 698890 42380 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 42444 698339 42472 703802
rect 43364 702506 43392 709786
rect 43456 706790 43484 709854
rect 43444 706784 43496 706790
rect 43444 706726 43496 706732
rect 43548 706246 43576 717470
rect 43640 708626 43668 721511
rect 43628 708620 43680 708626
rect 43628 708562 43680 708568
rect 43536 706240 43588 706246
rect 43536 706182 43588 706188
rect 43352 702500 43404 702506
rect 43352 702442 43404 702448
rect 42182 698311 42472 698339
rect 8588 688052 8616 688908
rect 9048 688052 9076 688908
rect 9508 688052 9536 688908
rect 9968 688052 9996 688908
rect 10428 688052 10456 688908
rect 10888 688052 10916 688908
rect 11348 688052 11376 688908
rect 11808 688052 11836 688908
rect 12268 688052 12296 688908
rect 12728 688052 12756 688908
rect 13188 688052 13216 688908
rect 13648 688052 13676 688908
rect 14108 688052 14136 688908
rect 41510 688392 41566 688401
rect 41510 688327 41512 688336
rect 41564 688327 41566 688336
rect 41512 688298 41564 688304
rect 41786 687712 41842 687721
rect 41786 687647 41788 687656
rect 41840 687647 41842 687656
rect 41788 687618 41840 687624
rect 41786 687304 41842 687313
rect 41786 687239 41788 687248
rect 41840 687239 41842 687248
rect 41788 687210 41840 687216
rect 43732 686089 43760 728855
rect 43810 726064 43866 726073
rect 43810 725999 43866 726008
rect 43824 712298 43852 725999
rect 43994 725656 44050 725665
rect 43994 725591 44050 725600
rect 43902 725248 43958 725257
rect 43902 725183 43958 725192
rect 43812 712292 43864 712298
rect 43812 712234 43864 712240
rect 43812 712156 43864 712162
rect 43812 712098 43864 712104
rect 43824 709442 43852 712098
rect 43916 709918 43944 725183
rect 43904 709912 43956 709918
rect 43904 709854 43956 709860
rect 44008 709850 44036 725591
rect 44086 724432 44142 724441
rect 44086 724367 44142 724376
rect 43996 709844 44048 709850
rect 43996 709786 44048 709792
rect 44100 709730 44128 724367
rect 44364 714196 44416 714202
rect 44364 714138 44416 714144
rect 44272 712292 44324 712298
rect 44272 712234 44324 712240
rect 43916 709702 44128 709730
rect 43812 709436 43864 709442
rect 43812 709378 43864 709384
rect 43916 709334 43944 709702
rect 44284 709646 44312 712234
rect 43996 709640 44048 709646
rect 43996 709582 44048 709588
rect 44272 709640 44324 709646
rect 44272 709582 44324 709588
rect 43824 709306 43944 709334
rect 43824 701962 43852 709306
rect 43812 701956 43864 701962
rect 43812 701898 43864 701904
rect 44008 699446 44036 709582
rect 44376 709578 44404 714138
rect 44088 709572 44140 709578
rect 44088 709514 44140 709520
rect 44364 709572 44416 709578
rect 44364 709514 44416 709520
rect 44100 701826 44128 709514
rect 44088 701820 44140 701826
rect 44088 701762 44140 701768
rect 43996 699440 44048 699446
rect 43996 699382 44048 699388
rect 44610 686924 44638 729660
rect 44702 728488 44730 771198
rect 44794 770897 44822 813607
rect 48332 786622 48360 817226
rect 48320 786616 48372 786622
rect 48320 786558 48372 786564
rect 51000 786554 51028 817634
rect 59266 814600 59322 814609
rect 59266 814535 59322 814544
rect 58256 800488 58308 800494
rect 58256 800430 58308 800436
rect 58268 790945 58296 800430
rect 58254 790936 58310 790945
rect 58254 790871 58310 790880
rect 58072 789404 58124 789410
rect 58072 789346 58124 789352
rect 58084 788497 58112 789346
rect 58532 789336 58584 789342
rect 58530 789304 58532 789313
rect 58584 789304 58586 789313
rect 58530 789239 58586 789248
rect 58070 788488 58126 788497
rect 58070 788423 58126 788432
rect 59280 787409 59308 814535
rect 62120 805996 62172 806002
rect 62120 805938 62172 805944
rect 59266 787400 59322 787409
rect 59266 787335 59322 787344
rect 58440 786616 58492 786622
rect 58440 786558 58492 786564
rect 50988 786548 51040 786554
rect 50988 786490 51040 786496
rect 58452 784961 58480 786558
rect 58532 786548 58584 786554
rect 58532 786490 58584 786496
rect 58544 786185 58572 786490
rect 58530 786176 58586 786185
rect 58530 786111 58586 786120
rect 58438 784952 58494 784961
rect 58438 784887 58494 784896
rect 53748 774784 53800 774790
rect 53748 774726 53800 774732
rect 50988 773900 51040 773906
rect 50988 773842 51040 773848
rect 45468 773492 45520 773498
rect 45468 773434 45520 773440
rect 44778 770888 44838 770897
rect 44778 770819 44838 770828
rect 44794 770796 44822 770819
rect 44794 770485 44822 770500
rect 44778 770476 44838 770485
rect 44778 770407 44838 770416
rect 44686 728478 44746 728488
rect 44686 728408 44746 728418
rect 44702 728388 44730 728408
rect 44702 728078 44730 728094
rect 44686 728068 44746 728078
rect 44686 727998 44746 728008
rect 44594 686914 44654 686924
rect 44594 686844 44654 686854
rect 44610 686836 44638 686844
rect 44610 686540 44638 686548
rect 44594 686530 44654 686540
rect 44594 686460 44654 686470
rect 43718 686080 43774 686089
rect 43718 686015 43774 686024
rect 43074 685672 43130 685681
rect 43074 685607 43130 685616
rect 42246 683224 42302 683233
rect 42246 683159 42302 683168
rect 41878 682000 41934 682009
rect 41878 681935 41934 681944
rect 41694 681456 41750 681465
rect 41694 681391 41750 681400
rect 41708 676546 41736 681391
rect 41786 678736 41842 678745
rect 41786 678671 41842 678680
rect 41800 678638 41828 678671
rect 41788 678632 41840 678638
rect 41788 678574 41840 678580
rect 41786 678328 41842 678337
rect 41786 678263 41842 678272
rect 41800 676666 41828 678263
rect 41788 676660 41840 676666
rect 41788 676602 41840 676608
rect 41708 676518 41828 676546
rect 5446 676288 5502 676297
rect 5446 676223 5502 676232
rect 5460 674830 5488 676223
rect 5538 676152 5594 676161
rect 5538 676087 5594 676096
rect 5552 675782 5580 676087
rect 30562 676016 30618 676025
rect 30562 675951 30618 675960
rect 30576 675782 30604 675951
rect 5540 675776 5592 675782
rect 5540 675718 5592 675724
rect 30564 675776 30616 675782
rect 30564 675718 30616 675724
rect 5448 674824 5500 674830
rect 5448 674766 5500 674772
rect 41800 670614 41828 676518
rect 41892 672450 41920 681935
rect 42062 680368 42118 680377
rect 42062 680303 42118 680312
rect 41880 672444 41932 672450
rect 41880 672386 41932 672392
rect 42076 670721 42104 680303
rect 42062 670712 42118 670721
rect 42062 670647 42118 670656
rect 41788 670608 41840 670614
rect 41788 670550 41840 670556
rect 41788 670404 41840 670410
rect 41788 670346 41840 670352
rect 41800 669868 41828 670346
rect 42168 667978 42196 668032
rect 42260 667978 42288 683159
rect 42338 681184 42394 681193
rect 42338 681119 42394 681128
rect 42352 671838 42380 681119
rect 42430 679552 42486 679561
rect 42430 679487 42486 679496
rect 42340 671832 42392 671838
rect 42340 671774 42392 671780
rect 42340 670812 42392 670818
rect 42340 670754 42392 670760
rect 42168 667950 42288 667978
rect 42248 667888 42300 667894
rect 42248 667830 42300 667836
rect 42156 667752 42208 667758
rect 42156 667694 42208 667700
rect 42168 667352 42196 667694
rect 42156 666732 42208 666738
rect 42156 666674 42208 666680
rect 42168 666165 42196 666674
rect 42260 666074 42288 667830
rect 42352 667758 42380 670754
rect 42444 670750 42472 679487
rect 43088 672586 43116 685607
rect 43258 683632 43314 683641
rect 43258 683567 43314 683576
rect 43168 676660 43220 676666
rect 43168 676602 43220 676608
rect 43076 672580 43128 672586
rect 43076 672522 43128 672528
rect 43076 672444 43128 672450
rect 43076 672386 43128 672392
rect 42432 670744 42484 670750
rect 42432 670686 42484 670692
rect 42340 667752 42392 667758
rect 42340 667694 42392 667700
rect 42260 666046 42380 666074
rect 42182 665502 42288 665530
rect 42156 665236 42208 665242
rect 42156 665178 42208 665184
rect 42168 664972 42196 665178
rect 42156 664692 42208 664698
rect 42156 664634 42208 664640
rect 42168 664325 42196 664634
rect 42156 664216 42208 664222
rect 42156 664158 42208 664164
rect 42168 663680 42196 664158
rect 42156 663400 42208 663406
rect 42156 663342 42208 663348
rect 42168 663136 42196 663342
rect 42156 661088 42208 661094
rect 42156 661030 42208 661036
rect 42168 660620 42196 661030
rect 42156 660544 42208 660550
rect 42156 660486 42208 660492
rect 42168 660008 42196 660486
rect 42260 659666 42288 665502
rect 42248 659660 42300 659666
rect 42248 659602 42300 659608
rect 42248 659524 42300 659530
rect 42248 659466 42300 659472
rect 42260 659371 42288 659466
rect 42182 659343 42288 659371
rect 42156 659252 42208 659258
rect 42156 659194 42208 659200
rect 42168 658784 42196 659194
rect 42156 657416 42208 657422
rect 42156 657358 42208 657364
rect 42168 656948 42196 657358
rect 42352 656350 42380 666046
rect 43088 663406 43116 672386
rect 43180 671922 43208 676602
rect 43272 672042 43300 683567
rect 43534 682816 43590 682825
rect 43534 682751 43590 682760
rect 43442 682408 43498 682417
rect 43442 682343 43498 682352
rect 43352 674824 43404 674830
rect 43352 674766 43404 674772
rect 43260 672036 43312 672042
rect 43260 671978 43312 671984
rect 43180 671894 43300 671922
rect 43168 671832 43220 671838
rect 43168 671774 43220 671780
rect 43180 667894 43208 671774
rect 43168 667888 43220 667894
rect 43168 667830 43220 667836
rect 43168 667752 43220 667758
rect 43168 667694 43220 667700
rect 43180 664222 43208 667694
rect 43272 665242 43300 671894
rect 43260 665236 43312 665242
rect 43260 665178 43312 665184
rect 43258 665136 43314 665145
rect 43258 665071 43314 665080
rect 43168 664216 43220 664222
rect 43168 664158 43220 664164
rect 43076 663400 43128 663406
rect 43076 663342 43128 663348
rect 43272 660550 43300 665071
rect 43364 661094 43392 674766
rect 43456 672178 43484 682343
rect 43548 680898 43576 682751
rect 43548 680870 43944 680898
rect 43718 680776 43774 680785
rect 43718 680711 43774 680720
rect 43626 679960 43682 679969
rect 43626 679895 43682 679904
rect 43536 672580 43588 672586
rect 43536 672522 43588 672528
rect 43444 672172 43496 672178
rect 43444 672114 43496 672120
rect 43444 672036 43496 672042
rect 43444 671978 43496 671984
rect 43456 662414 43484 671978
rect 43548 670886 43576 672522
rect 43536 670880 43588 670886
rect 43536 670822 43588 670828
rect 43536 670744 43588 670750
rect 43536 670686 43588 670692
rect 43548 664698 43576 670686
rect 43640 666738 43668 679895
rect 43732 670682 43760 680711
rect 43720 670676 43772 670682
rect 43720 670618 43772 670624
rect 43628 666732 43680 666738
rect 43628 666674 43680 666680
rect 43536 664692 43588 664698
rect 43536 664634 43588 664640
rect 43628 664556 43680 664562
rect 43628 664498 43680 664504
rect 43456 662386 43576 662414
rect 43352 661088 43404 661094
rect 43352 661030 43404 661036
rect 43260 660544 43312 660550
rect 43260 660486 43312 660492
rect 42432 659728 42484 659734
rect 42432 659670 42484 659676
rect 42182 656322 42380 656350
rect 42156 656056 42208 656062
rect 42156 655998 42208 656004
rect 42168 655656 42196 655998
rect 42444 655126 42472 659670
rect 43548 657422 43576 662386
rect 43640 659530 43668 664498
rect 43628 659524 43680 659530
rect 43628 659466 43680 659472
rect 43536 657416 43588 657422
rect 43536 657358 43588 657364
rect 43916 656062 43944 680870
rect 44088 678632 44140 678638
rect 44088 678574 44140 678580
rect 43996 672172 44048 672178
rect 43996 672114 44048 672120
rect 44008 670970 44036 672114
rect 44100 671106 44128 678574
rect 44100 671078 44220 671106
rect 44008 670942 44128 670970
rect 43996 670880 44048 670886
rect 43996 670822 44048 670828
rect 43904 656056 43956 656062
rect 43904 655998 43956 656004
rect 42182 655098 42472 655126
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 41512 645108 41564 645114
rect 41512 645050 41564 645056
rect 41524 644745 41552 645050
rect 41788 645040 41840 645046
rect 41788 644982 41840 644988
rect 41800 644949 41828 644982
rect 41786 644940 41842 644949
rect 41786 644875 41842 644884
rect 41510 644736 41566 644745
rect 41510 644671 41566 644680
rect 41786 644124 41842 644133
rect 41786 644059 41788 644068
rect 41840 644059 41842 644068
rect 41788 644030 41840 644036
rect 44008 643113 44036 670822
rect 44100 659258 44128 670942
rect 44192 667758 44220 671078
rect 44272 670676 44324 670682
rect 44272 670618 44324 670624
rect 44180 667752 44232 667758
rect 44180 667694 44232 667700
rect 44284 664562 44312 670618
rect 44272 664556 44324 664562
rect 44272 664498 44324 664504
rect 44088 659252 44140 659258
rect 44088 659194 44140 659200
rect 44610 643724 44638 686460
rect 44702 685288 44730 727998
rect 44794 727697 44822 770407
rect 45480 745210 45508 773434
rect 48228 767440 48280 767446
rect 48228 767382 48280 767388
rect 45468 745204 45520 745210
rect 45468 745146 45520 745152
rect 44778 727688 44838 727697
rect 44778 727619 44838 727628
rect 44794 727608 44822 727619
rect 44794 727285 44822 727312
rect 44778 727276 44838 727285
rect 44778 727207 44838 727216
rect 44686 685278 44746 685288
rect 44686 685208 44746 685218
rect 44702 685190 44730 685208
rect 44702 684878 44730 684900
rect 44686 684868 44746 684878
rect 44686 684798 44746 684808
rect 44594 643714 44654 643724
rect 44594 643644 44654 643654
rect 44610 643636 44638 643644
rect 44610 643340 44638 643342
rect 44594 643330 44654 643340
rect 44594 643260 44654 643270
rect 43994 643104 44050 643113
rect 43994 643039 44050 643048
rect 43902 642288 43958 642297
rect 43902 642223 43958 642232
rect 43074 640384 43130 640393
rect 43074 640319 43130 640328
rect 42338 639840 42394 639849
rect 42338 639775 42394 639784
rect 42246 638208 42302 638217
rect 42246 638143 42302 638152
rect 30194 637800 30250 637809
rect 30194 637735 30250 637744
rect 30102 637392 30158 637401
rect 30102 637327 30158 637336
rect 20628 632664 20680 632670
rect 30116 632641 30144 637327
rect 30208 632670 30236 637735
rect 38474 634944 38530 634953
rect 38474 634879 38530 634888
rect 30196 632664 30248 632670
rect 20628 632606 20680 632612
rect 24766 632632 24822 632641
rect 20640 630834 20668 632606
rect 24766 632567 24822 632576
rect 30102 632632 30158 632641
rect 30196 632606 30248 632612
rect 30102 632567 30158 632576
rect 20628 630828 20680 630834
rect 20628 630770 20680 630776
rect 24780 630766 24808 632567
rect 24768 630760 24820 630766
rect 24768 630702 24820 630708
rect 38488 629270 38516 634879
rect 41510 634536 41566 634545
rect 41510 634471 41566 634480
rect 41524 633321 41552 634471
rect 41510 633312 41566 633321
rect 41510 633247 41512 633256
rect 41564 633247 41566 633256
rect 41512 633218 41564 633224
rect 38476 629264 38528 629270
rect 38476 629206 38528 629212
rect 42260 627178 42288 638143
rect 42168 627150 42288 627178
rect 42168 626620 42196 627150
rect 42352 625326 42380 639775
rect 42706 636984 42762 636993
rect 42706 636919 42762 636928
rect 42432 630964 42484 630970
rect 42432 630906 42484 630912
rect 42444 627473 42472 630906
rect 42430 627464 42486 627473
rect 42430 627399 42486 627408
rect 42720 626754 42748 636919
rect 43088 629406 43116 640319
rect 43166 639024 43222 639033
rect 43166 638959 43222 638968
rect 43180 630902 43208 638959
rect 43626 638616 43682 638625
rect 43626 638551 43682 638560
rect 43258 636576 43314 636585
rect 43258 636511 43314 636520
rect 43168 630896 43220 630902
rect 43168 630838 43220 630844
rect 43168 630760 43220 630766
rect 43168 630702 43220 630708
rect 43076 629400 43128 629406
rect 43076 629342 43128 629348
rect 43076 629264 43128 629270
rect 43076 629206 43128 629212
rect 42708 626748 42760 626754
rect 42708 626690 42760 626696
rect 42708 626612 42760 626618
rect 42708 626554 42760 626560
rect 42156 625320 42208 625326
rect 42156 625262 42208 625268
rect 42340 625320 42392 625326
rect 42340 625262 42392 625268
rect 42168 624784 42196 625262
rect 42720 624510 42748 626554
rect 42340 624504 42392 624510
rect 42340 624446 42392 624452
rect 42708 624504 42760 624510
rect 42708 624446 42760 624452
rect 42182 624158 42288 624186
rect 42156 623484 42208 623490
rect 42156 623426 42208 623432
rect 42168 622948 42196 623426
rect 42260 622470 42288 624158
rect 42248 622464 42300 622470
rect 42248 622406 42300 622412
rect 42352 622350 42380 624446
rect 42708 622464 42760 622470
rect 42708 622406 42760 622412
rect 42182 622322 42380 622350
rect 42340 622260 42392 622266
rect 42340 622202 42392 622208
rect 42352 621806 42380 622202
rect 42168 621738 42196 621792
rect 42260 621778 42380 621806
rect 42260 621738 42288 621778
rect 42168 621710 42288 621738
rect 42340 621716 42392 621722
rect 42340 621658 42392 621664
rect 42352 621126 42380 621658
rect 42182 621098 42380 621126
rect 42338 620936 42394 620945
rect 42338 620871 42394 620880
rect 42064 620832 42116 620838
rect 42064 620774 42116 620780
rect 42076 620500 42104 620774
rect 42064 620220 42116 620226
rect 42064 620162 42116 620168
rect 42076 619956 42104 620162
rect 42352 617454 42380 620871
rect 42432 619200 42484 619206
rect 42432 619142 42484 619148
rect 42182 617426 42380 617454
rect 42064 617364 42116 617370
rect 42064 617306 42116 617312
rect 42076 616828 42104 617306
rect 42444 616162 42472 619142
rect 42720 618254 42748 622406
rect 43088 622266 43116 629206
rect 43076 622260 43128 622266
rect 43076 622202 43128 622208
rect 43074 622160 43130 622169
rect 43074 622095 43130 622104
rect 43088 620226 43116 622095
rect 43076 620220 43128 620226
rect 43076 620162 43128 620168
rect 43180 619206 43208 630702
rect 43272 623490 43300 636511
rect 43442 636168 43498 636177
rect 43442 636103 43498 636112
rect 43350 635352 43406 635361
rect 43350 635287 43406 635296
rect 43364 626890 43392 635287
rect 43352 626884 43404 626890
rect 43352 626826 43404 626832
rect 43352 626748 43404 626754
rect 43352 626690 43404 626696
rect 43260 623484 43312 623490
rect 43260 623426 43312 623432
rect 43168 619200 43220 619206
rect 43168 619142 43220 619148
rect 42708 618248 42760 618254
rect 42708 618190 42760 618196
rect 43364 617370 43392 626690
rect 43456 621722 43484 636103
rect 43640 627065 43668 638551
rect 43718 635760 43774 635769
rect 43718 635695 43774 635704
rect 43732 630970 43760 635695
rect 43720 630964 43772 630970
rect 43720 630906 43772 630912
rect 43812 630896 43864 630902
rect 43812 630838 43864 630844
rect 43720 630828 43772 630834
rect 43720 630770 43772 630776
rect 43626 627056 43682 627065
rect 43626 626991 43682 627000
rect 43628 626884 43680 626890
rect 43628 626826 43680 626832
rect 43444 621716 43496 621722
rect 43444 621658 43496 621664
rect 43640 620838 43668 626826
rect 43628 620832 43680 620838
rect 43628 620774 43680 620780
rect 43352 617364 43404 617370
rect 43352 617306 43404 617312
rect 42182 616134 42472 616162
rect 42340 616072 42392 616078
rect 42340 616014 42392 616020
rect 42248 616004 42300 616010
rect 42248 615946 42300 615952
rect 42156 615868 42208 615874
rect 42156 615810 42208 615816
rect 42168 615604 42196 615810
rect 42156 614236 42208 614242
rect 42156 614178 42208 614184
rect 42168 613768 42196 614178
rect 42260 613135 42288 615946
rect 42182 613107 42288 613135
rect 42352 612490 42380 616014
rect 43732 616010 43760 630770
rect 43720 616004 43772 616010
rect 43720 615946 43772 615952
rect 43824 615874 43852 630838
rect 43812 615868 43864 615874
rect 43812 615810 43864 615816
rect 42432 615528 42484 615534
rect 42432 615470 42484 615476
rect 42182 612462 42380 612490
rect 42444 611946 42472 615470
rect 42182 611918 42472 611946
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 41786 601760 41842 601769
rect 41786 601695 41788 601704
rect 41840 601695 41842 601704
rect 41788 601666 41840 601672
rect 43916 601497 43944 642223
rect 44086 639432 44142 639441
rect 44086 639367 44142 639376
rect 43996 629400 44048 629406
rect 43996 629342 44048 629348
rect 44008 614242 44036 629342
rect 44100 616078 44128 639367
rect 44088 616072 44140 616078
rect 44088 616014 44140 616020
rect 43996 614236 44048 614242
rect 43996 614178 44048 614184
rect 41510 601488 41566 601497
rect 41510 601423 41566 601432
rect 43902 601488 43958 601497
rect 43902 601423 43958 601432
rect 41524 599865 41552 601423
rect 42706 601080 42762 601089
rect 42706 601015 42762 601024
rect 41510 599856 41566 599865
rect 41510 599791 41566 599800
rect 42720 599185 42748 601015
rect 43074 600672 43130 600681
rect 43074 600607 43130 600616
rect 42706 599176 42762 599185
rect 42706 599111 42762 599120
rect 43088 599049 43116 600607
rect 44610 600524 44638 643260
rect 44702 642088 44730 684798
rect 44794 684497 44822 727207
rect 45744 687268 45796 687274
rect 45744 687210 45796 687216
rect 44778 684488 44838 684497
rect 44778 684419 44838 684428
rect 44794 684392 44822 684419
rect 44794 684085 44822 684096
rect 44778 684076 44838 684085
rect 44778 684007 44838 684016
rect 44686 642078 44746 642088
rect 44686 642008 44746 642018
rect 44702 641986 44730 642008
rect 44702 641678 44730 641694
rect 44686 641668 44746 641678
rect 44686 641598 44746 641608
rect 44594 600514 44654 600524
rect 44594 600444 44654 600454
rect 44610 600436 44638 600444
rect 44610 600140 44638 600152
rect 44594 600130 44654 600140
rect 44594 600060 44654 600070
rect 43902 599312 43958 599321
rect 43902 599247 43958 599256
rect 43074 599040 43130 599049
rect 43074 598975 43130 598984
rect 43166 596864 43222 596873
rect 43166 596799 43222 596808
rect 41786 595232 41842 595241
rect 41786 595167 41842 595176
rect 38566 593328 38622 593337
rect 38566 593263 38622 593272
rect 38580 587858 38608 593263
rect 41510 591288 41566 591297
rect 41510 591223 41566 591232
rect 41524 590073 41552 591223
rect 41510 590064 41566 590073
rect 41510 589999 41566 590008
rect 41524 589286 41552 589999
rect 41512 589280 41564 589286
rect 41512 589222 41564 589228
rect 38568 587852 38620 587858
rect 38568 587794 38620 587800
rect 41800 584202 41828 595167
rect 42430 594824 42486 594833
rect 42430 594759 42486 594768
rect 42340 587852 42392 587858
rect 42340 587794 42392 587800
rect 41800 584174 42288 584202
rect 42260 583454 42288 584174
rect 42182 583426 42288 583454
rect 42248 582616 42300 582622
rect 42248 582558 42300 582564
rect 42156 582140 42208 582146
rect 42156 582082 42208 582088
rect 42168 581604 42196 582082
rect 42156 581528 42208 581534
rect 42156 581470 42208 581476
rect 42168 580961 42196 581470
rect 42260 580378 42288 582558
rect 42248 580372 42300 580378
rect 42248 580314 42300 580320
rect 42352 580258 42380 587794
rect 42444 584254 42472 594759
rect 43076 593020 43128 593026
rect 43076 592962 43128 592968
rect 43088 585313 43116 592962
rect 43180 592090 43208 596799
rect 43718 596456 43774 596465
rect 43718 596391 43774 596400
rect 43350 595640 43406 595649
rect 43350 595575 43406 595584
rect 43364 593026 43392 595575
rect 43442 594416 43498 594425
rect 43442 594351 43498 594360
rect 43352 593020 43404 593026
rect 43352 592962 43404 592968
rect 43352 592884 43404 592890
rect 43352 592826 43404 592832
rect 43180 592062 43300 592090
rect 43166 591968 43222 591977
rect 43166 591903 43222 591912
rect 43074 585304 43130 585313
rect 43074 585239 43130 585248
rect 43076 585200 43128 585206
rect 43076 585142 43128 585148
rect 42432 584248 42484 584254
rect 42432 584190 42484 584196
rect 43088 581534 43116 585142
rect 43076 581528 43128 581534
rect 43076 581470 43128 581476
rect 43074 581360 43130 581369
rect 43074 581295 43130 581304
rect 42168 580230 42380 580258
rect 42168 579768 42196 580230
rect 42248 580168 42300 580174
rect 42248 580110 42300 580116
rect 42260 579850 42288 580110
rect 42260 579822 42380 579850
rect 42352 579135 42380 579822
rect 42182 579107 42380 579135
rect 42248 579012 42300 579018
rect 42248 578954 42300 578960
rect 42156 578808 42208 578814
rect 42156 578750 42208 578756
rect 42168 578544 42196 578750
rect 42156 578468 42208 578474
rect 42156 578410 42208 578416
rect 42168 577932 42196 578410
rect 42260 577295 42288 578954
rect 42182 577267 42288 577295
rect 42248 577176 42300 577182
rect 42248 577118 42300 577124
rect 42156 576972 42208 576978
rect 42156 576914 42208 576920
rect 42168 576708 42196 576914
rect 42260 574274 42288 577118
rect 43088 576978 43116 581295
rect 43180 578814 43208 591903
rect 43272 582146 43300 592062
rect 43364 583914 43392 592826
rect 43352 583908 43404 583914
rect 43352 583850 43404 583856
rect 43350 583808 43406 583817
rect 43350 583743 43406 583752
rect 43260 582140 43312 582146
rect 43260 582082 43312 582088
rect 43260 582004 43312 582010
rect 43260 581946 43312 581952
rect 43168 578808 43220 578814
rect 43168 578750 43220 578756
rect 43076 576972 43128 576978
rect 43076 576914 43128 576920
rect 42340 576020 42392 576026
rect 42340 575962 42392 575968
rect 42182 574246 42288 574274
rect 42156 573844 42208 573850
rect 42156 573786 42208 573792
rect 42168 573580 42196 573786
rect 42352 572982 42380 575962
rect 42432 574116 42484 574122
rect 42432 574058 42484 574064
rect 42182 572954 42380 572982
rect 42340 572892 42392 572898
rect 42340 572834 42392 572840
rect 42352 572438 42380 572834
rect 42168 572370 42196 572424
rect 42260 572410 42380 572438
rect 42260 572370 42288 572410
rect 42168 572342 42288 572370
rect 42248 572008 42300 572014
rect 42248 571950 42300 571956
rect 42064 570988 42116 570994
rect 42064 570930 42116 570936
rect 42076 570588 42104 570930
rect 42260 569922 42288 571950
rect 42340 571668 42392 571674
rect 42340 571610 42392 571616
rect 42182 569894 42288 569922
rect 42352 569310 42380 571610
rect 42168 569242 42196 569296
rect 42260 569282 42380 569310
rect 42260 569242 42288 569282
rect 42168 569214 42288 569242
rect 42444 568766 42472 574058
rect 43272 570994 43300 581946
rect 43364 573850 43392 583743
rect 43456 580530 43484 594351
rect 43534 594008 43590 594017
rect 43534 593943 43590 593952
rect 43548 583817 43576 593943
rect 43626 592376 43682 592385
rect 43626 592311 43682 592320
rect 43534 583808 43590 583817
rect 43534 583743 43590 583752
rect 43536 583704 43588 583710
rect 43536 583646 43588 583652
rect 43548 582010 43576 583646
rect 43536 582004 43588 582010
rect 43536 581946 43588 581952
rect 43456 580502 43576 580530
rect 43444 580440 43496 580446
rect 43444 580382 43496 580388
rect 43352 573844 43404 573850
rect 43352 573786 43404 573792
rect 43456 572898 43484 580382
rect 43548 576026 43576 580502
rect 43640 579018 43668 592311
rect 43628 579012 43680 579018
rect 43628 578954 43680 578960
rect 43536 576020 43588 576026
rect 43536 575962 43588 575968
rect 43444 572892 43496 572898
rect 43444 572834 43496 572840
rect 43732 571674 43760 596391
rect 43810 593192 43866 593201
rect 43810 593127 43866 593136
rect 43824 578474 43852 593127
rect 43916 578474 43944 599247
rect 44086 597272 44142 597281
rect 44086 597207 44142 597216
rect 43994 596048 44050 596057
rect 43994 595983 44050 595992
rect 44008 580446 44036 595983
rect 44100 592890 44128 597207
rect 44088 592884 44140 592890
rect 44088 592826 44140 592832
rect 44086 592784 44142 592793
rect 44086 592719 44142 592728
rect 43996 580440 44048 580446
rect 43996 580382 44048 580388
rect 44100 580378 44128 592719
rect 44272 584248 44324 584254
rect 44272 584190 44324 584196
rect 44088 580372 44140 580378
rect 44088 580314 44140 580320
rect 44088 580168 44140 580174
rect 44088 580110 44140 580116
rect 43812 578468 43864 578474
rect 43812 578410 43864 578416
rect 43904 578468 43956 578474
rect 43904 578410 43956 578416
rect 43904 578264 43956 578270
rect 43904 578206 43956 578212
rect 43720 571668 43772 571674
rect 43720 571610 43772 571616
rect 43260 570988 43312 570994
rect 43260 570930 43312 570936
rect 42168 568698 42196 568752
rect 42260 568738 42472 568766
rect 42260 568698 42288 568738
rect 42168 568670 42288 568698
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 41512 558816 41564 558822
rect 41510 558784 41512 558793
rect 41564 558784 41566 558793
rect 41510 558719 41566 558728
rect 41512 558680 41564 558686
rect 41512 558622 41564 558628
rect 41524 558385 41552 558622
rect 41510 558376 41566 558385
rect 41510 558311 41566 558320
rect 41512 557592 41564 557598
rect 41510 557560 41512 557569
rect 41564 557560 41566 557569
rect 41510 557495 41566 557504
rect 43916 556481 43944 578206
rect 44100 577182 44128 580110
rect 44088 577176 44140 577182
rect 44088 577118 44140 577124
rect 44284 576994 44312 584190
rect 44100 576966 44312 576994
rect 44100 572014 44128 576966
rect 44088 572008 44140 572014
rect 44088 571950 44140 571956
rect 44610 557324 44638 600060
rect 44702 598888 44730 641598
rect 44794 641297 44822 684007
rect 45756 659598 45784 687210
rect 45744 659592 45796 659598
rect 45744 659534 45796 659540
rect 44778 641288 44838 641297
rect 44778 641219 44838 641228
rect 44794 641188 44822 641219
rect 44794 640885 44822 640892
rect 44778 640876 44838 640885
rect 44778 640807 44838 640816
rect 44686 598878 44746 598888
rect 44686 598808 44746 598818
rect 44702 598790 44730 598808
rect 44702 598478 44730 598504
rect 44686 598468 44746 598478
rect 44686 598398 44746 598408
rect 44594 557314 44654 557324
rect 44594 557244 44654 557254
rect 44610 557236 44638 557244
rect 44610 556940 44638 556946
rect 44594 556930 44654 556940
rect 44594 556860 44654 556870
rect 43902 556472 43958 556481
rect 43902 556407 43958 556416
rect 38106 555520 38162 555529
rect 38106 555455 38162 555464
rect 38120 546417 38148 555455
rect 43350 553616 43406 553625
rect 43350 553551 43406 553560
rect 41786 551984 41842 551993
rect 41786 551919 41842 551928
rect 41602 549808 41658 549817
rect 41602 549743 41658 549752
rect 41418 549400 41474 549409
rect 41418 549335 41474 549344
rect 38106 546408 38162 546417
rect 41432 546378 41460 549335
rect 41510 548992 41566 549001
rect 41510 548927 41566 548936
rect 41524 548690 41552 548927
rect 41512 548684 41564 548690
rect 41512 548626 41564 548632
rect 41510 548584 41566 548593
rect 41510 548519 41566 548528
rect 41524 548486 41552 548519
rect 41512 548480 41564 548486
rect 41512 548422 41564 548428
rect 41510 548176 41566 548185
rect 41510 548111 41566 548120
rect 41524 546961 41552 548111
rect 41510 546952 41566 546961
rect 41510 546887 41512 546896
rect 41564 546887 41566 546896
rect 41512 546858 41564 546864
rect 41616 546446 41644 549743
rect 41604 546440 41656 546446
rect 41604 546382 41656 546388
rect 38106 546343 38162 546352
rect 41420 546372 41472 546378
rect 41420 546314 41472 546320
rect 41800 541074 41828 551919
rect 43166 550352 43222 550361
rect 43166 550287 43222 550296
rect 41788 541068 41840 541074
rect 41788 541010 41840 541016
rect 42248 541068 42300 541074
rect 42248 541010 42300 541016
rect 43076 541068 43128 541074
rect 43076 541010 43128 541016
rect 41788 540796 41840 540802
rect 41788 540738 41840 540744
rect 41800 540260 41828 540738
rect 42064 538960 42116 538966
rect 42064 538902 42116 538908
rect 42076 538424 42104 538902
rect 42260 538234 42288 541010
rect 42168 538206 42288 538234
rect 42168 537744 42196 538206
rect 43088 538150 43116 541010
rect 42248 538144 42300 538150
rect 42248 538086 42300 538092
rect 43076 538144 43128 538150
rect 43076 538086 43128 538092
rect 42064 537124 42116 537130
rect 42064 537066 42116 537072
rect 42076 536588 42104 537066
rect 42260 535922 42288 538086
rect 43180 537130 43208 550287
rect 43260 548480 43312 548486
rect 43260 548422 43312 548428
rect 43168 537124 43220 537130
rect 43168 537066 43220 537072
rect 42182 535894 42288 535922
rect 42246 535800 42302 535809
rect 42246 535735 42302 535744
rect 42156 535628 42208 535634
rect 42156 535570 42208 535576
rect 42168 535364 42196 535570
rect 42064 535084 42116 535090
rect 42064 535026 42116 535032
rect 42076 534752 42104 535026
rect 42156 534472 42208 534478
rect 42156 534414 42208 534420
rect 42168 534072 42196 534414
rect 42156 533996 42208 534002
rect 42156 533938 42208 533944
rect 42168 533528 42196 533938
rect 42154 532808 42210 532817
rect 42260 532794 42288 535735
rect 43272 535634 43300 548422
rect 43364 538966 43392 553551
rect 43628 548684 43680 548690
rect 43628 548626 43680 548632
rect 43444 546372 43496 546378
rect 43444 546314 43496 546320
rect 43352 538960 43404 538966
rect 43352 538902 43404 538908
rect 43350 538792 43406 538801
rect 43350 538727 43406 538736
rect 43260 535628 43312 535634
rect 43260 535570 43312 535576
rect 43364 534002 43392 538727
rect 43352 533996 43404 534002
rect 43352 533938 43404 533944
rect 43074 533080 43130 533089
rect 43074 533015 43130 533024
rect 42430 532808 42486 532817
rect 42260 532766 42380 532794
rect 42154 532743 42210 532752
rect 42168 532658 42196 532743
rect 42168 532630 42288 532658
rect 42156 531480 42208 531486
rect 42156 531422 42208 531428
rect 42168 531045 42196 531422
rect 42156 530732 42208 530738
rect 42156 530674 42208 530680
rect 42168 530400 42196 530674
rect 42260 530618 42288 532630
rect 42352 530738 42380 532766
rect 42430 532743 42486 532752
rect 42340 530732 42392 530738
rect 42340 530674 42392 530680
rect 42260 530590 42380 530618
rect 42352 530346 42380 530590
rect 42260 530318 42380 530346
rect 42260 529771 42288 530318
rect 42338 530224 42394 530233
rect 42338 530159 42394 530168
rect 42182 529743 42288 529771
rect 42352 529666 42380 530159
rect 42260 529638 42380 529666
rect 42156 529508 42208 529514
rect 42156 529450 42208 529456
rect 42168 529205 42196 529450
rect 42156 527808 42208 527814
rect 42156 527750 42208 527756
rect 42168 527340 42196 527750
rect 42260 527218 42288 529638
rect 42444 527814 42472 532743
rect 43088 529514 43116 533015
rect 43456 531486 43484 546314
rect 43640 534478 43668 548626
rect 43720 546440 43772 546446
rect 43720 546382 43772 546388
rect 43732 535090 43760 546382
rect 43720 535084 43772 535090
rect 43720 535026 43772 535032
rect 43628 534472 43680 534478
rect 43628 534414 43680 534420
rect 43444 531480 43496 531486
rect 43444 531422 43496 531428
rect 43166 530768 43222 530777
rect 43166 530703 43222 530712
rect 43076 529508 43128 529514
rect 43076 529450 43128 529456
rect 42432 527808 42484 527814
rect 42432 527750 42484 527756
rect 42168 527190 42288 527218
rect 42168 526728 42196 527190
rect 43180 526454 43208 530703
rect 43260 529984 43312 529990
rect 43260 529926 43312 529932
rect 42156 526448 42208 526454
rect 42156 526390 42208 526396
rect 43168 526448 43220 526454
rect 43168 526390 43220 526396
rect 42168 526077 42196 526390
rect 43272 525774 43300 529926
rect 42156 525768 42208 525774
rect 42156 525710 42208 525716
rect 43260 525768 43312 525774
rect 43260 525710 43312 525716
rect 42168 525504 42196 525710
rect 42430 455968 42486 455977
rect 42430 455903 42486 455912
rect 42444 450809 42472 455903
rect 42430 450800 42486 450809
rect 42430 450735 42486 450744
rect 42430 445904 42486 445913
rect 42430 445839 42486 445848
rect 42444 440745 42472 445839
rect 42430 440736 42486 440745
rect 42430 440671 42486 440680
rect 8588 431596 8616 431732
rect 9048 431596 9076 431732
rect 9508 431596 9536 431732
rect 9968 431596 9996 431732
rect 10428 431596 10456 431732
rect 10888 431596 10916 431732
rect 11348 431596 11376 431732
rect 11808 431596 11836 431732
rect 12268 431596 12296 431732
rect 12728 431596 12756 431732
rect 13188 431596 13216 431732
rect 13648 431596 13676 431732
rect 14108 431596 14136 431732
rect 30024 427689 30052 440316
rect 30116 428097 30144 440316
rect 41786 430944 41842 430953
rect 41786 430879 41788 430888
rect 41840 430879 41842 430888
rect 41788 430850 41840 430856
rect 41786 430536 41842 430545
rect 41786 430471 41842 430480
rect 30102 428088 30158 428097
rect 30102 428023 30158 428032
rect 41800 427881 41828 430471
rect 42062 430128 42118 430137
rect 42062 430063 42118 430072
rect 42076 428321 42104 430063
rect 44610 429724 44638 556860
rect 44702 555688 44730 598398
rect 44794 598097 44822 640807
rect 44778 598088 44838 598097
rect 44778 598019 44838 598028
rect 44794 597998 44822 598019
rect 44794 597685 44822 597702
rect 44778 597676 44838 597685
rect 44778 597607 44838 597616
rect 44686 555678 44746 555688
rect 44686 555608 44746 555618
rect 44702 555590 44730 555608
rect 44702 555278 44730 555294
rect 44686 555268 44746 555278
rect 44686 555198 44746 555208
rect 44594 429714 44654 429724
rect 44594 429644 44654 429654
rect 44610 429636 44638 429644
rect 44610 429340 44638 429348
rect 44594 429330 44654 429340
rect 44594 429260 44654 429270
rect 43718 428496 43774 428505
rect 43718 428431 43774 428440
rect 42054 428312 42110 428321
rect 42054 428247 42110 428256
rect 42076 428238 42104 428247
rect 41786 427872 41842 427881
rect 41786 427807 41842 427816
rect 30010 427680 30066 427689
rect 30010 427615 30066 427624
rect 43442 426456 43498 426465
rect 43442 426391 43498 426400
rect 42338 426048 42394 426057
rect 42338 425983 42394 425992
rect 42246 424416 42302 424425
rect 42246 424351 42302 424360
rect 41878 422784 41934 422793
rect 41878 422719 41934 422728
rect 41786 420744 41842 420753
rect 41786 420679 41842 420688
rect 41800 419529 41828 420679
rect 41786 419520 41842 419529
rect 41786 419455 41788 419464
rect 41840 419455 41842 419464
rect 41788 419426 41840 419432
rect 41892 416634 41920 422719
rect 41970 422376 42026 422385
rect 41970 422311 42026 422320
rect 41984 416702 42012 422311
rect 41972 416696 42024 416702
rect 41972 416638 42024 416644
rect 41880 416628 41932 416634
rect 41880 416570 41932 416576
rect 42260 413114 42288 424351
rect 42168 413086 42288 413114
rect 42168 412624 42196 413086
rect 42352 412978 42380 425983
rect 42706 425640 42762 425649
rect 42706 425575 42762 425584
rect 42260 412950 42380 412978
rect 42260 411254 42288 412950
rect 42168 411226 42288 411254
rect 42340 411256 42392 411262
rect 42168 410788 42196 411226
rect 42340 411198 42392 411204
rect 42182 410162 42288 410190
rect 42260 409562 42288 410162
rect 42248 409556 42300 409562
rect 42248 409498 42300 409504
rect 42352 409442 42380 411198
rect 42168 409414 42380 409442
rect 42168 408952 42196 409414
rect 42340 409352 42392 409358
rect 42340 409294 42392 409300
rect 42352 408898 42380 409294
rect 42260 408870 42380 408898
rect 42064 408060 42116 408066
rect 42064 408002 42116 408008
rect 42076 407796 42104 408002
rect 42168 407930 42196 408340
rect 42156 407924 42208 407930
rect 42156 407866 42208 407872
rect 42156 407652 42208 407658
rect 42156 407594 42208 407600
rect 42168 407116 42196 407594
rect 42064 406836 42116 406842
rect 42064 406778 42116 406784
rect 42076 406504 42104 406778
rect 42156 406224 42208 406230
rect 42156 406166 42208 406172
rect 42168 405929 42196 406166
rect 42260 405686 42288 408870
rect 42340 407924 42392 407930
rect 42340 407866 42392 407872
rect 42248 405680 42300 405686
rect 42248 405622 42300 405628
rect 42248 405544 42300 405550
rect 42248 405486 42300 405492
rect 42156 403912 42208 403918
rect 42156 403854 42208 403860
rect 42168 403444 42196 403854
rect 42156 403368 42208 403374
rect 42156 403310 42208 403316
rect 42168 402801 42196 403310
rect 42260 402166 42288 405486
rect 42352 402966 42380 407866
rect 42720 405210 42748 425575
rect 43350 421560 43406 421569
rect 43350 421495 43406 421504
rect 43258 421152 43314 421161
rect 43258 421087 43314 421096
rect 43168 416696 43220 416702
rect 43168 416638 43220 416644
rect 43076 416628 43128 416634
rect 43076 416570 43128 416576
rect 43088 411262 43116 416570
rect 43076 411256 43128 411262
rect 43076 411198 43128 411204
rect 43076 410848 43128 410854
rect 43076 410790 43128 410796
rect 43088 405550 43116 410790
rect 43180 407658 43208 416638
rect 43272 408066 43300 421087
rect 43260 408060 43312 408066
rect 43260 408002 43312 408008
rect 43168 407652 43220 407658
rect 43168 407594 43220 407600
rect 43364 406842 43392 421495
rect 43352 406836 43404 406842
rect 43352 406778 43404 406784
rect 43076 405544 43128 405550
rect 43076 405486 43128 405492
rect 42432 405204 42484 405210
rect 42432 405146 42484 405152
rect 42708 405204 42760 405210
rect 42708 405146 42760 405152
rect 42340 402960 42392 402966
rect 42340 402902 42392 402908
rect 42340 402824 42392 402830
rect 42340 402766 42392 402772
rect 42182 402138 42288 402166
rect 42352 401622 42380 402766
rect 42182 401594 42380 401622
rect 42340 400648 42392 400654
rect 42340 400590 42392 400596
rect 42352 399786 42380 400590
rect 42182 399758 42380 399786
rect 42340 399696 42392 399702
rect 42340 399638 42392 399644
rect 42352 399135 42380 399638
rect 42182 399107 42380 399135
rect 42444 398494 42472 405146
rect 43456 400654 43484 426391
rect 43534 425232 43590 425241
rect 43534 425167 43590 425176
rect 43548 402830 43576 425167
rect 43626 424824 43682 424833
rect 43626 424759 43682 424768
rect 43640 406230 43668 424759
rect 43628 406224 43680 406230
rect 43628 406166 43680 406172
rect 43536 402824 43588 402830
rect 43536 402766 43588 402772
rect 43444 400648 43496 400654
rect 43444 400590 43496 400596
rect 42182 398466 42472 398494
rect 42168 394670 42196 397936
rect 42156 394664 42208 394670
rect 42156 394606 42208 394612
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41512 387864 41564 387870
rect 41512 387806 41564 387812
rect 41524 387569 41552 387806
rect 41788 387796 41840 387802
rect 41788 387738 41840 387744
rect 41800 387705 41828 387738
rect 41786 387696 41842 387705
rect 41786 387631 41842 387640
rect 41510 387560 41566 387569
rect 41510 387495 41566 387504
rect 41510 386744 41566 386753
rect 41510 386679 41512 386688
rect 41564 386679 41566 386688
rect 41512 386650 41564 386656
rect 43732 385665 43760 428431
rect 43902 424008 43958 424017
rect 43902 423943 43958 423952
rect 43810 423600 43866 423609
rect 43810 423535 43866 423544
rect 43824 410854 43852 423535
rect 43916 417194 43944 423943
rect 43994 423192 44050 423201
rect 43994 423127 44050 423136
rect 44008 417330 44036 423127
rect 44086 421968 44142 421977
rect 44086 421903 44142 421912
rect 44100 417466 44128 421903
rect 44100 417438 44220 417466
rect 44008 417302 44128 417330
rect 43916 417166 44036 417194
rect 43812 410848 43864 410854
rect 43812 410790 43864 410796
rect 44008 409902 44036 417166
rect 43812 409896 43864 409902
rect 43812 409838 43864 409844
rect 43996 409896 44048 409902
rect 43996 409838 44048 409844
rect 43824 399702 43852 409838
rect 43996 409760 44048 409766
rect 43996 409702 44048 409708
rect 44008 403918 44036 409702
rect 43996 403912 44048 403918
rect 43996 403854 44048 403860
rect 44100 403374 44128 417302
rect 44192 409766 44220 417438
rect 44180 409760 44232 409766
rect 44180 409702 44232 409708
rect 44088 403368 44140 403374
rect 44088 403310 44140 403316
rect 43812 399696 43864 399702
rect 43812 399638 43864 399644
rect 44610 386524 44638 429260
rect 44702 428094 44730 555198
rect 44794 554897 44822 597607
rect 44778 554888 44838 554897
rect 44778 554819 44838 554828
rect 44794 554818 44822 554819
rect 44794 554485 44822 554490
rect 44778 554476 44838 554485
rect 44778 554407 44838 554416
rect 44686 428084 44746 428094
rect 44686 428014 44746 428024
rect 44702 427678 44730 427694
rect 44686 427668 44746 427678
rect 44686 427598 44746 427608
rect 44594 386514 44654 386524
rect 44594 386444 44654 386454
rect 44610 386436 44638 386444
rect 44610 386140 44638 386152
rect 44594 386130 44654 386140
rect 44594 386060 44654 386070
rect 43718 385656 43774 385665
rect 43718 385591 43774 385600
rect 43534 385248 43590 385257
rect 43534 385183 43590 385192
rect 43442 383208 43498 383217
rect 43442 383143 43498 383152
rect 42706 382800 42762 382809
rect 42706 382735 42762 382744
rect 38198 381032 38254 381041
rect 38198 380967 38254 380976
rect 38212 375358 38240 380967
rect 41970 379944 42026 379953
rect 41970 379879 42026 379888
rect 41602 378584 41658 378593
rect 41602 378519 41658 378528
rect 41418 378176 41474 378185
rect 41418 378111 41474 378120
rect 38200 375352 38252 375358
rect 38200 375294 38252 375300
rect 41432 375290 41460 378111
rect 41510 377768 41566 377777
rect 41510 377703 41566 377712
rect 41420 375284 41472 375290
rect 41420 375226 41472 375232
rect 41524 371482 41552 377703
rect 41616 372842 41644 378519
rect 41786 377496 41842 377505
rect 41786 377431 41842 377440
rect 41800 376281 41828 377431
rect 41786 376272 41842 376281
rect 41786 376207 41788 376216
rect 41840 376207 41842 376216
rect 41788 376178 41840 376184
rect 41604 372836 41656 372842
rect 41604 372778 41656 372784
rect 41512 371476 41564 371482
rect 41512 371418 41564 371424
rect 41984 370258 42012 379879
rect 42248 375352 42300 375358
rect 42248 375294 42300 375300
rect 41972 370252 42024 370258
rect 41972 370194 42024 370200
rect 42260 369458 42288 375294
rect 42720 374270 42748 382735
rect 43074 381984 43130 381993
rect 43074 381919 43130 381928
rect 42340 374264 42392 374270
rect 42340 374206 42392 374212
rect 42708 374264 42760 374270
rect 42708 374206 42760 374212
rect 42182 369430 42288 369458
rect 42248 369368 42300 369374
rect 42248 369310 42300 369316
rect 42156 368144 42208 368150
rect 42156 368086 42208 368092
rect 42168 367608 42196 368086
rect 42260 367554 42288 369310
rect 42352 368150 42380 374206
rect 42708 371476 42760 371482
rect 42708 371418 42760 371424
rect 42340 368144 42392 368150
rect 42340 368086 42392 368092
rect 42260 367526 42380 367554
rect 42182 366947 42288 366975
rect 42156 366308 42208 366314
rect 42156 366250 42208 366256
rect 42168 365772 42196 366250
rect 42260 365242 42288 366947
rect 42352 366178 42380 367526
rect 42340 366172 42392 366178
rect 42340 366114 42392 366120
rect 42260 365214 42380 365242
rect 42168 364970 42196 365121
rect 42352 365090 42380 365214
rect 42340 365084 42392 365090
rect 42340 365026 42392 365032
rect 42168 364942 42380 364970
rect 42156 364812 42208 364818
rect 42156 364754 42208 364760
rect 42168 364548 42196 364754
rect 42248 364132 42300 364138
rect 42248 364074 42300 364080
rect 42260 363950 42288 364074
rect 42182 363922 42288 363950
rect 42156 363860 42208 363866
rect 42156 363802 42208 363808
rect 42168 363256 42196 363802
rect 42156 363180 42208 363186
rect 42156 363122 42208 363128
rect 42168 362712 42196 363122
rect 42352 361622 42380 364942
rect 42720 364818 42748 371418
rect 42708 364812 42760 364818
rect 42708 364754 42760 364760
rect 42708 364676 42760 364682
rect 42708 364618 42760 364624
rect 42432 361956 42484 361962
rect 42432 361898 42484 361904
rect 42340 361616 42392 361622
rect 42340 361558 42392 361564
rect 42064 360664 42116 360670
rect 42064 360606 42116 360612
rect 42076 360264 42104 360606
rect 42340 360324 42392 360330
rect 42340 360266 42392 360272
rect 42156 359984 42208 359990
rect 42156 359926 42208 359932
rect 42168 359584 42196 359926
rect 42352 358986 42380 360266
rect 42182 358958 42380 358986
rect 42444 358442 42472 361898
rect 42720 361350 42748 364618
rect 43088 361962 43116 381919
rect 43258 381576 43314 381585
rect 43258 381511 43314 381520
rect 43166 379536 43222 379545
rect 43166 379471 43222 379480
rect 43180 366314 43208 379471
rect 43272 379386 43300 381511
rect 43456 379506 43484 383143
rect 43444 379500 43496 379506
rect 43444 379442 43496 379448
rect 43272 379358 43484 379386
rect 43548 379370 43576 385183
rect 43718 382392 43774 382401
rect 43718 382327 43774 382336
rect 43732 380894 43760 382327
rect 43640 380866 43760 380894
rect 43456 379250 43484 379358
rect 43536 379364 43588 379370
rect 43536 379306 43588 379312
rect 43352 379228 43404 379234
rect 43456 379222 43576 379250
rect 43352 379170 43404 379176
rect 43260 375284 43312 375290
rect 43260 375226 43312 375232
rect 43168 366308 43220 366314
rect 43168 366250 43220 366256
rect 43168 366172 43220 366178
rect 43168 366114 43220 366120
rect 43180 363798 43208 366114
rect 43272 363866 43300 375226
rect 43260 363860 43312 363866
rect 43260 363802 43312 363808
rect 43168 363792 43220 363798
rect 43168 363734 43220 363740
rect 43076 361956 43128 361962
rect 43076 361898 43128 361904
rect 42708 361344 42760 361350
rect 42708 361286 42760 361292
rect 42168 358306 42196 358428
rect 42260 358414 42472 358442
rect 42260 358306 42288 358414
rect 43364 358358 43392 379170
rect 43442 379128 43498 379137
rect 43442 379063 43498 379072
rect 43456 364138 43484 379063
rect 43444 364132 43496 364138
rect 43444 364074 43496 364080
rect 43444 363996 43496 364002
rect 43444 363938 43496 363944
rect 43456 360330 43484 363938
rect 43548 363186 43576 379222
rect 43536 363180 43588 363186
rect 43536 363122 43588 363128
rect 43444 360324 43496 360330
rect 43444 360266 43496 360272
rect 42168 358278 42288 358306
rect 42432 358352 42484 358358
rect 42432 358294 42484 358300
rect 43352 358352 43404 358358
rect 43352 358294 43404 358300
rect 42444 356606 42472 358294
rect 42168 356538 42196 356592
rect 42260 356578 42472 356606
rect 42260 356538 42288 356578
rect 42168 356510 42288 356538
rect 43640 356522 43668 380866
rect 43718 380760 43774 380769
rect 43718 380695 43774 380704
rect 43732 371346 43760 380695
rect 43902 380352 43958 380361
rect 43902 380287 43958 380296
rect 43720 371340 43772 371346
rect 43720 371282 43772 371288
rect 43812 371136 43864 371142
rect 43812 371078 43864 371084
rect 42432 356516 42484 356522
rect 42432 356458 42484 356464
rect 43628 356516 43680 356522
rect 43628 356458 43680 356464
rect 42340 356448 42392 356454
rect 42340 356390 42392 356396
rect 42352 355926 42380 356390
rect 42182 355898 42380 355926
rect 42444 355314 42472 356458
rect 43824 356454 43852 371078
rect 43916 364002 43944 380287
rect 44088 379364 44140 379370
rect 44088 379306 44140 379312
rect 43996 372836 44048 372842
rect 43996 372778 44048 372784
rect 43904 363996 43956 364002
rect 43904 363938 43956 363944
rect 44008 363882 44036 372778
rect 43916 363854 44036 363882
rect 43916 360670 43944 363854
rect 43996 363792 44048 363798
rect 43996 363734 44048 363740
rect 43904 360664 43956 360670
rect 43904 360606 43956 360612
rect 44008 359990 44036 363734
rect 43996 359984 44048 359990
rect 43996 359926 44048 359932
rect 43812 356448 43864 356454
rect 43812 356390 43864 356396
rect 42168 355178 42196 355300
rect 42260 355286 42472 355314
rect 42260 355178 42288 355286
rect 42168 355150 42288 355178
rect 42168 350538 42196 354725
rect 42156 350532 42208 350538
rect 42156 350474 42208 350480
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 41510 344312 41566 344321
rect 41510 344247 41512 344256
rect 41564 344247 41566 344256
rect 41512 344218 41564 344224
rect 41510 343904 41566 343913
rect 41510 343839 41512 343848
rect 41564 343839 41566 343848
rect 41512 343810 41564 343816
rect 41510 343496 41566 343505
rect 41510 343431 41512 343440
rect 41564 343431 41566 343440
rect 41512 343402 41564 343408
rect 44100 342922 44128 379306
rect 44610 343324 44638 386060
rect 44702 384888 44730 427598
rect 44794 427297 44822 554407
rect 45744 546916 45796 546922
rect 45744 546858 45796 546864
rect 44778 427288 44838 427297
rect 44778 427219 44838 427228
rect 44794 427208 44822 427219
rect 44794 426885 44822 426892
rect 44778 426876 44838 426885
rect 44778 426807 44838 426816
rect 44686 384878 44746 384888
rect 44686 384808 44746 384818
rect 44702 384790 44730 384808
rect 44702 384478 44730 384494
rect 44686 384468 44746 384478
rect 44686 384398 44746 384408
rect 44594 343314 44654 343324
rect 44594 343244 44654 343254
rect 44594 342930 44654 342940
rect 41512 342916 41564 342922
rect 41512 342858 41564 342864
rect 44088 342916 44140 342922
rect 44088 342858 44140 342864
rect 44594 342860 44654 342870
rect 41524 342689 41552 342858
rect 41510 342680 41566 342689
rect 41510 342615 41566 342624
rect 43350 342136 43406 342145
rect 43350 342071 43406 342080
rect 32862 339824 32918 339833
rect 32862 339759 32918 339768
rect 33046 339824 33102 339833
rect 33046 339759 33102 339768
rect 32876 329769 32904 339759
rect 33060 330002 33088 339759
rect 43166 338464 43222 338473
rect 43166 338399 43222 338408
rect 41786 338056 41842 338065
rect 41786 337991 41842 338000
rect 41510 336968 41566 336977
rect 41510 336903 41566 336912
rect 41418 336560 41474 336569
rect 41418 336495 41474 336504
rect 41432 331226 41460 336495
rect 41420 331220 41472 331226
rect 41420 331162 41472 331168
rect 41524 330138 41552 336903
rect 41602 334112 41658 334121
rect 41602 334047 41658 334056
rect 41616 332897 41644 334047
rect 41602 332888 41658 332897
rect 41602 332823 41604 332832
rect 41656 332823 41658 332832
rect 41604 332794 41656 332800
rect 41512 330132 41564 330138
rect 41512 330074 41564 330080
rect 33048 329996 33100 330002
rect 33048 329938 33100 329944
rect 32862 329760 32918 329769
rect 32862 329695 32918 329704
rect 41800 327010 41828 337991
rect 42338 336424 42394 336433
rect 42338 336359 42394 336368
rect 42248 329996 42300 330002
rect 42248 329938 42300 329944
rect 41788 327004 41840 327010
rect 41788 326946 41840 326952
rect 41788 326800 41840 326806
rect 41788 326742 41840 326748
rect 41800 326264 41828 326742
rect 42168 324306 42196 324428
rect 42260 324306 42288 329938
rect 42168 324278 42288 324306
rect 42182 323734 42288 323762
rect 42260 323202 42288 323734
rect 42248 323196 42300 323202
rect 42248 323138 42300 323144
rect 42352 323082 42380 336359
rect 42706 335608 42762 335617
rect 42706 335543 42762 335552
rect 42168 323054 42380 323082
rect 42168 322934 42196 323054
rect 42248 322992 42300 322998
rect 42248 322934 42300 322940
rect 42076 322906 42196 322934
rect 42076 322592 42104 322906
rect 42260 322046 42288 322934
rect 42248 322040 42300 322046
rect 42248 321982 42300 321988
rect 42182 321898 42380 321926
rect 42248 321836 42300 321842
rect 42248 321778 42300 321784
rect 42156 321632 42208 321638
rect 42156 321574 42208 321580
rect 42168 321368 42196 321574
rect 42260 320739 42288 321778
rect 42182 320711 42288 320739
rect 42248 320612 42300 320618
rect 42248 320554 42300 320560
rect 42156 320476 42208 320482
rect 42156 320418 42208 320424
rect 42168 320076 42196 320418
rect 42260 319546 42288 320554
rect 42182 319518 42288 319546
rect 42352 317422 42380 321898
rect 42720 318782 42748 335543
rect 43076 330132 43128 330138
rect 43076 330074 43128 330080
rect 42432 318776 42484 318782
rect 42432 318718 42484 318724
rect 42708 318776 42760 318782
rect 42708 318718 42760 318724
rect 42340 317416 42392 317422
rect 42340 317358 42392 317364
rect 42444 317059 42472 318718
rect 42182 317031 42472 317059
rect 43088 316946 43116 330074
rect 43180 320618 43208 338399
rect 43258 336016 43314 336025
rect 43258 335951 43314 335960
rect 43272 321842 43300 335951
rect 43260 321836 43312 321842
rect 43260 321778 43312 321784
rect 43168 320612 43220 320618
rect 43168 320554 43220 320560
rect 42432 316940 42484 316946
rect 42432 316882 42484 316888
rect 43076 316940 43128 316946
rect 43076 316882 43128 316888
rect 42340 316872 42392 316878
rect 42340 316814 42392 316820
rect 42352 316418 42380 316814
rect 42182 316390 42380 316418
rect 42444 315771 42472 316882
rect 42182 315743 42472 315771
rect 41970 315616 42026 315625
rect 41970 315551 42026 315560
rect 41984 315180 42012 315551
rect 42154 313848 42210 313857
rect 42154 313783 42210 313792
rect 42168 313344 42196 313783
rect 41786 313168 41842 313177
rect 41786 313103 41842 313112
rect 41800 312732 41828 313103
rect 41786 312352 41842 312361
rect 41786 312287 41842 312296
rect 41800 312052 41828 312287
rect 42076 306338 42104 311508
rect 42064 306332 42116 306338
rect 42064 306274 42116 306280
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41880 301436 41932 301442
rect 41880 301378 41932 301384
rect 41788 301368 41840 301374
rect 41786 301336 41788 301345
rect 41840 301336 41842 301345
rect 41786 301271 41842 301280
rect 41788 301232 41840 301238
rect 41788 301174 41840 301180
rect 41800 299305 41828 301174
rect 41892 300937 41920 301378
rect 43364 301238 43392 342071
rect 43626 335200 43682 335209
rect 43626 335135 43682 335144
rect 43442 334792 43498 334801
rect 43442 334727 43498 334736
rect 43456 321638 43484 334727
rect 43536 331220 43588 331226
rect 43536 331162 43588 331168
rect 43444 321632 43496 321638
rect 43444 321574 43496 321580
rect 43548 316878 43576 331162
rect 43640 320482 43668 335135
rect 43720 322040 43772 322046
rect 43720 321982 43772 321988
rect 43628 320476 43680 320482
rect 43628 320418 43680 320424
rect 43732 318782 43760 321982
rect 43720 318776 43772 318782
rect 43720 318718 43772 318724
rect 43536 316872 43588 316878
rect 43536 316814 43588 316820
rect 43352 301232 43404 301238
rect 43352 301174 43404 301180
rect 41878 300928 41934 300937
rect 41878 300863 41934 300872
rect 42706 300520 42762 300529
rect 42706 300455 42762 300464
rect 41786 299296 41842 299305
rect 41786 299231 41842 299240
rect 42720 298217 42748 300455
rect 44610 300124 44638 342860
rect 44702 341688 44730 384398
rect 44794 384097 44822 426807
rect 44778 384088 44838 384097
rect 44778 384019 44838 384028
rect 44794 384012 44822 384019
rect 44794 383685 44822 383692
rect 44778 383676 44838 383685
rect 44778 383607 44838 383616
rect 44686 341678 44746 341688
rect 44686 341608 44746 341618
rect 44686 341268 44746 341278
rect 44686 341198 44746 341208
rect 44594 300114 44654 300124
rect 44594 300044 44654 300054
rect 44610 299740 44638 299744
rect 44594 299730 44654 299740
rect 44594 299660 44654 299670
rect 43074 298888 43130 298897
rect 43074 298823 43130 298832
rect 42706 298208 42762 298217
rect 42706 298143 42762 298152
rect 42340 295384 42392 295390
rect 42340 295326 42392 295332
rect 41878 294808 41934 294817
rect 41878 294743 41934 294752
rect 30010 292768 30066 292777
rect 30010 292703 30066 292712
rect 30024 288862 30052 292703
rect 41786 291952 41842 291961
rect 41786 291887 41788 291896
rect 41840 291887 41842 291896
rect 41788 291858 41840 291864
rect 41786 291544 41842 291553
rect 41786 291479 41842 291488
rect 41800 289882 41828 291479
rect 41788 289876 41840 289882
rect 41788 289818 41840 289824
rect 30012 288856 30064 288862
rect 30012 288798 30064 288804
rect 41892 283830 41920 294743
rect 42248 288448 42300 288454
rect 42248 288390 42300 288396
rect 41880 283824 41932 283830
rect 41880 283766 41932 283772
rect 41880 283620 41932 283626
rect 41880 283562 41932 283568
rect 41892 283045 41920 283562
rect 42156 281784 42208 281790
rect 42156 281726 42208 281732
rect 42168 281180 42196 281726
rect 42156 281104 42208 281110
rect 42156 281046 42208 281052
rect 42168 280568 42196 281046
rect 42156 279880 42208 279886
rect 42156 279822 42208 279828
rect 42168 279344 42196 279822
rect 42156 279268 42208 279274
rect 42156 279210 42208 279216
rect 42168 278732 42196 279210
rect 42064 278656 42116 278662
rect 42064 278598 42116 278604
rect 42076 278188 42104 278598
rect 42260 277794 42288 288390
rect 42352 281110 42380 295326
rect 42430 293992 42486 294001
rect 42430 293927 42486 293936
rect 42444 285530 42472 293927
rect 42708 289876 42760 289882
rect 42708 289818 42760 289824
rect 42432 285524 42484 285530
rect 42432 285466 42484 285472
rect 42340 281104 42392 281110
rect 42340 281046 42392 281052
rect 42340 280492 42392 280498
rect 42340 280434 42392 280440
rect 42168 277766 42288 277794
rect 42168 277508 42196 277766
rect 42352 276910 42380 280434
rect 42720 278662 42748 289818
rect 43088 285666 43116 298823
rect 43626 296440 43682 296449
rect 43626 296375 43682 296384
rect 43258 296032 43314 296041
rect 43258 295967 43314 295976
rect 43166 293176 43222 293185
rect 43166 293111 43222 293120
rect 43076 285660 43128 285666
rect 43076 285602 43128 285608
rect 43076 285524 43128 285530
rect 43076 285466 43128 285472
rect 42708 278656 42760 278662
rect 42708 278598 42760 278604
rect 42708 278520 42760 278526
rect 42708 278462 42760 278468
rect 42182 276882 42380 276910
rect 42340 276820 42392 276826
rect 42340 276762 42392 276768
rect 42248 276752 42300 276758
rect 42248 276694 42300 276700
rect 42064 276616 42116 276622
rect 42064 276558 42116 276564
rect 42076 276352 42104 276558
rect 42156 274304 42208 274310
rect 42156 274246 42208 274252
rect 42168 273836 42196 274246
rect 42064 273556 42116 273562
rect 42064 273498 42116 273504
rect 42076 273224 42104 273498
rect 42260 272558 42288 276694
rect 42182 272530 42288 272558
rect 42352 272014 42380 276762
rect 42720 275602 42748 278462
rect 43088 276758 43116 285466
rect 43180 279886 43208 293111
rect 43168 279880 43220 279886
rect 43168 279822 43220 279828
rect 43076 276752 43128 276758
rect 43076 276694 43128 276700
rect 42432 275596 42484 275602
rect 42432 275538 42484 275544
rect 42708 275596 42760 275602
rect 42708 275538 42760 275544
rect 42182 271986 42380 272014
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 41800 270164 41828 270399
rect 42444 269535 42472 275538
rect 42182 269507 42472 269535
rect 43272 269414 43300 295967
rect 43534 295216 43590 295225
rect 43534 295151 43590 295160
rect 43352 292596 43404 292602
rect 43352 292538 43404 292544
rect 43364 279274 43392 292538
rect 43444 291916 43496 291922
rect 43444 291858 43496 291864
rect 43456 280498 43484 291858
rect 43444 280492 43496 280498
rect 43444 280434 43496 280440
rect 43352 279268 43404 279274
rect 43352 279210 43404 279216
rect 43548 276622 43576 295151
rect 43640 281790 43668 296375
rect 43718 295624 43774 295633
rect 43718 295559 43774 295568
rect 43732 295334 43760 295559
rect 43732 295306 43852 295334
rect 43720 285660 43772 285666
rect 43720 285602 43772 285608
rect 43628 281784 43680 281790
rect 43628 281726 43680 281732
rect 43628 281648 43680 281654
rect 43628 281590 43680 281596
rect 43536 276616 43588 276622
rect 43536 276558 43588 276564
rect 43640 273562 43668 281590
rect 43628 273556 43680 273562
rect 43628 273498 43680 273504
rect 42432 269408 42484 269414
rect 42432 269350 42484 269356
rect 43260 269408 43312 269414
rect 43260 269350 43312 269356
rect 42444 268886 42472 269350
rect 42182 268858 42472 268886
rect 42168 264790 42196 268328
rect 42156 264784 42208 264790
rect 42156 264726 42208 264732
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 41788 258120 41840 258126
rect 41786 258088 41788 258097
rect 41840 258088 41842 258097
rect 41786 258023 41842 258032
rect 41512 257984 41564 257990
rect 41510 257952 41512 257961
rect 41564 257952 41566 257961
rect 41510 257887 41566 257896
rect 41512 257576 41564 257582
rect 41510 257544 41512 257553
rect 41564 257544 41566 257553
rect 41510 257479 41566 257488
rect 43732 256057 43760 285602
rect 43824 276826 43852 295306
rect 43902 294400 43958 294409
rect 43902 294335 43958 294344
rect 43916 278526 43944 294335
rect 43994 293584 44050 293593
rect 43994 293519 44050 293528
rect 44008 284306 44036 293519
rect 44086 292360 44142 292369
rect 44086 292295 44142 292304
rect 44100 284458 44128 292295
rect 44100 284430 44220 284458
rect 43996 284300 44048 284306
rect 43996 284242 44048 284248
rect 44192 284186 44220 284430
rect 44272 284300 44324 284306
rect 44272 284242 44324 284248
rect 44100 284158 44220 284186
rect 43904 278520 43956 278526
rect 43904 278462 43956 278468
rect 43812 276820 43864 276826
rect 43812 276762 43864 276768
rect 44100 274310 44128 284158
rect 44284 281654 44312 284242
rect 44272 281648 44324 281654
rect 44272 281590 44324 281596
rect 44088 274304 44140 274310
rect 44088 274246 44140 274252
rect 44610 256923 44638 299660
rect 44702 298488 44730 341198
rect 44794 340897 44822 383607
rect 44778 340888 44838 340897
rect 44778 340819 44838 340828
rect 44794 340814 44822 340819
rect 44794 340485 44822 340494
rect 44778 340476 44838 340485
rect 44778 340407 44838 340416
rect 44686 298478 44746 298488
rect 44686 298408 44746 298418
rect 44702 298406 44730 298408
rect 44686 298068 44746 298078
rect 44686 297998 44746 298008
rect 44594 256914 44654 256923
rect 44594 256845 44654 256854
rect 44610 256840 44638 256845
rect 44610 256539 44638 256546
rect 44594 256530 44654 256539
rect 44594 256461 44654 256470
rect 43718 256048 43774 256057
rect 43718 255983 43774 255992
rect 42246 255640 42302 255649
rect 42246 255575 42302 255584
rect 30102 251424 30158 251433
rect 30102 251359 30158 251368
rect 30116 245886 30144 251359
rect 38106 248976 38162 248985
rect 38106 248911 38162 248920
rect 20720 245880 20772 245886
rect 20720 245822 20772 245828
rect 30104 245880 30156 245886
rect 30104 245822 30156 245828
rect 20732 244390 20760 245822
rect 38120 245478 38148 248911
rect 38198 248568 38254 248577
rect 38198 248503 38254 248512
rect 38108 245472 38160 245478
rect 38108 245414 38160 245420
rect 38212 245410 38240 248503
rect 41510 248160 41566 248169
rect 41510 248095 41566 248104
rect 41418 247752 41474 247761
rect 41418 247687 41420 247696
rect 41472 247687 41474 247696
rect 41420 247658 41472 247664
rect 41418 247344 41474 247353
rect 41418 247279 41474 247288
rect 41432 245682 41460 247279
rect 41524 246974 41552 248095
rect 41512 246968 41564 246974
rect 41512 246910 41564 246916
rect 41510 246528 41566 246537
rect 41510 246463 41566 246472
rect 41524 245750 41552 246463
rect 41512 245744 41564 245750
rect 41512 245686 41564 245692
rect 41420 245676 41472 245682
rect 41420 245618 41472 245624
rect 38200 245404 38252 245410
rect 38200 245346 38252 245352
rect 42260 244474 42288 255575
rect 42338 253600 42394 253609
rect 42338 253535 42394 253544
rect 42352 244594 42380 253535
rect 43810 253192 43866 253201
rect 43810 253127 43866 253136
rect 43258 252376 43314 252385
rect 43258 252311 43314 252320
rect 42706 249928 42762 249937
rect 42706 249863 42762 249872
rect 42340 244588 42392 244594
rect 42340 244530 42392 244536
rect 42260 244446 42380 244474
rect 20720 244384 20772 244390
rect 20720 244326 20772 244332
rect 42248 244384 42300 244390
rect 42248 244326 42300 244332
rect 42260 239850 42288 244326
rect 42182 239822 42288 239850
rect 42248 239760 42300 239766
rect 42248 239702 42300 239708
rect 42156 238536 42208 238542
rect 42156 238478 42208 238484
rect 42168 238000 42196 238478
rect 42260 236178 42288 239702
rect 42182 236150 42288 236178
rect 42248 236088 42300 236094
rect 42248 236030 42300 236036
rect 42156 235408 42208 235414
rect 42156 235350 42208 235356
rect 42168 234969 42196 235350
rect 42156 234660 42208 234666
rect 42156 234602 42208 234608
rect 42168 234328 42196 234602
rect 42260 233695 42288 236030
rect 42182 233667 42288 233695
rect 42248 233572 42300 233578
rect 42248 233514 42300 233520
rect 42156 233368 42208 233374
rect 42156 233310 42208 233316
rect 42168 233104 42196 233310
rect 42260 230670 42288 233514
rect 42182 230642 42288 230670
rect 42248 230580 42300 230586
rect 42248 230522 42300 230528
rect 42156 230376 42208 230382
rect 42156 230318 42208 230324
rect 42168 229976 42196 230318
rect 42156 229900 42208 229906
rect 42156 229842 42208 229848
rect 42168 229364 42196 229842
rect 42260 228834 42288 230522
rect 42182 228806 42288 228834
rect 42064 227384 42116 227390
rect 42064 227326 42116 227332
rect 42076 226984 42104 227326
rect 42156 226840 42208 226846
rect 42156 226782 42208 226788
rect 42168 226304 42196 226782
rect 41786 225992 41842 226001
rect 41786 225927 41842 225936
rect 41800 225692 41828 225927
rect 41696 222216 41748 222222
rect 41696 222158 41748 222164
rect 8208 217932 8260 217938
rect 8208 217874 8260 217880
rect 8220 202473 8248 217874
rect 41512 216708 41564 216714
rect 41512 216650 41564 216656
rect 41420 216640 41472 216646
rect 41420 216582 41472 216588
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 31668 215416 31720 215422
rect 31668 215358 31720 215364
rect 30102 204096 30158 204105
rect 30102 204031 30158 204040
rect 30116 202473 30144 204031
rect 31680 203697 31708 215358
rect 41432 214305 41460 216582
rect 41524 214713 41552 216650
rect 41708 215121 41736 222158
rect 42168 220794 42196 225148
rect 42156 220788 42208 220794
rect 42156 220730 42208 220736
rect 41694 215112 41750 215121
rect 41694 215047 41750 215056
rect 41510 214704 41566 214713
rect 41510 214639 41566 214648
rect 41418 214296 41474 214305
rect 41418 214231 41474 214240
rect 41512 213308 41564 213314
rect 41512 213250 41564 213256
rect 41524 212673 41552 213250
rect 42352 212945 42380 244446
rect 42720 239766 42748 249863
rect 43074 249520 43130 249529
rect 43074 249455 43130 249464
rect 43088 245562 43116 249455
rect 43272 245614 43300 252311
rect 43534 251968 43590 251977
rect 43534 251903 43590 251912
rect 43352 246968 43404 246974
rect 43352 246910 43404 246916
rect 43260 245608 43312 245614
rect 43088 245534 43208 245562
rect 43260 245550 43312 245556
rect 43076 245404 43128 245410
rect 43076 245346 43128 245352
rect 42708 239760 42760 239766
rect 42708 239702 42760 239708
rect 43088 236094 43116 245346
rect 43076 236088 43128 236094
rect 43076 236030 43128 236036
rect 43180 234666 43208 245534
rect 43260 245472 43312 245478
rect 43260 245414 43312 245420
rect 43168 234660 43220 234666
rect 43168 234602 43220 234608
rect 43272 233578 43300 245414
rect 43364 235414 43392 246910
rect 43444 245540 43496 245546
rect 43444 245482 43496 245488
rect 43456 244730 43484 245482
rect 43444 244724 43496 244730
rect 43444 244666 43496 244672
rect 43444 244588 43496 244594
rect 43444 244530 43496 244536
rect 43352 235408 43404 235414
rect 43352 235350 43404 235356
rect 43260 233572 43312 233578
rect 43260 233514 43312 233520
rect 43456 227390 43484 244530
rect 43548 233374 43576 251903
rect 43626 251152 43682 251161
rect 43626 251087 43682 251096
rect 43536 233368 43588 233374
rect 43536 233310 43588 233316
rect 43444 227384 43496 227390
rect 43444 227326 43496 227332
rect 43640 226846 43668 251087
rect 43718 250744 43774 250753
rect 43718 250679 43774 250688
rect 43732 244866 43760 250679
rect 43720 244860 43772 244866
rect 43720 244802 43772 244808
rect 43720 244724 43772 244730
rect 43720 244666 43772 244672
rect 43732 230586 43760 244666
rect 43824 238542 43852 253127
rect 43994 250336 44050 250345
rect 43994 250271 44050 250280
rect 43904 244860 43956 244866
rect 43904 244802 43956 244808
rect 43812 238536 43864 238542
rect 43812 238478 43864 238484
rect 43720 230580 43772 230586
rect 43720 230522 43772 230528
rect 43916 229906 43944 244802
rect 44008 230382 44036 250271
rect 43996 230376 44048 230382
rect 43996 230318 44048 230324
rect 43904 229900 43956 229906
rect 43904 229842 43956 229848
rect 43628 226840 43680 226846
rect 43628 226782 43680 226788
rect 44610 213719 44638 256461
rect 44702 255287 44730 297998
rect 44794 297697 44822 340407
rect 44778 297688 44838 297697
rect 44778 297619 44838 297628
rect 44794 297614 44822 297619
rect 44794 297285 44822 297286
rect 44778 297276 44838 297285
rect 44778 297207 44838 297216
rect 44686 255278 44746 255287
rect 44686 255209 44746 255218
rect 44702 255206 44730 255209
rect 44702 254877 44730 254888
rect 44686 254868 44746 254877
rect 44686 254799 44746 254808
rect 44592 213710 44648 213719
rect 44592 213645 44648 213654
rect 44610 213642 44638 213645
rect 42338 212936 42394 212945
rect 42338 212871 42394 212880
rect 41510 212664 41566 212673
rect 41510 212599 41566 212608
rect 44702 212085 44730 254799
rect 44794 254497 44822 297207
rect 44778 254488 44838 254497
rect 44778 254419 44838 254428
rect 44794 254412 44822 254419
rect 44794 254085 44822 254094
rect 44778 254076 44838 254085
rect 44778 254007 44838 254016
rect 44688 212076 44744 212085
rect 44688 212011 44744 212020
rect 44702 211996 44730 212011
rect 44794 211275 44822 254007
rect 45652 247716 45704 247722
rect 45652 247658 45704 247664
rect 45664 230518 45692 247658
rect 45652 230512 45704 230518
rect 45652 230454 45704 230460
rect 45756 219774 45784 546858
rect 45928 419484 45980 419490
rect 45928 419426 45980 419432
rect 45940 230722 45968 419426
rect 46020 376236 46072 376242
rect 46020 376178 46072 376184
rect 45928 230716 45980 230722
rect 45928 230658 45980 230664
rect 46032 230586 46060 376178
rect 46572 344276 46624 344282
rect 46572 344218 46624 344224
rect 46388 343868 46440 343874
rect 46388 343810 46440 343816
rect 46204 332852 46256 332858
rect 46204 332794 46256 332800
rect 46112 287088 46164 287094
rect 46112 287030 46164 287036
rect 46124 257582 46152 287030
rect 46112 257576 46164 257582
rect 46112 257518 46164 257524
rect 46216 230654 46244 332794
rect 46400 311846 46428 343810
rect 46480 343460 46532 343466
rect 46480 343402 46532 343408
rect 46492 314634 46520 343402
rect 46480 314628 46532 314634
rect 46480 314570 46532 314576
rect 46584 314566 46612 344218
rect 46572 314560 46624 314566
rect 46572 314502 46624 314508
rect 46388 311840 46440 311846
rect 46388 311782 46440 311788
rect 48240 277438 48268 767382
rect 48320 762884 48372 762890
rect 48320 762826 48372 762832
rect 48332 277642 48360 762826
rect 51000 742422 51028 773842
rect 50988 742416 51040 742422
rect 50988 742358 51040 742364
rect 53760 742354 53788 774726
rect 59268 756288 59320 756294
rect 59268 756230 59320 756236
rect 58440 747924 58492 747930
rect 58440 747866 58492 747872
rect 58452 747697 58480 747866
rect 58438 747688 58494 747697
rect 58438 747623 58494 747632
rect 59280 746473 59308 756230
rect 59266 746464 59322 746473
rect 59266 746399 59322 746408
rect 58440 745272 58492 745278
rect 58440 745214 58492 745220
rect 58452 744977 58480 745214
rect 58532 745204 58584 745210
rect 58532 745146 58584 745152
rect 58438 744968 58494 744977
rect 58438 744903 58494 744912
rect 58544 744161 58572 745146
rect 58530 744152 58586 744161
rect 58530 744087 58586 744096
rect 58440 742416 58492 742422
rect 57978 742384 58034 742393
rect 53748 742348 53800 742354
rect 58440 742358 58492 742364
rect 57978 742319 57980 742328
rect 53748 742290 53800 742296
rect 58032 742319 58034 742328
rect 57980 742290 58032 742296
rect 58452 741849 58480 742358
rect 58438 741840 58494 741849
rect 58438 741775 58494 741784
rect 59634 729192 59690 729201
rect 59634 729127 59690 729136
rect 59266 729056 59322 729065
rect 59266 728991 59322 729000
rect 59280 728654 59308 728991
rect 59450 728920 59506 728929
rect 59450 728855 59506 728864
rect 59188 728626 59308 728654
rect 53748 717664 53800 717670
rect 53748 717606 53800 717612
rect 50988 687676 51040 687682
rect 50988 687618 51040 687624
rect 51000 656878 51028 687618
rect 50988 656872 51040 656878
rect 50988 656814 51040 656820
rect 50988 644088 51040 644094
rect 50988 644030 51040 644036
rect 48412 633276 48464 633282
rect 48412 633218 48464 633224
rect 48320 277636 48372 277642
rect 48320 277578 48372 277584
rect 48424 277574 48452 633218
rect 51000 615466 51028 644030
rect 50988 615460 51040 615466
rect 50988 615402 51040 615408
rect 50988 557592 51040 557598
rect 50988 557534 51040 557540
rect 51000 529922 51028 557534
rect 50988 529916 51040 529922
rect 50988 529858 51040 529864
rect 50988 386708 51040 386714
rect 50988 386650 51040 386656
rect 51000 358766 51028 386650
rect 50988 358760 51040 358766
rect 50988 358702 51040 358708
rect 50986 290728 51042 290737
rect 50986 290663 51042 290672
rect 48594 289912 48650 289921
rect 48594 289847 48650 289856
rect 48504 281580 48556 281586
rect 48504 281522 48556 281528
rect 48412 277568 48464 277574
rect 48412 277510 48464 277516
rect 48228 277432 48280 277438
rect 48228 277374 48280 277380
rect 46204 230648 46256 230654
rect 46204 230590 46256 230596
rect 46020 230580 46072 230586
rect 46020 230522 46072 230528
rect 45744 219768 45796 219774
rect 45744 219710 45796 219716
rect 47314 217155 47342 217158
rect 47298 217146 47358 217155
rect 47298 217077 47358 217086
rect 47314 211689 47342 217077
rect 47406 216889 47434 216896
rect 47390 216880 47450 216889
rect 47390 216811 47450 216820
rect 47298 211680 47358 211689
rect 47298 211611 47358 211620
rect 47314 211608 47342 211611
rect 44778 211266 44834 211275
rect 44778 211201 44834 211210
rect 44794 211192 44822 211201
rect 47406 210875 47434 216811
rect 47498 216613 47526 216618
rect 47482 216604 47542 216613
rect 47482 216535 47542 216544
rect 47498 213317 47526 216535
rect 48228 215484 48280 215490
rect 48228 215426 48280 215432
rect 47482 213308 47542 213317
rect 47482 213239 47542 213248
rect 47498 213236 47526 213239
rect 47390 210866 47450 210875
rect 47390 210797 47450 210806
rect 37830 210216 37886 210225
rect 37830 210151 37886 210160
rect 31666 203688 31722 203697
rect 31666 203623 31722 203632
rect 8206 202464 8262 202473
rect 8206 202399 8262 202408
rect 30102 202464 30158 202473
rect 30102 202399 30158 202408
rect 37844 198801 37872 210151
rect 38014 209808 38070 209817
rect 38014 209743 38070 209752
rect 37922 206952 37978 206961
rect 37922 206887 37978 206896
rect 37936 201482 37964 206887
rect 37924 201476 37976 201482
rect 37924 201418 37976 201424
rect 38028 200938 38056 209743
rect 38290 209400 38346 209409
rect 38290 209335 38346 209344
rect 38198 208992 38254 209001
rect 38198 208927 38254 208936
rect 38106 208584 38162 208593
rect 38106 208519 38162 208528
rect 38120 204406 38148 208519
rect 38212 204474 38240 208927
rect 38304 204513 38332 209335
rect 38566 208176 38622 208185
rect 38566 208111 38622 208120
rect 38382 207768 38438 207777
rect 38382 207703 38438 207712
rect 38396 204921 38424 207703
rect 38474 207360 38530 207369
rect 38474 207295 38530 207304
rect 38488 205086 38516 207295
rect 38476 205080 38528 205086
rect 38476 205022 38528 205028
rect 38382 204912 38438 204921
rect 38382 204847 38438 204856
rect 38290 204504 38346 204513
rect 38200 204468 38252 204474
rect 38290 204439 38346 204448
rect 38200 204410 38252 204416
rect 38108 204400 38160 204406
rect 38108 204342 38160 204348
rect 38580 204338 38608 208111
rect 42706 206816 42762 206825
rect 42706 206751 42762 206760
rect 42338 205184 42394 205193
rect 42338 205119 42394 205128
rect 38568 204332 38620 204338
rect 38568 204274 38620 204280
rect 42248 204332 42300 204338
rect 42248 204274 42300 204280
rect 38016 200932 38068 200938
rect 38016 200874 38068 200880
rect 37830 198792 37886 198801
rect 37830 198727 37886 198736
rect 42260 196670 42288 204274
rect 42182 196642 42288 196670
rect 42248 196580 42300 196586
rect 42248 196522 42300 196528
rect 42260 194834 42288 196522
rect 42182 194806 42288 194834
rect 42064 193520 42116 193526
rect 42064 193462 42116 193468
rect 42076 192984 42104 193462
rect 42352 191774 42380 205119
rect 42720 193526 42748 206751
rect 43258 206408 43314 206417
rect 43258 206343 43314 206352
rect 43074 205592 43130 205601
rect 43074 205527 43130 205536
rect 42708 193520 42760 193526
rect 42708 193462 42760 193468
rect 42182 191746 42380 191774
rect 43088 191690 43116 205527
rect 43168 200932 43220 200938
rect 43168 200874 43220 200880
rect 43180 196586 43208 200874
rect 43168 196580 43220 196586
rect 43168 196522 43220 196528
rect 42340 191684 42392 191690
rect 42340 191626 42392 191632
rect 43076 191684 43128 191690
rect 43076 191626 43128 191632
rect 42064 191480 42116 191486
rect 42064 191422 42116 191428
rect 42076 191148 42104 191422
rect 42352 190482 42380 191626
rect 43272 191486 43300 206343
rect 43442 206000 43498 206009
rect 43442 205935 43498 205944
rect 43352 204400 43404 204406
rect 43352 204342 43404 204348
rect 43260 191480 43312 191486
rect 43260 191422 43312 191428
rect 42182 190454 42380 190482
rect 43364 190398 43392 204342
rect 42340 190392 42392 190398
rect 42340 190334 42392 190340
rect 43352 190392 43404 190398
rect 43352 190334 43404 190340
rect 42352 189938 42380 190334
rect 42182 189910 42380 189938
rect 43456 189854 43484 205935
rect 43536 205080 43588 205086
rect 43536 205022 43588 205028
rect 42248 189848 42300 189854
rect 42248 189790 42300 189796
rect 43444 189848 43496 189854
rect 43444 189790 43496 189796
rect 42260 187459 42288 189790
rect 42340 189780 42392 189786
rect 42340 189722 42392 189728
rect 42182 187431 42288 187459
rect 42352 186810 42380 189722
rect 42432 189168 42484 189174
rect 42432 189110 42484 189116
rect 42182 186782 42380 186810
rect 42340 186720 42392 186726
rect 42340 186662 42392 186668
rect 42352 186198 42380 186662
rect 42168 186130 42196 186184
rect 42260 186170 42380 186198
rect 42260 186130 42288 186170
rect 42168 186102 42288 186130
rect 42444 185619 42472 189110
rect 43548 186726 43576 205022
rect 48240 204785 48268 215426
rect 48226 204776 48282 204785
rect 48226 204711 48282 204720
rect 43628 204468 43680 204474
rect 43628 204410 43680 204416
rect 43640 189174 43668 204410
rect 43720 201476 43772 201482
rect 43720 201418 43772 201424
rect 43732 189786 43760 201418
rect 43720 189780 43772 189786
rect 43720 189722 43772 189728
rect 43628 189168 43680 189174
rect 43628 189110 43680 189116
rect 43536 186720 43588 186726
rect 43536 186662 43588 186668
rect 42182 185591 42472 185619
rect 41878 184240 41934 184249
rect 41878 184175 41934 184184
rect 41892 183765 41920 184175
rect 41786 183424 41842 183433
rect 41786 183359 41842 183368
rect 41800 183124 41828 183359
rect 41786 182744 41842 182753
rect 41786 182679 41842 182688
rect 41800 182477 41828 182679
rect 48516 182170 48544 281522
rect 48608 219502 48636 289847
rect 51000 219706 51028 290663
rect 51080 284368 51132 284374
rect 51080 284310 51132 284316
rect 51092 257990 51120 284310
rect 51080 257984 51132 257990
rect 51080 257926 51132 257932
rect 52276 256760 52328 256766
rect 52276 256702 52328 256708
rect 52184 245812 52236 245818
rect 52184 245754 52236 245760
rect 52092 230848 52144 230854
rect 52092 230790 52144 230796
rect 50988 219700 51040 219706
rect 50988 219642 51040 219648
rect 48596 219496 48648 219502
rect 48596 219438 48648 219444
rect 42156 182164 42208 182170
rect 42156 182106 42208 182112
rect 48504 182164 48556 182170
rect 48504 182106 48556 182112
rect 42168 181900 42196 182106
rect 52104 51134 52132 230790
rect 52092 51128 52144 51134
rect 52092 51070 52144 51076
rect 52196 42770 52224 245754
rect 52288 47122 52316 256702
rect 52736 227724 52788 227730
rect 52736 227666 52788 227672
rect 52748 217410 52776 227666
rect 53564 222284 53616 222290
rect 53564 222226 53616 222232
rect 53576 217410 53604 222226
rect 53760 220046 53788 717606
rect 58532 703860 58584 703866
rect 58532 703802 58584 703808
rect 58544 702137 58572 703802
rect 58530 702128 58586 702137
rect 58530 702063 58586 702072
rect 59188 698193 59216 728626
rect 59360 714876 59412 714882
rect 59360 714818 59412 714824
rect 59268 712156 59320 712162
rect 59268 712098 59320 712104
rect 59280 703361 59308 712098
rect 59372 704449 59400 714818
rect 59358 704440 59414 704449
rect 59358 704375 59414 704384
rect 59266 703352 59322 703361
rect 59266 703287 59322 703296
rect 59464 700913 59492 728855
rect 59450 700904 59506 700913
rect 59450 700839 59506 700848
rect 59648 699689 59676 729127
rect 59634 699680 59690 699689
rect 59634 699615 59690 699624
rect 59174 698184 59230 698193
rect 59174 698119 59230 698128
rect 53840 688356 53892 688362
rect 53840 688298 53892 688304
rect 53852 656810 53880 688298
rect 60648 670812 60700 670818
rect 60648 670754 60700 670760
rect 60660 661201 60688 670754
rect 60646 661192 60702 661201
rect 60646 661127 60702 661136
rect 58440 659728 58492 659734
rect 58440 659670 58492 659676
rect 58452 658889 58480 659670
rect 58532 659660 58584 659666
rect 58532 659602 58584 659608
rect 58544 659569 58572 659602
rect 58624 659592 58676 659598
rect 58530 659560 58586 659569
rect 58624 659534 58676 659540
rect 58530 659495 58586 659504
rect 58438 658880 58494 658889
rect 58438 658815 58494 658824
rect 58636 657665 58664 659534
rect 58622 657656 58678 657665
rect 58622 657591 58678 657600
rect 58440 656872 58492 656878
rect 58440 656814 58492 656820
rect 53840 656804 53892 656810
rect 53840 656746 53892 656752
rect 58452 655353 58480 656814
rect 58992 656804 59044 656810
rect 58992 656746 59044 656752
rect 59004 656577 59032 656746
rect 58990 656568 59046 656577
rect 58990 656503 59046 656512
rect 58438 655344 58494 655353
rect 58438 655279 58494 655288
rect 53840 645108 53892 645114
rect 53840 645050 53892 645056
rect 53852 612134 53880 645050
rect 56508 645040 56560 645046
rect 56508 644982 56560 644988
rect 56520 612746 56548 644982
rect 58532 626612 58584 626618
rect 58532 626554 58584 626560
rect 58164 618248 58216 618254
rect 58164 618190 58216 618196
rect 58176 617817 58204 618190
rect 58162 617808 58218 617817
rect 58162 617743 58218 617752
rect 58544 616865 58572 626554
rect 58530 616856 58586 616865
rect 58530 616791 58586 616800
rect 58532 615528 58584 615534
rect 58530 615496 58532 615505
rect 58584 615496 58586 615505
rect 58164 615460 58216 615466
rect 58530 615431 58586 615440
rect 58164 615402 58216 615408
rect 58176 614553 58204 615402
rect 58162 614544 58218 614553
rect 58162 614479 58218 614488
rect 56508 612740 56560 612746
rect 56508 612682 56560 612688
rect 57980 612740 58032 612746
rect 57980 612682 58032 612688
rect 57992 612649 58020 612682
rect 57978 612640 58034 612649
rect 57978 612575 58034 612584
rect 53840 612128 53892 612134
rect 57980 612128 58032 612134
rect 53840 612070 53892 612076
rect 57978 612096 57980 612105
rect 58032 612096 58034 612105
rect 57978 612031 58034 612040
rect 56508 601724 56560 601730
rect 56508 601666 56560 601672
rect 53840 589280 53892 589286
rect 53840 589222 53892 589228
rect 53748 220040 53800 220046
rect 53748 219982 53800 219988
rect 53852 219978 53880 589222
rect 56520 571334 56548 601666
rect 59266 599176 59322 599185
rect 59266 599111 59322 599120
rect 58532 585200 58584 585206
rect 58532 585142 58584 585148
rect 58544 574841 58572 585142
rect 58530 574832 58586 574841
rect 58530 574767 58586 574776
rect 56508 571328 56560 571334
rect 56508 571270 56560 571276
rect 58716 571328 58768 571334
rect 58716 571270 58768 571276
rect 58728 570081 58756 571270
rect 58714 570072 58770 570081
rect 58714 570007 58770 570016
rect 59280 568585 59308 599111
rect 59450 599040 59506 599049
rect 59450 598975 59506 598984
rect 59360 582616 59412 582622
rect 59360 582558 59412 582564
rect 59372 573617 59400 582558
rect 59358 573608 59414 573617
rect 59358 573543 59414 573552
rect 59464 571305 59492 598975
rect 60648 574116 60700 574122
rect 60648 574058 60700 574064
rect 60660 572393 60688 574058
rect 60646 572384 60702 572393
rect 60646 572319 60702 572328
rect 59450 571296 59506 571305
rect 59450 571231 59506 571240
rect 59266 568576 59322 568585
rect 59266 568511 59322 568520
rect 56508 558816 56560 558822
rect 56508 558758 56560 558764
rect 53932 558680 53984 558686
rect 53932 558622 53984 558628
rect 53944 527066 53972 558622
rect 56520 527134 56548 558758
rect 59268 541068 59320 541074
rect 59268 541010 59320 541016
rect 59280 530641 59308 541010
rect 59452 541000 59504 541006
rect 59452 540942 59504 540948
rect 59464 531729 59492 540942
rect 59450 531720 59506 531729
rect 59450 531655 59506 531664
rect 59266 530632 59322 530641
rect 59266 530567 59322 530576
rect 58532 529984 58584 529990
rect 58532 529926 58584 529932
rect 58348 529916 58400 529922
rect 58348 529858 58400 529864
rect 58360 528193 58388 529858
rect 58544 529417 58572 529926
rect 58530 529408 58586 529417
rect 58530 529343 58586 529352
rect 58346 528184 58402 528193
rect 58346 528119 58402 528128
rect 56508 527128 56560 527134
rect 60648 527128 60700 527134
rect 56508 527070 56560 527076
rect 60646 527096 60648 527105
rect 60700 527096 60702 527105
rect 53932 527060 53984 527066
rect 53932 527002 53984 527008
rect 59360 527060 59412 527066
rect 60646 527031 60702 527040
rect 59360 527002 59412 527008
rect 59372 525881 59400 527002
rect 59358 525872 59414 525881
rect 59358 525807 59414 525816
rect 56508 430908 56560 430914
rect 56508 430850 56560 430856
rect 56520 399702 56548 430850
rect 59266 428088 59322 428097
rect 59266 428023 59322 428032
rect 58164 405680 58216 405686
rect 58164 405622 58216 405628
rect 58176 404161 58204 405622
rect 58162 404152 58218 404161
rect 58162 404087 58218 404096
rect 58164 402960 58216 402966
rect 58162 402928 58164 402937
rect 58216 402928 58218 402937
rect 58162 402863 58218 402872
rect 58898 400752 58954 400761
rect 58898 400687 58954 400696
rect 56508 399696 56560 399702
rect 56508 399638 56560 399644
rect 58164 399696 58216 399702
rect 58164 399638 58216 399644
rect 58176 399401 58204 399638
rect 58162 399392 58218 399401
rect 58162 399327 58218 399336
rect 58912 394670 58940 400687
rect 59280 400081 59308 428023
rect 59450 427952 59506 427961
rect 59450 427887 59506 427896
rect 59266 400072 59322 400081
rect 59266 400007 59322 400016
rect 59464 398313 59492 427887
rect 59450 398304 59506 398313
rect 59450 398239 59506 398248
rect 58900 394664 58952 394670
rect 58900 394606 58952 394612
rect 53932 387864 53984 387870
rect 53932 387806 53984 387812
rect 53944 355978 53972 387806
rect 56508 387796 56560 387802
rect 56508 387738 56560 387744
rect 56520 356046 56548 387738
rect 58348 361548 58400 361554
rect 58348 361490 58400 361496
rect 58164 361344 58216 361350
rect 58164 361286 58216 361292
rect 58176 360913 58204 361286
rect 58162 360904 58218 360913
rect 58162 360839 58218 360848
rect 58360 359825 58388 361490
rect 58346 359816 58402 359825
rect 58346 359751 58402 359760
rect 58532 358760 58584 358766
rect 58532 358702 58584 358708
rect 58544 357377 58572 358702
rect 58622 357504 58678 357513
rect 58622 357439 58678 357448
rect 58530 357368 58586 357377
rect 58530 357303 58586 357312
rect 56508 356040 56560 356046
rect 58072 356040 58124 356046
rect 56508 355982 56560 355988
rect 58070 356008 58072 356017
rect 58124 356008 58126 356017
rect 53932 355972 53984 355978
rect 58070 355943 58126 355952
rect 53932 355914 53984 355920
rect 58636 350538 58664 357439
rect 59360 355972 59412 355978
rect 59360 355914 59412 355920
rect 59372 355065 59400 355914
rect 59358 355056 59414 355065
rect 59358 354991 59414 355000
rect 58624 350532 58676 350538
rect 58624 350474 58676 350480
rect 58440 318776 58492 318782
rect 58440 318718 58492 318724
rect 58164 317416 58216 317422
rect 58452 317393 58480 318718
rect 58164 317358 58216 317364
rect 58438 317384 58494 317393
rect 58176 316577 58204 317358
rect 58438 317319 58494 317328
rect 58162 316568 58218 316577
rect 58162 316503 58218 316512
rect 58346 314800 58402 314809
rect 58346 314735 58402 314744
rect 58164 314560 58216 314566
rect 58164 314502 58216 314508
rect 58176 313041 58204 314502
rect 58162 313032 58218 313041
rect 58162 312967 58218 312976
rect 58360 306338 58388 314735
rect 58532 314628 58584 314634
rect 58532 314570 58584 314576
rect 58544 314129 58572 314570
rect 58530 314120 58586 314129
rect 58530 314055 58586 314064
rect 58532 311840 58584 311846
rect 58530 311808 58532 311817
rect 58584 311808 58586 311817
rect 58530 311743 58586 311752
rect 58348 306332 58400 306338
rect 58348 306274 58400 306280
rect 54024 301436 54076 301442
rect 54024 301378 54076 301384
rect 54036 289814 54064 301378
rect 57888 301368 57940 301374
rect 57888 301310 57940 301316
rect 57900 291553 57928 301310
rect 58438 298208 58494 298217
rect 58438 298143 58494 298152
rect 58346 293992 58402 294001
rect 58346 293927 58402 293936
rect 58360 292602 58388 293927
rect 58348 292596 58400 292602
rect 58348 292538 58400 292544
rect 58452 292505 58480 298143
rect 58530 295488 58586 295497
rect 58530 295423 58586 295432
rect 58544 295390 58572 295423
rect 58532 295384 58584 295390
rect 58532 295326 58584 295332
rect 59450 292768 59506 292777
rect 59450 292703 59506 292712
rect 58438 292496 58494 292505
rect 58438 292431 58494 292440
rect 57886 291544 57942 291553
rect 57886 291479 57942 291488
rect 54024 289808 54076 289814
rect 58532 289808 58584 289814
rect 54024 289750 54076 289756
rect 58530 289776 58532 289785
rect 58584 289776 58586 289785
rect 58530 289711 58586 289720
rect 57978 288008 58034 288017
rect 57978 287943 58034 287952
rect 57992 287162 58020 287943
rect 58530 287192 58586 287201
rect 56508 287156 56560 287162
rect 56508 287098 56560 287104
rect 57980 287156 58032 287162
rect 58530 287127 58586 287136
rect 57980 287098 58032 287104
rect 53932 285184 53984 285190
rect 53932 285126 53984 285132
rect 53944 258126 53972 285126
rect 53932 258120 53984 258126
rect 53932 258062 53984 258068
rect 56046 227624 56102 227633
rect 56046 227559 56102 227568
rect 55128 224936 55180 224942
rect 55128 224878 55180 224884
rect 54390 222184 54446 222193
rect 54390 222119 54446 222128
rect 53840 219972 53892 219978
rect 53840 219914 53892 219920
rect 54404 217410 54432 222119
rect 55140 217410 55168 224878
rect 56060 217410 56088 227559
rect 56520 220794 56548 287098
rect 58544 287094 58572 287127
rect 58532 287088 58584 287094
rect 58532 287030 58584 287036
rect 57978 285696 58034 285705
rect 57978 285631 58034 285640
rect 57992 285190 58020 285631
rect 57980 285184 58032 285190
rect 57980 285126 58032 285132
rect 58530 284472 58586 284481
rect 58530 284407 58586 284416
rect 58544 284374 58572 284407
rect 58532 284368 58584 284374
rect 58532 284310 58584 284316
rect 57978 283248 58034 283257
rect 57978 283183 58034 283192
rect 57992 281586 58020 283183
rect 59266 282160 59322 282169
rect 59266 282095 59322 282104
rect 57980 281580 58032 281586
rect 57980 281522 58032 281528
rect 56692 245744 56744 245750
rect 56692 245686 56744 245692
rect 56600 245676 56652 245682
rect 56600 245618 56652 245624
rect 56508 220788 56560 220794
rect 56508 220730 56560 220736
rect 56612 219910 56640 245618
rect 56600 219904 56652 219910
rect 56600 219846 56652 219852
rect 56704 219842 56732 245686
rect 57610 227760 57666 227769
rect 57610 227695 57666 227704
rect 56874 224904 56930 224913
rect 56874 224839 56930 224848
rect 56692 219836 56744 219842
rect 56692 219778 56744 219784
rect 56888 217410 56916 224839
rect 57624 217410 57652 227695
rect 58622 225040 58678 225049
rect 58622 224975 58678 224984
rect 58636 217410 58664 224975
rect 59174 222320 59230 222329
rect 59174 222255 59230 222264
rect 59188 217410 59216 222255
rect 52440 217382 52776 217410
rect 53268 217382 53604 217410
rect 54096 217382 54432 217410
rect 54924 217382 55168 217410
rect 55752 217382 56088 217410
rect 56580 217382 56916 217410
rect 57408 217382 57652 217410
rect 58328 217382 58664 217410
rect 59156 217382 59216 217410
rect 59280 216646 59308 282095
rect 59358 279712 59414 279721
rect 59358 279647 59414 279656
rect 59372 216714 59400 279647
rect 59464 264790 59492 292703
rect 61842 291136 61898 291145
rect 61842 291071 61898 291080
rect 59542 280936 59598 280945
rect 59542 280871 59598 280880
rect 59452 264784 59504 264790
rect 59452 264726 59504 264732
rect 59556 222222 59584 280871
rect 60280 225004 60332 225010
rect 60280 224946 60332 224952
rect 59544 222216 59596 222222
rect 59544 222158 59596 222164
rect 60292 217410 60320 224946
rect 61106 222456 61162 222465
rect 61106 222391 61162 222400
rect 61120 217410 61148 222391
rect 61856 217870 61884 291071
rect 61936 222216 61988 222222
rect 61936 222158 61988 222164
rect 61844 217864 61896 217870
rect 61844 217806 61896 217812
rect 61948 217410 61976 222158
rect 62132 221490 62160 805938
rect 655520 792192 655572 792198
rect 655520 792134 655572 792140
rect 655426 778424 655482 778433
rect 655426 778359 655482 778368
rect 654968 775532 655020 775538
rect 654968 775474 655020 775480
rect 654980 773537 655008 775474
rect 654966 773528 655022 773537
rect 654966 773463 655022 773472
rect 655152 737044 655204 737050
rect 655152 736986 655204 736992
rect 655164 730289 655192 736986
rect 655150 730280 655206 730289
rect 655150 730215 655206 730224
rect 655440 715018 655468 778359
rect 655532 775577 655560 792134
rect 656532 783896 656584 783902
rect 656532 783838 656584 783844
rect 655610 777064 655666 777073
rect 655610 776999 655666 777008
rect 655518 775568 655574 775577
rect 655518 775503 655574 775512
rect 655518 731504 655574 731513
rect 655518 731439 655574 731448
rect 655428 715012 655480 715018
rect 655428 714954 655480 714960
rect 654232 692912 654284 692918
rect 654232 692854 654284 692860
rect 654140 690056 654192 690062
rect 654140 689998 654192 690004
rect 654152 684457 654180 689998
rect 654244 685817 654272 692854
rect 655426 687304 655482 687313
rect 655426 687239 655482 687248
rect 654230 685808 654286 685817
rect 654230 685743 654286 685752
rect 654138 684448 654194 684457
rect 654138 684383 654194 684392
rect 654416 648644 654468 648650
rect 654416 648586 654468 648592
rect 654428 639441 654456 648586
rect 654414 639432 654470 639441
rect 654414 639367 654470 639376
rect 655440 623898 655468 687239
rect 655532 668098 655560 731439
rect 655624 715154 655652 776999
rect 655794 775976 655850 775985
rect 655794 775911 655850 775920
rect 655702 734360 655758 734369
rect 655702 734295 655758 734304
rect 655612 715148 655664 715154
rect 655612 715090 655664 715096
rect 655610 689480 655666 689489
rect 655610 689415 655666 689424
rect 655520 668092 655572 668098
rect 655520 668034 655572 668040
rect 655518 643240 655574 643249
rect 655518 643175 655574 643184
rect 655428 623892 655480 623898
rect 655428 623834 655480 623840
rect 655428 612876 655480 612882
rect 655428 612818 655480 612824
rect 655440 595377 655468 612818
rect 655426 595368 655482 595377
rect 655426 595303 655482 595312
rect 655532 579834 655560 643175
rect 655624 624034 655652 689415
rect 655716 670818 655744 734295
rect 655808 715290 655836 775911
rect 656544 774761 656572 783838
rect 656530 774752 656586 774761
rect 656530 774687 656586 774696
rect 655980 747992 656032 747998
rect 655980 747934 656032 747940
rect 655886 732728 655942 732737
rect 655886 732663 655942 732672
rect 655796 715284 655848 715290
rect 655796 715226 655848 715232
rect 655794 688256 655850 688265
rect 655794 688191 655850 688200
rect 655704 670812 655756 670818
rect 655704 670754 655756 670760
rect 655704 656940 655756 656946
rect 655704 656882 655756 656888
rect 655716 640257 655744 656882
rect 655702 640248 655758 640257
rect 655702 640183 655758 640192
rect 655808 624170 655836 688191
rect 655900 670954 655928 732663
rect 655992 731377 656020 747934
rect 656072 736976 656124 736982
rect 656072 736918 656124 736924
rect 655978 731368 656034 731377
rect 655978 731303 656034 731312
rect 656084 728657 656112 736918
rect 656070 728648 656126 728657
rect 656070 728583 656126 728592
rect 670436 713454 670464 892978
rect 670528 715426 670556 894406
rect 670608 893852 670660 893858
rect 670608 893794 670660 893800
rect 670516 715420 670568 715426
rect 670516 715362 670568 715368
rect 670516 714876 670568 714882
rect 670516 714818 670568 714824
rect 669872 713448 669924 713454
rect 669872 713390 669924 713396
rect 670424 713448 670476 713454
rect 670424 713390 670476 713396
rect 669884 712366 669912 713390
rect 669872 712360 669924 712366
rect 669872 712302 669924 712308
rect 670332 712292 670384 712298
rect 670332 712234 670384 712240
rect 655980 703860 656032 703866
rect 655980 703802 656032 703808
rect 655992 687041 656020 703802
rect 655978 687032 656034 687041
rect 655978 686967 656034 686976
rect 655888 670948 655940 670954
rect 655888 670890 655940 670896
rect 669596 669316 669648 669322
rect 669596 669258 669648 669264
rect 669608 668234 669636 669258
rect 669596 668228 669648 668234
rect 669596 668170 669648 668176
rect 670240 665304 670292 665310
rect 670240 665246 670292 665252
rect 656440 645924 656492 645930
rect 656440 645866 656492 645872
rect 655978 641880 656034 641889
rect 655978 641815 656034 641824
rect 655796 624164 655848 624170
rect 655796 624106 655848 624112
rect 655612 624028 655664 624034
rect 655612 623970 655664 623976
rect 655612 601724 655664 601730
rect 655612 601666 655664 601672
rect 655624 593065 655652 601666
rect 655886 597816 655942 597825
rect 655886 597751 655942 597760
rect 655702 596592 655758 596601
rect 655702 596527 655758 596536
rect 655610 593056 655666 593065
rect 655610 592991 655666 593000
rect 655520 579828 655572 579834
rect 655520 579770 655572 579776
rect 654232 557592 654284 557598
rect 654232 557534 654284 557540
rect 654140 554804 654192 554810
rect 654140 554746 654192 554752
rect 654152 548593 654180 554746
rect 654244 549273 654272 557534
rect 655610 553344 655666 553353
rect 655610 553279 655666 553288
rect 655426 552120 655482 552129
rect 655426 552055 655482 552064
rect 654230 549264 654286 549273
rect 654230 549199 654286 549208
rect 654138 548584 654194 548593
rect 654138 548519 654194 548528
rect 655440 491434 655468 552055
rect 655518 551032 655574 551041
rect 655518 550967 655574 550976
rect 655532 491570 655560 550967
rect 655624 491706 655652 553279
rect 655716 535634 655744 596527
rect 655794 595504 655850 595513
rect 655794 595439 655850 595448
rect 655704 535628 655756 535634
rect 655704 535570 655756 535576
rect 655808 532914 655836 595439
rect 655900 535770 655928 597751
rect 655992 579970 656020 641815
rect 656162 640656 656218 640665
rect 656162 640591 656218 640600
rect 656176 580106 656204 640591
rect 656452 638217 656480 645866
rect 656438 638208 656494 638217
rect 656438 638143 656494 638152
rect 670252 621042 670280 665246
rect 670344 665242 670372 712234
rect 670424 712224 670476 712230
rect 670424 712166 670476 712172
rect 670436 668166 670464 712166
rect 670528 669322 670556 714818
rect 670620 712434 670648 893794
rect 671988 883244 672040 883250
rect 671988 883186 672040 883192
rect 670608 712428 670660 712434
rect 670608 712370 670660 712376
rect 670516 669316 670568 669322
rect 670516 669258 670568 669264
rect 670424 668160 670476 668166
rect 670424 668102 670476 668108
rect 670608 668024 670660 668030
rect 670608 667966 670660 667972
rect 670332 665236 670384 665242
rect 670332 665178 670384 665184
rect 670620 624102 670648 667966
rect 670608 624096 670660 624102
rect 670608 624038 670660 624044
rect 670516 623960 670568 623966
rect 670516 623902 670568 623908
rect 670424 621104 670476 621110
rect 670424 621046 670476 621052
rect 670240 621036 670292 621042
rect 670240 620978 670292 620984
rect 656808 601792 656860 601798
rect 656808 601734 656860 601740
rect 656820 594289 656848 601734
rect 656806 594280 656862 594289
rect 656806 594215 656862 594224
rect 656164 580100 656216 580106
rect 656164 580042 656216 580048
rect 655980 579964 656032 579970
rect 655980 579906 656032 579912
rect 670436 576978 670464 621046
rect 670528 579698 670556 623902
rect 670608 621172 670660 621178
rect 670608 621114 670660 621120
rect 670516 579692 670568 579698
rect 670516 579634 670568 579640
rect 670424 576972 670476 576978
rect 670424 576914 670476 576920
rect 670620 576910 670648 621114
rect 670608 576904 670660 576910
rect 670608 576846 670660 576852
rect 655980 568676 656032 568682
rect 655980 568618 656032 568624
rect 655992 550905 656020 568618
rect 655978 550896 656034 550905
rect 655978 550831 656034 550840
rect 655888 535764 655940 535770
rect 655888 535706 655940 535712
rect 655796 532908 655848 532914
rect 655796 532850 655848 532856
rect 655612 491700 655664 491706
rect 655612 491642 655664 491648
rect 655520 491564 655572 491570
rect 655520 491506 655572 491512
rect 655428 491428 655480 491434
rect 655428 491370 655480 491376
rect 655704 403164 655756 403170
rect 655704 403106 655756 403112
rect 655520 403096 655572 403102
rect 655520 403038 655572 403044
rect 655428 403028 655480 403034
rect 655428 402970 655480 402976
rect 654508 372564 654560 372570
rect 654508 372506 654560 372512
rect 654520 370977 654548 372506
rect 655440 372201 655468 402970
rect 655532 373289 655560 403038
rect 655716 374513 655744 403106
rect 655702 374504 655758 374513
rect 655702 374439 655758 374448
rect 655518 373280 655574 373289
rect 655518 373215 655574 373224
rect 655426 372192 655482 372201
rect 655426 372127 655482 372136
rect 654506 370968 654562 370977
rect 654506 370903 654562 370912
rect 655520 356516 655572 356522
rect 655520 356458 655572 356464
rect 655428 356380 655480 356386
rect 655428 356322 655480 356328
rect 655440 327457 655468 356322
rect 655532 329905 655560 356458
rect 655612 356244 655664 356250
rect 655612 356186 655664 356192
rect 655518 329896 655574 329905
rect 655518 329831 655574 329840
rect 655624 328273 655652 356186
rect 655980 335368 656032 335374
rect 655980 335310 656032 335316
rect 655610 328264 655666 328273
rect 655610 328199 655666 328208
rect 655426 327448 655482 327457
rect 655426 327383 655482 327392
rect 655992 325689 656020 335310
rect 655978 325680 656034 325689
rect 655978 325615 656034 325624
rect 655428 312180 655480 312186
rect 655428 312122 655480 312128
rect 655440 300801 655468 312122
rect 655704 312044 655756 312050
rect 655704 311986 655756 311992
rect 655520 311976 655572 311982
rect 655520 311918 655572 311924
rect 655532 303385 655560 311918
rect 655518 303376 655574 303385
rect 655518 303311 655574 303320
rect 655716 302161 655744 311986
rect 671620 311908 671672 311914
rect 671620 311850 671672 311856
rect 655702 302152 655758 302161
rect 655702 302087 655758 302096
rect 655426 300792 655482 300801
rect 655426 300727 655482 300736
rect 655058 298752 655114 298761
rect 655058 298687 655114 298696
rect 655072 298178 655100 298687
rect 655060 298172 655112 298178
rect 655060 298114 655112 298120
rect 656162 297528 656218 297537
rect 656162 297463 656218 297472
rect 655794 296304 655850 296313
rect 655794 296239 655850 296248
rect 655610 293992 655666 294001
rect 655610 293927 655666 293936
rect 655426 292768 655482 292777
rect 655426 292703 655482 292712
rect 654138 289232 654194 289241
rect 654138 289167 654194 289176
rect 654152 289134 654180 289167
rect 654140 289128 654192 289134
rect 654140 289070 654192 289076
rect 654138 288008 654194 288017
rect 654138 287943 654194 287952
rect 654152 287094 654180 287943
rect 654140 287088 654192 287094
rect 654140 287030 654192 287036
rect 655242 285696 655298 285705
rect 655242 285631 655298 285640
rect 655256 284986 655284 285631
rect 655244 284980 655296 284986
rect 655244 284922 655296 284928
rect 654506 284744 654562 284753
rect 654506 284679 654508 284688
rect 654560 284679 654562 284688
rect 654508 284650 654560 284656
rect 654230 283656 654286 283665
rect 654230 283591 654286 283600
rect 654244 283218 654272 283591
rect 654232 283212 654284 283218
rect 654232 283154 654284 283160
rect 655242 282160 655298 282169
rect 655242 282095 655298 282104
rect 655256 281586 655284 282095
rect 655244 281580 655296 281586
rect 655244 281522 655296 281528
rect 654138 280936 654194 280945
rect 654138 280871 654194 280880
rect 654152 280430 654180 280871
rect 654140 280424 654192 280430
rect 654140 280366 654192 280372
rect 654874 279712 654930 279721
rect 654874 279647 654930 279656
rect 654888 278798 654916 279647
rect 654876 278792 654928 278798
rect 654876 278734 654928 278740
rect 63406 276040 63462 276049
rect 63406 275975 63462 275984
rect 62670 227896 62726 227905
rect 62670 227831 62726 227840
rect 59984 217382 60320 217410
rect 60812 217382 61148 217410
rect 61640 217382 61976 217410
rect 62040 221462 62160 221490
rect 62040 216782 62068 221462
rect 62684 217410 62712 227831
rect 63314 225176 63370 225185
rect 63314 225111 63370 225120
rect 62948 217864 63000 217870
rect 62948 217806 63000 217812
rect 62468 217382 62712 217410
rect 62028 216776 62080 216782
rect 62028 216718 62080 216724
rect 62960 216714 62988 217806
rect 63328 217410 63356 225111
rect 63296 217382 63356 217410
rect 63420 217297 63448 275975
rect 65904 271862 65932 278052
rect 65892 271856 65944 271862
rect 65892 271798 65944 271804
rect 67100 269142 67128 278052
rect 67088 269136 67140 269142
rect 67088 269078 67140 269084
rect 68204 266354 68232 278052
rect 69400 271833 69428 278052
rect 70596 271969 70624 278052
rect 70582 271960 70638 271969
rect 70582 271895 70638 271904
rect 69386 271824 69442 271833
rect 69386 271759 69442 271768
rect 71792 269113 71820 278052
rect 72988 269278 73016 278052
rect 72976 269272 73028 269278
rect 72976 269214 73028 269220
rect 71778 269104 71834 269113
rect 71778 269039 71834 269048
rect 74184 267918 74212 278052
rect 75380 269346 75408 278052
rect 75368 269340 75420 269346
rect 75368 269282 75420 269288
rect 76484 269249 76512 278052
rect 77680 269385 77708 278052
rect 78876 269521 78904 278052
rect 80072 272377 80100 278052
rect 80058 272368 80114 272377
rect 80058 272303 80114 272312
rect 81268 272105 81296 278052
rect 81254 272096 81310 272105
rect 81254 272031 81310 272040
rect 82464 271930 82492 278052
rect 83660 272241 83688 278052
rect 83646 272232 83702 272241
rect 83646 272167 83702 272176
rect 82452 271924 82504 271930
rect 82452 271866 82504 271872
rect 84764 269657 84792 278052
rect 85960 269793 85988 278052
rect 85946 269784 86002 269793
rect 85946 269719 86002 269728
rect 84750 269648 84806 269657
rect 84750 269583 84806 269592
rect 78862 269512 78918 269521
rect 78862 269447 78918 269456
rect 87156 269414 87184 278052
rect 88352 272649 88380 278052
rect 88338 272640 88394 272649
rect 88338 272575 88394 272584
rect 89548 271998 89576 278052
rect 90744 272513 90772 278052
rect 90730 272504 90786 272513
rect 90730 272439 90786 272448
rect 91848 272066 91876 278052
rect 91836 272060 91888 272066
rect 91836 272002 91888 272008
rect 89536 271992 89588 271998
rect 89536 271934 89588 271940
rect 93044 269929 93072 278052
rect 93030 269920 93086 269929
rect 93030 269855 93086 269864
rect 94240 269550 94268 278052
rect 94228 269544 94280 269550
rect 94228 269486 94280 269492
rect 95436 269482 95464 278052
rect 96632 272921 96660 278052
rect 96618 272912 96674 272921
rect 96618 272847 96674 272856
rect 97828 272134 97856 278052
rect 99024 272785 99052 278052
rect 99010 272776 99066 272785
rect 99010 272711 99066 272720
rect 97816 272128 97868 272134
rect 97816 272070 97868 272076
rect 100128 270065 100156 278052
rect 101324 270201 101352 278052
rect 101310 270192 101366 270201
rect 101310 270127 101366 270136
rect 100114 270056 100170 270065
rect 100114 269991 100170 270000
rect 102520 269618 102548 278052
rect 103716 273057 103744 278052
rect 103702 273048 103758 273057
rect 103702 272983 103758 272992
rect 104912 272202 104940 278052
rect 106108 273193 106136 278052
rect 106094 273184 106150 273193
rect 106094 273119 106150 273128
rect 104900 272196 104952 272202
rect 104900 272138 104952 272144
rect 107212 270337 107240 278052
rect 107198 270328 107254 270337
rect 107198 270263 107254 270272
rect 108408 269686 108436 278052
rect 109604 269754 109632 278052
rect 110800 271425 110828 278052
rect 111996 271697 112024 278052
rect 111982 271688 112038 271697
rect 111982 271623 112038 271632
rect 110786 271416 110842 271425
rect 110786 271351 110842 271360
rect 113192 269822 113220 278052
rect 114388 269890 114416 278052
rect 115492 271561 115520 278052
rect 115478 271552 115534 271561
rect 115478 271487 115534 271496
rect 114376 269884 114428 269890
rect 114376 269826 114428 269832
rect 113180 269816 113232 269822
rect 113180 269758 113232 269764
rect 109592 269748 109644 269754
rect 109592 269690 109644 269696
rect 108396 269680 108448 269686
rect 108396 269622 108448 269628
rect 102508 269612 102560 269618
rect 102508 269554 102560 269560
rect 95424 269476 95476 269482
rect 95424 269418 95476 269424
rect 87144 269408 87196 269414
rect 77666 269376 77722 269385
rect 87144 269350 87196 269356
rect 77666 269311 77722 269320
rect 76470 269240 76526 269249
rect 76470 269175 76526 269184
rect 74172 267912 74224 267918
rect 74172 267854 74224 267860
rect 116688 266422 116716 278052
rect 117884 271289 117912 278052
rect 117870 271280 117926 271289
rect 117870 271215 117926 271224
rect 119080 269958 119108 278052
rect 120276 270473 120304 278052
rect 120262 270464 120318 270473
rect 120262 270399 120318 270408
rect 121472 270026 121500 278052
rect 122576 271153 122604 278052
rect 123772 272270 123800 278052
rect 124968 272338 124996 278052
rect 124956 272332 125008 272338
rect 124956 272274 125008 272280
rect 123760 272264 123812 272270
rect 123760 272206 123812 272212
rect 122562 271144 122618 271153
rect 122562 271079 122618 271088
rect 126164 270162 126192 278052
rect 126152 270156 126204 270162
rect 126152 270098 126204 270104
rect 127360 270094 127388 278052
rect 127348 270088 127400 270094
rect 127348 270030 127400 270036
rect 121460 270020 121512 270026
rect 121460 269962 121512 269968
rect 119068 269952 119120 269958
rect 119068 269894 119120 269900
rect 128556 268977 128584 278052
rect 129660 272406 129688 278052
rect 130856 272542 130884 278052
rect 130844 272536 130896 272542
rect 130844 272478 130896 272484
rect 132052 272474 132080 278052
rect 132040 272468 132092 272474
rect 132040 272410 132092 272416
rect 129648 272400 129700 272406
rect 129648 272342 129700 272348
rect 133248 270570 133276 278052
rect 134444 271454 134472 278052
rect 134432 271448 134484 271454
rect 134432 271390 134484 271396
rect 133236 270564 133288 270570
rect 133236 270506 133288 270512
rect 135640 270230 135668 278052
rect 136836 272610 136864 278052
rect 137940 272678 137968 278052
rect 139136 272746 139164 278052
rect 139124 272740 139176 272746
rect 139124 272682 139176 272688
rect 137928 272672 137980 272678
rect 137928 272614 137980 272620
rect 136824 272604 136876 272610
rect 136824 272546 136876 272552
rect 140332 270366 140360 278052
rect 141528 270434 141556 278052
rect 142724 270842 142752 278052
rect 143920 273018 143948 278052
rect 143908 273012 143960 273018
rect 143908 272954 143960 272960
rect 145116 272882 145144 278052
rect 145104 272876 145156 272882
rect 145104 272818 145156 272824
rect 146220 272814 146248 278052
rect 146208 272808 146260 272814
rect 146208 272750 146260 272756
rect 142712 270836 142764 270842
rect 142712 270778 142764 270784
rect 146208 270836 146260 270842
rect 146208 270778 146260 270784
rect 141516 270428 141568 270434
rect 141516 270370 141568 270376
rect 140320 270360 140372 270366
rect 140320 270302 140372 270308
rect 135628 270224 135680 270230
rect 135628 270166 135680 270172
rect 128542 268968 128598 268977
rect 128542 268903 128598 268912
rect 146220 268841 146248 270778
rect 147416 270502 147444 278052
rect 148612 272950 148640 278052
rect 149808 273086 149836 278052
rect 149796 273080 149848 273086
rect 149796 273022 149848 273028
rect 148600 272944 148652 272950
rect 148600 272886 148652 272892
rect 147404 270496 147456 270502
rect 147404 270438 147456 270444
rect 146206 268832 146262 268841
rect 146206 268767 146262 268776
rect 151004 268705 151032 278052
rect 152200 269006 152228 278052
rect 153396 269074 153424 278052
rect 154500 273222 154528 278052
rect 154488 273216 154540 273222
rect 154488 273158 154540 273164
rect 155696 271794 155724 278052
rect 156892 273154 156920 278052
rect 156880 273148 156932 273154
rect 156880 273090 156932 273096
rect 155684 271788 155736 271794
rect 155684 271730 155736 271736
rect 153384 269068 153436 269074
rect 153384 269010 153436 269016
rect 152188 269000 152240 269006
rect 152188 268942 152240 268948
rect 150990 268696 151046 268705
rect 150990 268631 151046 268640
rect 158088 268569 158116 278052
rect 158074 268560 158130 268569
rect 158074 268495 158130 268504
rect 159284 268433 159312 278052
rect 160480 268870 160508 278052
rect 161584 271726 161612 278052
rect 161572 271720 161624 271726
rect 161572 271662 161624 271668
rect 162780 271590 162808 278052
rect 163976 271658 164004 278052
rect 163964 271652 164016 271658
rect 163964 271594 164016 271600
rect 162768 271584 162820 271590
rect 162768 271526 162820 271532
rect 165172 268938 165200 278052
rect 165160 268932 165212 268938
rect 165160 268874 165212 268880
rect 160468 268864 160520 268870
rect 160468 268806 160520 268812
rect 166368 268734 166396 278052
rect 167564 268802 167592 278052
rect 168760 271386 168788 278052
rect 168748 271380 168800 271386
rect 168748 271322 168800 271328
rect 169864 271318 169892 278052
rect 171060 271522 171088 278052
rect 171048 271516 171100 271522
rect 171048 271458 171100 271464
rect 169852 271312 169904 271318
rect 169852 271254 169904 271260
rect 167552 268796 167604 268802
rect 167552 268738 167604 268744
rect 166356 268728 166408 268734
rect 166356 268670 166408 268676
rect 172256 268666 172284 278052
rect 172244 268660 172296 268666
rect 172244 268602 172296 268608
rect 173452 268598 173480 278052
rect 173440 268592 173492 268598
rect 173440 268534 173492 268540
rect 174648 268530 174676 278052
rect 175844 271114 175872 278052
rect 176844 271856 176896 271862
rect 176844 271798 176896 271804
rect 176856 271250 176884 271798
rect 176844 271244 176896 271250
rect 176844 271186 176896 271192
rect 175832 271108 175884 271114
rect 175832 271050 175884 271056
rect 176948 270774 176976 278052
rect 178144 271182 178172 278052
rect 178132 271176 178184 271182
rect 178132 271118 178184 271124
rect 176936 270768 176988 270774
rect 176936 270710 176988 270716
rect 174636 268524 174688 268530
rect 174636 268466 174688 268472
rect 179340 268462 179368 278052
rect 179328 268456 179380 268462
rect 159270 268424 159326 268433
rect 179328 268398 179380 268404
rect 159270 268359 159326 268368
rect 180536 268326 180564 278052
rect 181732 268394 181760 278052
rect 182928 271046 182956 278052
rect 182916 271040 182968 271046
rect 182916 270982 182968 270988
rect 181720 268388 181772 268394
rect 181720 268330 181772 268336
rect 180524 268320 180576 268326
rect 180524 268262 180576 268268
rect 184124 268258 184152 278052
rect 184112 268252 184164 268258
rect 184112 268194 184164 268200
rect 185228 268190 185256 278052
rect 186424 270910 186452 278052
rect 187620 270978 187648 278052
rect 187608 270972 187660 270978
rect 187608 270914 187660 270920
rect 186412 270904 186464 270910
rect 186412 270846 186464 270852
rect 188816 270842 188844 278052
rect 188804 270836 188856 270842
rect 188804 270778 188856 270784
rect 185216 268184 185268 268190
rect 185216 268126 185268 268132
rect 190012 268122 190040 278052
rect 191208 270570 191236 278052
rect 192116 271244 192168 271250
rect 192116 271186 192168 271192
rect 191196 270564 191248 270570
rect 191196 270506 191248 270512
rect 190000 268116 190052 268122
rect 190000 268058 190052 268064
rect 116676 266416 116728 266422
rect 116676 266358 116728 266364
rect 68192 266348 68244 266354
rect 68192 266290 68244 266296
rect 192128 264330 192156 271186
rect 192404 268054 192432 278052
rect 193508 269142 193536 278052
rect 194138 271960 194194 271969
rect 194138 271895 194194 271904
rect 193678 271824 193734 271833
rect 193678 271759 193734 271768
rect 192760 269136 192812 269142
rect 192760 269078 192812 269084
rect 193496 269136 193548 269142
rect 193496 269078 193548 269084
rect 192392 268048 192444 268054
rect 192392 267990 192444 267996
rect 192128 264302 192418 264330
rect 192772 264316 192800 269078
rect 193220 266348 193272 266354
rect 193220 266290 193272 266296
rect 193232 264316 193260 266290
rect 193692 264316 193720 271759
rect 194152 264316 194180 271895
rect 194704 271862 194732 278052
rect 194692 271856 194744 271862
rect 194692 271798 194744 271804
rect 195796 271448 195848 271454
rect 195796 271390 195848 271396
rect 195428 269340 195480 269346
rect 195428 269282 195480 269288
rect 195060 269272 195112 269278
rect 195060 269214 195112 269220
rect 194598 269104 194654 269113
rect 194598 269039 194654 269048
rect 194612 264316 194640 269039
rect 195072 264316 195100 269214
rect 195440 264316 195468 269282
rect 195808 267986 195836 271390
rect 195900 269210 195928 278052
rect 196898 272368 196954 272377
rect 196898 272303 196954 272312
rect 195980 272060 196032 272066
rect 195980 272002 196032 272008
rect 195888 269204 195940 269210
rect 195888 269146 195940 269152
rect 195992 268297 196020 272002
rect 196806 269376 196862 269385
rect 196806 269311 196862 269320
rect 196346 269240 196402 269249
rect 196346 269175 196402 269184
rect 195978 268288 196034 268297
rect 195978 268223 196034 268232
rect 195796 267980 195848 267986
rect 195796 267922 195848 267928
rect 195888 267912 195940 267918
rect 195888 267854 195940 267860
rect 195900 264316 195928 267854
rect 196360 264316 196388 269175
rect 196820 264316 196848 269311
rect 196912 264330 196940 272303
rect 197096 271454 197124 278052
rect 198094 272096 198150 272105
rect 198094 272031 198150 272040
rect 197084 271448 197136 271454
rect 197084 271390 197136 271396
rect 197188 271250 197400 271266
rect 197188 271244 197412 271250
rect 197188 271238 197360 271244
rect 197188 271114 197216 271238
rect 197360 271186 197412 271192
rect 197176 271108 197228 271114
rect 197176 271050 197228 271056
rect 197268 271108 197320 271114
rect 197268 271050 197320 271056
rect 197280 270774 197308 271050
rect 197268 270768 197320 270774
rect 197268 270710 197320 270716
rect 197726 269512 197782 269521
rect 197726 269447 197782 269456
rect 196912 264302 197294 264330
rect 197740 264316 197768 269447
rect 198108 264316 198136 272031
rect 198292 270638 198320 278052
rect 199488 276014 199516 278052
rect 199488 275986 199608 276014
rect 199106 272232 199162 272241
rect 199106 272167 199162 272176
rect 198556 271924 198608 271930
rect 198556 271866 198608 271872
rect 198280 270632 198332 270638
rect 198280 270574 198332 270580
rect 198568 264316 198596 271866
rect 199014 269648 199070 269657
rect 199014 269583 199070 269592
rect 199028 264316 199056 269583
rect 199120 264330 199148 272167
rect 199580 270706 199608 275986
rect 199568 270700 199620 270706
rect 199568 270642 199620 270648
rect 199934 269784 199990 269793
rect 199934 269719 199990 269728
rect 199120 264302 199502 264330
rect 199948 264316 199976 269719
rect 200396 269408 200448 269414
rect 200396 269350 200448 269356
rect 200408 264316 200436 269350
rect 200592 269278 200620 278052
rect 201222 272640 201278 272649
rect 201222 272575 201278 272584
rect 200764 271992 200816 271998
rect 200764 271934 200816 271940
rect 200580 269272 200632 269278
rect 200580 269214 200632 269220
rect 200776 264316 200804 271934
rect 201236 264316 201264 272575
rect 201682 272504 201738 272513
rect 201682 272439 201738 272448
rect 201696 264316 201724 272439
rect 201788 272066 201816 278052
rect 201776 272060 201828 272066
rect 201776 272002 201828 272008
rect 202604 269544 202656 269550
rect 202604 269486 202656 269492
rect 202142 268288 202198 268297
rect 202142 268223 202198 268232
rect 202156 264316 202184 268223
rect 202616 264316 202644 269486
rect 202984 269414 203012 278052
rect 203892 272128 203944 272134
rect 203892 272070 203944 272076
rect 203062 269920 203118 269929
rect 203062 269855 203118 269864
rect 202972 269408 203024 269414
rect 202972 269350 203024 269356
rect 203076 264316 203104 269855
rect 203524 269476 203576 269482
rect 203524 269418 203576 269424
rect 203536 264316 203564 269418
rect 203904 264316 203932 272070
rect 204180 269346 204208 278052
rect 204350 272912 204406 272921
rect 204350 272847 204406 272856
rect 204168 269340 204220 269346
rect 204168 269282 204220 269288
rect 204364 264316 204392 272847
rect 204810 272776 204866 272785
rect 204810 272711 204866 272720
rect 204824 264316 204852 272711
rect 205376 272134 205404 278052
rect 206284 272196 206336 272202
rect 206284 272138 206336 272144
rect 205364 272128 205416 272134
rect 205364 272070 205416 272076
rect 205270 270192 205326 270201
rect 205270 270127 205326 270136
rect 205284 264316 205312 270127
rect 205730 270056 205786 270065
rect 205730 269991 205786 270000
rect 205744 264316 205772 269991
rect 206192 269612 206244 269618
rect 206192 269554 206244 269560
rect 206204 264316 206232 269554
rect 206296 264330 206324 272138
rect 206572 269482 206600 278052
rect 207782 278038 208072 278066
rect 208886 278038 209176 278066
rect 207478 273184 207534 273193
rect 207478 273119 207534 273128
rect 207018 273048 207074 273057
rect 207018 272983 207074 272992
rect 206560 269476 206612 269482
rect 206560 269418 206612 269424
rect 206296 264302 206586 264330
rect 207032 264316 207060 272983
rect 207492 264316 207520 273119
rect 207848 270292 207900 270298
rect 207848 270234 207900 270240
rect 207940 270292 207992 270298
rect 207940 270234 207992 270240
rect 207860 267918 207888 270234
rect 207952 270094 207980 270234
rect 207940 270088 207992 270094
rect 207940 270030 207992 270036
rect 208044 269686 208072 278038
rect 208308 273148 208360 273154
rect 208308 273090 208360 273096
rect 208320 271998 208348 273090
rect 208308 271992 208360 271998
rect 208308 271934 208360 271940
rect 208124 270496 208176 270502
rect 208124 270438 208176 270444
rect 208136 270094 208164 270438
rect 208398 270328 208454 270337
rect 208398 270263 208454 270272
rect 208124 270088 208176 270094
rect 208124 270030 208176 270036
rect 207940 269680 207992 269686
rect 207940 269622 207992 269628
rect 208032 269680 208084 269686
rect 208032 269622 208084 269628
rect 207848 267912 207900 267918
rect 207848 267854 207900 267860
rect 207952 264316 207980 269622
rect 208412 264316 208440 270263
rect 208860 269748 208912 269754
rect 208860 269690 208912 269696
rect 208872 264316 208900 269690
rect 209148 269550 209176 278038
rect 209226 271688 209282 271697
rect 209226 271623 209282 271632
rect 209136 269544 209188 269550
rect 209136 269486 209188 269492
rect 209240 264316 209268 271623
rect 209686 271416 209742 271425
rect 209686 271351 209742 271360
rect 209700 264316 209728 271351
rect 210068 269618 210096 278052
rect 210606 271552 210662 271561
rect 210606 271487 210662 271496
rect 210148 269816 210200 269822
rect 210148 269758 210200 269764
rect 210056 269612 210108 269618
rect 210056 269554 210108 269560
rect 210160 264316 210188 269758
rect 210620 264316 210648 271487
rect 211068 269884 211120 269890
rect 211068 269826 211120 269832
rect 211080 264316 211108 269826
rect 211264 269754 211292 278052
rect 212354 271280 212410 271289
rect 212354 271215 212410 271224
rect 211896 269952 211948 269958
rect 211896 269894 211948 269900
rect 211252 269748 211304 269754
rect 211252 269690 211304 269696
rect 211528 266416 211580 266422
rect 211528 266358 211580 266364
rect 211540 264316 211568 266358
rect 211908 264316 211936 269894
rect 212368 264316 212396 271215
rect 212460 269890 212488 278052
rect 213274 271144 213330 271153
rect 213274 271079 213330 271088
rect 212814 270464 212870 270473
rect 212814 270399 212870 270408
rect 212448 269884 212500 269890
rect 212448 269826 212500 269832
rect 212828 264316 212856 270399
rect 213288 264316 213316 271079
rect 213656 270162 213684 278052
rect 214196 272264 214248 272270
rect 214196 272206 214248 272212
rect 213460 270156 213512 270162
rect 213460 270098 213512 270104
rect 213644 270156 213696 270162
rect 213644 270098 213696 270104
rect 213472 267782 213500 270098
rect 213736 270020 213788 270026
rect 213736 269962 213788 269968
rect 213460 267776 213512 267782
rect 213460 267718 213512 267724
rect 213748 264316 213776 269962
rect 214208 264316 214236 272206
rect 214852 269822 214880 278052
rect 215668 272400 215720 272406
rect 215668 272342 215720 272348
rect 215024 272332 215076 272338
rect 215024 272274 215076 272280
rect 214840 269816 214892 269822
rect 214840 269758 214892 269764
rect 214656 267776 214708 267782
rect 214656 267718 214708 267724
rect 214668 264316 214696 267718
rect 215036 264316 215064 272274
rect 215484 270292 215536 270298
rect 215484 270234 215536 270240
rect 215496 264316 215524 270234
rect 215680 264330 215708 272342
rect 215956 270026 215984 278052
rect 216864 272536 216916 272542
rect 216864 272478 216916 272484
rect 215944 270020 215996 270026
rect 215944 269962 215996 269968
rect 216402 268968 216458 268977
rect 216402 268903 216458 268912
rect 215680 264302 215970 264330
rect 216416 264316 216444 268903
rect 216876 264316 216904 272478
rect 217152 269958 217180 278052
rect 217692 272468 217744 272474
rect 217692 272410 217744 272416
rect 217140 269952 217192 269958
rect 217140 269894 217192 269900
rect 217324 267912 217376 267918
rect 217324 267854 217376 267860
rect 217336 264316 217364 267854
rect 217704 264316 217732 272410
rect 218348 270298 218376 278052
rect 219440 272672 219492 272678
rect 219440 272614 219492 272620
rect 218612 272604 218664 272610
rect 218612 272546 218664 272552
rect 218336 270292 218388 270298
rect 218336 270234 218388 270240
rect 218152 267980 218204 267986
rect 218152 267922 218204 267928
rect 218164 264316 218192 267922
rect 218624 264316 218652 272546
rect 219072 270360 219124 270366
rect 219072 270302 219124 270308
rect 219084 264316 219112 270302
rect 219452 264330 219480 272614
rect 219544 267986 219572 278052
rect 220360 272740 220412 272746
rect 220360 272682 220412 272688
rect 219992 270428 220044 270434
rect 219992 270370 220044 270376
rect 219532 267980 219584 267986
rect 219532 267922 219584 267928
rect 219452 264302 219558 264330
rect 220004 264316 220032 270370
rect 220372 264316 220400 272682
rect 220740 270230 220768 278052
rect 221280 273012 221332 273018
rect 221280 272954 221332 272960
rect 220820 270496 220872 270502
rect 220820 270438 220872 270444
rect 220728 270224 220780 270230
rect 220728 270166 220780 270172
rect 220832 264316 220860 270438
rect 221292 264316 221320 272954
rect 221936 270366 221964 278052
rect 222200 272876 222252 272882
rect 222200 272818 222252 272824
rect 221924 270360 221976 270366
rect 221924 270302 221976 270308
rect 221738 268832 221794 268841
rect 221738 268767 221794 268776
rect 221752 264316 221780 268767
rect 222212 264316 222240 272818
rect 223028 272808 223080 272814
rect 223028 272750 223080 272756
rect 222660 270088 222712 270094
rect 222660 270030 222712 270036
rect 222672 264316 222700 270030
rect 223040 264316 223068 272750
rect 223132 270094 223160 278052
rect 223212 272944 223264 272950
rect 223212 272886 223264 272892
rect 223120 270088 223172 270094
rect 223120 270030 223172 270036
rect 223224 264330 223252 272886
rect 224236 270434 224264 278052
rect 225328 273216 225380 273222
rect 225328 273158 225380 273164
rect 224408 273080 224460 273086
rect 224408 273022 224460 273028
rect 224224 270428 224276 270434
rect 224224 270370 224276 270376
rect 223946 268696 224002 268705
rect 223946 268631 224002 268640
rect 223224 264302 223514 264330
rect 223960 264316 223988 268631
rect 224420 264316 224448 273022
rect 224868 269000 224920 269006
rect 224868 268942 224920 268948
rect 224880 264316 224908 268942
rect 225340 264316 225368 273158
rect 225432 270502 225460 278052
rect 226628 272202 226656 278052
rect 227824 272474 227852 278052
rect 227812 272468 227864 272474
rect 227812 272410 227864 272416
rect 229020 272338 229048 278052
rect 229008 272332 229060 272338
rect 229008 272274 229060 272280
rect 230216 272270 230244 278052
rect 231320 272406 231348 278052
rect 232516 272678 232544 278052
rect 232504 272672 232556 272678
rect 232504 272614 232556 272620
rect 233712 272542 233740 278052
rect 234908 272882 234936 278052
rect 236104 272950 236132 278052
rect 236092 272944 236144 272950
rect 236092 272886 236144 272892
rect 234896 272876 234948 272882
rect 234896 272818 234948 272824
rect 237300 272610 237328 278052
rect 238496 272814 238524 278052
rect 238484 272808 238536 272814
rect 238484 272750 238536 272756
rect 239600 272746 239628 278052
rect 239588 272740 239640 272746
rect 239588 272682 239640 272688
rect 237288 272604 237340 272610
rect 237288 272546 237340 272552
rect 233700 272536 233752 272542
rect 233700 272478 233752 272484
rect 231308 272400 231360 272406
rect 231308 272342 231360 272348
rect 230204 272264 230256 272270
rect 230204 272206 230256 272212
rect 226616 272196 226668 272202
rect 226616 272138 226668 272144
rect 240140 272060 240192 272066
rect 240140 272002 240192 272008
rect 227076 271992 227128 271998
rect 227076 271934 227128 271940
rect 225880 271788 225932 271794
rect 225880 271730 225932 271736
rect 225420 270496 225472 270502
rect 225420 270438 225472 270444
rect 225788 269068 225840 269074
rect 225788 269010 225840 269016
rect 225800 264316 225828 269010
rect 225892 264330 225920 271730
rect 226614 268560 226670 268569
rect 226614 268495 226670 268504
rect 225892 264302 226182 264330
rect 226628 264316 226656 268495
rect 227088 264316 227116 271934
rect 227996 271720 228048 271726
rect 227996 271662 228048 271668
rect 227534 268424 227590 268433
rect 227534 268359 227590 268368
rect 227548 264316 227576 268359
rect 228008 264316 228036 271662
rect 229744 271652 229796 271658
rect 229744 271594 229796 271600
rect 228824 271584 228876 271590
rect 228824 271526 228876 271532
rect 228456 268864 228508 268870
rect 228456 268806 228508 268812
rect 228468 264316 228496 268806
rect 228836 264316 228864 271526
rect 229284 268932 229336 268938
rect 229284 268874 229336 268880
rect 229296 264316 229324 268874
rect 229756 264316 229784 271594
rect 232412 271516 232464 271522
rect 232412 271458 232464 271464
rect 230664 271380 230716 271386
rect 230664 271322 230716 271328
rect 230204 268728 230256 268734
rect 230204 268670 230256 268676
rect 230216 264316 230244 268670
rect 230676 264316 230704 271322
rect 231492 271312 231544 271318
rect 231492 271254 231544 271260
rect 231124 268796 231176 268802
rect 231124 268738 231176 268744
rect 231136 264316 231164 268738
rect 231504 264316 231532 271254
rect 231860 271176 231912 271182
rect 231860 271118 231912 271124
rect 231872 267918 231900 271118
rect 231952 268660 232004 268666
rect 231952 268602 232004 268608
rect 231860 267912 231912 267918
rect 231860 267854 231912 267860
rect 231964 264316 231992 268602
rect 232424 264316 232452 271458
rect 233332 271244 233384 271250
rect 233332 271186 233384 271192
rect 232872 268592 232924 268598
rect 232872 268534 232924 268540
rect 232884 264316 232912 268534
rect 233344 264316 233372 271186
rect 234160 271108 234212 271114
rect 234160 271050 234212 271056
rect 233792 268524 233844 268530
rect 233792 268466 233844 268472
rect 233804 264316 233832 268466
rect 234172 264316 234200 271050
rect 236000 271040 236052 271046
rect 236000 270982 236052 270988
rect 234620 270768 234672 270774
rect 234620 270710 234672 270716
rect 234632 269074 234660 270710
rect 234620 269068 234672 269074
rect 234620 269010 234672 269016
rect 234620 268456 234672 268462
rect 234620 268398 234672 268404
rect 234632 264316 234660 268398
rect 235540 268320 235592 268326
rect 235540 268262 235592 268268
rect 235080 267912 235132 267918
rect 235080 267854 235132 267860
rect 235092 264316 235120 267854
rect 235552 264316 235580 268262
rect 236012 264316 236040 270982
rect 238208 270972 238260 270978
rect 238208 270914 238260 270920
rect 237288 270904 237340 270910
rect 237288 270846 237340 270852
rect 236460 268388 236512 268394
rect 236460 268330 236512 268336
rect 236472 264316 236500 268330
rect 236920 268252 236972 268258
rect 236920 268194 236972 268200
rect 236932 264316 236960 268194
rect 237300 264316 237328 270846
rect 237748 268184 237800 268190
rect 237748 268126 237800 268132
rect 237760 264316 237788 268126
rect 238220 264316 238248 270914
rect 239128 270836 239180 270842
rect 239128 270778 239180 270784
rect 238668 268116 238720 268122
rect 238668 268058 238720 268064
rect 238680 264316 238708 268058
rect 239140 264316 239168 270778
rect 239588 269068 239640 269074
rect 239588 269010 239640 269016
rect 239600 264316 239628 269010
rect 240152 268530 240180 272002
rect 240796 271998 240824 278052
rect 241992 273018 242020 278052
rect 243188 273086 243216 278052
rect 243176 273080 243228 273086
rect 243176 273022 243228 273028
rect 241980 273012 242032 273018
rect 241980 272954 242032 272960
rect 240784 271992 240836 271998
rect 240784 271934 240836 271940
rect 244384 271862 244412 278052
rect 244924 272128 244976 272134
rect 244924 272070 244976 272076
rect 240876 271856 240928 271862
rect 240876 271798 240928 271804
rect 244372 271856 244424 271862
rect 244372 271798 244424 271804
rect 240416 269136 240468 269142
rect 240416 269078 240468 269084
rect 240140 268524 240192 268530
rect 240140 268466 240192 268472
rect 239956 268048 240008 268054
rect 239956 267990 240008 267996
rect 239968 264316 239996 267990
rect 240428 264316 240456 269078
rect 240888 264316 240916 271798
rect 241796 271448 241848 271454
rect 241796 271390 241848 271396
rect 241336 269204 241388 269210
rect 241336 269146 241388 269152
rect 241348 264316 241376 269146
rect 241808 264316 241836 271390
rect 242624 270700 242676 270706
rect 242624 270642 242676 270648
rect 242256 270632 242308 270638
rect 242256 270574 242308 270580
rect 242268 264316 242296 270574
rect 242636 264316 242664 270642
rect 244004 269408 244056 269414
rect 244004 269350 244056 269356
rect 243084 269272 243136 269278
rect 243084 269214 243136 269220
rect 243096 264316 243124 269214
rect 243544 268524 243596 268530
rect 243544 268466 243596 268472
rect 243556 264316 243584 268466
rect 244016 264316 244044 269350
rect 244464 269340 244516 269346
rect 244464 269282 244516 269288
rect 244476 264316 244504 269282
rect 244936 264316 244964 272070
rect 245580 271930 245608 278052
rect 245568 271924 245620 271930
rect 245568 271866 245620 271872
rect 246776 271862 246804 278052
rect 246764 271856 246816 271862
rect 246764 271798 246816 271804
rect 247880 271114 247908 278052
rect 249076 271794 249104 278052
rect 249064 271788 249116 271794
rect 249064 271730 249116 271736
rect 250272 271318 250300 278052
rect 251468 271726 251496 278052
rect 251456 271720 251508 271726
rect 251456 271662 251508 271668
rect 252664 271386 252692 278052
rect 253388 272468 253440 272474
rect 253388 272410 253440 272416
rect 252928 272196 252980 272202
rect 252928 272138 252980 272144
rect 252652 271380 252704 271386
rect 252652 271322 252704 271328
rect 250260 271312 250312 271318
rect 250260 271254 250312 271260
rect 247868 271108 247920 271114
rect 247868 271050 247920 271056
rect 252468 270496 252520 270502
rect 252468 270438 252520 270444
rect 252008 270428 252060 270434
rect 252008 270370 252060 270376
rect 251088 270360 251140 270366
rect 251088 270302 251140 270308
rect 249800 270292 249852 270298
rect 249800 270234 249852 270240
rect 248052 270156 248104 270162
rect 248052 270098 248104 270104
rect 247592 269884 247644 269890
rect 247592 269826 247644 269832
rect 247132 269748 247184 269754
rect 247132 269690 247184 269696
rect 245752 269680 245804 269686
rect 245752 269622 245804 269628
rect 245292 269476 245344 269482
rect 245292 269418 245344 269424
rect 245304 264316 245332 269418
rect 245764 264316 245792 269622
rect 246672 269612 246724 269618
rect 246672 269554 246724 269560
rect 246212 269544 246264 269550
rect 246212 269486 246264 269492
rect 246224 264316 246252 269486
rect 246684 264316 246712 269554
rect 247144 264316 247172 269690
rect 247604 264316 247632 269826
rect 248064 264316 248092 270098
rect 248880 270020 248932 270026
rect 248880 269962 248932 269968
rect 248420 269816 248472 269822
rect 248420 269758 248472 269764
rect 248432 264316 248460 269758
rect 248892 264316 248920 269962
rect 249340 269952 249392 269958
rect 249340 269894 249392 269900
rect 249352 264316 249380 269894
rect 249812 264316 249840 270234
rect 250720 270224 250772 270230
rect 250720 270166 250772 270172
rect 250260 267980 250312 267986
rect 250260 267922 250312 267928
rect 250272 264316 250300 267922
rect 250732 264316 250760 270166
rect 251100 264316 251128 270302
rect 251548 270088 251600 270094
rect 251548 270030 251600 270036
rect 251560 264316 251588 270030
rect 252020 264316 252048 270370
rect 252480 264316 252508 270438
rect 252940 264316 252968 272138
rect 253400 264316 253428 272410
rect 253756 272332 253808 272338
rect 253756 272274 253808 272280
rect 253768 264316 253796 272274
rect 253860 271658 253888 278052
rect 254676 272400 254728 272406
rect 254676 272342 254728 272348
rect 254216 272264 254268 272270
rect 254216 272206 254268 272212
rect 253848 271652 253900 271658
rect 253848 271594 253900 271600
rect 254228 264316 254256 272206
rect 254688 264316 254716 272342
rect 254964 271454 254992 278052
rect 256056 272876 256108 272882
rect 256056 272818 256108 272824
rect 255136 272672 255188 272678
rect 255136 272614 255188 272620
rect 254952 271448 255004 271454
rect 254952 271390 255004 271396
rect 255148 264316 255176 272614
rect 255596 272536 255648 272542
rect 255596 272478 255648 272484
rect 255608 264316 255636 272478
rect 256068 264316 256096 272818
rect 256160 270706 256188 278052
rect 256424 272944 256476 272950
rect 256424 272886 256476 272892
rect 256148 270700 256200 270706
rect 256148 270642 256200 270648
rect 256436 264316 256464 272886
rect 257252 272604 257304 272610
rect 257252 272546 257304 272552
rect 257264 264330 257292 272546
rect 257356 271590 257384 278052
rect 257436 272808 257488 272814
rect 257436 272750 257488 272756
rect 257344 271584 257396 271590
rect 257344 271526 257396 271532
rect 257448 264330 257476 272750
rect 257804 272740 257856 272746
rect 257804 272682 257856 272688
rect 256910 264302 257292 264330
rect 257370 264302 257476 264330
rect 257816 264316 257844 272682
rect 258264 272128 258316 272134
rect 258264 272070 258316 272076
rect 258276 264316 258304 272070
rect 258552 271522 258580 278052
rect 259748 273086 259776 278052
rect 260944 273154 260972 278052
rect 260932 273148 260984 273154
rect 260932 273090 260984 273096
rect 259184 273080 259236 273086
rect 259184 273022 259236 273028
rect 259736 273080 259788 273086
rect 259736 273022 259788 273028
rect 258724 273012 258776 273018
rect 258724 272954 258776 272960
rect 258540 271516 258592 271522
rect 258540 271458 258592 271464
rect 258736 264316 258764 272954
rect 259196 264316 259224 273022
rect 260012 272060 260064 272066
rect 260012 272002 260064 272008
rect 259552 271924 259604 271930
rect 259552 271866 259604 271872
rect 259564 264316 259592 271866
rect 260024 264316 260052 272002
rect 262140 271998 262168 278052
rect 263244 273222 263272 278052
rect 263232 273216 263284 273222
rect 263232 273158 263284 273164
rect 262128 271992 262180 271998
rect 262128 271934 262180 271940
rect 264440 271862 264468 278052
rect 265348 273080 265400 273086
rect 265348 273022 265400 273028
rect 260472 271856 260524 271862
rect 260472 271798 260524 271804
rect 264428 271856 264480 271862
rect 264428 271798 264480 271804
rect 260484 264316 260512 271798
rect 261392 271788 261444 271794
rect 261392 271730 261444 271736
rect 260932 271108 260984 271114
rect 260932 271050 260984 271056
rect 260944 264316 260972 271050
rect 261404 264316 261432 271730
rect 262220 271720 262272 271726
rect 262220 271662 262272 271668
rect 261852 271312 261904 271318
rect 261852 271254 261904 271260
rect 261864 264316 261892 271254
rect 262232 264316 262260 271662
rect 263140 271652 263192 271658
rect 263140 271594 263192 271600
rect 262864 271380 262916 271386
rect 262864 271322 262916 271328
rect 262876 264330 262904 271322
rect 262706 264302 262904 264330
rect 263152 264316 263180 271594
rect 264520 271584 264572 271590
rect 264520 271526 264572 271532
rect 263600 271448 263652 271454
rect 263600 271390 263652 271396
rect 263612 264316 263640 271390
rect 264060 270700 264112 270706
rect 264060 270642 264112 270648
rect 264072 264316 264100 270642
rect 264532 264316 264560 271526
rect 264888 271516 264940 271522
rect 264888 271458 264940 271464
rect 264900 264316 264928 271458
rect 265360 264316 265388 273022
rect 265636 270502 265664 278052
rect 266728 273216 266780 273222
rect 266728 273158 266780 273164
rect 265808 273148 265860 273154
rect 265808 273090 265860 273096
rect 265624 270496 265676 270502
rect 265624 270438 265676 270444
rect 265820 264316 265848 273090
rect 266268 271992 266320 271998
rect 266268 271934 266320 271940
rect 266280 264316 266308 271934
rect 266740 264316 266768 273158
rect 266832 271522 266860 278052
rect 268042 278038 268516 278066
rect 267188 271856 267240 271862
rect 267188 271798 267240 271804
rect 266820 271516 266872 271522
rect 266820 271458 266872 271464
rect 267200 264316 267228 271798
rect 268016 271516 268068 271522
rect 268016 271458 268068 271464
rect 267556 270496 267608 270502
rect 267556 270438 267608 270444
rect 267568 264316 267596 270438
rect 268028 264316 268056 271458
rect 268488 264316 268516 278038
rect 268948 278038 269146 278066
rect 268948 264316 268976 278038
rect 270328 270502 270356 278052
rect 269396 270496 269448 270502
rect 269396 270438 269448 270444
rect 270316 270496 270368 270502
rect 270316 270438 270368 270444
rect 271144 270496 271196 270502
rect 271144 270438 271196 270444
rect 269408 264316 269436 270438
rect 269856 270428 269908 270434
rect 269856 270370 269908 270376
rect 269868 264316 269896 270370
rect 270684 270224 270736 270230
rect 270684 270166 270736 270172
rect 270316 269136 270368 269142
rect 270316 269078 270368 269084
rect 270328 264316 270356 269078
rect 270696 264316 270724 270166
rect 271156 264316 271184 270438
rect 271524 270434 271552 278052
rect 271512 270428 271564 270434
rect 271512 270370 271564 270376
rect 271604 270428 271656 270434
rect 271604 270370 271656 270376
rect 271616 264316 271644 270370
rect 272064 270360 272116 270366
rect 272064 270302 272116 270308
rect 272076 264316 272104 270302
rect 272524 270020 272576 270026
rect 272524 269962 272576 269968
rect 272536 264316 272564 269962
rect 272720 269142 272748 278052
rect 273916 270230 273944 278052
rect 275112 270502 275140 278052
rect 275100 270496 275152 270502
rect 275100 270438 275152 270444
rect 276216 270434 276244 278052
rect 276940 270496 276992 270502
rect 276940 270438 276992 270444
rect 276204 270428 276256 270434
rect 276204 270370 276256 270376
rect 273904 270224 273956 270230
rect 273904 270166 273956 270172
rect 272984 270156 273036 270162
rect 272984 270098 273036 270104
rect 272708 269136 272760 269142
rect 272708 269078 272760 269084
rect 272996 264316 273024 270098
rect 273720 270088 273772 270094
rect 273720 270030 273772 270036
rect 273732 264330 273760 270030
rect 274732 269680 274784 269686
rect 274732 269622 274784 269628
rect 273812 268728 273864 268734
rect 273812 268670 273864 268676
rect 273378 264302 273760 264330
rect 273824 264316 273852 268670
rect 274272 268660 274324 268666
rect 274272 268602 274324 268608
rect 274284 264316 274312 268602
rect 274744 264316 274772 269622
rect 275192 268320 275244 268326
rect 275192 268262 275244 268268
rect 275204 264316 275232 268262
rect 275652 268252 275704 268258
rect 275652 268194 275704 268200
rect 275664 264316 275692 268194
rect 276480 267980 276532 267986
rect 276480 267922 276532 267928
rect 276296 267912 276348 267918
rect 276296 267854 276348 267860
rect 276308 264330 276336 267854
rect 276046 264302 276336 264330
rect 276492 264316 276520 267922
rect 276952 264316 276980 270438
rect 277412 270366 277440 278052
rect 277492 270428 277544 270434
rect 277492 270370 277544 270376
rect 277400 270360 277452 270366
rect 277400 270302 277452 270308
rect 277504 264330 277532 270370
rect 277860 270360 277912 270366
rect 277860 270302 277912 270308
rect 277426 264302 277532 264330
rect 277872 264316 277900 270302
rect 278608 270026 278636 278052
rect 278688 270224 278740 270230
rect 278688 270166 278740 270172
rect 278596 270020 278648 270026
rect 278596 269962 278648 269968
rect 278320 269748 278372 269754
rect 278320 269690 278372 269696
rect 278332 264316 278360 269690
rect 278700 264316 278728 270166
rect 279804 270162 279832 278052
rect 279792 270156 279844 270162
rect 279792 270098 279844 270104
rect 281000 270094 281028 278052
rect 280988 270088 281040 270094
rect 280988 270030 281040 270036
rect 281080 270088 281132 270094
rect 281080 270030 281132 270036
rect 279148 270020 279200 270026
rect 279148 269962 279200 269968
rect 279160 264316 279188 269962
rect 279608 269952 279660 269958
rect 279608 269894 279660 269900
rect 279620 264316 279648 269894
rect 280068 269884 280120 269890
rect 280068 269826 280120 269832
rect 280080 264316 280108 269826
rect 280528 269816 280580 269822
rect 280528 269758 280580 269764
rect 280540 264316 280568 269758
rect 281092 269754 281120 270030
rect 281080 269748 281132 269754
rect 281080 269690 281132 269696
rect 281816 269680 281868 269686
rect 281816 269622 281868 269628
rect 281448 269612 281500 269618
rect 281448 269554 281500 269560
rect 280988 269544 281040 269550
rect 280988 269486 281040 269492
rect 281000 264316 281028 269486
rect 281460 264316 281488 269554
rect 281828 264316 281856 269622
rect 282196 268734 282224 278052
rect 282736 269476 282788 269482
rect 282736 269418 282788 269424
rect 282276 269408 282328 269414
rect 282276 269350 282328 269356
rect 282184 268728 282236 268734
rect 282184 268670 282236 268676
rect 282288 264316 282316 269350
rect 282748 264316 282776 269418
rect 283196 269272 283248 269278
rect 283196 269214 283248 269220
rect 283208 264316 283236 269214
rect 283392 268666 283420 278052
rect 284208 271380 284260 271386
rect 284208 271322 284260 271328
rect 283656 269340 283708 269346
rect 283656 269282 283708 269288
rect 283380 268660 283432 268666
rect 283380 268602 283432 268608
rect 283668 264316 283696 269282
rect 284220 264330 284248 271322
rect 284496 269754 284524 278052
rect 285404 271720 285456 271726
rect 285404 271662 285456 271668
rect 284484 269748 284536 269754
rect 284484 269690 284536 269696
rect 284944 269204 284996 269210
rect 284944 269146 284996 269152
rect 284484 269136 284536 269142
rect 284484 269078 284536 269084
rect 284142 264302 284248 264330
rect 284496 264316 284524 269078
rect 284956 264316 284984 269146
rect 285416 264316 285444 271662
rect 285692 268326 285720 278052
rect 286692 272196 286744 272202
rect 286692 272138 286744 272144
rect 285864 271448 285916 271454
rect 285864 271390 285916 271396
rect 285680 268320 285732 268326
rect 285680 268262 285732 268268
rect 285876 264316 285904 271390
rect 286704 264330 286732 272138
rect 286888 268258 286916 278052
rect 287612 272332 287664 272338
rect 287612 272274 287664 272280
rect 287152 272060 287204 272066
rect 287152 272002 287204 272008
rect 286968 271992 287020 271998
rect 286968 271934 287020 271940
rect 286876 268252 286928 268258
rect 286876 268194 286928 268200
rect 286980 264330 287008 271934
rect 286350 264302 286732 264330
rect 286810 264302 287008 264330
rect 287164 264316 287192 272002
rect 287624 264316 287652 272274
rect 288084 267918 288112 278052
rect 288164 272536 288216 272542
rect 288164 272478 288216 272484
rect 288072 267912 288124 267918
rect 288072 267854 288124 267860
rect 288176 264330 288204 272478
rect 288900 272264 288952 272270
rect 288900 272206 288952 272212
rect 288912 264330 288940 272206
rect 289280 267986 289308 278052
rect 289544 271924 289596 271930
rect 289544 271866 289596 271872
rect 289268 267980 289320 267986
rect 289268 267922 289320 267928
rect 289556 264974 289584 271866
rect 289636 271856 289688 271862
rect 289636 271798 289688 271804
rect 289372 264946 289584 264974
rect 289372 264330 289400 264946
rect 289648 264330 289676 271798
rect 289820 271584 289872 271590
rect 289820 271526 289872 271532
rect 288098 264302 288204 264330
rect 288558 264302 288940 264330
rect 289018 264302 289400 264330
rect 289478 264302 289676 264330
rect 289832 264316 289860 271526
rect 290280 271516 290332 271522
rect 290280 271458 290332 271464
rect 290292 264316 290320 271458
rect 290476 270502 290504 278052
rect 291200 273216 291252 273222
rect 291200 273158 291252 273164
rect 290740 271652 290792 271658
rect 290740 271594 290792 271600
rect 290464 270496 290516 270502
rect 290464 270438 290516 270444
rect 290752 264316 290780 271594
rect 291212 264316 291240 273158
rect 291580 270366 291608 278052
rect 292120 273148 292172 273154
rect 292120 273090 292172 273096
rect 291660 271788 291712 271794
rect 291660 271730 291712 271736
rect 291568 270360 291620 270366
rect 291568 270302 291620 270308
rect 291672 264316 291700 271730
rect 292132 264316 292160 273090
rect 292580 272128 292632 272134
rect 292580 272070 292632 272076
rect 292592 264316 292620 272070
rect 292776 270230 292804 278052
rect 293868 273080 293920 273086
rect 293868 273022 293920 273028
rect 293408 272468 293460 272474
rect 293408 272410 293460 272416
rect 292764 270224 292816 270230
rect 292764 270166 292816 270172
rect 292948 269000 293000 269006
rect 292948 268942 293000 268948
rect 292960 264316 292988 268942
rect 293420 264316 293448 272410
rect 293880 264316 293908 273022
rect 293972 270094 294000 278052
rect 294880 272944 294932 272950
rect 294880 272886 294932 272892
rect 293960 270088 294012 270094
rect 293960 270030 294012 270036
rect 294328 269068 294380 269074
rect 294328 269010 294380 269016
rect 294340 264316 294368 269010
rect 294892 264330 294920 272886
rect 295168 270162 295196 278052
rect 296076 273012 296128 273018
rect 296076 272954 296128 272960
rect 295248 272740 295300 272746
rect 295248 272682 295300 272688
rect 295156 270156 295208 270162
rect 295156 270098 295208 270104
rect 294814 264302 294920 264330
rect 295260 264316 295288 272682
rect 295616 270496 295668 270502
rect 295616 270438 295668 270444
rect 295628 264316 295656 270438
rect 296088 264316 296116 272954
rect 296364 270026 296392 278052
rect 296996 270428 297048 270434
rect 296996 270370 297048 270376
rect 296352 270020 296404 270026
rect 296352 269962 296404 269968
rect 296536 268796 296588 268802
rect 296536 268738 296588 268744
rect 296548 264316 296576 268738
rect 297008 264316 297036 270370
rect 297560 269958 297588 278052
rect 298480 278038 298770 278066
rect 298284 270360 298336 270366
rect 298284 270302 298336 270308
rect 297916 270292 297968 270298
rect 297916 270234 297968 270240
rect 297548 269952 297600 269958
rect 297548 269894 297600 269900
rect 297456 268932 297508 268938
rect 297456 268874 297508 268880
rect 297468 264316 297496 268874
rect 297928 264316 297956 270234
rect 298296 264316 298324 270302
rect 298480 269890 298508 278038
rect 298744 270156 298796 270162
rect 298744 270098 298796 270104
rect 298468 269884 298520 269890
rect 298468 269826 298520 269832
rect 298756 264316 298784 270098
rect 299860 269822 299888 278052
rect 300124 270224 300176 270230
rect 300124 270166 300176 270172
rect 299848 269816 299900 269822
rect 299848 269758 299900 269764
rect 299204 268660 299256 268666
rect 299204 268602 299256 268608
rect 299216 264316 299244 268602
rect 299664 267164 299716 267170
rect 299664 267106 299716 267112
rect 299676 264316 299704 267106
rect 300136 264316 300164 270166
rect 300584 270088 300636 270094
rect 300584 270030 300636 270036
rect 300596 264316 300624 270030
rect 301056 269550 301084 278052
rect 301412 272876 301464 272882
rect 301412 272818 301464 272824
rect 301044 269544 301096 269550
rect 301044 269486 301096 269492
rect 300952 267096 301004 267102
rect 300952 267038 301004 267044
rect 300964 264316 300992 267038
rect 301424 264316 301452 272818
rect 301872 272808 301924 272814
rect 301872 272750 301924 272756
rect 301884 264316 301912 272750
rect 302252 269618 302280 278052
rect 303252 270020 303304 270026
rect 303252 269962 303304 269968
rect 302792 269952 302844 269958
rect 302792 269894 302844 269900
rect 302240 269612 302292 269618
rect 302240 269554 302292 269560
rect 302332 267028 302384 267034
rect 302332 266970 302384 266976
rect 302344 264316 302372 266970
rect 302804 264316 302832 269894
rect 303264 264316 303292 269962
rect 303448 269686 303476 278052
rect 304080 272672 304132 272678
rect 304080 272614 304132 272620
rect 303436 269680 303488 269686
rect 303436 269622 303488 269628
rect 303712 266960 303764 266966
rect 303712 266902 303764 266908
rect 303724 264316 303752 266902
rect 304092 264316 304120 272614
rect 304540 272604 304592 272610
rect 304540 272546 304592 272552
rect 304552 264316 304580 272546
rect 304644 269414 304672 278052
rect 305460 269884 305512 269890
rect 305460 269826 305512 269832
rect 304632 269408 304684 269414
rect 304632 269350 304684 269356
rect 305000 266892 305052 266898
rect 305000 266834 305052 266840
rect 305012 264316 305040 266834
rect 305472 264316 305500 269826
rect 305840 269482 305868 278052
rect 306748 269816 306800 269822
rect 306748 269758 306800 269764
rect 305920 269748 305972 269754
rect 305920 269690 305972 269696
rect 305828 269476 305880 269482
rect 305828 269418 305880 269424
rect 305932 264316 305960 269690
rect 306380 266824 306432 266830
rect 306380 266766 306432 266772
rect 306392 264316 306420 266766
rect 306760 264316 306788 269758
rect 307036 269278 307064 278052
rect 307208 272400 307260 272406
rect 307208 272342 307260 272348
rect 307024 269272 307076 269278
rect 307024 269214 307076 269220
rect 307220 264316 307248 272342
rect 308140 269346 308168 278052
rect 309336 271386 309364 278052
rect 309324 271380 309376 271386
rect 309324 271322 309376 271328
rect 308220 269680 308272 269686
rect 308220 269622 308272 269628
rect 308128 269340 308180 269346
rect 308128 269282 308180 269288
rect 307668 266756 307720 266762
rect 307668 266698 307720 266704
rect 307680 264316 307708 266698
rect 308232 264330 308260 269622
rect 310532 269142 310560 278052
rect 310796 269612 310848 269618
rect 310796 269554 310848 269560
rect 310520 269136 310572 269142
rect 310520 269078 310572 269084
rect 309876 268728 309928 268734
rect 309876 268670 309928 268676
rect 309416 268252 309468 268258
rect 309416 268194 309468 268200
rect 308588 267844 308640 267850
rect 308588 267786 308640 267792
rect 308154 264302 308260 264330
rect 308600 264316 308628 267786
rect 309048 266688 309100 266694
rect 309048 266630 309100 266636
rect 309060 264316 309088 266630
rect 309428 264316 309456 268194
rect 309888 264316 309916 268670
rect 310336 266620 310388 266626
rect 310336 266562 310388 266568
rect 310348 264316 310376 266562
rect 310808 264316 310836 269554
rect 311728 269210 311756 278052
rect 312924 271726 312952 278052
rect 313556 271856 313608 271862
rect 313384 271804 313556 271810
rect 313384 271798 313608 271804
rect 313384 271794 313596 271798
rect 313372 271788 313596 271794
rect 313424 271782 313596 271788
rect 313372 271730 313424 271736
rect 312912 271720 312964 271726
rect 312912 271662 312964 271668
rect 313556 271720 313608 271726
rect 313556 271662 313608 271668
rect 313280 271652 313332 271658
rect 313280 271594 313332 271600
rect 313292 271522 313320 271594
rect 313280 271516 313332 271522
rect 313280 271458 313332 271464
rect 312544 270564 312596 270570
rect 312544 270506 312596 270512
rect 311716 269204 311768 269210
rect 311716 269146 311768 269152
rect 312556 268802 312584 270506
rect 313464 269544 313516 269550
rect 313464 269486 313516 269492
rect 312544 268796 312596 268802
rect 312544 268738 312596 268744
rect 312544 268592 312596 268598
rect 312544 268534 312596 268540
rect 312084 268184 312136 268190
rect 312084 268126 312136 268132
rect 311256 267980 311308 267986
rect 311256 267922 311308 267928
rect 311268 264316 311296 267922
rect 311716 266552 311768 266558
rect 311716 266494 311768 266500
rect 311728 264316 311756 266494
rect 312096 264316 312124 268126
rect 312556 264316 312584 268534
rect 313004 266484 313056 266490
rect 313004 266426 313056 266432
rect 313016 264316 313044 266426
rect 313476 264316 313504 269486
rect 313568 268666 313596 271662
rect 314120 271318 314148 278052
rect 315224 272202 315252 278052
rect 315212 272196 315264 272202
rect 315212 272138 315264 272144
rect 315304 272196 315356 272202
rect 315304 272138 315356 272144
rect 314660 271448 314712 271454
rect 314660 271390 314712 271396
rect 314108 271312 314160 271318
rect 314108 271254 314160 271260
rect 314672 268938 314700 271390
rect 314660 268932 314712 268938
rect 314660 268874 314712 268880
rect 313556 268660 313608 268666
rect 313556 268602 313608 268608
rect 313924 268116 313976 268122
rect 313924 268058 313976 268064
rect 313936 264316 313964 268058
rect 314844 268048 314896 268054
rect 314844 267990 314896 267996
rect 314384 265328 314436 265334
rect 314384 265270 314436 265276
rect 314396 264316 314424 265270
rect 314856 264316 314884 267990
rect 315316 264330 315344 272138
rect 316420 271998 316448 278052
rect 317616 272066 317644 278052
rect 318812 272338 318840 278052
rect 319904 274780 319956 274786
rect 319904 274722 319956 274728
rect 318800 272332 318852 272338
rect 318800 272274 318852 272280
rect 318892 272332 318944 272338
rect 318892 272274 318944 272280
rect 317604 272060 317656 272066
rect 317604 272002 317656 272008
rect 317880 272060 317932 272066
rect 317880 272002 317932 272008
rect 316408 271992 316460 271998
rect 316408 271934 316460 271940
rect 316132 269476 316184 269482
rect 316132 269418 316184 269424
rect 315672 266348 315724 266354
rect 315672 266290 315724 266296
rect 315238 264302 315344 264330
rect 315684 264316 315712 266290
rect 316144 264316 316172 269418
rect 316592 269408 316644 269414
rect 316592 269350 316644 269356
rect 316604 264316 316632 269350
rect 317512 269340 317564 269346
rect 317512 269282 317564 269288
rect 317052 265600 317104 265606
rect 317052 265542 317104 265548
rect 317064 264316 317092 265542
rect 317524 264316 317552 269282
rect 317892 264316 317920 272002
rect 318800 271992 318852 271998
rect 318800 271934 318852 271940
rect 318340 265260 318392 265266
rect 318340 265202 318392 265208
rect 318352 264316 318380 265202
rect 318812 264316 318840 271934
rect 318904 268598 318932 272274
rect 319260 269272 319312 269278
rect 319260 269214 319312 269220
rect 318892 268592 318944 268598
rect 318892 268534 318944 268540
rect 319272 264316 319300 269214
rect 319916 264330 319944 274722
rect 320008 272542 320036 278052
rect 320272 274916 320324 274922
rect 320272 274858 320324 274864
rect 319996 272536 320048 272542
rect 319996 272478 320048 272484
rect 320088 272536 320140 272542
rect 320088 272478 320140 272484
rect 320100 268734 320128 272478
rect 320180 270700 320232 270706
rect 320180 270642 320232 270648
rect 320088 268728 320140 268734
rect 320088 268670 320140 268676
rect 320192 267850 320220 270642
rect 320180 267844 320232 267850
rect 320180 267786 320232 267792
rect 320284 264330 320312 274858
rect 321008 274712 321060 274718
rect 321008 274654 321060 274660
rect 320548 271856 320600 271862
rect 320548 271798 320600 271804
rect 319746 264302 319944 264330
rect 320206 264302 320312 264330
rect 320560 264316 320588 271798
rect 321020 264316 321048 274654
rect 321204 272270 321232 278052
rect 321192 272264 321244 272270
rect 321192 272206 321244 272212
rect 322400 271930 322428 278052
rect 322756 274644 322808 274650
rect 322756 274586 322808 274592
rect 322388 271924 322440 271930
rect 322388 271866 322440 271872
rect 321928 269204 321980 269210
rect 321928 269146 321980 269152
rect 321468 265396 321520 265402
rect 321468 265338 321520 265344
rect 321480 264316 321508 265338
rect 321940 264316 321968 269146
rect 322768 264330 322796 274586
rect 323216 271856 323268 271862
rect 323216 271798 323268 271804
rect 322848 269136 322900 269142
rect 322848 269078 322900 269084
rect 322414 264302 322796 264330
rect 322860 264316 322888 269078
rect 323228 264316 323256 271798
rect 323504 271658 323532 278052
rect 323676 273624 323728 273630
rect 323676 273566 323728 273572
rect 323492 271652 323544 271658
rect 323492 271594 323544 271600
rect 323688 264316 323716 273566
rect 324700 271590 324728 278052
rect 325516 273760 325568 273766
rect 325516 273702 325568 273708
rect 325332 272264 325384 272270
rect 325332 272206 325384 272212
rect 324688 271584 324740 271590
rect 324688 271526 324740 271532
rect 324136 270836 324188 270842
rect 324136 270778 324188 270784
rect 324148 264316 324176 270778
rect 325344 268054 325372 272206
rect 325332 268048 325384 268054
rect 325332 267990 325384 267996
rect 324596 267912 324648 267918
rect 324596 267854 324648 267860
rect 324608 264316 324636 267854
rect 325528 264974 325556 273702
rect 325896 271386 325924 278052
rect 326344 273692 326396 273698
rect 326344 273634 326396 273640
rect 325884 271380 325936 271386
rect 325884 271322 325936 271328
rect 325976 270904 326028 270910
rect 325976 270846 326028 270852
rect 325608 265464 325660 265470
rect 325608 265406 325660 265412
rect 325436 264946 325556 264974
rect 325436 264330 325464 264946
rect 325620 264330 325648 265406
rect 325082 264302 325464 264330
rect 325542 264302 325648 264330
rect 325988 264316 326016 270846
rect 326356 264316 326384 273634
rect 327092 271522 327120 278052
rect 327724 273828 327776 273834
rect 327724 273770 327776 273776
rect 327080 271516 327132 271522
rect 327080 271458 327132 271464
rect 327172 270768 327224 270774
rect 327172 270710 327224 270716
rect 327184 268190 327212 270710
rect 327540 270632 327592 270638
rect 327540 270574 327592 270580
rect 327552 268258 327580 270574
rect 327540 268252 327592 268258
rect 327540 268194 327592 268200
rect 327172 268184 327224 268190
rect 327172 268126 327224 268132
rect 327264 268184 327316 268190
rect 327264 268126 327316 268132
rect 326804 265532 326856 265538
rect 326804 265474 326856 265480
rect 326816 264316 326844 265474
rect 327276 264316 327304 268126
rect 327736 264316 327764 273770
rect 328288 273222 328316 278052
rect 329012 273896 329064 273902
rect 329012 273838 329064 273844
rect 328276 273216 328328 273222
rect 328276 273158 328328 273164
rect 328644 270972 328696 270978
rect 328644 270914 328696 270920
rect 328184 268252 328236 268258
rect 328184 268194 328236 268200
rect 328196 264316 328224 268194
rect 328656 264316 328684 270914
rect 329024 264316 329052 273838
rect 329484 271794 329512 278052
rect 330588 273154 330616 278052
rect 331680 274032 331732 274038
rect 331680 273974 331732 273980
rect 330760 273964 330812 273970
rect 330760 273906 330812 273912
rect 330576 273148 330628 273154
rect 330576 273090 330628 273096
rect 329472 271788 329524 271794
rect 329472 271730 329524 271736
rect 329932 268320 329984 268326
rect 329932 268262 329984 268268
rect 329472 268048 329524 268054
rect 329472 267990 329524 267996
rect 329484 264316 329512 267990
rect 329944 264316 329972 268262
rect 330772 264330 330800 273906
rect 331312 268524 331364 268530
rect 331312 268466 331364 268472
rect 330852 268388 330904 268394
rect 330852 268330 330904 268336
rect 330418 264302 330800 264330
rect 330864 264316 330892 268330
rect 331324 264316 331352 268466
rect 331692 264316 331720 273974
rect 331784 272134 331812 278052
rect 331772 272128 331824 272134
rect 331772 272070 331824 272076
rect 331864 272128 331916 272134
rect 331864 272070 331916 272076
rect 331876 268530 331904 272070
rect 332140 271108 332192 271114
rect 332140 271050 332192 271056
rect 331864 268524 331916 268530
rect 331864 268466 331916 268472
rect 332152 264316 332180 271050
rect 332416 271040 332468 271046
rect 332416 270982 332468 270988
rect 332428 268054 332456 270982
rect 332980 269006 333008 278052
rect 333428 274100 333480 274106
rect 333428 274042 333480 274048
rect 332968 269000 333020 269006
rect 332968 268942 333020 268948
rect 332600 268456 332652 268462
rect 332600 268398 332652 268404
rect 332416 268048 332468 268054
rect 332416 267990 332468 267996
rect 332612 264316 332640 268398
rect 332692 268116 332744 268122
rect 332692 268058 332744 268064
rect 332704 267918 332732 268058
rect 332692 267912 332744 267918
rect 332692 267854 332744 267860
rect 333440 264330 333468 274042
rect 334176 272474 334204 278052
rect 334348 274168 334400 274174
rect 334348 274110 334400 274116
rect 334164 272468 334216 272474
rect 334164 272410 334216 272416
rect 334256 272468 334308 272474
rect 334256 272410 334308 272416
rect 333520 268524 333572 268530
rect 333520 268466 333572 268472
rect 333086 264302 333468 264330
rect 333532 264316 333560 268466
rect 334268 264330 334296 272410
rect 334006 264302 334296 264330
rect 334360 264316 334388 274110
rect 335372 273086 335400 278052
rect 335728 274236 335780 274242
rect 335728 274178 335780 274184
rect 335360 273080 335412 273086
rect 335360 273022 335412 273028
rect 334808 271176 334860 271182
rect 334808 271118 334860 271124
rect 334820 264316 334848 271118
rect 335268 268592 335320 268598
rect 335268 268534 335320 268540
rect 335280 264316 335308 268534
rect 335740 264316 335768 274178
rect 336464 271312 336516 271318
rect 336464 271254 336516 271260
rect 336188 268660 336240 268666
rect 336188 268602 336240 268608
rect 336200 264316 336228 268602
rect 336476 264330 336504 271254
rect 336568 269074 336596 278052
rect 337108 274304 337160 274310
rect 337108 274246 337160 274252
rect 336556 269068 336608 269074
rect 336556 269010 336608 269016
rect 336476 264302 336674 264330
rect 337120 264316 337148 274246
rect 337764 272950 337792 278052
rect 337752 272944 337804 272950
rect 337752 272886 337804 272892
rect 338868 272746 338896 278052
rect 339776 274372 339828 274378
rect 339776 274314 339828 274320
rect 338856 272740 338908 272746
rect 338856 272682 338908 272688
rect 339408 272740 339460 272746
rect 339408 272682 339460 272688
rect 337476 271244 337528 271250
rect 337476 271186 337528 271192
rect 337488 264316 337516 271186
rect 338856 268796 338908 268802
rect 338856 268738 338908 268744
rect 337936 268728 337988 268734
rect 337936 268670 337988 268676
rect 337948 264316 337976 268670
rect 338396 265668 338448 265674
rect 338396 265610 338448 265616
rect 338408 264316 338436 265610
rect 338868 264316 338896 268738
rect 339420 264330 339448 272682
rect 339342 264302 339448 264330
rect 339788 264316 339816 274314
rect 340064 270502 340092 278052
rect 341260 273018 341288 278052
rect 341248 273012 341300 273018
rect 341248 272954 341300 272960
rect 342168 271448 342220 271454
rect 342168 271390 342220 271396
rect 340144 271380 340196 271386
rect 340144 271322 340196 271328
rect 340052 270496 340104 270502
rect 340052 270438 340104 270444
rect 340156 264316 340184 271322
rect 341524 268932 341576 268938
rect 341524 268874 341576 268880
rect 340604 268864 340656 268870
rect 340604 268806 340656 268812
rect 340616 264316 340644 268806
rect 341064 265736 341116 265742
rect 341064 265678 341116 265684
rect 341076 264316 341104 265678
rect 341536 264316 341564 268874
rect 342180 264330 342208 271390
rect 342456 270570 342484 278052
rect 342536 274440 342588 274446
rect 342536 274382 342588 274388
rect 342444 270564 342496 270570
rect 342444 270506 342496 270512
rect 342548 264330 342576 274382
rect 342812 273080 342864 273086
rect 342812 273022 342864 273028
rect 342010 264302 342208 264330
rect 342470 264302 342576 264330
rect 342824 264316 342852 273022
rect 343652 270434 343680 278052
rect 343732 274576 343784 274582
rect 343732 274518 343784 274524
rect 343640 270428 343692 270434
rect 343640 270370 343692 270376
rect 343272 269068 343324 269074
rect 343272 269010 343324 269016
rect 343284 264316 343312 269010
rect 343744 264316 343772 274518
rect 344848 271522 344876 278052
rect 345112 274508 345164 274514
rect 345112 274450 345164 274456
rect 344836 271516 344888 271522
rect 344836 271458 344888 271464
rect 344928 271516 344980 271522
rect 344928 271458 344980 271464
rect 344192 269000 344244 269006
rect 344192 268942 344244 268948
rect 344204 264316 344232 268942
rect 344940 264330 344968 271458
rect 344678 264302 344968 264330
rect 345124 264316 345152 274450
rect 345480 273216 345532 273222
rect 345480 273158 345532 273164
rect 345492 264316 345520 273158
rect 345952 270298 345980 278052
rect 347148 270570 347176 278052
rect 347780 276004 347832 276010
rect 347780 275946 347832 275952
rect 347596 271584 347648 271590
rect 347596 271526 347648 271532
rect 347136 270564 347188 270570
rect 347136 270506 347188 270512
rect 346032 270496 346084 270502
rect 346032 270438 346084 270444
rect 345940 270292 345992 270298
rect 345940 270234 345992 270240
rect 346044 264330 346072 270438
rect 346860 270428 346912 270434
rect 346860 270370 346912 270376
rect 346400 265804 346452 265810
rect 346400 265746 346452 265752
rect 345966 264302 346072 264330
rect 346412 264316 346440 265746
rect 346872 264316 346900 270370
rect 347608 264330 347636 271526
rect 347346 264302 347636 264330
rect 347792 264316 347820 275946
rect 347872 273012 347924 273018
rect 347872 272954 347924 272960
rect 347884 270230 347912 272954
rect 348240 271652 348292 271658
rect 348240 271594 348292 271600
rect 347872 270224 347924 270230
rect 347872 270166 347924 270172
rect 348252 264316 348280 271594
rect 348344 270162 348372 278052
rect 349540 271726 349568 278052
rect 350172 275936 350224 275942
rect 350172 275878 350224 275884
rect 350080 272944 350132 272950
rect 350080 272886 350132 272892
rect 349528 271720 349580 271726
rect 349528 271662 349580 271668
rect 348608 270360 348660 270366
rect 348608 270302 348660 270308
rect 348332 270156 348384 270162
rect 348332 270098 348384 270104
rect 348620 264316 348648 270302
rect 349528 270292 349580 270298
rect 349528 270234 349580 270240
rect 349068 265872 349120 265878
rect 349068 265814 349120 265820
rect 349080 264316 349108 265814
rect 349540 264316 349568 270234
rect 350092 264330 350120 272886
rect 350014 264302 350120 264330
rect 350184 264330 350212 275878
rect 350736 267170 350764 278052
rect 351932 273018 351960 278052
rect 351920 273012 351972 273018
rect 351920 272954 351972 272960
rect 350908 271720 350960 271726
rect 350908 271662 350960 271668
rect 350724 267164 350776 267170
rect 350724 267106 350776 267112
rect 350184 264302 350474 264330
rect 350920 264316 350948 271662
rect 353022 271144 353078 271153
rect 353022 271079 353078 271088
rect 351276 270224 351328 270230
rect 351276 270166 351328 270172
rect 351288 264316 351316 270166
rect 352194 268424 352250 268433
rect 352194 268359 352250 268368
rect 351736 265940 351788 265946
rect 351736 265882 351788 265888
rect 351748 264316 351776 265882
rect 352208 264316 352236 268359
rect 353036 264330 353064 271079
rect 353128 270094 353156 278052
rect 353208 275868 353260 275874
rect 353208 275810 353260 275816
rect 353116 270088 353168 270094
rect 353116 270030 353168 270036
rect 353220 264330 353248 275810
rect 353576 271788 353628 271794
rect 353576 271730 353628 271736
rect 352682 264302 353064 264330
rect 353142 264302 353248 264330
rect 353588 264316 353616 271730
rect 353942 268560 353998 268569
rect 353942 268495 353998 268504
rect 353956 264316 353984 268495
rect 354232 267102 354260 278052
rect 355428 272882 355456 278052
rect 355784 275800 355836 275806
rect 355784 275742 355836 275748
rect 355416 272876 355468 272882
rect 355416 272818 355468 272824
rect 355322 271280 355378 271289
rect 355322 271215 355378 271224
rect 354862 268696 354918 268705
rect 354862 268631 354918 268640
rect 354220 267096 354272 267102
rect 354220 267038 354272 267044
rect 354404 266008 354456 266014
rect 354404 265950 354456 265956
rect 354416 264316 354444 265950
rect 354876 264316 354904 268631
rect 355336 264316 355364 271215
rect 355796 264316 355824 275742
rect 356244 273148 356296 273154
rect 356244 273090 356296 273096
rect 356256 264316 356284 273090
rect 356624 272814 356652 278052
rect 356612 272808 356664 272814
rect 356612 272750 356664 272756
rect 357530 268968 357586 268977
rect 357530 268903 357586 268912
rect 356610 268832 356666 268841
rect 356610 268767 356666 268776
rect 356624 264316 356652 268767
rect 357072 266076 357124 266082
rect 357072 266018 357124 266024
rect 357084 264316 357112 266018
rect 357544 264316 357572 268903
rect 357820 267034 357848 278052
rect 358544 275732 358596 275738
rect 358544 275674 358596 275680
rect 357990 271416 358046 271425
rect 357990 271351 358046 271360
rect 357808 267028 357860 267034
rect 357808 266970 357860 266976
rect 358004 264316 358032 271351
rect 358556 264330 358584 275674
rect 358910 271552 358966 271561
rect 358910 271487 358966 271496
rect 358478 264302 358584 264330
rect 358924 264316 358952 271487
rect 359016 269958 359044 278052
rect 359936 278038 360226 278066
rect 359372 270156 359424 270162
rect 359372 270098 359424 270104
rect 359004 269952 359056 269958
rect 359004 269894 359056 269900
rect 359384 264316 359412 270098
rect 359936 270026 359964 278038
rect 361026 271688 361082 271697
rect 361026 271623 361082 271632
rect 360200 270088 360252 270094
rect 360200 270030 360252 270036
rect 359924 270020 359976 270026
rect 359924 269962 359976 269968
rect 359740 266144 359792 266150
rect 359740 266086 359792 266092
rect 359752 264316 359780 266086
rect 360212 264316 360240 270030
rect 361040 264330 361068 271623
rect 361408 266966 361436 278052
rect 361488 275664 361540 275670
rect 361488 275606 361540 275612
rect 361396 266960 361448 266966
rect 361396 266902 361448 266908
rect 361500 264330 361528 275606
rect 361580 273012 361632 273018
rect 361580 272954 361632 272960
rect 360686 264302 361068 264330
rect 361146 264302 361528 264330
rect 361592 264316 361620 272954
rect 362512 272678 362540 278052
rect 362500 272672 362552 272678
rect 362500 272614 362552 272620
rect 363708 272610 363736 278052
rect 363972 275596 364024 275602
rect 363972 275538 364024 275544
rect 363880 272808 363932 272814
rect 363880 272750 363932 272756
rect 363696 272604 363748 272610
rect 363696 272546 363748 272552
rect 362866 270464 362922 270473
rect 362866 270399 362922 270408
rect 362038 270328 362094 270337
rect 362038 270263 362094 270272
rect 362052 264316 362080 270263
rect 362408 266212 362460 266218
rect 362408 266154 362460 266160
rect 362420 264316 362448 266154
rect 362880 264316 362908 270399
rect 363892 264974 363920 272750
rect 363708 264946 363920 264974
rect 363708 264330 363736 264946
rect 363984 264330 364012 275538
rect 364062 273184 364118 273193
rect 364062 273119 364118 273128
rect 363354 264302 363736 264330
rect 363814 264302 364012 264330
rect 364076 264330 364104 273119
rect 364708 270020 364760 270026
rect 364708 269962 364760 269968
rect 364076 264302 364274 264330
rect 364720 264316 364748 269962
rect 364904 266898 364932 278052
rect 365534 270192 365590 270201
rect 365534 270127 365590 270136
rect 364892 266892 364944 266898
rect 364892 266834 364944 266840
rect 365076 266280 365128 266286
rect 365076 266222 365128 266228
rect 365088 264316 365116 266222
rect 365548 264316 365576 270127
rect 366100 269890 366128 278052
rect 366456 275528 366508 275534
rect 366456 275470 366508 275476
rect 366088 269884 366140 269890
rect 366088 269826 366140 269832
rect 365994 268288 366050 268297
rect 365994 268223 366050 268232
rect 366008 264316 366036 268223
rect 366468 264316 366496 275470
rect 366914 273048 366970 273057
rect 366914 272983 366970 272992
rect 366928 264316 366956 272983
rect 367296 269754 367324 278052
rect 367376 269952 367428 269958
rect 367376 269894 367428 269900
rect 367284 269748 367336 269754
rect 367284 269690 367336 269696
rect 367388 264316 367416 269894
rect 368204 269884 368256 269890
rect 368204 269826 368256 269832
rect 367744 267708 367796 267714
rect 367744 267650 367796 267656
rect 367756 264316 367784 267650
rect 368216 264316 368244 269826
rect 368492 266830 368520 278052
rect 369124 275460 369176 275466
rect 369124 275402 369176 275408
rect 368662 272912 368718 272921
rect 368662 272847 368718 272856
rect 368480 266824 368532 266830
rect 368480 266766 368532 266772
rect 368676 264316 368704 272847
rect 369136 264316 369164 275402
rect 369596 269822 369624 278052
rect 369674 272776 369730 272785
rect 369674 272711 369730 272720
rect 369584 269816 369636 269822
rect 369584 269758 369636 269764
rect 369688 264330 369716 272711
rect 370792 272406 370820 278052
rect 371792 275392 371844 275398
rect 371792 275334 371844 275340
rect 370780 272400 370832 272406
rect 370780 272342 370832 272348
rect 370042 270056 370098 270065
rect 370042 269991 370098 270000
rect 369610 264302 369716 264330
rect 370056 264316 370084 269991
rect 370870 269920 370926 269929
rect 370870 269855 370926 269864
rect 370504 267640 370556 267646
rect 370504 267582 370556 267588
rect 370516 264316 370544 267582
rect 370884 264316 370912 269855
rect 371332 267980 371384 267986
rect 371332 267922 371384 267928
rect 371344 264316 371372 267922
rect 371804 264316 371832 275334
rect 371988 266762 372016 278052
rect 372804 272876 372856 272882
rect 372804 272818 372856 272824
rect 372618 272640 372674 272649
rect 372618 272575 372674 272584
rect 372434 272504 372490 272513
rect 372434 272439 372490 272448
rect 372068 272400 372120 272406
rect 372068 272342 372120 272348
rect 372080 268297 372108 272342
rect 372066 268288 372122 268297
rect 372066 268223 372122 268232
rect 371976 266756 372028 266762
rect 371976 266698 372028 266704
rect 372448 264330 372476 272439
rect 372632 268002 372660 272575
rect 372712 269816 372764 269822
rect 372712 269758 372764 269764
rect 372540 267986 372660 268002
rect 372528 267980 372660 267986
rect 372580 267974 372660 267980
rect 372528 267922 372580 267928
rect 372278 264302 372476 264330
rect 372724 264316 372752 269758
rect 372816 267918 372844 272818
rect 373184 269686 373212 278052
rect 374380 270706 374408 278052
rect 375288 275324 375340 275330
rect 375288 275266 375340 275272
rect 374368 270700 374420 270706
rect 374368 270642 374420 270648
rect 374000 269748 374052 269754
rect 374000 269690 374052 269696
rect 373172 269680 373224 269686
rect 373172 269622 373224 269628
rect 372804 267912 372856 267918
rect 372804 267854 372856 267860
rect 373172 267572 373224 267578
rect 373172 267514 373224 267520
rect 373184 264316 373212 267514
rect 373540 267504 373592 267510
rect 373540 267446 373592 267452
rect 373552 264316 373580 267446
rect 374012 264316 374040 269690
rect 374460 267436 374512 267442
rect 374460 267378 374512 267384
rect 374472 264316 374500 267378
rect 375300 264330 375328 275266
rect 375380 272672 375432 272678
rect 375380 272614 375432 272620
rect 374946 264302 375328 264330
rect 375392 264316 375420 272614
rect 375576 266694 375604 278052
rect 376772 270638 376800 278052
rect 377876 272542 377904 278052
rect 377956 275256 378008 275262
rect 377956 275198 378008 275204
rect 377864 272536 377916 272542
rect 377864 272478 377916 272484
rect 376760 270632 376812 270638
rect 376760 270574 376812 270580
rect 376666 269784 376722 269793
rect 376666 269719 376722 269728
rect 376208 267368 376260 267374
rect 376208 267310 376260 267316
rect 375840 267300 375892 267306
rect 375840 267242 375892 267248
rect 375564 266688 375616 266694
rect 375564 266630 375616 266636
rect 375852 264316 375880 267242
rect 376220 264316 376248 267310
rect 376680 264316 376708 269719
rect 377128 267232 377180 267238
rect 377128 267174 377180 267180
rect 377140 264316 377168 267174
rect 377968 264330 377996 275198
rect 378048 272604 378100 272610
rect 378048 272546 378100 272552
rect 377614 264302 377996 264330
rect 378060 264316 378088 272546
rect 378508 267164 378560 267170
rect 378508 267106 378560 267112
rect 378520 264316 378548 267106
rect 378876 267096 378928 267102
rect 378876 267038 378928 267044
rect 378888 264316 378916 267038
rect 379072 266626 379100 278052
rect 379336 269680 379388 269686
rect 379336 269622 379388 269628
rect 379060 266620 379112 266626
rect 379060 266562 379112 266568
rect 379348 264316 379376 269622
rect 380268 269618 380296 278052
rect 380348 275188 380400 275194
rect 380348 275130 380400 275136
rect 380256 269612 380308 269618
rect 380256 269554 380308 269560
rect 379796 267028 379848 267034
rect 379796 266970 379848 266976
rect 379808 264316 379836 266970
rect 380360 264330 380388 275130
rect 381464 272882 381492 278052
rect 381452 272876 381504 272882
rect 381452 272818 381504 272824
rect 380714 272368 380770 272377
rect 380714 272303 380770 272312
rect 380282 264302 380388 264330
rect 380728 264316 380756 272303
rect 382002 269648 382058 269657
rect 382002 269583 382058 269592
rect 381636 266960 381688 266966
rect 381636 266902 381688 266908
rect 381176 266892 381228 266898
rect 381176 266834 381228 266840
rect 381188 264316 381216 266834
rect 381648 264316 381676 266902
rect 382016 264316 382044 269583
rect 382464 266824 382516 266830
rect 382464 266766 382516 266772
rect 382476 264316 382504 266766
rect 382660 266558 382688 278052
rect 382924 275120 382976 275126
rect 382924 275062 382976 275068
rect 382648 266552 382700 266558
rect 382648 266494 382700 266500
rect 382936 264316 382964 275062
rect 383660 272876 383712 272882
rect 383660 272818 383712 272824
rect 383476 270700 383528 270706
rect 383476 270642 383528 270648
rect 383488 264330 383516 270642
rect 383672 268054 383700 272818
rect 383856 270774 383884 278052
rect 384960 272338 384988 278052
rect 385592 275052 385644 275058
rect 385592 274994 385644 275000
rect 384948 272332 385000 272338
rect 384948 272274 385000 272280
rect 383844 270768 383896 270774
rect 383844 270710 383896 270716
rect 384672 269612 384724 269618
rect 384672 269554 384724 269560
rect 383660 268048 383712 268054
rect 383660 267990 383712 267996
rect 384304 266756 384356 266762
rect 384304 266698 384356 266704
rect 383844 266688 383896 266694
rect 383844 266630 383896 266636
rect 383410 264302 383516 264330
rect 383856 264316 383884 266630
rect 384316 264316 384344 266698
rect 384684 264316 384712 269554
rect 385132 266620 385184 266626
rect 385132 266562 385184 266568
rect 385144 264316 385172 266562
rect 385604 264316 385632 274994
rect 386156 266490 386184 278052
rect 386984 278038 387366 278066
rect 386236 270768 386288 270774
rect 386236 270710 386288 270716
rect 386144 266484 386196 266490
rect 386144 266426 386196 266432
rect 386248 264330 386276 270710
rect 386984 269550 387012 278038
rect 387248 276072 387300 276078
rect 387248 276014 387300 276020
rect 387260 274922 387288 276014
rect 387248 274916 387300 274922
rect 387248 274858 387300 274864
rect 388260 273556 388312 273562
rect 388260 273498 388312 273504
rect 386972 269544 387024 269550
rect 386972 269486 387024 269492
rect 387340 269544 387392 269550
rect 387340 269486 387392 269492
rect 386970 267200 387026 267209
rect 386970 267135 387026 267144
rect 386512 266552 386564 266558
rect 386512 266494 386564 266500
rect 386078 264302 386276 264330
rect 386524 264316 386552 266494
rect 386984 264316 387012 267135
rect 387352 264316 387380 269486
rect 387432 269340 387484 269346
rect 387432 269282 387484 269288
rect 387444 268054 387472 269282
rect 387432 268048 387484 268054
rect 387432 267990 387484 267996
rect 387800 266484 387852 266490
rect 387800 266426 387852 266432
rect 387812 264316 387840 266426
rect 388272 264316 388300 273498
rect 388548 272882 388576 278052
rect 388536 272876 388588 272882
rect 388536 272818 388588 272824
rect 388996 270632 389048 270638
rect 388996 270574 389048 270580
rect 389008 264330 389036 270574
rect 389638 267064 389694 267073
rect 389638 266999 389694 267008
rect 389180 266416 389232 266422
rect 389180 266358 389232 266364
rect 388746 264302 389036 264330
rect 389192 264316 389220 266358
rect 389652 264316 389680 266999
rect 389744 265334 389772 278052
rect 390468 272876 390520 272882
rect 390468 272818 390520 272824
rect 390480 272406 390508 272818
rect 390468 272400 390520 272406
rect 390468 272342 390520 272348
rect 390008 272332 390060 272338
rect 390008 272274 390060 272280
rect 389732 265328 389784 265334
rect 389732 265270 389784 265276
rect 390020 264316 390048 272274
rect 390940 272270 390968 278052
rect 391020 273284 391072 273290
rect 391020 273226 391072 273232
rect 390928 272264 390980 272270
rect 390928 272206 390980 272212
rect 390466 266928 390522 266937
rect 390466 266863 390522 266872
rect 390480 264316 390508 266863
rect 391032 264330 391060 273226
rect 391572 272536 391624 272542
rect 391572 272478 391624 272484
rect 391204 272400 391256 272406
rect 391204 272342 391256 272348
rect 391112 272332 391164 272338
rect 391112 272274 391164 272280
rect 391124 270638 391152 272274
rect 391216 270774 391244 272342
rect 391204 270768 391256 270774
rect 391204 270710 391256 270716
rect 391584 270706 391612 272478
rect 392136 272202 392164 278052
rect 392228 278038 393254 278066
rect 392124 272196 392176 272202
rect 392124 272138 392176 272144
rect 391572 270700 391624 270706
rect 391572 270642 391624 270648
rect 391112 270632 391164 270638
rect 391112 270574 391164 270580
rect 391386 269512 391442 269521
rect 391386 269447 391442 269456
rect 390954 264302 391060 264330
rect 391400 264316 391428 269447
rect 391846 266792 391902 266801
rect 391846 266727 391902 266736
rect 391860 264316 391888 266727
rect 392228 266354 392256 278038
rect 393594 274272 393650 274281
rect 393594 274207 393650 274216
rect 392768 269476 392820 269482
rect 392768 269418 392820 269424
rect 392216 266348 392268 266354
rect 392216 266290 392268 266296
rect 392308 266348 392360 266354
rect 392308 266290 392360 266296
rect 392320 264316 392348 266290
rect 392780 264316 392808 269418
rect 393134 266656 393190 266665
rect 393134 266591 393190 266600
rect 393148 264316 393176 266591
rect 393608 264316 393636 274207
rect 394056 272196 394108 272202
rect 394056 272138 394108 272144
rect 394068 264316 394096 272138
rect 394436 269414 394464 278052
rect 395434 272232 395490 272241
rect 395434 272167 395490 272176
rect 394424 269408 394476 269414
rect 394424 269350 394476 269356
rect 394514 266520 394570 266529
rect 394514 266455 394570 266464
rect 394528 264316 394556 266455
rect 394700 265600 394752 265606
rect 394700 265542 394752 265548
rect 394976 265600 395028 265606
rect 394976 265542 395028 265548
rect 394712 265402 394740 265542
rect 394700 265396 394752 265402
rect 394700 265338 394752 265344
rect 394988 264316 395016 265542
rect 395448 264316 395476 272167
rect 395632 269346 395660 278052
rect 396262 275768 396318 275777
rect 396262 275703 396318 275712
rect 395802 274408 395858 274417
rect 395802 274343 395858 274352
rect 395620 269340 395672 269346
rect 395620 269282 395672 269288
rect 395816 264316 395844 274343
rect 396276 264316 396304 275703
rect 396724 269408 396776 269414
rect 396724 269350 396776 269356
rect 396736 264316 396764 269350
rect 396828 265402 396856 278052
rect 397366 275904 397422 275913
rect 397366 275839 397422 275848
rect 397184 269204 397236 269210
rect 397184 269146 397236 269152
rect 397196 267986 397224 269146
rect 397184 267980 397236 267986
rect 397184 267922 397236 267928
rect 396816 265396 396868 265402
rect 396816 265338 396868 265344
rect 397380 264330 397408 275839
rect 398024 268054 398052 278052
rect 398930 275632 398986 275641
rect 398930 275567 398986 275576
rect 398470 275496 398526 275505
rect 398470 275431 398526 275440
rect 398012 268048 398064 268054
rect 398012 267990 398064 267996
rect 398104 267776 398156 267782
rect 398104 267718 398156 267724
rect 397642 267472 397698 267481
rect 397642 267407 397698 267416
rect 397210 264302 397408 264330
rect 397656 264316 397684 267407
rect 398116 264316 398144 267718
rect 398484 264316 398512 275431
rect 398944 264316 398972 275567
rect 399220 272066 399248 278052
rect 400232 278038 400338 278066
rect 399850 275224 399906 275233
rect 399850 275159 399906 275168
rect 399208 272060 399260 272066
rect 399208 272002 399260 272008
rect 399576 272060 399628 272066
rect 399576 272002 399628 272008
rect 399392 269340 399444 269346
rect 399392 269282 399444 269288
rect 399404 264316 399432 269282
rect 399588 267782 399616 272002
rect 399576 267776 399628 267782
rect 399576 267718 399628 267724
rect 399864 264316 399892 275159
rect 400232 265266 400260 278038
rect 401138 275360 401194 275369
rect 401138 275295 401194 275304
rect 400772 269272 400824 269278
rect 400772 269214 400824 269220
rect 400312 265328 400364 265334
rect 400312 265270 400364 265276
rect 400220 265260 400272 265266
rect 400220 265202 400272 265208
rect 400324 264316 400352 265270
rect 400784 264316 400812 269214
rect 401152 264316 401180 275295
rect 401520 271998 401548 278052
rect 401966 275088 402022 275097
rect 401966 275023 402022 275032
rect 401600 274984 401652 274990
rect 401600 274926 401652 274932
rect 401612 273562 401640 274926
rect 401692 274848 401744 274854
rect 401692 274790 401744 274796
rect 401600 273556 401652 273562
rect 401600 273498 401652 273504
rect 401704 273290 401732 274790
rect 401692 273284 401744 273290
rect 401692 273226 401744 273232
rect 401508 271992 401560 271998
rect 401508 271934 401560 271940
rect 401600 269136 401652 269142
rect 401600 269078 401652 269084
rect 401612 268122 401640 269078
rect 401600 268116 401652 268122
rect 401600 268058 401652 268064
rect 401980 264330 402008 275023
rect 402518 274952 402574 274961
rect 402518 274887 402574 274896
rect 402060 270768 402112 270774
rect 402060 270710 402112 270716
rect 401626 264302 402008 264330
rect 402072 264316 402100 270710
rect 402532 264316 402560 274887
rect 402716 269210 402744 278052
rect 403912 274786 403940 278052
rect 405108 276078 405136 278052
rect 405096 276072 405148 276078
rect 405096 276014 405148 276020
rect 405372 274916 405424 274922
rect 405372 274858 405424 274864
rect 405186 274816 405242 274825
rect 403900 274780 403952 274786
rect 403900 274722 403952 274728
rect 404268 274780 404320 274786
rect 405186 274751 405242 274760
rect 404268 274722 404320 274728
rect 403438 269376 403494 269385
rect 403438 269311 403494 269320
rect 402704 269204 402756 269210
rect 402704 269146 402756 269152
rect 402978 267608 403034 267617
rect 402978 267543 403034 267552
rect 402992 264316 403020 267543
rect 403452 264316 403480 269311
rect 403900 269136 403952 269142
rect 403900 269078 403952 269084
rect 403912 264316 403940 269078
rect 404280 264316 404308 274722
rect 404726 272096 404782 272105
rect 404726 272031 404782 272040
rect 404740 264316 404768 272031
rect 405200 264316 405228 274751
rect 405384 269142 405412 274858
rect 406304 271930 406332 278052
rect 407500 274718 407528 278052
rect 407488 274712 407540 274718
rect 407488 274654 407540 274660
rect 408314 274680 408370 274689
rect 408314 274615 408370 274624
rect 407854 274544 407910 274553
rect 407854 274479 407910 274488
rect 406568 273488 406620 273494
rect 406568 273430 406620 273436
rect 406292 271924 406344 271930
rect 406292 271866 406344 271872
rect 406106 269240 406162 269249
rect 406106 269175 406162 269184
rect 405372 269136 405424 269142
rect 405372 269078 405424 269084
rect 405646 267744 405702 267753
rect 405646 267679 405702 267688
rect 405660 264316 405688 267679
rect 406120 264316 406148 269175
rect 406580 264316 406608 273430
rect 407396 271992 407448 271998
rect 407396 271934 407448 271940
rect 406934 267336 406990 267345
rect 406934 267271 406990 267280
rect 406948 264316 406976 267271
rect 407408 264316 407436 271934
rect 407868 264316 407896 274479
rect 408328 264316 408356 274615
rect 408604 265402 408632 278052
rect 409236 274712 409288 274718
rect 409236 274654 409288 274660
rect 408776 269204 408828 269210
rect 408776 269146 408828 269152
rect 408592 265396 408644 265402
rect 408592 265338 408644 265344
rect 408788 264316 408816 269146
rect 409248 264316 409276 274654
rect 409800 267986 409828 278052
rect 410996 274650 411024 278052
rect 410984 274644 411036 274650
rect 410984 274586 411036 274592
rect 410522 271960 410578 271969
rect 410522 271895 410578 271904
rect 411444 271924 411496 271930
rect 410062 271824 410118 271833
rect 410062 271759 410118 271768
rect 409788 267980 409840 267986
rect 409788 267922 409840 267928
rect 409604 265396 409656 265402
rect 409604 265338 409656 265344
rect 409616 264316 409644 265338
rect 410076 264316 410104 271759
rect 410536 264316 410564 271895
rect 411444 271866 411496 271872
rect 410982 269104 411038 269113
rect 410982 269039 411038 269048
rect 410996 264316 411024 269039
rect 411456 264316 411484 271866
rect 411904 269136 411956 269142
rect 411904 269078 411956 269084
rect 411916 264316 411944 269078
rect 412192 268122 412220 278052
rect 413388 271862 413416 278052
rect 414584 273630 414612 278052
rect 414572 273624 414624 273630
rect 414572 273566 414624 273572
rect 413652 271992 413704 271998
rect 413652 271934 413704 271940
rect 413376 271856 413428 271862
rect 413376 271798 413428 271804
rect 413664 270774 413692 271934
rect 415780 270842 415808 278052
rect 415768 270836 415820 270842
rect 415768 270778 415820 270784
rect 413652 270768 413704 270774
rect 413652 270710 413704 270716
rect 412180 268116 412232 268122
rect 412180 268058 412232 268064
rect 416884 268054 416912 278052
rect 418080 273766 418108 278052
rect 418068 273760 418120 273766
rect 418068 273702 418120 273708
rect 416872 268048 416924 268054
rect 416872 267990 416924 267996
rect 419276 265470 419304 278052
rect 420472 270910 420500 278052
rect 421668 273698 421696 278052
rect 421656 273692 421708 273698
rect 421656 273634 421708 273640
rect 420460 270904 420512 270910
rect 420460 270846 420512 270852
rect 422864 265538 422892 278052
rect 423968 268190 423996 278052
rect 425164 273834 425192 278052
rect 425152 273828 425204 273834
rect 425152 273770 425204 273776
rect 426360 268258 426388 278052
rect 427556 270978 427584 278052
rect 428752 273902 428780 278052
rect 429108 274712 429160 274718
rect 429108 274654 429160 274660
rect 428740 273896 428792 273902
rect 428740 273838 428792 273844
rect 429120 273562 429148 274654
rect 429108 273556 429160 273562
rect 429108 273498 429160 273504
rect 429948 271046 429976 278052
rect 429936 271040 429988 271046
rect 429936 270982 429988 270988
rect 427544 270972 427596 270978
rect 427544 270914 427596 270920
rect 431144 268326 431172 278052
rect 432248 273970 432276 278052
rect 432236 273964 432288 273970
rect 432236 273906 432288 273912
rect 433444 268394 433472 278052
rect 434640 272134 434668 278052
rect 435836 274038 435864 278052
rect 435824 274032 435876 274038
rect 435824 273974 435876 273980
rect 434628 272128 434680 272134
rect 434628 272070 434680 272076
rect 435732 272128 435784 272134
rect 435732 272070 435784 272076
rect 433432 268388 433484 268394
rect 433432 268330 433484 268336
rect 431132 268320 431184 268326
rect 431132 268262 431184 268268
rect 426348 268252 426400 268258
rect 426348 268194 426400 268200
rect 423956 268184 424008 268190
rect 423956 268126 424008 268132
rect 422852 265532 422904 265538
rect 422852 265474 422904 265480
rect 419264 265464 419316 265470
rect 419264 265406 419316 265412
rect 435744 265402 435772 272070
rect 437032 271114 437060 278052
rect 437020 271108 437072 271114
rect 437020 271050 437072 271056
rect 438228 268462 438256 278052
rect 439332 274106 439360 278052
rect 439320 274100 439372 274106
rect 439320 274042 439372 274048
rect 440528 268530 440556 278052
rect 441724 272474 441752 278052
rect 442920 274174 442948 278052
rect 442908 274168 442960 274174
rect 442908 274110 442960 274116
rect 441712 272468 441764 272474
rect 441712 272410 441764 272416
rect 441804 272468 441856 272474
rect 441804 272410 441856 272416
rect 440516 268524 440568 268530
rect 440516 268466 440568 268472
rect 438216 268456 438268 268462
rect 438216 268398 438268 268404
rect 441816 267753 441844 272410
rect 444116 271182 444144 278052
rect 444104 271176 444156 271182
rect 444104 271118 444156 271124
rect 445312 268598 445340 278052
rect 446508 274242 446536 278052
rect 446496 274236 446548 274242
rect 446496 274178 446548 274184
rect 447612 268666 447640 278052
rect 448808 271318 448836 278052
rect 450004 274310 450032 278052
rect 449992 274304 450044 274310
rect 449992 274246 450044 274252
rect 448796 271312 448848 271318
rect 448796 271254 448848 271260
rect 451200 271250 451228 278052
rect 451188 271244 451240 271250
rect 451188 271186 451240 271192
rect 452396 268734 452424 278052
rect 452384 268728 452436 268734
rect 452384 268670 452436 268676
rect 447600 268660 447652 268666
rect 447600 268602 447652 268608
rect 445300 268592 445352 268598
rect 445300 268534 445352 268540
rect 441802 267744 441858 267753
rect 441802 267679 441858 267688
rect 453592 265674 453620 278052
rect 454696 268802 454724 278052
rect 455892 272746 455920 278052
rect 457088 274378 457116 278052
rect 457076 274372 457128 274378
rect 457076 274314 457128 274320
rect 455880 272740 455932 272746
rect 455880 272682 455932 272688
rect 455972 272740 456024 272746
rect 455972 272682 456024 272688
rect 454684 268796 454736 268802
rect 454684 268738 454736 268744
rect 455984 267617 456012 272682
rect 458284 271386 458312 278052
rect 458272 271380 458324 271386
rect 458272 271322 458324 271328
rect 459480 268870 459508 278052
rect 459468 268864 459520 268870
rect 459468 268806 459520 268812
rect 455970 267608 456026 267617
rect 455970 267543 456026 267552
rect 460676 265742 460704 278052
rect 461872 268938 461900 278052
rect 462976 271454 463004 278052
rect 464172 274446 464200 278052
rect 464160 274440 464212 274446
rect 464160 274382 464212 274388
rect 465368 273086 465396 278052
rect 465356 273080 465408 273086
rect 465356 273022 465408 273028
rect 462964 271448 463016 271454
rect 462964 271390 463016 271396
rect 466564 269074 466592 278052
rect 467760 274582 467788 278052
rect 467748 274576 467800 274582
rect 467748 274518 467800 274524
rect 467748 273080 467800 273086
rect 467748 273022 467800 273028
rect 466552 269068 466604 269074
rect 466552 269010 466604 269016
rect 461860 268932 461912 268938
rect 461860 268874 461912 268880
rect 460664 265736 460716 265742
rect 460664 265678 460716 265684
rect 453580 265668 453632 265674
rect 453580 265610 453632 265616
rect 435732 265396 435784 265402
rect 435732 265338 435784 265344
rect 467760 265334 467788 273022
rect 468956 269006 468984 278052
rect 470152 271522 470180 278052
rect 471256 274514 471284 278052
rect 471244 274508 471296 274514
rect 471244 274450 471296 274456
rect 472452 273222 472480 278052
rect 472440 273216 472492 273222
rect 472440 273158 472492 273164
rect 472532 273216 472584 273222
rect 472532 273158 472584 273164
rect 470140 271516 470192 271522
rect 470140 271458 470192 271464
rect 468944 269000 468996 269006
rect 468944 268942 468996 268948
rect 472544 267481 472572 273158
rect 473648 270502 473676 278052
rect 473636 270496 473688 270502
rect 473636 270438 473688 270444
rect 472530 267472 472586 267481
rect 472530 267407 472586 267416
rect 474844 265810 474872 278052
rect 476040 270434 476068 278052
rect 477236 271590 477264 278052
rect 478340 276010 478368 278052
rect 478328 276004 478380 276010
rect 478328 275946 478380 275952
rect 479536 271658 479564 278052
rect 479524 271652 479576 271658
rect 479524 271594 479576 271600
rect 477224 271584 477276 271590
rect 477224 271526 477276 271532
rect 476028 270428 476080 270434
rect 476028 270370 476080 270376
rect 480732 270366 480760 278052
rect 480720 270360 480772 270366
rect 480720 270302 480772 270308
rect 481928 265878 481956 278052
rect 483124 270298 483152 278052
rect 484320 272950 484348 278052
rect 485516 275942 485544 278052
rect 485504 275936 485556 275942
rect 485504 275878 485556 275884
rect 484308 272944 484360 272950
rect 484308 272886 484360 272892
rect 485044 272944 485096 272950
rect 485044 272886 485096 272892
rect 483112 270292 483164 270298
rect 483112 270234 483164 270240
rect 485056 267345 485084 272886
rect 486620 271726 486648 278052
rect 486608 271720 486660 271726
rect 486608 271662 486660 271668
rect 487816 270230 487844 278052
rect 487804 270224 487856 270230
rect 487804 270166 487856 270172
rect 485042 267336 485098 267345
rect 485042 267271 485098 267280
rect 489012 265946 489040 278052
rect 490208 268433 490236 278052
rect 491404 271153 491432 278052
rect 492600 275874 492628 278052
rect 492588 275868 492640 275874
rect 492588 275810 492640 275816
rect 493704 271794 493732 278052
rect 493692 271788 493744 271794
rect 493692 271730 493744 271736
rect 491390 271144 491446 271153
rect 491390 271079 491446 271088
rect 494900 268569 494928 278052
rect 494886 268560 494942 268569
rect 494886 268495 494942 268504
rect 490194 268424 490250 268433
rect 490194 268359 490250 268368
rect 496096 266014 496124 278052
rect 497292 268705 497320 278052
rect 498488 271289 498516 278052
rect 499684 275806 499712 278052
rect 499672 275800 499724 275806
rect 499672 275742 499724 275748
rect 500880 273154 500908 278052
rect 500868 273148 500920 273154
rect 500868 273090 500920 273096
rect 498660 271788 498712 271794
rect 498660 271730 498712 271736
rect 498474 271280 498530 271289
rect 498474 271215 498530 271224
rect 497278 268696 497334 268705
rect 497278 268631 497334 268640
rect 496084 266008 496136 266014
rect 496084 265950 496136 265956
rect 489000 265940 489052 265946
rect 489000 265882 489052 265888
rect 481916 265872 481968 265878
rect 481916 265814 481968 265820
rect 474832 265804 474884 265810
rect 474832 265746 474884 265752
rect 498672 265606 498700 271730
rect 501984 268841 502012 278052
rect 501970 268832 502026 268841
rect 501970 268767 502026 268776
rect 503180 266082 503208 278052
rect 504376 268977 504404 278052
rect 505572 271425 505600 278052
rect 506768 275738 506796 278052
rect 506756 275732 506808 275738
rect 506756 275674 506808 275680
rect 507964 271561 507992 278052
rect 507950 271552 508006 271561
rect 507950 271487 508006 271496
rect 505558 271416 505614 271425
rect 505558 271351 505614 271360
rect 509068 270162 509096 278052
rect 509056 270156 509108 270162
rect 509056 270098 509108 270104
rect 504362 268968 504418 268977
rect 504362 268903 504418 268912
rect 510264 266150 510292 278052
rect 511460 270094 511488 278052
rect 512656 271697 512684 278052
rect 513852 275670 513880 278052
rect 513840 275664 513892 275670
rect 513840 275606 513892 275612
rect 515048 273018 515076 278052
rect 515036 273012 515088 273018
rect 515036 272954 515088 272960
rect 512642 271688 512698 271697
rect 512642 271623 512698 271632
rect 516244 270337 516272 278052
rect 516230 270328 516286 270337
rect 516230 270263 516286 270272
rect 511448 270088 511500 270094
rect 511448 270030 511500 270036
rect 517348 266218 517376 278052
rect 518544 270473 518572 278052
rect 519740 272814 519768 278052
rect 520936 275602 520964 278052
rect 520924 275596 520976 275602
rect 520924 275538 520976 275544
rect 522132 273193 522160 278052
rect 522118 273184 522174 273193
rect 522118 273119 522174 273128
rect 519728 272808 519780 272814
rect 519728 272750 519780 272756
rect 518530 270464 518586 270473
rect 518530 270399 518586 270408
rect 523328 270026 523356 278052
rect 523316 270020 523368 270026
rect 523316 269962 523368 269968
rect 524524 266286 524552 278052
rect 525628 270201 525656 278052
rect 526824 272882 526852 278052
rect 528020 275534 528048 278052
rect 528008 275528 528060 275534
rect 528008 275470 528060 275476
rect 529216 273057 529244 278052
rect 529202 273048 529258 273057
rect 529202 272983 529258 272992
rect 526812 272876 526864 272882
rect 526812 272818 526864 272824
rect 525614 270192 525670 270201
rect 525614 270127 525670 270136
rect 530412 269958 530440 278052
rect 530400 269952 530452 269958
rect 530400 269894 530452 269900
rect 531608 267714 531636 278052
rect 532712 269890 532740 278052
rect 533908 272921 533936 278052
rect 535104 275466 535132 278052
rect 535092 275460 535144 275466
rect 535092 275402 535144 275408
rect 533894 272912 533950 272921
rect 533894 272847 533950 272856
rect 536300 272785 536328 278052
rect 536286 272776 536342 272785
rect 536286 272711 536342 272720
rect 537496 270065 537524 278052
rect 537482 270056 537538 270065
rect 537482 269991 537538 270000
rect 532700 269884 532752 269890
rect 532700 269826 532752 269832
rect 531596 267708 531648 267714
rect 531596 267650 531648 267656
rect 538692 267646 538720 278052
rect 539888 269929 539916 278052
rect 540992 272649 541020 278052
rect 542188 275398 542216 278052
rect 542176 275392 542228 275398
rect 542176 275334 542228 275340
rect 540978 272640 541034 272649
rect 540978 272575 541034 272584
rect 543384 272513 543412 278052
rect 543370 272504 543426 272513
rect 543370 272439 543426 272448
rect 539874 269920 539930 269929
rect 539874 269855 539930 269864
rect 544580 269822 544608 278052
rect 544568 269816 544620 269822
rect 544568 269758 544620 269764
rect 538680 267640 538732 267646
rect 538680 267582 538732 267588
rect 545776 267578 545804 278052
rect 545764 267572 545816 267578
rect 545764 267514 545816 267520
rect 546972 267510 547000 278052
rect 548076 269754 548104 278052
rect 548064 269748 548116 269754
rect 548064 269690 548116 269696
rect 546960 267504 547012 267510
rect 546960 267446 547012 267452
rect 549272 267442 549300 278052
rect 550468 275330 550496 278052
rect 550456 275324 550508 275330
rect 550456 275266 550508 275272
rect 551664 272678 551692 278052
rect 551652 272672 551704 272678
rect 551652 272614 551704 272620
rect 549260 267436 549312 267442
rect 549260 267378 549312 267384
rect 552860 267306 552888 278052
rect 554056 267374 554084 278052
rect 555252 269793 555280 278052
rect 555238 269784 555294 269793
rect 555238 269719 555294 269728
rect 554044 267368 554096 267374
rect 554044 267310 554096 267316
rect 552848 267300 552900 267306
rect 552848 267242 552900 267248
rect 556356 267238 556384 278052
rect 557552 275262 557580 278052
rect 557540 275256 557592 275262
rect 557540 275198 557592 275204
rect 558748 272610 558776 278052
rect 558736 272604 558788 272610
rect 558736 272546 558788 272552
rect 556344 267232 556396 267238
rect 556344 267174 556396 267180
rect 559944 267170 559972 278052
rect 559932 267164 559984 267170
rect 559932 267106 559984 267112
rect 561140 267102 561168 278052
rect 562336 269686 562364 278052
rect 562324 269680 562376 269686
rect 562324 269622 562376 269628
rect 561128 267096 561180 267102
rect 561128 267038 561180 267044
rect 563440 267034 563468 278052
rect 564636 275194 564664 278052
rect 564624 275188 564676 275194
rect 564624 275130 564676 275136
rect 565832 272377 565860 278052
rect 565818 272368 565874 272377
rect 565818 272303 565874 272312
rect 563428 267028 563480 267034
rect 563428 266970 563480 266976
rect 567028 266898 567056 278052
rect 568224 266966 568252 278052
rect 569420 269657 569448 278052
rect 569406 269648 569462 269657
rect 569406 269583 569462 269592
rect 568212 266960 568264 266966
rect 568212 266902 568264 266908
rect 567016 266892 567068 266898
rect 567016 266834 567068 266840
rect 570616 266830 570644 278052
rect 571720 275126 571748 278052
rect 571708 275120 571760 275126
rect 571708 275062 571760 275068
rect 572916 272542 572944 278052
rect 572904 272536 572956 272542
rect 572904 272478 572956 272484
rect 570604 266824 570656 266830
rect 570604 266766 570656 266772
rect 574112 266694 574140 278052
rect 575308 266762 575336 278052
rect 576504 269618 576532 278052
rect 576492 269612 576544 269618
rect 576492 269554 576544 269560
rect 575296 266756 575348 266762
rect 575296 266698 575348 266704
rect 574100 266688 574152 266694
rect 574100 266630 574152 266636
rect 577700 266626 577728 278052
rect 578896 275058 578924 278052
rect 578884 275052 578936 275058
rect 578884 274994 578936 275000
rect 580000 272406 580028 278052
rect 579988 272400 580040 272406
rect 579988 272342 580040 272348
rect 577688 266620 577740 266626
rect 577688 266562 577740 266568
rect 581196 266558 581224 278052
rect 582392 267209 582420 278052
rect 583588 269550 583616 278052
rect 583576 269544 583628 269550
rect 583576 269486 583628 269492
rect 582378 267200 582434 267209
rect 582378 267135 582434 267144
rect 581184 266552 581236 266558
rect 581184 266494 581236 266500
rect 584784 266490 584812 278052
rect 585980 274990 586008 278052
rect 585968 274984 586020 274990
rect 585968 274926 586020 274932
rect 587084 272338 587112 278052
rect 587072 272332 587124 272338
rect 587072 272274 587124 272280
rect 584772 266484 584824 266490
rect 584772 266426 584824 266432
rect 588280 266422 588308 278052
rect 589476 267073 589504 278052
rect 590672 272270 590700 278052
rect 590660 272264 590712 272270
rect 590660 272206 590712 272212
rect 589462 267064 589518 267073
rect 589462 266999 589518 267008
rect 591868 266937 591896 278052
rect 593064 274854 593092 278052
rect 593052 274848 593104 274854
rect 593052 274790 593104 274796
rect 594260 269521 594288 278052
rect 594246 269512 594302 269521
rect 594246 269447 594302 269456
rect 591854 266928 591910 266937
rect 591854 266863 591910 266872
rect 595364 266801 595392 278052
rect 595350 266792 595406 266801
rect 595350 266727 595406 266736
rect 588268 266416 588320 266422
rect 588268 266358 588320 266364
rect 596560 266354 596588 278052
rect 597756 269482 597784 278052
rect 597744 269476 597796 269482
rect 597744 269418 597796 269424
rect 598952 266665 598980 278052
rect 600148 274281 600176 278052
rect 600134 274272 600190 274281
rect 600134 274207 600190 274216
rect 601344 272202 601372 278052
rect 601332 272196 601384 272202
rect 601332 272138 601384 272144
rect 598938 266656 598994 266665
rect 598938 266591 598994 266600
rect 602448 266529 602476 278052
rect 603644 271794 603672 278052
rect 604840 272241 604868 278052
rect 606036 274417 606064 278052
rect 607232 275777 607260 278052
rect 607218 275768 607274 275777
rect 607218 275703 607274 275712
rect 606022 274408 606078 274417
rect 606022 274343 606078 274352
rect 604826 272232 604882 272241
rect 604826 272167 604882 272176
rect 603632 271788 603684 271794
rect 603632 271730 603684 271736
rect 608428 269414 608456 278052
rect 609624 275913 609652 278052
rect 609610 275904 609666 275913
rect 609610 275839 609666 275848
rect 610728 273222 610756 278052
rect 610716 273216 610768 273222
rect 610716 273158 610768 273164
rect 611924 272066 611952 278052
rect 613120 275505 613148 278052
rect 614316 275641 614344 278052
rect 614302 275632 614358 275641
rect 614302 275567 614358 275576
rect 613106 275496 613162 275505
rect 613106 275431 613162 275440
rect 611912 272060 611964 272066
rect 611912 272002 611964 272008
rect 608416 269408 608468 269414
rect 608416 269350 608468 269356
rect 615512 269346 615540 278052
rect 616708 275233 616736 278052
rect 616694 275224 616750 275233
rect 616694 275159 616750 275168
rect 617812 273086 617840 278052
rect 617800 273080 617852 273086
rect 617800 273022 617852 273028
rect 615500 269340 615552 269346
rect 615500 269282 615552 269288
rect 619008 269278 619036 278052
rect 620204 275369 620232 278052
rect 620190 275360 620246 275369
rect 620190 275295 620246 275304
rect 621400 275097 621428 278052
rect 621386 275088 621442 275097
rect 621386 275023 621442 275032
rect 622596 271998 622624 278052
rect 623792 274961 623820 278052
rect 623778 274952 623834 274961
rect 623778 274887 623834 274896
rect 624988 272746 625016 278052
rect 624976 272740 625028 272746
rect 624976 272682 625028 272688
rect 622584 271992 622636 271998
rect 622584 271934 622636 271940
rect 626092 269385 626120 278052
rect 627288 274922 627316 278052
rect 627276 274916 627328 274922
rect 627276 274858 627328 274864
rect 628484 274786 628512 278052
rect 628472 274780 628524 274786
rect 628472 274722 628524 274728
rect 629680 272105 629708 278052
rect 630876 274825 630904 278052
rect 630862 274816 630918 274825
rect 630862 274751 630918 274760
rect 632072 272474 632100 278052
rect 632060 272468 632112 272474
rect 632060 272410 632112 272416
rect 629666 272096 629722 272105
rect 629666 272031 629722 272040
rect 626078 269376 626134 269385
rect 626078 269311 626134 269320
rect 618996 269272 619048 269278
rect 633268 269249 633296 278052
rect 634372 274718 634400 278052
rect 634360 274712 634412 274718
rect 634360 274654 634412 274660
rect 635568 272950 635596 278052
rect 635556 272944 635608 272950
rect 635556 272886 635608 272892
rect 636764 271930 636792 278052
rect 637960 274553 637988 278052
rect 639156 274689 639184 278052
rect 639142 274680 639198 274689
rect 639142 274615 639198 274624
rect 637946 274544 638002 274553
rect 637946 274479 638002 274488
rect 636752 271924 636804 271930
rect 636752 271866 636804 271872
rect 618996 269214 619048 269220
rect 633254 269240 633310 269249
rect 640352 269210 640380 278052
rect 641456 274650 641484 278052
rect 641444 274644 641496 274650
rect 641444 274586 641496 274592
rect 642652 272134 642680 278052
rect 642640 272128 642692 272134
rect 642640 272070 642692 272076
rect 643848 271833 643876 278052
rect 645044 271969 645072 278052
rect 645030 271960 645086 271969
rect 645030 271895 645086 271904
rect 643834 271824 643890 271833
rect 643834 271759 643890 271768
rect 633254 269175 633310 269184
rect 640340 269204 640392 269210
rect 640340 269146 640392 269152
rect 646240 269113 646268 278052
rect 647436 271862 647464 278052
rect 648646 278038 648752 278066
rect 648620 277636 648672 277642
rect 648620 277578 648672 277584
rect 647424 271856 647476 271862
rect 647424 271798 647476 271804
rect 646226 269104 646282 269113
rect 646226 269039 646282 269048
rect 602434 266520 602490 266529
rect 602434 266455 602490 266464
rect 596548 266348 596600 266354
rect 596548 266290 596600 266296
rect 524512 266280 524564 266286
rect 524512 266222 524564 266228
rect 517336 266212 517388 266218
rect 517336 266154 517388 266160
rect 510252 266144 510304 266150
rect 510252 266086 510304 266092
rect 503168 266076 503220 266082
rect 503168 266018 503220 266024
rect 498660 265600 498712 265606
rect 498660 265542 498712 265548
rect 467748 265328 467800 265334
rect 467748 265270 467800 265276
rect 184938 258632 184994 258641
rect 184938 258567 184994 258576
rect 184952 256766 184980 258567
rect 184940 256760 184992 256766
rect 184940 256702 184992 256708
rect 416778 252784 416834 252793
rect 416778 252719 416834 252728
rect 416792 251258 416820 252719
rect 416780 251252 416832 251258
rect 416780 251194 416832 251200
rect 567108 251252 567160 251258
rect 567108 251194 567160 251200
rect 416778 249520 416834 249529
rect 416778 249455 416834 249464
rect 416792 248470 416820 249455
rect 416780 248464 416832 248470
rect 416780 248406 416832 248412
rect 564348 248464 564400 248470
rect 564348 248406 564400 248412
rect 184938 248024 184994 248033
rect 184938 247959 184994 247968
rect 184952 245818 184980 247959
rect 416778 246392 416834 246401
rect 416778 246327 416834 246336
rect 184940 245812 184992 245818
rect 184940 245754 184992 245760
rect 416792 245682 416820 246327
rect 416780 245676 416832 245682
rect 416780 245618 416832 245624
rect 418066 243128 418122 243137
rect 418066 243063 418122 243072
rect 184940 237448 184992 237454
rect 184938 237416 184940 237425
rect 184992 237416 184994 237425
rect 184938 237351 184994 237360
rect 158720 229084 158772 229090
rect 158720 229026 158772 229032
rect 152832 229016 152884 229022
rect 84658 228984 84714 228993
rect 152832 228958 152884 228964
rect 84658 228919 84714 228928
rect 82726 228576 82782 228585
rect 82726 228511 82782 228520
rect 77942 228440 77998 228449
rect 77942 228375 77998 228384
rect 76286 228304 76342 228313
rect 76286 228239 76342 228248
rect 71226 228168 71282 228177
rect 71226 228103 71282 228112
rect 64510 228032 64566 228041
rect 64510 227967 64566 227976
rect 64524 217410 64552 227967
rect 69480 227860 69532 227866
rect 69480 227802 69532 227808
rect 65340 227792 65392 227798
rect 65340 227734 65392 227740
rect 65352 217410 65380 227734
rect 66996 222828 67048 222834
rect 66996 222770 67048 222776
rect 66166 222728 66222 222737
rect 66166 222663 66222 222672
rect 66180 217410 66208 222663
rect 67008 217410 67036 222770
rect 67822 222592 67878 222601
rect 67822 222527 67878 222536
rect 67836 217410 67864 222527
rect 68652 222352 68704 222358
rect 68652 222294 68704 222300
rect 68664 217410 68692 222294
rect 69492 217410 69520 227802
rect 70398 225312 70454 225321
rect 70398 225247 70454 225256
rect 70412 217410 70440 225247
rect 71240 217410 71268 228103
rect 72056 227996 72108 228002
rect 72056 227938 72108 227944
rect 72068 217410 72096 227938
rect 73712 225072 73764 225078
rect 73712 225014 73764 225020
rect 72882 223000 72938 223009
rect 72882 222935 72938 222944
rect 72896 217410 72924 222935
rect 73724 217410 73752 225014
rect 74446 222864 74502 222873
rect 74446 222799 74502 222808
rect 74460 217410 74488 222799
rect 75368 222420 75420 222426
rect 75368 222362 75420 222368
rect 75380 217410 75408 222362
rect 76300 217410 76328 228239
rect 77114 225448 77170 225457
rect 77114 225383 77170 225392
rect 77128 217410 77156 225383
rect 77956 217410 77984 228375
rect 78772 227928 78824 227934
rect 78772 227870 78824 227876
rect 78784 217410 78812 227870
rect 80426 225584 80482 225593
rect 80426 225519 80482 225528
rect 79598 223136 79654 223145
rect 79598 223071 79654 223080
rect 79612 217410 79640 223071
rect 80440 217410 80468 225519
rect 82176 222624 82228 222630
rect 82176 222566 82228 222572
rect 81256 222488 81308 222494
rect 81256 222430 81308 222436
rect 81268 217410 81296 222430
rect 82188 217410 82216 222566
rect 82740 217410 82768 228511
rect 83830 225720 83886 225729
rect 83830 225655 83886 225664
rect 83844 217410 83872 225655
rect 84672 217410 84700 228919
rect 150256 228880 150308 228886
rect 88062 228848 88118 228857
rect 150256 228822 150308 228828
rect 88062 228783 88118 228792
rect 86314 228712 86370 228721
rect 86314 228647 86370 228656
rect 85488 222556 85540 222562
rect 85488 222498 85540 222504
rect 85500 217410 85528 222498
rect 86328 217410 86356 228647
rect 87144 223304 87196 223310
rect 87144 223246 87196 223252
rect 87156 217410 87184 223246
rect 88076 217410 88104 228783
rect 146024 228744 146076 228750
rect 146024 228686 146076 228692
rect 138480 228676 138532 228682
rect 138480 228618 138532 228624
rect 136824 228472 136876 228478
rect 136824 228414 136876 228420
rect 131764 228404 131816 228410
rect 131764 228346 131816 228352
rect 125048 228336 125100 228342
rect 125048 228278 125100 228284
rect 123392 228200 123444 228206
rect 123392 228142 123444 228148
rect 114928 228132 114980 228138
rect 114928 228074 114980 228080
rect 108212 228064 108264 228070
rect 108212 228006 108264 228012
rect 93030 227488 93086 227497
rect 93030 227423 93086 227432
rect 88892 225208 88944 225214
rect 88892 225150 88944 225156
rect 88904 217410 88932 225150
rect 92204 225140 92256 225146
rect 92204 225082 92256 225088
rect 91376 222760 91428 222766
rect 91376 222702 91428 222708
rect 89720 222692 89772 222698
rect 89720 222634 89772 222640
rect 89732 217410 89760 222634
rect 90548 222012 90600 222018
rect 90548 221954 90600 221960
rect 90560 217410 90588 221954
rect 91388 217410 91416 222702
rect 92216 217410 92244 225082
rect 93044 217410 93072 227423
rect 94778 227352 94834 227361
rect 94778 227287 94834 227296
rect 93768 223508 93820 223514
rect 93768 223450 93820 223456
rect 93780 217410 93808 223450
rect 94792 217410 94820 227287
rect 101494 227216 101550 227225
rect 101494 227151 101550 227160
rect 99838 227080 99894 227089
rect 99838 227015 99894 227024
rect 98918 225992 98974 226001
rect 98918 225927 98974 225936
rect 97264 225344 97316 225350
rect 97264 225286 97316 225292
rect 95608 225276 95660 225282
rect 95608 225218 95660 225224
rect 95620 217410 95648 225218
rect 96434 223272 96490 223281
rect 96434 223207 96490 223216
rect 96448 217410 96476 223207
rect 97276 217410 97304 225286
rect 98090 223408 98146 223417
rect 98090 223343 98146 223352
rect 98104 217410 98132 223343
rect 98932 217410 98960 225927
rect 99852 217410 99880 227015
rect 100668 225412 100720 225418
rect 100668 225354 100720 225360
rect 100680 217410 100708 225354
rect 101508 217410 101536 227151
rect 106554 226944 106610 226953
rect 106554 226879 106610 226888
rect 103978 226128 104034 226137
rect 103978 226063 104034 226072
rect 102046 225856 102102 225865
rect 102046 225791 102102 225800
rect 102060 217410 102088 225791
rect 103150 223544 103206 223553
rect 103150 223479 103206 223488
rect 103164 217410 103192 223479
rect 103992 217410 104020 226063
rect 105728 225548 105780 225554
rect 105728 225490 105780 225496
rect 104806 222048 104862 222057
rect 104806 221983 104862 221992
rect 104820 217410 104848 221983
rect 105740 217410 105768 225490
rect 106568 217410 106596 226879
rect 107384 225480 107436 225486
rect 107384 225422 107436 225428
rect 107396 217410 107424 225422
rect 108224 217410 108252 228006
rect 113086 226808 113142 226817
rect 113086 226743 113142 226752
rect 109038 226264 109094 226273
rect 109038 226199 109094 226208
rect 109052 217410 109080 226199
rect 110696 225616 110748 225622
rect 110696 225558 110748 225564
rect 109866 221912 109922 221921
rect 109866 221847 109922 221856
rect 109880 217410 109908 221847
rect 110708 217410 110736 225558
rect 112442 224768 112498 224777
rect 112442 224703 112498 224712
rect 111614 221776 111670 221785
rect 111614 221711 111670 221720
rect 111628 217410 111656 221711
rect 112456 217410 112484 224703
rect 113100 217410 113128 226743
rect 114100 225684 114152 225690
rect 114100 225626 114152 225632
rect 114112 217410 114140 225626
rect 114284 224868 114336 224874
rect 114284 224810 114336 224816
rect 114296 222834 114324 224810
rect 114284 222828 114336 222834
rect 114284 222770 114336 222776
rect 114940 217410 114968 228074
rect 119160 225820 119212 225826
rect 119160 225762 119212 225768
rect 115754 224632 115810 224641
rect 115754 224567 115810 224576
rect 115768 217410 115796 224567
rect 117502 224496 117558 224505
rect 117502 224431 117558 224440
rect 116584 222828 116636 222834
rect 116584 222770 116636 222776
rect 116596 217410 116624 222770
rect 117516 217410 117544 224431
rect 118330 221368 118386 221377
rect 118330 221303 118386 221312
rect 118344 217410 118372 221303
rect 119172 217410 119200 225762
rect 120814 224360 120870 224369
rect 120814 224295 120870 224304
rect 119986 221640 120042 221649
rect 119986 221575 120042 221584
rect 120000 217410 120028 221575
rect 120828 217410 120856 224295
rect 121366 221504 121422 221513
rect 121366 221439 121422 221448
rect 121380 217410 121408 221439
rect 122472 220108 122524 220114
rect 122472 220050 122524 220056
rect 122484 217410 122512 220050
rect 123404 217410 123432 228142
rect 124128 225752 124180 225758
rect 124128 225694 124180 225700
rect 124140 217410 124168 225694
rect 125060 217410 125088 228278
rect 130108 228268 130160 228274
rect 130108 228210 130160 228216
rect 127532 225888 127584 225894
rect 127532 225830 127584 225836
rect 126704 222896 126756 222902
rect 126704 222838 126756 222844
rect 125876 220176 125928 220182
rect 125876 220118 125928 220124
rect 125888 217410 125916 220118
rect 126716 217410 126744 222838
rect 127544 217410 127572 225830
rect 128360 222964 128412 222970
rect 128360 222906 128412 222912
rect 128372 217410 128400 222906
rect 129280 220244 129332 220250
rect 129280 220186 129332 220192
rect 129292 217410 129320 220186
rect 130120 217410 130148 228210
rect 130936 225956 130988 225962
rect 130936 225898 130988 225904
rect 130948 217410 130976 225898
rect 131776 217410 131804 228346
rect 134248 226024 134300 226030
rect 134248 225966 134300 225972
rect 133420 223032 133472 223038
rect 133420 222974 133472 222980
rect 132408 220312 132460 220318
rect 132408 220254 132460 220260
rect 132420 217410 132448 220254
rect 133432 217410 133460 222974
rect 134260 217410 134288 225966
rect 135168 223100 135220 223106
rect 135168 223042 135220 223048
rect 135180 217410 135208 223042
rect 135996 220380 136048 220386
rect 135996 220322 136048 220328
rect 136008 217410 136036 220322
rect 136836 217410 136864 228414
rect 137652 226092 137704 226098
rect 137652 226034 137704 226040
rect 137664 217410 137692 226034
rect 138492 217410 138520 228618
rect 143448 228608 143500 228614
rect 143448 228550 143500 228556
rect 141056 226160 141108 226166
rect 141056 226102 141108 226108
rect 140136 223168 140188 223174
rect 140136 223110 140188 223116
rect 139308 220448 139360 220454
rect 139308 220390 139360 220396
rect 139320 217410 139348 220390
rect 140148 217410 140176 223110
rect 141068 217410 141096 226102
rect 141884 223236 141936 223242
rect 141884 223178 141936 223184
rect 141896 217410 141924 223178
rect 142712 220516 142764 220522
rect 142712 220458 142764 220464
rect 142724 217410 142752 220458
rect 143460 217410 143488 228550
rect 145196 228540 145248 228546
rect 145196 228482 145248 228488
rect 144368 226296 144420 226302
rect 144368 226238 144420 226244
rect 144380 217410 144408 226238
rect 145208 217410 145236 228482
rect 146036 217410 146064 228686
rect 147772 226228 147824 226234
rect 147772 226170 147824 226176
rect 146300 224052 146352 224058
rect 146300 223994 146352 224000
rect 146312 223514 146340 223994
rect 146300 223508 146352 223514
rect 146300 223450 146352 223456
rect 146944 223440 146996 223446
rect 146944 223382 146996 223388
rect 146956 217410 146984 223382
rect 147784 217410 147812 226170
rect 148600 223372 148652 223378
rect 148600 223314 148652 223320
rect 148612 217410 148640 223314
rect 149428 221468 149480 221474
rect 149428 221410 149480 221416
rect 149440 217410 149468 221410
rect 150268 217410 150296 228822
rect 151728 228812 151780 228818
rect 151728 228754 151780 228760
rect 151084 224732 151136 224738
rect 151084 224674 151136 224680
rect 151096 217410 151124 224674
rect 151740 217410 151768 228754
rect 152844 217410 152872 228958
rect 156972 228948 157024 228954
rect 156972 228890 157024 228896
rect 156144 227656 156196 227662
rect 156144 227598 156196 227604
rect 154488 224800 154540 224806
rect 154488 224742 154540 224748
rect 153660 223508 153712 223514
rect 153660 223450 153712 223456
rect 153672 217410 153700 223450
rect 154500 217410 154528 224742
rect 155316 223576 155368 223582
rect 155316 223518 155368 223524
rect 155328 217410 155356 223518
rect 156156 217410 156184 227598
rect 156984 217410 157012 228890
rect 157800 224596 157852 224602
rect 157800 224538 157852 224544
rect 157812 217410 157840 224538
rect 158732 217410 158760 229026
rect 162768 227588 162820 227594
rect 162768 227530 162820 227536
rect 161204 224664 161256 224670
rect 161204 224606 161256 224612
rect 160098 224224 160154 224233
rect 160098 224159 160154 224168
rect 160112 222018 160140 224159
rect 160376 222080 160428 222086
rect 160376 222022 160428 222028
rect 160100 222012 160152 222018
rect 160100 221954 160152 221960
rect 159548 221536 159600 221542
rect 159548 221478 159600 221484
rect 159560 217410 159588 221478
rect 160388 217410 160416 222022
rect 161216 217410 161244 224606
rect 162032 222148 162084 222154
rect 162032 222090 162084 222096
rect 162044 217410 162072 222090
rect 162780 217410 162808 227530
rect 165436 227520 165488 227526
rect 165436 227462 165488 227468
rect 163688 227452 163740 227458
rect 163688 227394 163740 227400
rect 163700 217410 163728 227394
rect 164608 220856 164660 220862
rect 164608 220798 164660 220804
rect 164620 217410 164648 220798
rect 165448 217410 165476 227462
rect 167092 227384 167144 227390
rect 167092 227326 167144 227332
rect 166356 224460 166408 224466
rect 166356 224402 166408 224408
rect 166264 221332 166316 221338
rect 166264 221274 166316 221280
rect 166276 217410 166304 221274
rect 166368 220862 166396 224402
rect 166356 220856 166408 220862
rect 166356 220798 166408 220804
rect 167104 217410 167132 227326
rect 173624 227316 173676 227322
rect 173624 227258 173676 227264
rect 169576 227248 169628 227254
rect 169576 227190 169628 227196
rect 169116 224528 169168 224534
rect 169116 224470 169168 224476
rect 168748 221944 168800 221950
rect 168748 221886 168800 221892
rect 167920 220856 167972 220862
rect 167920 220798 167972 220804
rect 167932 217410 167960 220798
rect 168760 217410 168788 221886
rect 169128 220862 169156 224470
rect 169116 220856 169168 220862
rect 169116 220798 169168 220804
rect 169588 217410 169616 227190
rect 172152 227180 172204 227186
rect 172152 227122 172204 227128
rect 171048 224392 171100 224398
rect 171048 224334 171100 224340
rect 170496 222012 170548 222018
rect 170496 221954 170548 221960
rect 170508 217410 170536 221954
rect 171060 217410 171088 224334
rect 172164 217410 172192 227122
rect 172426 224088 172482 224097
rect 172426 224023 172482 224032
rect 172440 223310 172468 224023
rect 172428 223304 172480 223310
rect 172428 223246 172480 223252
rect 172980 221264 173032 221270
rect 172980 221206 173032 221212
rect 172992 217410 173020 221206
rect 173636 217410 173664 227258
rect 181904 227112 181956 227118
rect 181904 227054 181956 227060
rect 176384 227044 176436 227050
rect 176384 226986 176436 226992
rect 175464 223304 175516 223310
rect 175464 223246 175516 223252
rect 174636 220856 174688 220862
rect 174636 220798 174688 220804
rect 174648 217410 174676 220798
rect 175476 217410 175504 223246
rect 176396 217410 176424 226986
rect 180524 226976 180576 226982
rect 180524 226918 180576 226924
rect 176660 224324 176712 224330
rect 176660 224266 176712 224272
rect 176672 220862 176700 224266
rect 178040 224188 178092 224194
rect 178040 224130 178092 224136
rect 177212 221876 177264 221882
rect 177212 221818 177264 221824
rect 176660 220856 176712 220862
rect 176660 220798 176712 220804
rect 177224 217410 177252 221818
rect 178052 217410 178080 224130
rect 179696 221672 179748 221678
rect 179696 221614 179748 221620
rect 178868 221196 178920 221202
rect 178868 221138 178920 221144
rect 178880 217410 178908 221138
rect 179708 217410 179736 221614
rect 180536 217410 180564 226918
rect 181352 224256 181404 224262
rect 181352 224198 181404 224204
rect 181364 217410 181392 224198
rect 181916 221202 181944 227054
rect 190368 226908 190420 226914
rect 190368 226850 190420 226856
rect 189264 226840 189316 226846
rect 189264 226782 189316 226788
rect 186412 226772 186464 226778
rect 186412 226714 186464 226720
rect 183008 226364 183060 226370
rect 183008 226306 183060 226312
rect 183020 222290 183048 226306
rect 184756 224120 184808 224126
rect 184756 224062 184808 224068
rect 183008 222284 183060 222290
rect 183008 222226 183060 222232
rect 183928 221808 183980 221814
rect 183928 221750 183980 221756
rect 182088 221740 182140 221746
rect 182088 221682 182140 221688
rect 181904 221196 181956 221202
rect 181904 221138 181956 221144
rect 182100 217410 182128 221682
rect 183100 221128 183152 221134
rect 183100 221070 183152 221076
rect 183112 217410 183140 221070
rect 183940 217410 183968 221750
rect 184768 217410 184796 224062
rect 185584 223644 185636 223650
rect 185584 223586 185636 223592
rect 185596 217410 185624 223586
rect 186424 217410 186452 226714
rect 188160 223984 188212 223990
rect 188160 223926 188212 223932
rect 187240 222284 187292 222290
rect 187240 222226 187292 222232
rect 187252 217410 187280 222226
rect 188172 217410 188200 223926
rect 188436 223848 188488 223854
rect 188436 223790 188488 223796
rect 188448 221474 188476 223790
rect 189276 223650 189304 226782
rect 189264 223644 189316 223650
rect 189264 223586 189316 223592
rect 188436 221468 188488 221474
rect 188436 221410 188488 221416
rect 189816 221196 189868 221202
rect 189816 221138 189868 221144
rect 188988 221060 189040 221066
rect 188988 221002 189040 221008
rect 189000 217410 189028 221002
rect 189828 217410 189856 221138
rect 190380 217410 190408 226850
rect 192312 226370 192340 231676
rect 192300 226364 192352 226370
rect 192300 226306 192352 226312
rect 192588 224942 192616 231676
rect 192956 227730 192984 231676
rect 192944 227724 192996 227730
rect 192944 227666 192996 227672
rect 193036 226636 193088 226642
rect 193036 226578 193088 226584
rect 192760 225412 192812 225418
rect 192760 225354 192812 225360
rect 192772 225214 192800 225354
rect 192668 225208 192720 225214
rect 192668 225150 192720 225156
rect 192760 225208 192812 225214
rect 192760 225150 192812 225156
rect 192680 224942 192708 225150
rect 192576 224936 192628 224942
rect 192576 224878 192628 224884
rect 192668 224936 192720 224942
rect 192668 224878 192720 224884
rect 191472 223780 191524 223786
rect 191472 223722 191524 223728
rect 191484 217410 191512 223722
rect 193048 221406 193076 226578
rect 193324 222193 193352 231676
rect 193692 224913 193720 231676
rect 193772 227928 193824 227934
rect 193772 227870 193824 227876
rect 193784 226574 193812 227870
rect 193772 226568 193824 226574
rect 193772 226510 193824 226516
rect 194060 225049 194088 231676
rect 194428 227633 194456 231676
rect 194796 227769 194824 231676
rect 194782 227760 194838 227769
rect 194782 227695 194838 227704
rect 194414 227624 194470 227633
rect 194414 227559 194470 227568
rect 194046 225040 194102 225049
rect 195164 225010 195192 231676
rect 194046 224975 194102 224984
rect 195152 225004 195204 225010
rect 195152 224946 195204 224952
rect 195244 225004 195296 225010
rect 195244 224946 195296 224952
rect 193678 224904 193734 224913
rect 193678 224839 193734 224848
rect 193310 222184 193366 222193
rect 193310 222119 193366 222128
rect 194048 221604 194100 221610
rect 194048 221546 194100 221552
rect 192300 221400 192352 221406
rect 192300 221342 192352 221348
rect 193036 221400 193088 221406
rect 193036 221342 193088 221348
rect 193128 221400 193180 221406
rect 193128 221342 193180 221348
rect 192312 217410 192340 221342
rect 193140 217410 193168 221342
rect 194060 217410 194088 221546
rect 195256 217546 195284 224946
rect 195440 222222 195468 231676
rect 195808 222329 195836 231676
rect 195888 226704 195940 226710
rect 195888 226646 195940 226652
rect 195794 222320 195850 222329
rect 195794 222255 195850 222264
rect 195428 222216 195480 222222
rect 195428 222158 195480 222164
rect 195704 221468 195756 221474
rect 195704 221410 195756 221416
rect 194980 217518 195284 217546
rect 194980 217410 195008 217518
rect 195716 217410 195744 221410
rect 195900 221406 195928 226646
rect 196176 222465 196204 231676
rect 196544 225185 196572 231676
rect 196912 227798 196940 231676
rect 197280 227905 197308 231676
rect 197648 228041 197676 231676
rect 197634 228032 197690 228041
rect 197634 227967 197690 227976
rect 197266 227896 197322 227905
rect 197266 227831 197322 227840
rect 196900 227792 196952 227798
rect 196900 227734 196952 227740
rect 197360 227724 197412 227730
rect 197360 227666 197412 227672
rect 196530 225176 196586 225185
rect 196530 225111 196586 225120
rect 196162 222456 196218 222465
rect 196162 222391 196218 222400
rect 196072 221604 196124 221610
rect 196072 221546 196124 221552
rect 196164 221604 196216 221610
rect 196164 221546 196216 221552
rect 196084 221474 196112 221546
rect 196072 221468 196124 221474
rect 196072 221410 196124 221416
rect 195888 221400 195940 221406
rect 195888 221342 195940 221348
rect 196176 221066 196204 221546
rect 196164 221060 196216 221066
rect 196164 221002 196216 221008
rect 196532 220924 196584 220930
rect 196532 220866 196584 220872
rect 196544 217410 196572 220866
rect 197372 217410 197400 227666
rect 197452 225208 197504 225214
rect 197452 225150 197504 225156
rect 197464 224058 197492 225150
rect 198016 224874 198044 231676
rect 198004 224868 198056 224874
rect 198004 224810 198056 224816
rect 198188 224868 198240 224874
rect 198188 224810 198240 224816
rect 197452 224052 197504 224058
rect 197452 223994 197504 224000
rect 198200 217410 198228 224810
rect 198292 222358 198320 231676
rect 198660 222737 198688 231676
rect 198740 227860 198792 227866
rect 198740 227802 198792 227808
rect 198646 222728 198702 222737
rect 198646 222663 198702 222672
rect 198752 222630 198780 227802
rect 198924 227792 198976 227798
rect 198924 227734 198976 227740
rect 198740 222624 198792 222630
rect 198740 222566 198792 222572
rect 198280 222352 198332 222358
rect 198280 222294 198332 222300
rect 198936 217410 198964 227734
rect 199028 222601 199056 231676
rect 199396 225321 199424 231676
rect 199764 228002 199792 231676
rect 199752 227996 199804 228002
rect 199752 227938 199804 227944
rect 200132 227934 200160 231676
rect 200500 228177 200528 231676
rect 200486 228168 200542 228177
rect 200486 228103 200542 228112
rect 200120 227928 200172 227934
rect 200120 227870 200172 227876
rect 199382 225312 199438 225321
rect 199382 225247 199438 225256
rect 200868 225078 200896 231676
rect 200856 225072 200908 225078
rect 200856 225014 200908 225020
rect 199014 222592 199070 222601
rect 199014 222527 199070 222536
rect 201144 222426 201172 231676
rect 201408 225072 201460 225078
rect 201408 225014 201460 225020
rect 201132 222420 201184 222426
rect 201132 222362 201184 222368
rect 200764 222216 200816 222222
rect 200764 222158 200816 222164
rect 199936 221060 199988 221066
rect 199936 221002 199988 221008
rect 199948 217410 199976 221002
rect 200776 217410 200804 222158
rect 201420 217410 201448 225014
rect 201512 223009 201540 231676
rect 201682 226536 201738 226545
rect 201682 226471 201738 226480
rect 201592 226432 201644 226438
rect 201592 226374 201644 226380
rect 201498 223000 201554 223009
rect 201498 222935 201554 222944
rect 201604 222766 201632 226374
rect 201592 222760 201644 222766
rect 201592 222702 201644 222708
rect 201696 222698 201724 226471
rect 201880 222873 201908 231676
rect 202248 225457 202276 231676
rect 202616 226574 202644 231676
rect 202984 228313 203012 231676
rect 203352 228449 203380 231676
rect 203338 228440 203394 228449
rect 203338 228375 203394 228384
rect 202970 228304 203026 228313
rect 202970 228239 203026 228248
rect 203248 227996 203300 228002
rect 203248 227938 203300 227944
rect 202604 226568 202656 226574
rect 202604 226510 202656 226516
rect 202234 225448 202290 225457
rect 202234 225383 202290 225392
rect 201866 222864 201922 222873
rect 201866 222799 201922 222808
rect 201684 222692 201736 222698
rect 201684 222634 201736 222640
rect 202420 222352 202472 222358
rect 202420 222294 202472 222300
rect 202432 217410 202460 222294
rect 203260 217410 203288 227938
rect 203720 225593 203748 231676
rect 203996 227866 204024 231676
rect 203984 227860 204036 227866
rect 203984 227802 204036 227808
rect 204260 227724 204312 227730
rect 204260 227666 204312 227672
rect 204272 226642 204300 227666
rect 204260 226636 204312 226642
rect 204260 226578 204312 226584
rect 203706 225584 203762 225593
rect 203706 225519 203762 225528
rect 204364 223145 204392 231676
rect 204350 223136 204406 223145
rect 204350 223071 204406 223080
rect 204732 222494 204760 231676
rect 205100 225729 205128 231676
rect 205086 225720 205142 225729
rect 205086 225655 205142 225664
rect 204904 223916 204956 223922
rect 204904 223858 204956 223864
rect 204720 222488 204772 222494
rect 204720 222430 204772 222436
rect 204076 220856 204128 220862
rect 204076 220798 204128 220804
rect 204088 217410 204116 220798
rect 204916 217410 204944 223858
rect 205468 222562 205496 231676
rect 205836 228585 205864 231676
rect 206204 228993 206232 231676
rect 206190 228984 206246 228993
rect 206190 228919 206246 228928
rect 205822 228576 205878 228585
rect 205822 228511 205878 228520
rect 206572 224097 206600 231676
rect 206848 224942 206876 231676
rect 207018 228984 207074 228993
rect 207018 228919 207074 228928
rect 207032 225418 207060 228919
rect 207216 228721 207244 231676
rect 207584 228857 207612 231676
rect 207570 228848 207626 228857
rect 207570 228783 207626 228792
rect 207202 228712 207258 228721
rect 207202 228647 207258 228656
rect 207020 225412 207072 225418
rect 207020 225354 207072 225360
rect 206836 224936 206888 224942
rect 206836 224878 206888 224884
rect 206928 224936 206980 224942
rect 206928 224878 206980 224884
rect 206558 224088 206614 224097
rect 206558 224023 206614 224032
rect 206940 223786 206968 224878
rect 207952 224233 207980 231676
rect 208044 231662 208334 231690
rect 208044 225146 208072 231662
rect 208688 226545 208716 231676
rect 208674 226536 208730 226545
rect 208674 226471 208730 226480
rect 209056 226438 209084 231676
rect 209044 226432 209096 226438
rect 209044 226374 209096 226380
rect 208308 225208 208360 225214
rect 208308 225150 208360 225156
rect 208032 225140 208084 225146
rect 208032 225082 208084 225088
rect 207938 224224 207994 224233
rect 207938 224159 207994 224168
rect 206928 223780 206980 223786
rect 206928 223722 206980 223728
rect 207480 222624 207532 222630
rect 207480 222566 207532 222572
rect 205456 222556 205508 222562
rect 205456 222498 205508 222504
rect 205824 222420 205876 222426
rect 205824 222362 205876 222368
rect 205836 217410 205864 222362
rect 206652 220992 206704 220998
rect 206652 220934 206704 220940
rect 206664 217410 206692 220934
rect 207492 217410 207520 222566
rect 208320 217410 208348 225150
rect 209228 225140 209280 225146
rect 209228 225082 209280 225088
rect 208952 223780 209004 223786
rect 208952 223722 209004 223728
rect 208964 221338 208992 223722
rect 209136 222488 209188 222494
rect 209136 222430 209188 222436
rect 208952 221332 209004 221338
rect 208952 221274 209004 221280
rect 209148 217410 209176 222430
rect 209240 220862 209268 225082
rect 209424 223650 209452 231676
rect 209596 227928 209648 227934
rect 209596 227870 209648 227876
rect 209412 223644 209464 223650
rect 209412 223586 209464 223592
rect 209228 220856 209280 220862
rect 209228 220798 209280 220804
rect 64216 217382 64552 217410
rect 65044 217382 65380 217410
rect 65872 217382 66208 217410
rect 66700 217382 67036 217410
rect 67528 217382 67864 217410
rect 68356 217382 68692 217410
rect 69184 217382 69520 217410
rect 70104 217382 70440 217410
rect 70932 217382 71268 217410
rect 71760 217382 72096 217410
rect 72588 217382 72924 217410
rect 73416 217382 73752 217410
rect 74244 217382 74488 217410
rect 75072 217382 75408 217410
rect 75992 217382 76328 217410
rect 76820 217382 77156 217410
rect 77648 217382 77984 217410
rect 78476 217382 78812 217410
rect 79304 217382 79640 217410
rect 80132 217382 80468 217410
rect 80960 217382 81296 217410
rect 81880 217382 82216 217410
rect 82708 217382 82768 217410
rect 83536 217382 83872 217410
rect 84364 217382 84700 217410
rect 85192 217382 85528 217410
rect 86020 217382 86356 217410
rect 86848 217382 87184 217410
rect 87768 217382 88104 217410
rect 88596 217382 88932 217410
rect 89424 217382 89760 217410
rect 90252 217382 90588 217410
rect 91080 217382 91416 217410
rect 91908 217382 92244 217410
rect 92736 217382 93072 217410
rect 93656 217382 93808 217410
rect 94484 217382 94820 217410
rect 95312 217382 95648 217410
rect 96140 217382 96476 217410
rect 96968 217382 97304 217410
rect 97796 217382 98132 217410
rect 98624 217382 98960 217410
rect 99544 217382 99880 217410
rect 100372 217382 100708 217410
rect 101200 217382 101536 217410
rect 102028 217382 102088 217410
rect 102856 217382 103192 217410
rect 103684 217382 104020 217410
rect 104512 217382 104848 217410
rect 105432 217382 105768 217410
rect 106260 217382 106596 217410
rect 107088 217382 107424 217410
rect 107916 217382 108252 217410
rect 108744 217382 109080 217410
rect 109572 217382 109908 217410
rect 110400 217382 110736 217410
rect 111320 217382 111656 217410
rect 112148 217382 112484 217410
rect 112976 217382 113128 217410
rect 113804 217382 114140 217410
rect 114632 217382 114968 217410
rect 115460 217382 115796 217410
rect 116288 217382 116624 217410
rect 117208 217382 117544 217410
rect 118036 217382 118372 217410
rect 118864 217382 119200 217410
rect 119692 217382 120028 217410
rect 120520 217382 120856 217410
rect 121348 217382 121408 217410
rect 122176 217382 122512 217410
rect 123096 217382 123432 217410
rect 123924 217382 124168 217410
rect 124752 217382 125088 217410
rect 125580 217382 125916 217410
rect 126408 217382 126744 217410
rect 127236 217382 127572 217410
rect 128064 217382 128400 217410
rect 128984 217382 129320 217410
rect 129812 217382 130148 217410
rect 130640 217382 130976 217410
rect 131468 217382 131804 217410
rect 132296 217382 132448 217410
rect 133124 217382 133460 217410
rect 133952 217382 134288 217410
rect 134872 217382 135208 217410
rect 135700 217382 136036 217410
rect 136528 217382 136864 217410
rect 137356 217382 137692 217410
rect 138184 217382 138520 217410
rect 139012 217382 139348 217410
rect 139840 217382 140176 217410
rect 140760 217382 141096 217410
rect 141588 217382 141924 217410
rect 142416 217382 142752 217410
rect 143244 217382 143488 217410
rect 144072 217382 144408 217410
rect 144900 217382 145236 217410
rect 145728 217382 146064 217410
rect 146648 217382 146984 217410
rect 147476 217382 147812 217410
rect 148304 217382 148640 217410
rect 149132 217382 149468 217410
rect 149960 217382 150296 217410
rect 150788 217382 151124 217410
rect 151616 217382 151768 217410
rect 152536 217382 152872 217410
rect 153364 217382 153700 217410
rect 154192 217382 154528 217410
rect 155020 217382 155356 217410
rect 155848 217382 156184 217410
rect 156676 217382 157012 217410
rect 157504 217382 157840 217410
rect 158424 217382 158760 217410
rect 159252 217382 159588 217410
rect 160080 217382 160416 217410
rect 160908 217382 161244 217410
rect 161736 217382 162072 217410
rect 162564 217382 162808 217410
rect 163392 217382 163728 217410
rect 164312 217382 164648 217410
rect 165140 217382 165476 217410
rect 165968 217382 166304 217410
rect 166796 217382 167132 217410
rect 167624 217382 167960 217410
rect 168452 217382 168788 217410
rect 169280 217382 169616 217410
rect 170200 217382 170536 217410
rect 171028 217382 171088 217410
rect 171856 217382 172192 217410
rect 172684 217382 173020 217410
rect 173512 217382 173664 217410
rect 174340 217382 174676 217410
rect 175168 217382 175504 217410
rect 176088 217382 176424 217410
rect 176916 217382 177252 217410
rect 177744 217382 178080 217410
rect 178572 217382 178908 217410
rect 179400 217382 179736 217410
rect 180228 217382 180564 217410
rect 181056 217382 181392 217410
rect 181976 217382 182128 217410
rect 182804 217382 183140 217410
rect 183632 217382 183968 217410
rect 184460 217382 184796 217410
rect 185288 217382 185624 217410
rect 186116 217382 186452 217410
rect 186944 217382 187280 217410
rect 187864 217382 188200 217410
rect 188692 217382 189028 217410
rect 189520 217382 189856 217410
rect 190348 217382 190408 217410
rect 191176 217382 191512 217410
rect 192004 217382 192340 217410
rect 192832 217382 193168 217410
rect 193752 217382 194088 217410
rect 194580 217382 195008 217410
rect 195408 217382 195744 217410
rect 196236 217382 196572 217410
rect 197064 217382 197400 217410
rect 197892 217382 198228 217410
rect 198720 217382 198964 217410
rect 199640 217382 199976 217410
rect 200468 217382 200804 217410
rect 201296 217382 201448 217410
rect 202124 217382 202460 217410
rect 202952 217382 203288 217410
rect 203780 217382 204116 217410
rect 204608 217382 204944 217410
rect 205528 217382 205864 217410
rect 206356 217382 206692 217410
rect 207184 217382 207520 217410
rect 208012 217382 208348 217410
rect 208840 217382 209176 217410
rect 209608 217410 209636 227870
rect 209700 225350 209728 231676
rect 210068 227497 210096 231676
rect 210054 227488 210110 227497
rect 210054 227423 210110 227432
rect 210436 227361 210464 231676
rect 210804 228993 210832 231676
rect 210790 228984 210846 228993
rect 210790 228919 210846 228928
rect 210790 227624 210846 227633
rect 210790 227559 210846 227568
rect 210422 227352 210478 227361
rect 210422 227287 210478 227296
rect 209688 225344 209740 225350
rect 209688 225286 209740 225292
rect 209688 223712 209740 223718
rect 209688 223654 209740 223660
rect 209700 221542 209728 223654
rect 209688 221536 209740 221542
rect 209688 221478 209740 221484
rect 210804 217410 210832 227559
rect 211172 226001 211200 231676
rect 211158 225992 211214 226001
rect 211158 225927 211214 225936
rect 211540 223281 211568 231676
rect 211712 225276 211764 225282
rect 211712 225218 211764 225224
rect 211526 223272 211582 223281
rect 211526 223207 211582 223216
rect 211724 217410 211752 225218
rect 211908 223417 211936 231676
rect 212276 224058 212304 231676
rect 212354 227760 212410 227769
rect 212354 227695 212410 227704
rect 212264 224052 212316 224058
rect 212264 223994 212316 224000
rect 211894 223408 211950 223417
rect 211894 223343 211950 223352
rect 212368 217410 212396 227695
rect 212552 225865 212580 231676
rect 212920 227089 212948 231676
rect 213288 227225 213316 231676
rect 213274 227216 213330 227225
rect 213274 227151 213330 227160
rect 212906 227080 212962 227089
rect 212906 227015 212962 227024
rect 213656 226137 213684 231676
rect 213642 226128 213698 226137
rect 213642 226063 213698 226072
rect 212538 225856 212594 225865
rect 212538 225791 212594 225800
rect 214024 225554 214052 231676
rect 214012 225548 214064 225554
rect 214012 225490 214064 225496
rect 214392 223553 214420 231676
rect 214378 223544 214434 223553
rect 214378 223479 214434 223488
rect 214196 222760 214248 222766
rect 214196 222702 214248 222708
rect 213368 221536 213420 221542
rect 213368 221478 213420 221484
rect 213380 217410 213408 221478
rect 214208 217410 214236 222702
rect 214760 222057 214788 231676
rect 215128 225486 215156 231676
rect 215404 226273 215432 231676
rect 215772 226953 215800 231676
rect 216140 228070 216168 231676
rect 216128 228064 216180 228070
rect 216128 228006 216180 228012
rect 215758 226944 215814 226953
rect 215758 226879 215814 226888
rect 215390 226264 215446 226273
rect 215390 226199 215446 226208
rect 216508 225622 216536 231676
rect 216680 228064 216732 228070
rect 216680 228006 216732 228012
rect 216496 225616 216548 225622
rect 216496 225558 216548 225564
rect 216588 225616 216640 225622
rect 216588 225558 216640 225564
rect 215116 225480 215168 225486
rect 215116 225422 215168 225428
rect 215024 225344 215076 225350
rect 215024 225286 215076 225292
rect 214932 223644 214984 223650
rect 214932 223586 214984 223592
rect 214746 222048 214802 222057
rect 214746 221983 214802 221992
rect 214944 221270 214972 223586
rect 214932 221264 214984 221270
rect 214932 221206 214984 221212
rect 215036 217410 215064 225286
rect 216128 224052 216180 224058
rect 216128 223994 216180 224000
rect 215852 222556 215904 222562
rect 215852 222498 215904 222504
rect 215864 217410 215892 222498
rect 216140 221134 216168 223994
rect 216128 221128 216180 221134
rect 216128 221070 216180 221076
rect 216600 220930 216628 225558
rect 216588 220924 216640 220930
rect 216588 220866 216640 220872
rect 216692 217410 216720 228006
rect 216876 224777 216904 231676
rect 216862 224768 216918 224777
rect 216862 224703 216918 224712
rect 217244 221921 217272 231676
rect 217336 231662 217626 231690
rect 217230 221912 217286 221921
rect 217230 221847 217286 221856
rect 217336 221785 217364 231662
rect 217598 227896 217654 227905
rect 217598 227831 217654 227840
rect 217322 221776 217378 221785
rect 217322 221711 217378 221720
rect 217612 217410 217640 227831
rect 217980 225690 218008 231676
rect 217968 225684 218020 225690
rect 217968 225626 218020 225632
rect 218256 224641 218284 231676
rect 218624 226817 218652 231676
rect 218992 228138 219020 231676
rect 219254 228168 219310 228177
rect 218980 228132 219032 228138
rect 219254 228103 219310 228112
rect 218980 228074 219032 228080
rect 218610 226808 218666 226817
rect 218610 226743 218666 226752
rect 218428 225548 218480 225554
rect 218428 225490 218480 225496
rect 218242 224632 218298 224641
rect 218242 224567 218298 224576
rect 218440 217410 218468 225490
rect 219268 217410 219296 228103
rect 219360 224505 219388 231676
rect 219728 225826 219756 231676
rect 219716 225820 219768 225826
rect 219716 225762 219768 225768
rect 219346 224496 219402 224505
rect 219346 224431 219402 224440
rect 220096 222834 220124 231676
rect 220084 222828 220136 222834
rect 220084 222770 220136 222776
rect 220464 221377 220492 231676
rect 220726 228032 220782 228041
rect 220726 227967 220782 227976
rect 220450 221368 220506 221377
rect 220084 221332 220136 221338
rect 220450 221303 220506 221312
rect 220084 221274 220136 221280
rect 220096 217410 220124 221274
rect 220740 217410 220768 227967
rect 220832 224369 220860 231676
rect 220818 224360 220874 224369
rect 220818 224295 220874 224304
rect 221108 220114 221136 231676
rect 221476 221649 221504 231676
rect 221740 225480 221792 225486
rect 221740 225422 221792 225428
rect 221462 221640 221518 221649
rect 221462 221575 221518 221584
rect 221096 220108 221148 220114
rect 221096 220050 221148 220056
rect 221752 217410 221780 225422
rect 221844 221513 221872 231676
rect 222212 225758 222240 231676
rect 222304 231662 222594 231690
rect 222200 225752 222252 225758
rect 222200 225694 222252 225700
rect 221830 221504 221886 221513
rect 221830 221439 221886 221448
rect 222304 220182 222332 231662
rect 222948 228206 222976 231676
rect 223316 228342 223344 231676
rect 223304 228336 223356 228342
rect 223304 228278 223356 228284
rect 222936 228200 222988 228206
rect 222936 228142 222988 228148
rect 223488 228132 223540 228138
rect 223488 228074 223540 228080
rect 222568 222692 222620 222698
rect 222568 222634 222620 222640
rect 222292 220176 222344 220182
rect 222292 220118 222344 220124
rect 222580 217410 222608 222634
rect 223500 217410 223528 228074
rect 223684 225894 223712 231676
rect 223672 225888 223724 225894
rect 223672 225830 223724 225836
rect 223960 220250 223988 231676
rect 224052 231662 224342 231690
rect 224052 222902 224080 231662
rect 224696 222970 224724 231676
rect 225064 225962 225092 231676
rect 225052 225956 225104 225962
rect 225052 225898 225104 225904
rect 225144 225412 225196 225418
rect 225144 225354 225196 225360
rect 224684 222964 224736 222970
rect 224684 222906 224736 222912
rect 224040 222896 224092 222902
rect 224040 222838 224092 222844
rect 224316 222828 224368 222834
rect 224316 222770 224368 222776
rect 223948 220244 224000 220250
rect 223948 220186 224000 220192
rect 224328 217410 224356 222770
rect 225156 217410 225184 225354
rect 225432 220318 225460 231676
rect 225800 228274 225828 231676
rect 226168 228410 226196 231676
rect 226156 228404 226208 228410
rect 226156 228346 226208 228352
rect 225970 228304 226026 228313
rect 225788 228268 225840 228274
rect 225970 228239 226026 228248
rect 225788 228210 225840 228216
rect 225420 220312 225472 220318
rect 225420 220254 225472 220260
rect 225984 217410 226012 228239
rect 226536 226030 226564 231676
rect 226628 231662 226826 231690
rect 226524 226024 226576 226030
rect 226524 225966 226576 225972
rect 226628 220386 226656 231662
rect 227180 223038 227208 231676
rect 227548 223106 227576 231676
rect 227628 228268 227680 228274
rect 227628 228210 227680 228216
rect 227536 223100 227588 223106
rect 227536 223042 227588 223048
rect 227168 223032 227220 223038
rect 227168 222974 227220 222980
rect 226800 221060 226852 221066
rect 226800 221002 226852 221008
rect 226616 220380 226668 220386
rect 226616 220322 226668 220328
rect 226812 217410 226840 221002
rect 227640 217410 227668 228210
rect 227916 226098 227944 231676
rect 227904 226092 227956 226098
rect 227904 226034 227956 226040
rect 228284 220454 228312 231676
rect 228652 228478 228680 231676
rect 229020 228682 229048 231676
rect 229008 228676 229060 228682
rect 229008 228618 229060 228624
rect 228640 228472 228692 228478
rect 228640 228414 228692 228420
rect 229284 228336 229336 228342
rect 229284 228278 229336 228284
rect 228456 225616 228508 225622
rect 228456 225558 228508 225564
rect 228272 220448 228324 220454
rect 228272 220390 228324 220396
rect 228468 217410 228496 225558
rect 229296 217410 229324 228278
rect 229388 226166 229416 231676
rect 229376 226160 229428 226166
rect 229376 226102 229428 226108
rect 229664 220522 229692 231676
rect 230032 223174 230060 231676
rect 230400 223242 230428 231676
rect 230768 226302 230796 231676
rect 231136 228750 231164 231676
rect 231124 228744 231176 228750
rect 231124 228686 231176 228692
rect 231504 228614 231532 231676
rect 231492 228608 231544 228614
rect 231492 228550 231544 228556
rect 231872 228546 231900 231676
rect 231860 228540 231912 228546
rect 231860 228482 231912 228488
rect 231676 228200 231728 228206
rect 231676 228142 231728 228148
rect 230756 226296 230808 226302
rect 230756 226238 230808 226244
rect 231308 225820 231360 225826
rect 231308 225762 231360 225768
rect 230388 223236 230440 223242
rect 230388 223178 230440 223184
rect 230020 223168 230072 223174
rect 230020 223110 230072 223116
rect 231032 223032 231084 223038
rect 231032 222974 231084 222980
rect 230112 221128 230164 221134
rect 230112 221070 230164 221076
rect 230204 221128 230256 221134
rect 230204 221070 230256 221076
rect 230124 220930 230152 221070
rect 230112 220924 230164 220930
rect 230112 220866 230164 220872
rect 229652 220516 229704 220522
rect 229652 220458 229704 220464
rect 230216 217410 230244 221070
rect 231044 217410 231072 222974
rect 231216 221332 231268 221338
rect 231216 221274 231268 221280
rect 231228 220862 231256 221274
rect 231320 221202 231348 225762
rect 231308 221196 231360 221202
rect 231308 221138 231360 221144
rect 231216 220856 231268 220862
rect 231216 220798 231268 220804
rect 231688 217410 231716 228142
rect 232240 226234 232268 231676
rect 232228 226228 232280 226234
rect 232228 226170 232280 226176
rect 232044 225752 232096 225758
rect 232044 225694 232096 225700
rect 232056 220930 232084 225694
rect 232516 223854 232544 231676
rect 232504 223848 232556 223854
rect 232504 223790 232556 223796
rect 232884 223446 232912 231676
rect 232872 223440 232924 223446
rect 232872 223382 232924 223388
rect 233252 223378 233280 231676
rect 233516 226432 233568 226438
rect 233516 226374 233568 226380
rect 233240 223372 233292 223378
rect 233240 223314 233292 223320
rect 232596 223100 232648 223106
rect 232596 223042 232648 223048
rect 232608 222018 232636 223042
rect 232688 222896 232740 222902
rect 232688 222838 232740 222844
rect 232596 222012 232648 222018
rect 232596 221954 232648 221960
rect 232044 220924 232096 220930
rect 232044 220866 232096 220872
rect 232700 217410 232728 222838
rect 233528 221746 233556 226374
rect 233620 224738 233648 231676
rect 233988 229022 234016 231676
rect 233976 229016 234028 229022
rect 233976 228958 234028 228964
rect 234356 228886 234384 231676
rect 234344 228880 234396 228886
rect 234344 228822 234396 228828
rect 234724 228818 234752 231676
rect 234712 228812 234764 228818
rect 234712 228754 234764 228760
rect 235092 224806 235120 231676
rect 235264 228404 235316 228410
rect 235264 228346 235316 228352
rect 235080 224800 235132 224806
rect 235080 224742 235132 224748
rect 233608 224732 233660 224738
rect 233608 224674 233660 224680
rect 234344 221944 234396 221950
rect 234344 221886 234396 221892
rect 233516 221740 233568 221746
rect 233516 221682 233568 221688
rect 233516 221332 233568 221338
rect 233516 221274 233568 221280
rect 233528 217410 233556 221274
rect 234356 217410 234384 221886
rect 235276 217410 235304 228346
rect 235368 227662 235396 231676
rect 235356 227656 235408 227662
rect 235356 227598 235408 227604
rect 235736 223514 235764 231676
rect 236104 223582 236132 231676
rect 236276 226636 236328 226642
rect 236276 226578 236328 226584
rect 236092 223576 236144 223582
rect 236092 223518 236144 223524
rect 235724 223508 235776 223514
rect 235724 223450 235776 223456
rect 235908 223168 235960 223174
rect 235908 223110 235960 223116
rect 235920 222290 235948 223110
rect 236092 222964 236144 222970
rect 236092 222906 236144 222912
rect 235908 222284 235960 222290
rect 235908 222226 235960 222232
rect 235632 221672 235684 221678
rect 235684 221620 236040 221626
rect 235632 221614 236040 221620
rect 235644 221610 236040 221614
rect 235644 221604 236052 221610
rect 235644 221598 236000 221604
rect 236000 221546 236052 221552
rect 236104 217410 236132 222906
rect 236288 220998 236316 226578
rect 236472 224602 236500 231676
rect 236734 228440 236790 228449
rect 236734 228375 236790 228384
rect 236460 224596 236512 224602
rect 236460 224538 236512 224544
rect 236276 220992 236328 220998
rect 236276 220934 236328 220940
rect 236748 220862 236776 228375
rect 236840 223718 236868 231676
rect 237208 228954 237236 231676
rect 237576 229090 237604 231676
rect 237564 229084 237616 229090
rect 237564 229026 237616 229032
rect 237196 228948 237248 228954
rect 237196 228890 237248 228896
rect 237010 228576 237066 228585
rect 237010 228511 237066 228520
rect 236828 223712 236880 223718
rect 236828 223654 236880 223660
rect 237024 221474 237052 228511
rect 237944 224670 237972 231676
rect 238220 227594 238248 231676
rect 238312 231662 238602 231690
rect 238208 227588 238260 227594
rect 238208 227530 238260 227536
rect 237932 224664 237984 224670
rect 237932 224606 237984 224612
rect 237748 223372 237800 223378
rect 237748 223314 237800 223320
rect 237012 221468 237064 221474
rect 237012 221410 237064 221416
rect 236920 221400 236972 221406
rect 236920 221342 236972 221348
rect 236736 220856 236788 220862
rect 236736 220798 236788 220804
rect 236932 217410 236960 221342
rect 237760 217410 237788 223314
rect 238312 222086 238340 231662
rect 238576 228472 238628 228478
rect 238576 228414 238628 228420
rect 238300 222080 238352 222086
rect 238300 222022 238352 222028
rect 238588 217410 238616 228414
rect 238956 222154 238984 231676
rect 239324 224466 239352 231676
rect 239312 224460 239364 224466
rect 239312 224402 239364 224408
rect 239692 223786 239720 231676
rect 239772 228880 239824 228886
rect 239772 228822 239824 228828
rect 239680 223780 239732 223786
rect 239680 223722 239732 223728
rect 239404 223236 239456 223242
rect 239404 223178 239456 223184
rect 238944 222148 238996 222154
rect 238944 222090 238996 222096
rect 239416 217410 239444 223178
rect 239784 221134 239812 228822
rect 239956 228812 240008 228818
rect 239956 228754 240008 228760
rect 239864 228608 239916 228614
rect 239864 228550 239916 228556
rect 239876 221338 239904 228550
rect 239864 221332 239916 221338
rect 239864 221274 239916 221280
rect 239772 221128 239824 221134
rect 239772 221070 239824 221076
rect 239968 221066 239996 228754
rect 240060 227458 240088 231676
rect 240140 228540 240192 228546
rect 240140 228482 240192 228488
rect 240048 227452 240100 227458
rect 240048 227394 240100 227400
rect 239956 221060 240008 221066
rect 239956 221002 240008 221008
rect 240152 220946 240180 228482
rect 240428 227526 240456 231676
rect 240416 227520 240468 227526
rect 240416 227462 240468 227468
rect 240796 224534 240824 231676
rect 241072 227254 241100 231676
rect 241244 228948 241296 228954
rect 241244 228890 241296 228896
rect 241060 227248 241112 227254
rect 241060 227190 241112 227196
rect 240784 224528 240836 224534
rect 240784 224470 240836 224476
rect 241152 223508 241204 223514
rect 241152 223450 241204 223456
rect 240060 220918 240180 220946
rect 240060 217410 240088 220918
rect 241164 217410 241192 223450
rect 241256 221406 241284 228890
rect 241440 227390 241468 231676
rect 241428 227384 241480 227390
rect 241428 227326 241480 227332
rect 241808 222018 241836 231676
rect 241980 228744 242032 228750
rect 241980 228686 242032 228692
rect 241796 222012 241848 222018
rect 241796 221954 241848 221960
rect 241244 221400 241296 221406
rect 241244 221342 241296 221348
rect 241992 217410 242020 228686
rect 242176 224398 242204 231676
rect 242164 224392 242216 224398
rect 242164 224334 242216 224340
rect 242544 223650 242572 231676
rect 242926 231662 243124 231690
rect 243096 226334 243124 231662
rect 243280 227186 243308 231676
rect 243544 229016 243596 229022
rect 243544 228958 243596 228964
rect 243268 227180 243320 227186
rect 243268 227122 243320 227128
rect 242912 226306 243124 226334
rect 242532 223644 242584 223650
rect 242532 223586 242584 223592
rect 242912 223258 242940 226306
rect 243084 225956 243136 225962
rect 243084 225898 243136 225904
rect 242992 225888 243044 225894
rect 242992 225830 243044 225836
rect 242728 223230 242940 223258
rect 242728 223106 242756 223230
rect 242716 223100 242768 223106
rect 242716 223042 242768 223048
rect 242808 223100 242860 223106
rect 242808 223042 242860 223048
rect 242820 217410 242848 223042
rect 243004 221270 243032 225830
rect 242992 221264 243044 221270
rect 242992 221206 243044 221212
rect 243096 221202 243124 225898
rect 243084 221196 243136 221202
rect 243084 221138 243136 221144
rect 243556 217410 243584 228958
rect 243648 224330 243676 231676
rect 243924 227050 243952 231676
rect 244292 227322 244320 231676
rect 244280 227316 244332 227322
rect 244280 227258 244332 227264
rect 243912 227044 243964 227050
rect 243912 226986 243964 226992
rect 243636 224324 243688 224330
rect 243636 224266 243688 224272
rect 244660 223310 244688 231676
rect 245028 224194 245056 231676
rect 245292 228676 245344 228682
rect 245292 228618 245344 228624
rect 245016 224188 245068 224194
rect 245016 224130 245068 224136
rect 244648 223304 244700 223310
rect 244648 223246 244700 223252
rect 244464 222148 244516 222154
rect 244464 222090 244516 222096
rect 244476 217410 244504 222090
rect 245304 217410 245332 228618
rect 245396 221610 245424 231676
rect 245658 228848 245714 228857
rect 245658 228783 245714 228792
rect 245672 222766 245700 228783
rect 245660 222760 245712 222766
rect 245660 222702 245712 222708
rect 245764 221814 245792 231676
rect 246132 227118 246160 231676
rect 246212 229084 246264 229090
rect 246212 229026 246264 229032
rect 246120 227112 246172 227118
rect 246120 227054 246172 227060
rect 246120 222760 246172 222766
rect 246120 222702 246172 222708
rect 245752 221808 245804 221814
rect 245752 221750 245804 221756
rect 245384 221604 245436 221610
rect 245384 221546 245436 221552
rect 246132 217410 246160 222702
rect 246224 222630 246252 229026
rect 246500 224262 246528 231676
rect 246488 224256 246540 224262
rect 246488 224198 246540 224204
rect 246776 224058 246804 231676
rect 247040 227112 247092 227118
rect 247040 227054 247092 227060
rect 246764 224052 246816 224058
rect 246764 223994 246816 224000
rect 246212 222624 246264 222630
rect 246212 222566 246264 222572
rect 247052 217410 247080 227054
rect 247144 226982 247172 231676
rect 247132 226976 247184 226982
rect 247132 226918 247184 226924
rect 247512 226438 247540 231676
rect 247500 226432 247552 226438
rect 247500 226374 247552 226380
rect 247880 224126 247908 231676
rect 248248 226778 248276 231676
rect 248340 231662 248630 231690
rect 248236 226772 248288 226778
rect 248236 226714 248288 226720
rect 247868 224120 247920 224126
rect 247868 224062 247920 224068
rect 248340 221678 248368 231662
rect 248696 227656 248748 227662
rect 248696 227598 248748 227604
rect 248512 227248 248564 227254
rect 248512 227190 248564 227196
rect 248420 226772 248472 226778
rect 248420 226714 248472 226720
rect 248432 222834 248460 226714
rect 248524 223038 248552 227190
rect 248604 226908 248656 226914
rect 248604 226850 248656 226856
rect 248512 223032 248564 223038
rect 248512 222974 248564 222980
rect 248420 222828 248472 222834
rect 248420 222770 248472 222776
rect 248616 221950 248644 226850
rect 248604 221944 248656 221950
rect 248604 221886 248656 221892
rect 248328 221672 248380 221678
rect 248328 221614 248380 221620
rect 247868 221400 247920 221406
rect 247868 221342 247920 221348
rect 247880 217410 247908 221342
rect 248708 217410 248736 227598
rect 248984 226846 249012 231676
rect 248972 226840 249024 226846
rect 248972 226782 249024 226788
rect 249352 223990 249380 231676
rect 249628 225826 249656 231676
rect 249616 225820 249668 225826
rect 249616 225762 249668 225768
rect 249340 223984 249392 223990
rect 249340 223926 249392 223932
rect 249996 223174 250024 231676
rect 250088 231662 250378 231690
rect 249984 223168 250036 223174
rect 249984 223110 250036 223116
rect 250088 221542 250116 231662
rect 250352 227588 250404 227594
rect 250352 227530 250404 227536
rect 250076 221536 250128 221542
rect 250076 221478 250128 221484
rect 249524 221468 249576 221474
rect 249524 221410 249576 221416
rect 249536 217410 249564 221410
rect 250364 217410 250392 227530
rect 250732 224942 250760 231676
rect 251100 226710 251128 231676
rect 251468 226982 251496 231676
rect 251836 227730 251864 231676
rect 251824 227724 251876 227730
rect 251824 227666 251876 227672
rect 252008 227520 252060 227526
rect 252008 227462 252060 227468
rect 251456 226976 251508 226982
rect 251456 226918 251508 226924
rect 251088 226704 251140 226710
rect 251088 226646 251140 226652
rect 250720 224936 250772 224942
rect 250720 224878 250772 224884
rect 251088 221332 251140 221338
rect 251088 221274 251140 221280
rect 251100 217410 251128 221274
rect 252020 217410 252048 227462
rect 252204 225010 252232 231676
rect 252480 225690 252508 231676
rect 252848 225894 252876 231676
rect 252940 231662 253230 231690
rect 253308 231662 253598 231690
rect 252940 225962 252968 231662
rect 253204 227316 253256 227322
rect 253204 227258 253256 227264
rect 252928 225956 252980 225962
rect 252928 225898 252980 225904
rect 252836 225888 252888 225894
rect 252836 225830 252888 225836
rect 252468 225684 252520 225690
rect 252468 225626 252520 225632
rect 252192 225004 252244 225010
rect 252192 224946 252244 224952
rect 253216 223378 253244 227258
rect 253308 224874 253336 231662
rect 253756 227724 253808 227730
rect 253756 227666 253808 227672
rect 253572 227384 253624 227390
rect 253572 227326 253624 227332
rect 253296 224868 253348 224874
rect 253296 224810 253348 224816
rect 253584 223514 253612 227326
rect 253572 223508 253624 223514
rect 253572 223450 253624 223456
rect 253204 223372 253256 223378
rect 253204 223314 253256 223320
rect 252928 221264 252980 221270
rect 252928 221206 252980 221212
rect 252940 217410 252968 221206
rect 253768 217410 253796 227666
rect 253952 225758 253980 231676
rect 254320 227798 254348 231676
rect 254688 227866 254716 231676
rect 254676 227860 254728 227866
rect 254676 227802 254728 227808
rect 254308 227792 254360 227798
rect 254308 227734 254360 227740
rect 253940 225752 253992 225758
rect 253940 225694 253992 225700
rect 255056 225078 255084 231676
rect 255332 228002 255360 231676
rect 255320 227996 255372 228002
rect 255320 227938 255372 227944
rect 255504 227044 255556 227050
rect 255504 226986 255556 226992
rect 255320 226500 255372 226506
rect 255320 226442 255372 226448
rect 255044 225072 255096 225078
rect 255044 225014 255096 225020
rect 255332 222970 255360 226442
rect 255516 223242 255544 226986
rect 255504 223236 255556 223242
rect 255504 223178 255556 223184
rect 255320 222964 255372 222970
rect 255320 222906 255372 222912
rect 254584 222284 254636 222290
rect 254584 222226 254636 222232
rect 254596 217410 254624 222226
rect 255700 222222 255728 231676
rect 255964 227996 256016 228002
rect 255964 227938 256016 227944
rect 255780 226772 255832 226778
rect 255780 226714 255832 226720
rect 255792 222902 255820 226714
rect 255780 222896 255832 222902
rect 255780 222838 255832 222844
rect 255688 222216 255740 222222
rect 255688 222158 255740 222164
rect 255412 221672 255464 221678
rect 255412 221614 255464 221620
rect 255424 217410 255452 221614
rect 255976 221406 256004 227938
rect 256068 222358 256096 231676
rect 256436 223922 256464 231676
rect 256516 227792 256568 227798
rect 256516 227734 256568 227740
rect 256424 223916 256476 223922
rect 256424 223858 256476 223864
rect 256056 222352 256108 222358
rect 256056 222294 256108 222300
rect 255964 221400 256016 221406
rect 255964 221342 256016 221348
rect 256240 221400 256292 221406
rect 256240 221342 256292 221348
rect 256252 217410 256280 221342
rect 256528 221338 256556 227734
rect 256608 227180 256660 227186
rect 256608 227122 256660 227128
rect 256620 222154 256648 227122
rect 256804 226642 256832 231676
rect 256792 226636 256844 226642
rect 256792 226578 256844 226584
rect 257172 225146 257200 231676
rect 257160 225140 257212 225146
rect 257160 225082 257212 225088
rect 257068 222896 257120 222902
rect 257068 222838 257120 222844
rect 256608 222148 256660 222154
rect 256608 222090 256660 222096
rect 256516 221332 256568 221338
rect 256516 221274 256568 221280
rect 257080 217410 257108 222838
rect 257540 222426 257568 231676
rect 257908 225214 257936 231676
rect 258184 227934 258212 231676
rect 258552 229090 258580 231676
rect 258644 231662 258934 231690
rect 258540 229084 258592 229090
rect 258540 229026 258592 229032
rect 258172 227928 258224 227934
rect 258172 227870 258224 227876
rect 258356 227928 258408 227934
rect 258356 227870 258408 227876
rect 258172 226364 258224 226370
rect 258172 226306 258224 226312
rect 257896 225208 257948 225214
rect 257896 225150 257948 225156
rect 258184 222698 258212 226306
rect 258172 222692 258224 222698
rect 258172 222634 258224 222640
rect 257528 222420 257580 222426
rect 257528 222362 257580 222368
rect 257896 221740 257948 221746
rect 257896 221682 257948 221688
rect 257908 217410 257936 221682
rect 258368 221270 258396 227870
rect 258644 222494 258672 231662
rect 258724 227452 258776 227458
rect 258724 227394 258776 227400
rect 258736 227186 258764 227394
rect 258724 227180 258776 227186
rect 258724 227122 258776 227128
rect 258908 227112 258960 227118
rect 258908 227054 258960 227060
rect 259182 227080 259238 227089
rect 258724 226976 258776 226982
rect 258724 226918 258776 226924
rect 258736 222766 258764 226918
rect 258816 226704 258868 226710
rect 258816 226646 258868 226652
rect 258828 223106 258856 226646
rect 258816 223100 258868 223106
rect 258816 223042 258868 223048
rect 258724 222760 258776 222766
rect 258724 222702 258776 222708
rect 258632 222488 258684 222494
rect 258632 222430 258684 222436
rect 258816 222216 258868 222222
rect 258816 222158 258868 222164
rect 258356 221264 258408 221270
rect 258356 221206 258408 221212
rect 258828 217410 258856 222158
rect 258920 221474 258948 227054
rect 259182 227015 259238 227024
rect 259196 222562 259224 227015
rect 259288 225282 259316 231676
rect 259656 228585 259684 231676
rect 259642 228576 259698 228585
rect 259642 228511 259698 228520
rect 259552 227860 259604 227866
rect 259552 227802 259604 227808
rect 259276 225276 259328 225282
rect 259276 225218 259328 225224
rect 259368 222624 259420 222630
rect 259368 222566 259420 222572
rect 259184 222556 259236 222562
rect 259184 222498 259236 222504
rect 258908 221468 258960 221474
rect 258908 221410 258960 221416
rect 259380 217410 259408 222566
rect 259564 221406 259592 227802
rect 260024 227633 260052 231676
rect 260392 227769 260420 231676
rect 260378 227760 260434 227769
rect 260378 227695 260434 227704
rect 260010 227624 260066 227633
rect 260010 227559 260066 227568
rect 260760 225350 260788 231676
rect 261036 228070 261064 231676
rect 261404 228857 261432 231676
rect 261390 228848 261446 228857
rect 261390 228783 261446 228792
rect 261024 228064 261076 228070
rect 261024 228006 261076 228012
rect 261772 227089 261800 231676
rect 261758 227080 261814 227089
rect 261758 227015 261814 227024
rect 262140 225554 262168 231676
rect 262508 228449 262536 231676
rect 262494 228440 262550 228449
rect 262494 228375 262550 228384
rect 262876 227905 262904 231676
rect 263244 228177 263272 231676
rect 263230 228168 263286 228177
rect 263230 228103 263286 228112
rect 262862 227896 262918 227905
rect 262862 227831 262918 227840
rect 262128 225548 262180 225554
rect 262128 225490 262180 225496
rect 263612 225486 263640 231676
rect 263888 228138 263916 231676
rect 263876 228132 263928 228138
rect 263876 228074 263928 228080
rect 264256 228041 264284 231676
rect 264242 228032 264298 228041
rect 264242 227967 264298 227976
rect 264624 226370 264652 231676
rect 264612 226364 264664 226370
rect 264612 226306 264664 226312
rect 263600 225480 263652 225486
rect 263600 225422 263652 225428
rect 264992 225418 265020 231676
rect 265360 228818 265388 231676
rect 265348 228812 265400 228818
rect 265348 228754 265400 228760
rect 265728 226846 265756 231676
rect 266096 228313 266124 231676
rect 266082 228304 266138 228313
rect 266082 228239 266138 228248
rect 265716 226840 265768 226846
rect 265716 226782 265768 226788
rect 266464 225622 266492 231676
rect 266740 228886 266768 231676
rect 266728 228880 266780 228886
rect 266728 228822 266780 228828
rect 267108 228274 267136 231676
rect 267476 228342 267504 231676
rect 267464 228336 267516 228342
rect 267464 228278 267516 228284
rect 267096 228268 267148 228274
rect 267096 228210 267148 228216
rect 267844 228206 267872 231676
rect 268212 228614 268240 231676
rect 268200 228608 268252 228614
rect 268200 228550 268252 228556
rect 267832 228200 267884 228206
rect 267832 228142 267884 228148
rect 268580 227254 268608 231676
rect 268568 227248 268620 227254
rect 268568 227190 268620 227196
rect 268948 226778 268976 231676
rect 269316 228410 269344 231676
rect 269592 228954 269620 231676
rect 269580 228948 269632 228954
rect 269580 228890 269632 228896
rect 269304 228404 269356 228410
rect 269304 228346 269356 228352
rect 269960 226914 269988 231676
rect 269948 226908 270000 226914
rect 269948 226850 270000 226856
rect 268936 226772 268988 226778
rect 268936 226714 268988 226720
rect 270328 226506 270356 231676
rect 270696 228478 270724 231676
rect 271064 228546 271092 231676
rect 271052 228540 271104 228546
rect 271052 228482 271104 228488
rect 270684 228472 270736 228478
rect 270684 228414 270736 228420
rect 271432 227322 271460 231676
rect 271420 227316 271472 227322
rect 271420 227258 271472 227264
rect 271800 227050 271828 231676
rect 272168 228750 272196 231676
rect 272444 229022 272472 231676
rect 272432 229016 272484 229022
rect 272432 228958 272484 228964
rect 272156 228744 272208 228750
rect 272156 228686 272208 228692
rect 272812 227390 272840 231676
rect 272800 227384 272852 227390
rect 272800 227326 272852 227332
rect 271788 227044 271840 227050
rect 271788 226986 271840 226992
rect 273180 226710 273208 231676
rect 273548 228682 273576 231676
rect 273536 228676 273588 228682
rect 273536 228618 273588 228624
rect 273916 227186 273944 231676
rect 274284 227458 274312 231676
rect 274272 227452 274324 227458
rect 274272 227394 274324 227400
rect 273904 227180 273956 227186
rect 273904 227122 273956 227128
rect 274652 226982 274680 231676
rect 275020 227662 275048 231676
rect 275008 227656 275060 227662
rect 275008 227598 275060 227604
rect 275296 227594 275324 231676
rect 275664 228002 275692 231676
rect 275652 227996 275704 228002
rect 275652 227938 275704 227944
rect 275284 227588 275336 227594
rect 275284 227530 275336 227536
rect 276032 227118 276060 231676
rect 276400 227526 276428 231676
rect 276768 227730 276796 231676
rect 277136 227798 277164 231676
rect 277504 227934 277532 231676
rect 277492 227928 277544 227934
rect 277492 227870 277544 227876
rect 277124 227792 277176 227798
rect 277124 227734 277176 227740
rect 276756 227724 276808 227730
rect 276756 227666 276808 227672
rect 276388 227520 276440 227526
rect 276388 227462 276440 227468
rect 276020 227112 276072 227118
rect 276020 227054 276072 227060
rect 274640 226976 274692 226982
rect 274640 226918 274692 226924
rect 273168 226704 273220 226710
rect 273168 226646 273220 226652
rect 270316 226500 270368 226506
rect 270316 226442 270368 226448
rect 266452 225616 266504 225622
rect 266452 225558 266504 225564
rect 264980 225412 265032 225418
rect 264980 225354 265032 225360
rect 260748 225344 260800 225350
rect 260748 225286 260800 225292
rect 271420 223100 271472 223106
rect 271420 223042 271472 223048
rect 263784 222964 263836 222970
rect 263784 222906 263836 222912
rect 262956 222760 263008 222766
rect 262956 222702 263008 222708
rect 260472 222692 260524 222698
rect 260472 222634 260524 222640
rect 259552 221400 259604 221406
rect 259552 221342 259604 221348
rect 260484 217410 260512 222634
rect 261300 222556 261352 222562
rect 261300 222498 261352 222504
rect 261312 217410 261340 222498
rect 262128 222488 262180 222494
rect 262128 222430 262180 222436
rect 262140 217410 262168 222430
rect 262968 217410 262996 222702
rect 263796 217410 263824 222906
rect 264612 222828 264664 222834
rect 264612 222770 264664 222776
rect 264624 217410 264652 222770
rect 269672 222352 269724 222358
rect 269672 222294 269724 222300
rect 268016 221808 268068 221814
rect 268016 221750 268068 221756
rect 266360 221536 266412 221542
rect 266360 221478 266412 221484
rect 265532 221468 265584 221474
rect 265532 221410 265584 221416
rect 265544 217410 265572 221410
rect 266372 217410 266400 221478
rect 267188 221400 267240 221406
rect 267188 221342 267240 221348
rect 267200 217410 267228 221342
rect 268028 217410 268056 221750
rect 268844 221264 268896 221270
rect 268844 221206 268896 221212
rect 268856 217410 268884 221206
rect 269684 217410 269712 222294
rect 270408 221332 270460 221338
rect 270408 221274 270460 221280
rect 270420 217410 270448 221274
rect 271432 217410 271460 223042
rect 272248 222420 272300 222426
rect 272248 222362 272300 222368
rect 272260 217410 272288 222362
rect 273076 222148 273128 222154
rect 273076 222090 273128 222096
rect 273088 217410 273116 222090
rect 274732 222080 274784 222086
rect 274732 222022 274784 222028
rect 273904 221944 273956 221950
rect 273904 221886 273956 221892
rect 273916 217410 273944 221886
rect 274744 217410 274772 222022
rect 277872 221678 277900 231676
rect 278148 222902 278176 231676
rect 278136 222896 278188 222902
rect 278136 222838 278188 222844
rect 278516 222290 278544 231676
rect 278884 227866 278912 231676
rect 278872 227860 278924 227866
rect 278872 227802 278924 227808
rect 278688 223576 278740 223582
rect 278688 223518 278740 223524
rect 278504 222284 278556 222290
rect 278504 222226 278556 222232
rect 277860 221672 277912 221678
rect 277860 221614 277912 221620
rect 275560 221604 275612 221610
rect 275560 221546 275612 221552
rect 278136 221604 278188 221610
rect 278136 221546 278188 221552
rect 275572 217410 275600 221546
rect 277308 221196 277360 221202
rect 277308 221138 277360 221144
rect 276480 220992 276532 220998
rect 276480 220934 276532 220940
rect 276492 217410 276520 220934
rect 277320 217410 277348 221138
rect 278148 217410 278176 221546
rect 278700 217410 278728 223518
rect 279252 222222 279280 231676
rect 279620 222698 279648 231676
rect 279608 222692 279660 222698
rect 279608 222634 279660 222640
rect 279240 222216 279292 222222
rect 279240 222158 279292 222164
rect 279988 221746 280016 231676
rect 280356 222630 280384 231676
rect 280344 222624 280396 222630
rect 280344 222566 280396 222572
rect 280724 222494 280752 231676
rect 281000 222970 281028 231676
rect 280988 222964 281040 222970
rect 280988 222906 281040 222912
rect 281368 222562 281396 231676
rect 281736 222766 281764 231676
rect 281724 222760 281776 222766
rect 281724 222702 281776 222708
rect 281356 222556 281408 222562
rect 281356 222498 281408 222504
rect 280712 222488 280764 222494
rect 280712 222430 280764 222436
rect 281448 221876 281500 221882
rect 281448 221818 281500 221824
rect 279976 221740 280028 221746
rect 279976 221682 280028 221688
rect 279792 221060 279844 221066
rect 279792 221002 279844 221008
rect 279804 217410 279832 221002
rect 280620 220924 280672 220930
rect 280620 220866 280672 220872
rect 280632 217410 280660 220866
rect 281460 217410 281488 221818
rect 282104 221474 282132 231676
rect 282092 221468 282144 221474
rect 282092 221410 282144 221416
rect 282472 221406 282500 231676
rect 282840 222834 282868 231676
rect 282828 222828 282880 222834
rect 282828 222770 282880 222776
rect 283104 222488 283156 222494
rect 283104 222430 283156 222436
rect 282460 221400 282512 221406
rect 282460 221342 282512 221348
rect 282368 221128 282420 221134
rect 282368 221070 282420 221076
rect 282380 217410 282408 221070
rect 283116 217410 283144 222430
rect 283208 221542 283236 231676
rect 283196 221536 283248 221542
rect 283196 221478 283248 221484
rect 283576 221270 283604 231676
rect 283852 221338 283880 231676
rect 284220 221814 284248 231676
rect 284588 222358 284616 231676
rect 284956 222562 284984 231676
rect 284944 222556 284996 222562
rect 284944 222498 284996 222504
rect 284576 222352 284628 222358
rect 284576 222294 284628 222300
rect 285324 221950 285352 231676
rect 285692 223106 285720 231676
rect 285680 223100 285732 223106
rect 285680 223042 285732 223048
rect 286060 222154 286088 231676
rect 286048 222148 286100 222154
rect 286048 222090 286100 222096
rect 285312 221944 285364 221950
rect 285312 221886 285364 221892
rect 284208 221808 284260 221814
rect 284208 221750 284260 221756
rect 284852 221740 284904 221746
rect 284852 221682 284904 221688
rect 283932 221468 283984 221474
rect 283932 221410 283984 221416
rect 283840 221332 283892 221338
rect 283840 221274 283892 221280
rect 283564 221264 283616 221270
rect 283564 221206 283616 221212
rect 283748 221196 283800 221202
rect 283748 221138 283800 221144
rect 283760 220998 283788 221138
rect 283748 220992 283800 220998
rect 283748 220934 283800 220940
rect 283944 217410 283972 221410
rect 284864 217410 284892 221682
rect 286428 221678 286456 231676
rect 286416 221672 286468 221678
rect 286416 221614 286468 221620
rect 286508 221536 286560 221542
rect 286508 221478 286560 221484
rect 285680 220992 285732 220998
rect 285680 220934 285732 220940
rect 285692 217410 285720 220934
rect 286520 217410 286548 221478
rect 286704 221270 286732 231676
rect 287072 222086 287100 231676
rect 287060 222080 287112 222086
rect 287060 222022 287112 222028
rect 287060 221944 287112 221950
rect 287060 221886 287112 221892
rect 286692 221264 286744 221270
rect 286692 221206 286744 221212
rect 287072 221134 287100 221886
rect 287440 221202 287468 231676
rect 287808 223582 287836 231676
rect 287796 223576 287848 223582
rect 287796 223518 287848 223524
rect 287428 221196 287480 221202
rect 287428 221138 287480 221144
rect 287060 221128 287112 221134
rect 287060 221070 287112 221076
rect 287336 221128 287388 221134
rect 287336 221070 287388 221076
rect 287348 217410 287376 221070
rect 288176 220930 288204 231676
rect 288544 221610 288572 231676
rect 288532 221604 288584 221610
rect 288532 221546 288584 221552
rect 288256 221468 288308 221474
rect 288256 221410 288308 221416
rect 288164 220924 288216 220930
rect 288164 220866 288216 220872
rect 288268 217410 288296 221410
rect 288912 221066 288940 231676
rect 289280 221950 289308 231676
rect 289268 221944 289320 221950
rect 289268 221886 289320 221892
rect 289084 221400 289136 221406
rect 289084 221342 289136 221348
rect 288900 221060 288952 221066
rect 288900 221002 288952 221008
rect 289096 217410 289124 221342
rect 289556 221338 289584 231676
rect 289924 221882 289952 231676
rect 290292 222494 290320 231676
rect 290280 222488 290332 222494
rect 290280 222430 290332 222436
rect 289912 221876 289964 221882
rect 289912 221818 289964 221824
rect 289544 221332 289596 221338
rect 289544 221274 289596 221280
rect 289728 221264 289780 221270
rect 289728 221206 289780 221212
rect 289740 217410 289768 221206
rect 290660 220998 290688 231676
rect 290740 226908 290792 226914
rect 290740 226850 290792 226856
rect 290648 220992 290700 220998
rect 290648 220934 290700 220940
rect 290752 217410 290780 226850
rect 291028 221134 291056 231676
rect 291396 221746 291424 231676
rect 291384 221740 291436 221746
rect 291384 221682 291436 221688
rect 291764 221542 291792 231676
rect 291752 221536 291804 221542
rect 291752 221478 291804 221484
rect 292132 221406 292160 231676
rect 292408 226914 292436 231676
rect 292396 226908 292448 226914
rect 292396 226850 292448 226856
rect 292776 221474 292804 231676
rect 292764 221468 292816 221474
rect 292764 221410 292816 221416
rect 292120 221400 292172 221406
rect 292120 221342 292172 221348
rect 292396 221400 292448 221406
rect 292396 221342 292448 221348
rect 291568 221332 291620 221338
rect 291568 221274 291620 221280
rect 291016 221128 291068 221134
rect 291016 221070 291068 221076
rect 291580 217410 291608 221274
rect 292408 217410 292436 221342
rect 293144 221270 293172 231676
rect 293224 229016 293276 229022
rect 293224 228958 293276 228964
rect 293132 221264 293184 221270
rect 293132 221206 293184 221212
rect 293236 217410 293264 228958
rect 293512 221406 293540 231676
rect 293500 221400 293552 221406
rect 293500 221342 293552 221348
rect 293880 217410 293908 231676
rect 294248 221338 294276 231676
rect 294616 229022 294644 231676
rect 294998 231662 295196 231690
rect 294604 229016 294656 229022
rect 294604 228958 294656 228964
rect 295168 226334 295196 231662
rect 295260 227322 295288 231676
rect 295248 227316 295300 227322
rect 295248 227258 295300 227264
rect 295168 226306 295380 226334
rect 294236 221332 294288 221338
rect 294236 221274 294288 221280
rect 294972 221332 295024 221338
rect 294972 221274 295024 221280
rect 294984 217410 295012 221274
rect 209608 217382 209668 217410
rect 210496 217382 210832 217410
rect 211416 217382 211752 217410
rect 212244 217382 212396 217410
rect 213072 217382 213408 217410
rect 213900 217382 214236 217410
rect 214728 217382 215064 217410
rect 215556 217382 215892 217410
rect 216384 217382 216720 217410
rect 217304 217382 217640 217410
rect 218132 217382 218468 217410
rect 218960 217382 219296 217410
rect 219788 217382 220124 217410
rect 220616 217382 220768 217410
rect 221444 217382 221780 217410
rect 222272 217382 222608 217410
rect 223192 217382 223528 217410
rect 224020 217382 224356 217410
rect 224848 217382 225184 217410
rect 225676 217382 226012 217410
rect 226504 217382 226840 217410
rect 227332 217382 227668 217410
rect 228160 217382 228496 217410
rect 229080 217382 229324 217410
rect 229908 217382 230244 217410
rect 230736 217382 231072 217410
rect 231564 217382 231716 217410
rect 232392 217382 232728 217410
rect 233220 217382 233556 217410
rect 234048 217382 234384 217410
rect 234968 217382 235304 217410
rect 235796 217382 236132 217410
rect 236624 217382 236960 217410
rect 237452 217382 237788 217410
rect 238280 217382 238616 217410
rect 239108 217382 239444 217410
rect 239936 217382 240088 217410
rect 240856 217382 241192 217410
rect 241684 217382 242020 217410
rect 242512 217382 242848 217410
rect 243340 217382 243584 217410
rect 244168 217382 244504 217410
rect 244996 217382 245332 217410
rect 245824 217382 246160 217410
rect 246744 217382 247080 217410
rect 247572 217382 247908 217410
rect 248400 217382 248736 217410
rect 249228 217382 249564 217410
rect 250056 217382 250392 217410
rect 250884 217382 251128 217410
rect 251712 217382 252048 217410
rect 252632 217382 252968 217410
rect 253460 217382 253796 217410
rect 254288 217382 254624 217410
rect 255116 217382 255452 217410
rect 255944 217382 256280 217410
rect 256772 217382 257108 217410
rect 257600 217382 257936 217410
rect 258520 217382 258856 217410
rect 259348 217382 259408 217410
rect 260176 217382 260512 217410
rect 261004 217382 261340 217410
rect 261832 217382 262168 217410
rect 262660 217382 262996 217410
rect 263488 217382 263824 217410
rect 264408 217382 264652 217410
rect 265236 217382 265572 217410
rect 266064 217382 266400 217410
rect 266892 217382 267228 217410
rect 267720 217382 268056 217410
rect 268548 217382 268884 217410
rect 269376 217382 269712 217410
rect 270296 217382 270448 217410
rect 271124 217382 271460 217410
rect 271952 217382 272288 217410
rect 272780 217382 273116 217410
rect 273608 217382 273944 217410
rect 274436 217382 274772 217410
rect 275264 217382 275600 217410
rect 276184 217382 276520 217410
rect 277012 217382 277348 217410
rect 277840 217382 278176 217410
rect 278668 217382 278728 217410
rect 279496 217382 279832 217410
rect 280324 217382 280660 217410
rect 281152 217382 281488 217410
rect 282072 217382 282408 217410
rect 282900 217382 283144 217410
rect 283728 217382 283972 217410
rect 284556 217382 284892 217410
rect 285384 217382 285720 217410
rect 286212 217382 286548 217410
rect 287040 217382 287376 217410
rect 287960 217382 288296 217410
rect 288788 217382 289124 217410
rect 289616 217382 289768 217410
rect 290444 217382 290780 217410
rect 291272 217382 291608 217410
rect 292100 217382 292436 217410
rect 292928 217382 293264 217410
rect 293848 217382 293908 217410
rect 294676 217382 295012 217410
rect 295352 217410 295380 226306
rect 295628 221338 295656 231676
rect 295616 221332 295668 221338
rect 295616 221274 295668 221280
rect 295996 217410 296024 231676
rect 296364 229090 296392 231676
rect 296352 229084 296404 229090
rect 296352 229026 296404 229032
rect 296732 228954 296760 231676
rect 297114 231662 297404 231690
rect 296720 228948 296772 228954
rect 296720 228890 296772 228896
rect 296812 227316 296864 227322
rect 296812 227258 296864 227264
rect 296824 217410 296852 227258
rect 297376 226334 297404 231662
rect 297468 229022 297496 231676
rect 297456 229016 297508 229022
rect 297456 228958 297508 228964
rect 297836 226710 297864 231676
rect 298112 226982 298140 231676
rect 298494 231662 298784 231690
rect 298468 229084 298520 229090
rect 298468 229026 298520 229032
rect 298100 226976 298152 226982
rect 298100 226918 298152 226924
rect 297824 226704 297876 226710
rect 297824 226646 297876 226652
rect 297376 226306 297588 226334
rect 297560 217410 297588 226306
rect 298480 217410 298508 229026
rect 298756 227322 298784 231662
rect 298848 229090 298876 231676
rect 298836 229084 298888 229090
rect 298836 229026 298888 229032
rect 298744 227316 298796 227322
rect 298744 227258 298796 227264
rect 299216 226778 299244 231676
rect 299388 229016 299440 229022
rect 299388 228958 299440 228964
rect 299204 226772 299256 226778
rect 299204 226714 299256 226720
rect 299400 217410 299428 228958
rect 299584 226846 299612 231676
rect 299572 226840 299624 226846
rect 299572 226782 299624 226788
rect 299952 226370 299980 231676
rect 300216 228948 300268 228954
rect 300216 228890 300268 228896
rect 299940 226364 299992 226370
rect 299940 226306 299992 226312
rect 300228 217410 300256 228890
rect 300320 226642 300348 231676
rect 300688 226914 300716 231676
rect 300964 228274 300992 231676
rect 300952 228268 301004 228274
rect 300952 228210 301004 228216
rect 301044 227316 301096 227322
rect 301044 227258 301096 227264
rect 300676 226908 300728 226914
rect 300676 226850 300728 226856
rect 300308 226636 300360 226642
rect 300308 226578 300360 226584
rect 301056 217410 301084 227258
rect 301332 226574 301360 231676
rect 301700 227934 301728 231676
rect 301688 227928 301740 227934
rect 301688 227870 301740 227876
rect 302068 227254 302096 231676
rect 302436 227322 302464 231676
rect 302700 229084 302752 229090
rect 302700 229026 302752 229032
rect 302424 227316 302476 227322
rect 302424 227258 302476 227264
rect 302056 227248 302108 227254
rect 302056 227190 302108 227196
rect 301964 226976 302016 226982
rect 301964 226918 302016 226924
rect 301976 226710 302004 226918
rect 301872 226704 301924 226710
rect 301872 226646 301924 226652
rect 301964 226704 302016 226710
rect 301964 226646 302016 226652
rect 301320 226568 301372 226574
rect 301320 226510 301372 226516
rect 301884 217410 301912 226646
rect 302712 217410 302740 229026
rect 302804 228410 302832 231676
rect 302792 228404 302844 228410
rect 302792 228346 302844 228352
rect 303172 227390 303200 231676
rect 303540 229022 303568 231676
rect 303528 229016 303580 229022
rect 303528 228958 303580 228964
rect 303816 227458 303844 231676
rect 304184 229090 304212 231676
rect 304172 229084 304224 229090
rect 304172 229026 304224 229032
rect 304552 228954 304580 231676
rect 304540 228948 304592 228954
rect 304540 228890 304592 228896
rect 304920 228682 304948 231676
rect 304908 228676 304960 228682
rect 304908 228618 304960 228624
rect 305288 227526 305316 231676
rect 305656 228818 305684 231676
rect 305644 228812 305696 228818
rect 305644 228754 305696 228760
rect 306024 227662 306052 231676
rect 306012 227656 306064 227662
rect 306012 227598 306064 227604
rect 305276 227520 305328 227526
rect 305276 227462 305328 227468
rect 303804 227452 303856 227458
rect 303804 227394 303856 227400
rect 303160 227384 303212 227390
rect 303160 227326 303212 227332
rect 306392 227118 306420 231676
rect 306668 228750 306696 231676
rect 306656 228744 306708 228750
rect 306656 228686 306708 228692
rect 307036 228206 307064 231676
rect 307404 228614 307432 231676
rect 307392 228608 307444 228614
rect 307392 228550 307444 228556
rect 307772 228478 307800 231676
rect 307760 228472 307812 228478
rect 307760 228414 307812 228420
rect 308140 228342 308168 231676
rect 308508 228886 308536 231676
rect 308496 228880 308548 228886
rect 308496 228822 308548 228828
rect 308876 228546 308904 231676
rect 308864 228540 308916 228546
rect 308864 228482 308916 228488
rect 308128 228336 308180 228342
rect 308128 228278 308180 228284
rect 307024 228200 307076 228206
rect 307024 228142 307076 228148
rect 309244 227186 309272 231676
rect 309520 228138 309548 231676
rect 309508 228132 309560 228138
rect 309508 228074 309560 228080
rect 309416 227928 309468 227934
rect 309416 227870 309468 227876
rect 309232 227180 309284 227186
rect 309232 227122 309284 227128
rect 306380 227112 306432 227118
rect 306380 227054 306432 227060
rect 308588 226908 308640 226914
rect 308588 226850 308640 226856
rect 306932 226840 306984 226846
rect 306932 226782 306984 226788
rect 305276 226772 305328 226778
rect 305276 226714 305328 226720
rect 303620 226704 303672 226710
rect 303620 226646 303672 226652
rect 303632 217410 303660 226646
rect 304356 226364 304408 226370
rect 304356 226306 304408 226312
rect 304368 217410 304396 226306
rect 305288 217410 305316 226714
rect 306380 226636 306432 226642
rect 306380 226578 306432 226584
rect 306392 217410 306420 226578
rect 306944 217410 306972 226782
rect 307760 226568 307812 226574
rect 307760 226510 307812 226516
rect 307772 217410 307800 226510
rect 308600 217410 308628 226850
rect 309428 217410 309456 227870
rect 309888 226370 309916 231676
rect 310270 231662 310560 231690
rect 310244 228268 310296 228274
rect 310244 228210 310296 228216
rect 309876 226364 309928 226370
rect 309876 226306 309928 226312
rect 310256 217410 310284 228210
rect 310532 226982 310560 231662
rect 310624 227934 310652 231676
rect 310612 227928 310664 227934
rect 310612 227870 310664 227876
rect 310520 226976 310572 226982
rect 310520 226918 310572 226924
rect 310992 222290 311020 231676
rect 311164 228404 311216 228410
rect 311164 228346 311216 228352
rect 310980 222284 311032 222290
rect 310980 222226 311032 222232
rect 311176 217410 311204 228346
rect 311360 228002 311388 231676
rect 311728 228070 311756 231676
rect 311716 228064 311768 228070
rect 311716 228006 311768 228012
rect 311348 227996 311400 228002
rect 311348 227938 311400 227944
rect 312096 227866 312124 231676
rect 312084 227860 312136 227866
rect 312084 227802 312136 227808
rect 311992 227248 312044 227254
rect 311992 227190 312044 227196
rect 312004 217410 312032 227190
rect 312372 222222 312400 231676
rect 312740 227798 312768 231676
rect 312728 227792 312780 227798
rect 312728 227734 312780 227740
rect 312820 227384 312872 227390
rect 312820 227326 312872 227332
rect 312360 222216 312412 222222
rect 312360 222158 312412 222164
rect 312832 217410 312860 227326
rect 313108 221202 313136 231676
rect 313476 225214 313504 231676
rect 313648 227316 313700 227322
rect 313648 227258 313700 227264
rect 313464 225208 313516 225214
rect 313464 225150 313516 225156
rect 313096 221196 313148 221202
rect 313096 221138 313148 221144
rect 313660 217410 313688 227258
rect 313844 221338 313872 231676
rect 314212 221406 314240 231676
rect 314580 221474 314608 231676
rect 314660 229084 314712 229090
rect 314660 229026 314712 229032
rect 314568 221468 314620 221474
rect 314568 221410 314620 221416
rect 314200 221400 314252 221406
rect 314200 221342 314252 221348
rect 313832 221332 313884 221338
rect 313832 221274 313884 221280
rect 314672 217410 314700 229026
rect 314948 225146 314976 231676
rect 314936 225140 314988 225146
rect 314936 225082 314988 225088
rect 315224 221542 315252 231676
rect 315304 229016 315356 229022
rect 315304 228958 315356 228964
rect 315212 221536 315264 221542
rect 315212 221478 315264 221484
rect 315316 217410 315344 228958
rect 315592 221270 315620 231676
rect 315960 227730 315988 231676
rect 316132 228948 316184 228954
rect 316132 228890 316184 228896
rect 315948 227724 316000 227730
rect 315948 227666 316000 227672
rect 315580 221264 315632 221270
rect 315580 221206 315632 221212
rect 316144 217410 316172 228890
rect 316328 224942 316356 231676
rect 316316 224936 316368 224942
rect 316316 224878 316368 224884
rect 316696 221746 316724 231676
rect 316684 221740 316736 221746
rect 316684 221682 316736 221688
rect 317064 221678 317092 231676
rect 317432 228410 317460 231676
rect 317420 228404 317472 228410
rect 317420 228346 317472 228352
rect 317420 227452 317472 227458
rect 317420 227394 317472 227400
rect 317052 221672 317104 221678
rect 317052 221614 317104 221620
rect 317432 217410 317460 227394
rect 317800 225078 317828 231676
rect 317880 228812 317932 228818
rect 317880 228754 317932 228760
rect 317788 225072 317840 225078
rect 317788 225014 317840 225020
rect 295352 217382 295504 217410
rect 295996 217382 296332 217410
rect 296824 217382 297160 217410
rect 297560 217382 297988 217410
rect 298480 217382 298816 217410
rect 299400 217382 299736 217410
rect 300228 217382 300564 217410
rect 301056 217382 301392 217410
rect 301884 217382 302220 217410
rect 302712 217382 303048 217410
rect 303632 217382 303876 217410
rect 304368 217382 304704 217410
rect 305288 217382 305624 217410
rect 306392 217382 306452 217410
rect 306944 217382 307280 217410
rect 307772 217382 308108 217410
rect 308600 217382 308936 217410
rect 309428 217382 309764 217410
rect 310256 217382 310592 217410
rect 311176 217382 311512 217410
rect 312004 217382 312340 217410
rect 312832 217382 313168 217410
rect 313660 217382 313996 217410
rect 314672 217382 314824 217410
rect 315316 217382 315652 217410
rect 316144 217382 316480 217410
rect 317400 217382 317460 217410
rect 317892 217410 317920 228754
rect 318076 221950 318104 231676
rect 318064 221944 318116 221950
rect 318064 221886 318116 221892
rect 318444 221610 318472 231676
rect 318812 229022 318840 231676
rect 318800 229016 318852 229022
rect 318800 228958 318852 228964
rect 318708 228676 318760 228682
rect 318708 228618 318760 228624
rect 318432 221604 318484 221610
rect 318432 221546 318484 221552
rect 318720 217410 318748 228618
rect 319180 225010 319208 231676
rect 319562 231662 319852 231690
rect 319536 227656 319588 227662
rect 319536 227598 319588 227604
rect 319168 225004 319220 225010
rect 319168 224946 319220 224952
rect 319548 217410 319576 227598
rect 319824 222018 319852 231662
rect 319812 222012 319864 222018
rect 319812 221954 319864 221960
rect 319916 221882 319944 231676
rect 320284 227594 320312 231676
rect 320272 227588 320324 227594
rect 320272 227530 320324 227536
rect 320652 227526 320680 231676
rect 320364 227520 320416 227526
rect 320364 227462 320416 227468
rect 320640 227520 320692 227526
rect 320640 227462 320692 227468
rect 319904 221876 319956 221882
rect 319904 221818 319956 221824
rect 320376 217410 320404 227462
rect 320928 222086 320956 231676
rect 321192 228200 321244 228206
rect 321192 228142 321244 228148
rect 320916 222080 320968 222086
rect 320916 222022 320968 222028
rect 321204 217410 321232 228142
rect 321296 221814 321324 231676
rect 321664 227458 321692 231676
rect 322032 227662 322060 231676
rect 322020 227656 322072 227662
rect 322020 227598 322072 227604
rect 321652 227452 321704 227458
rect 321652 227394 321704 227400
rect 322020 227112 322072 227118
rect 322020 227054 322072 227060
rect 321284 221808 321336 221814
rect 321284 221750 321336 221756
rect 322032 217410 322060 227054
rect 322400 223514 322428 231676
rect 322388 223508 322440 223514
rect 322388 223450 322440 223456
rect 322768 222154 322796 231676
rect 322940 228608 322992 228614
rect 322940 228550 322992 228556
rect 322756 222148 322808 222154
rect 322756 222090 322808 222096
rect 322952 217410 322980 228550
rect 323136 227390 323164 231676
rect 323504 228682 323532 231676
rect 323492 228676 323544 228682
rect 323492 228618 323544 228624
rect 323124 227384 323176 227390
rect 323124 227326 323176 227332
rect 323780 223038 323808 231676
rect 323860 228744 323912 228750
rect 323860 228686 323912 228692
rect 323768 223032 323820 223038
rect 323768 222974 323820 222980
rect 323872 217410 323900 228686
rect 324148 223446 324176 231676
rect 324516 223582 324544 231676
rect 324596 228880 324648 228886
rect 324596 228822 324648 228828
rect 324504 223576 324556 223582
rect 324504 223518 324556 223524
rect 324136 223440 324188 223446
rect 324136 223382 324188 223388
rect 324608 217410 324636 228822
rect 324884 223378 324912 231676
rect 324872 223372 324924 223378
rect 324872 223314 324924 223320
rect 325252 222902 325280 231676
rect 325620 223174 325648 231676
rect 325700 228472 325752 228478
rect 325700 228414 325752 228420
rect 325608 223168 325660 223174
rect 325608 223110 325660 223116
rect 325240 222896 325292 222902
rect 325240 222838 325292 222844
rect 325712 217410 325740 228414
rect 325988 227322 326016 231676
rect 326252 228540 326304 228546
rect 326252 228482 326304 228488
rect 325976 227316 326028 227322
rect 325976 227258 326028 227264
rect 326264 217410 326292 228482
rect 326356 223242 326384 231676
rect 326344 223236 326396 223242
rect 326344 223178 326396 223184
rect 326632 222834 326660 231676
rect 327000 223310 327028 231676
rect 327080 228336 327132 228342
rect 327080 228278 327132 228284
rect 326988 223304 327040 223310
rect 326988 223246 327040 223252
rect 326620 222828 326672 222834
rect 326620 222770 326672 222776
rect 327092 217410 327120 228278
rect 327368 222970 327396 231676
rect 327356 222964 327408 222970
rect 327356 222906 327408 222912
rect 327736 222766 327764 231676
rect 327908 226364 327960 226370
rect 327908 226306 327960 226312
rect 327724 222760 327776 222766
rect 327724 222702 327776 222708
rect 327920 217410 327948 226306
rect 328104 222426 328132 231676
rect 328472 223106 328500 231676
rect 328854 231662 329144 231690
rect 328828 227180 328880 227186
rect 328828 227122 328880 227128
rect 328460 223100 328512 223106
rect 328460 223042 328512 223048
rect 328092 222420 328144 222426
rect 328092 222362 328144 222368
rect 328840 217410 328868 227122
rect 329116 226710 329144 231662
rect 329208 228410 329236 231676
rect 329196 228404 329248 228410
rect 329196 228346 329248 228352
rect 329104 226704 329156 226710
rect 329104 226646 329156 226652
rect 329484 222698 329512 231676
rect 329656 226976 329708 226982
rect 329656 226918 329708 226924
rect 329472 222692 329524 222698
rect 329472 222634 329524 222640
rect 329668 217410 329696 226918
rect 329852 222630 329880 231676
rect 329840 222624 329892 222630
rect 329840 222566 329892 222572
rect 330220 221134 330248 231676
rect 330588 228274 330616 231676
rect 330576 228268 330628 228274
rect 330576 228210 330628 228216
rect 330484 228132 330536 228138
rect 330484 228074 330536 228080
rect 330208 221128 330260 221134
rect 330208 221070 330260 221076
rect 330496 217410 330524 228074
rect 330956 222737 330984 231676
rect 331338 231662 331628 231690
rect 331312 227996 331364 228002
rect 331312 227938 331364 227944
rect 330942 222728 330998 222737
rect 330942 222663 330998 222672
rect 331324 217410 331352 227938
rect 331600 222562 331628 231662
rect 331692 227186 331720 231676
rect 332060 228478 332088 231676
rect 332048 228472 332100 228478
rect 332048 228414 332100 228420
rect 332140 227928 332192 227934
rect 332140 227870 332192 227876
rect 331680 227180 331732 227186
rect 331680 227122 331732 227128
rect 331588 222556 331640 222562
rect 331588 222498 331640 222504
rect 332152 217410 332180 227870
rect 332336 222601 332364 231676
rect 332322 222592 332378 222601
rect 332322 222527 332378 222536
rect 332704 222358 332732 231676
rect 332968 228064 333020 228070
rect 332968 228006 333020 228012
rect 332692 222352 332744 222358
rect 332692 222294 332744 222300
rect 332980 217410 333008 228006
rect 333072 222465 333100 231676
rect 333440 228138 333468 231676
rect 333428 228132 333480 228138
rect 333428 228074 333480 228080
rect 333058 222456 333114 222465
rect 333058 222391 333114 222400
rect 333808 222329 333836 231676
rect 333794 222320 333850 222329
rect 333794 222255 333850 222264
rect 333980 222284 334032 222290
rect 333980 222226 334032 222232
rect 333992 217410 334020 222226
rect 334176 220998 334204 231676
rect 334544 221649 334572 231676
rect 334912 228342 334940 231676
rect 335188 228546 335216 231676
rect 335570 231662 335860 231690
rect 335176 228540 335228 228546
rect 335176 228482 335228 228488
rect 334900 228336 334952 228342
rect 334900 228278 334952 228284
rect 335544 227860 335596 227866
rect 335544 227802 335596 227808
rect 334716 227792 334768 227798
rect 334716 227734 334768 227740
rect 334530 221640 334586 221649
rect 334530 221575 334586 221584
rect 334164 220992 334216 220998
rect 334164 220934 334216 220940
rect 334728 217410 334756 227734
rect 335556 217410 335584 227802
rect 335832 221785 335860 231662
rect 335924 222193 335952 231676
rect 336292 228954 336320 231676
rect 336280 228948 336332 228954
rect 336280 228890 336332 228896
rect 336660 228614 336688 231676
rect 336648 228608 336700 228614
rect 336648 228550 336700 228556
rect 337028 228070 337056 231676
rect 337016 228064 337068 228070
rect 337016 228006 337068 228012
rect 337200 222216 337252 222222
rect 335910 222184 335966 222193
rect 337200 222158 337252 222164
rect 335910 222119 335966 222128
rect 335818 221776 335874 221785
rect 335818 221711 335874 221720
rect 336740 221196 336792 221202
rect 336740 221138 336792 221144
rect 336752 217410 336780 221138
rect 317892 217382 318228 217410
rect 318720 217382 319056 217410
rect 319548 217382 319884 217410
rect 320376 217382 320712 217410
rect 321204 217382 321540 217410
rect 322032 217382 322368 217410
rect 322952 217382 323288 217410
rect 323872 217382 324116 217410
rect 324608 217382 324944 217410
rect 325712 217382 325772 217410
rect 326264 217382 326600 217410
rect 327092 217382 327428 217410
rect 327920 217382 328256 217410
rect 328840 217382 329176 217410
rect 329668 217382 330004 217410
rect 330496 217382 330832 217410
rect 331324 217382 331660 217410
rect 332152 217382 332488 217410
rect 332980 217382 333316 217410
rect 333992 217382 334144 217410
rect 334728 217382 335064 217410
rect 335556 217382 335892 217410
rect 336720 217382 336780 217410
rect 337212 217410 337240 222158
rect 337396 221202 337424 231676
rect 337764 228750 337792 231676
rect 337752 228744 337804 228750
rect 337752 228686 337804 228692
rect 337660 228200 337712 228206
rect 337660 228142 337712 228148
rect 337672 222290 337700 228142
rect 338040 227050 338068 231676
rect 338408 227934 338436 231676
rect 338396 227928 338448 227934
rect 338396 227870 338448 227876
rect 338304 227724 338356 227730
rect 338304 227666 338356 227672
rect 338028 227044 338080 227050
rect 338028 226986 338080 226992
rect 338316 222494 338344 227666
rect 338304 222488 338356 222494
rect 338304 222430 338356 222436
rect 338028 222420 338080 222426
rect 338212 222420 338264 222426
rect 338080 222380 338212 222408
rect 338028 222362 338080 222368
rect 338212 222362 338264 222368
rect 337660 222284 337712 222290
rect 337660 222226 337712 222232
rect 338776 221921 338804 231676
rect 339144 229090 339172 231676
rect 339132 229084 339184 229090
rect 339132 229026 339184 229032
rect 339512 228206 339540 231676
rect 339500 228200 339552 228206
rect 339500 228142 339552 228148
rect 339880 225214 339908 231676
rect 338856 225208 338908 225214
rect 338856 225150 338908 225156
rect 339868 225208 339920 225214
rect 339868 225150 339920 225156
rect 338762 221912 338818 221921
rect 338762 221847 338818 221856
rect 338028 221400 338080 221406
rect 338028 221342 338080 221348
rect 337384 221196 337436 221202
rect 337384 221138 337436 221144
rect 338040 217410 338068 221342
rect 338868 217410 338896 225150
rect 340248 224126 340276 231676
rect 340616 228818 340644 231676
rect 340892 228886 340920 231676
rect 340972 229016 341024 229022
rect 340972 228958 341024 228964
rect 340880 228880 340932 228886
rect 340880 228822 340932 228828
rect 340604 228812 340656 228818
rect 340604 228754 340656 228760
rect 340236 224120 340288 224126
rect 340236 224062 340288 224068
rect 340984 222222 341012 228958
rect 341260 228002 341288 231676
rect 341248 227996 341300 228002
rect 341248 227938 341300 227944
rect 341628 227866 341656 231676
rect 341616 227860 341668 227866
rect 341616 227802 341668 227808
rect 341996 227798 342024 231676
rect 342364 229022 342392 231676
rect 342352 229016 342404 229022
rect 342352 228958 342404 228964
rect 341984 227792 342036 227798
rect 341984 227734 342036 227740
rect 342076 227588 342128 227594
rect 342076 227530 342128 227536
rect 340972 222216 341024 222222
rect 340972 222158 341024 222164
rect 339684 221468 339736 221474
rect 339684 221410 339736 221416
rect 339696 217410 339724 221410
rect 342088 221338 342116 227530
rect 342536 225140 342588 225146
rect 342536 225082 342588 225088
rect 340604 221332 340656 221338
rect 340604 221274 340656 221280
rect 342076 221332 342128 221338
rect 342076 221274 342128 221280
rect 340616 217410 340644 221274
rect 341432 221264 341484 221270
rect 341432 221206 341484 221212
rect 341444 217410 341472 221206
rect 342548 217410 342576 225082
rect 342732 224602 342760 231676
rect 342904 227452 342956 227458
rect 342904 227394 342956 227400
rect 342720 224596 342772 224602
rect 342720 224538 342772 224544
rect 342916 221406 342944 227394
rect 342996 227384 343048 227390
rect 342996 227326 343048 227332
rect 342904 221400 342956 221406
rect 342904 221342 342956 221348
rect 343008 221066 343036 227326
rect 343100 225282 343128 231676
rect 343088 225276 343140 225282
rect 343088 225218 343140 225224
rect 343088 222488 343140 222494
rect 343088 222430 343140 222436
rect 342996 221060 343048 221066
rect 342996 221002 343048 221008
rect 343100 217410 343128 222430
rect 343468 219298 343496 231676
rect 343744 227594 343772 231676
rect 343732 227588 343784 227594
rect 343732 227530 343784 227536
rect 344112 224194 344140 231676
rect 344480 227730 344508 231676
rect 344468 227724 344520 227730
rect 344468 227666 344520 227672
rect 344100 224188 344152 224194
rect 344100 224130 344152 224136
rect 343548 222488 343600 222494
rect 343548 222430 343600 222436
rect 343560 221134 343588 222430
rect 343916 221536 343968 221542
rect 343916 221478 343968 221484
rect 343548 221128 343600 221134
rect 343548 221070 343600 221076
rect 343456 219292 343508 219298
rect 343456 219234 343508 219240
rect 343928 217410 343956 221478
rect 344848 220794 344876 231676
rect 345112 226704 345164 226710
rect 345112 226646 345164 226652
rect 345124 221678 345152 226646
rect 345216 224330 345244 231676
rect 345296 227316 345348 227322
rect 345296 227258 345348 227264
rect 345204 224324 345256 224330
rect 345204 224266 345256 224272
rect 345020 221672 345072 221678
rect 345020 221614 345072 221620
rect 345112 221672 345164 221678
rect 345112 221614 345164 221620
rect 344836 220788 344888 220794
rect 344836 220730 344888 220736
rect 345032 217410 345060 221614
rect 345308 221542 345336 227258
rect 345584 224262 345612 231676
rect 345952 231198 345980 231676
rect 345940 231192 345992 231198
rect 345940 231134 345992 231140
rect 345664 224936 345716 224942
rect 345664 224878 345716 224884
rect 345572 224256 345624 224262
rect 345572 224198 345624 224204
rect 345296 221536 345348 221542
rect 345296 221478 345348 221484
rect 345676 217410 345704 224878
rect 346320 219366 346348 231676
rect 346596 224942 346624 231676
rect 346584 224936 346636 224942
rect 346584 224878 346636 224884
rect 346964 224466 346992 231676
rect 347332 231062 347360 231676
rect 347320 231056 347372 231062
rect 347320 230998 347372 231004
rect 346952 224460 347004 224466
rect 346952 224402 347004 224408
rect 346492 222284 346544 222290
rect 346492 222226 346544 222232
rect 346584 222284 346636 222290
rect 346584 222226 346636 222232
rect 346308 219360 346360 219366
rect 346308 219302 346360 219308
rect 346504 217410 346532 222226
rect 346596 220998 346624 222226
rect 347320 221740 347372 221746
rect 347320 221682 347372 221688
rect 346584 220992 346636 220998
rect 346584 220934 346636 220940
rect 347332 217410 347360 221682
rect 347700 220658 347728 231676
rect 347780 227180 347832 227186
rect 347780 227122 347832 227128
rect 347792 221746 347820 227122
rect 348068 224534 348096 231676
rect 348056 224528 348108 224534
rect 348056 224470 348108 224476
rect 348436 224398 348464 231676
rect 348804 230926 348832 231676
rect 348792 230920 348844 230926
rect 348792 230862 348844 230868
rect 348976 225072 349028 225078
rect 348976 225014 349028 225020
rect 348424 224392 348476 224398
rect 348424 224334 348476 224340
rect 347780 221740 347832 221746
rect 347780 221682 347832 221688
rect 348148 221604 348200 221610
rect 348148 221546 348200 221552
rect 347688 220652 347740 220658
rect 347688 220594 347740 220600
rect 348160 217410 348188 221546
rect 348988 217410 349016 225014
rect 349172 220726 349200 231676
rect 349448 226302 349476 231676
rect 349436 226296 349488 226302
rect 349436 226238 349488 226244
rect 349816 224670 349844 231676
rect 350184 227322 350212 231676
rect 350172 227316 350224 227322
rect 350172 227258 350224 227264
rect 349804 224664 349856 224670
rect 349804 224606 349856 224612
rect 349804 222216 349856 222222
rect 349804 222158 349856 222164
rect 349896 222216 349948 222222
rect 349896 222158 349948 222164
rect 349160 220720 349212 220726
rect 349160 220662 349212 220668
rect 349816 217410 349844 222158
rect 349908 221202 349936 222158
rect 349896 221196 349948 221202
rect 349896 221138 349948 221144
rect 350552 220590 350580 231676
rect 350920 224874 350948 231676
rect 350908 224868 350960 224874
rect 350908 224810 350960 224816
rect 351288 224738 351316 231676
rect 351656 230858 351684 231676
rect 351644 230852 351696 230858
rect 351644 230794 351696 230800
rect 351276 224732 351328 224738
rect 351276 224674 351328 224680
rect 350632 221944 350684 221950
rect 350632 221886 350684 221892
rect 350540 220584 350592 220590
rect 350540 220526 350592 220532
rect 350644 217410 350672 221886
rect 351460 221876 351512 221882
rect 351460 221818 351512 221824
rect 351472 217410 351500 221818
rect 352024 220522 352052 231676
rect 352300 226098 352328 231676
rect 352668 226234 352696 231676
rect 353036 227186 353064 231676
rect 353024 227180 353076 227186
rect 353024 227122 353076 227128
rect 352656 226228 352708 226234
rect 352656 226170 352708 226176
rect 352288 226092 352340 226098
rect 352288 226034 352340 226040
rect 352380 225004 352432 225010
rect 352380 224946 352432 224952
rect 352012 220516 352064 220522
rect 352012 220458 352064 220464
rect 352392 217410 352420 224946
rect 353300 221332 353352 221338
rect 353300 221274 353352 221280
rect 353312 217410 353340 221274
rect 353404 220454 353432 231676
rect 353772 226166 353800 231676
rect 353760 226160 353812 226166
rect 353760 226102 353812 226108
rect 354140 224806 354168 231676
rect 354508 230790 354536 231676
rect 354890 231662 355088 231690
rect 354496 230784 354548 230790
rect 354496 230726 354548 230732
rect 354128 224800 354180 224806
rect 354128 224742 354180 224748
rect 354036 222012 354088 222018
rect 354036 221954 354088 221960
rect 353392 220448 353444 220454
rect 353392 220390 353444 220396
rect 354048 217410 354076 221954
rect 354864 221808 354916 221814
rect 354864 221750 354916 221756
rect 354876 217410 354904 221750
rect 355060 220318 355088 231662
rect 355152 225418 355180 231676
rect 355520 225962 355548 231676
rect 355888 231130 355916 231676
rect 355876 231124 355928 231130
rect 355876 231066 355928 231072
rect 356256 230994 356284 231676
rect 356244 230988 356296 230994
rect 356244 230930 356296 230936
rect 356060 227520 356112 227526
rect 356060 227462 356112 227468
rect 355508 225956 355560 225962
rect 355508 225898 355560 225904
rect 355140 225412 355192 225418
rect 355140 225354 355192 225360
rect 355048 220312 355100 220318
rect 355048 220254 355100 220260
rect 356072 217410 356100 227462
rect 356624 225894 356652 231676
rect 356992 226030 357020 231676
rect 357374 231662 357664 231690
rect 356980 226024 357032 226030
rect 356980 225966 357032 225972
rect 356612 225888 356664 225894
rect 356612 225830 356664 225836
rect 357348 222080 357400 222086
rect 357348 222022 357400 222028
rect 356520 221400 356572 221406
rect 356520 221342 356572 221348
rect 337212 217382 337548 217410
rect 338040 217382 338376 217410
rect 338868 217382 339204 217410
rect 339696 217382 340032 217410
rect 340616 217382 340952 217410
rect 341444 217382 341780 217410
rect 342548 217382 342608 217410
rect 343100 217382 343436 217410
rect 343928 217382 344264 217410
rect 345032 217382 345092 217410
rect 345676 217382 345920 217410
rect 346504 217382 346840 217410
rect 347332 217382 347668 217410
rect 348160 217382 348496 217410
rect 348988 217382 349324 217410
rect 349816 217382 350152 217410
rect 350644 217382 350980 217410
rect 351472 217382 351808 217410
rect 352392 217382 352728 217410
rect 353312 217382 353556 217410
rect 354048 217382 354384 217410
rect 354876 217382 355212 217410
rect 356040 217382 356100 217410
rect 356532 217410 356560 221342
rect 357360 217410 357388 222022
rect 357636 220386 357664 231662
rect 357728 230314 357756 231676
rect 357716 230308 357768 230314
rect 357716 230250 357768 230256
rect 358004 225078 358032 231676
rect 358372 225146 358400 231676
rect 358740 227118 358768 231676
rect 359108 230382 359136 231676
rect 359096 230376 359148 230382
rect 359096 230318 359148 230324
rect 359096 227656 359148 227662
rect 359096 227598 359148 227604
rect 358728 227112 358780 227118
rect 358728 227054 358780 227060
rect 358360 225140 358412 225146
rect 358360 225082 358412 225088
rect 357992 225072 358044 225078
rect 357992 225014 358044 225020
rect 358268 222148 358320 222154
rect 358268 222090 358320 222096
rect 357624 220380 357676 220386
rect 357624 220322 357676 220328
rect 358280 217410 358308 222090
rect 359108 217410 359136 227598
rect 359476 225826 359504 231676
rect 359844 226846 359872 231676
rect 359832 226840 359884 226846
rect 359832 226782 359884 226788
rect 359464 225820 359516 225826
rect 359464 225762 359516 225768
rect 359924 221060 359976 221066
rect 359924 221002 359976 221008
rect 359936 217410 359964 221002
rect 360212 220250 360240 231676
rect 360580 230110 360608 231676
rect 360568 230104 360620 230110
rect 360568 230046 360620 230052
rect 360856 225690 360884 231676
rect 360844 225684 360896 225690
rect 360844 225626 360896 225632
rect 361224 225010 361252 231676
rect 361592 226914 361620 231676
rect 361960 230178 361988 231676
rect 361948 230172 362000 230178
rect 361948 230114 362000 230120
rect 361580 226908 361632 226914
rect 361580 226850 361632 226856
rect 362328 225758 362356 231676
rect 362408 228676 362460 228682
rect 362408 228618 362460 228624
rect 362316 225752 362368 225758
rect 362316 225694 362368 225700
rect 361212 225004 361264 225010
rect 361212 224946 361264 224952
rect 360752 223508 360804 223514
rect 360752 223450 360804 223456
rect 360200 220244 360252 220250
rect 360200 220186 360252 220192
rect 360764 217410 360792 223450
rect 361764 223440 361816 223446
rect 361764 223382 361816 223388
rect 361776 217410 361804 223382
rect 362420 217410 362448 228618
rect 362696 225622 362724 231676
rect 363064 230246 363092 231676
rect 363052 230240 363104 230246
rect 363052 230182 363104 230188
rect 363432 229974 363460 231676
rect 363420 229968 363472 229974
rect 363420 229910 363472 229916
rect 362684 225616 362736 225622
rect 362684 225558 362736 225564
rect 363708 225486 363736 231676
rect 364076 229906 364104 231676
rect 364064 229900 364116 229906
rect 364064 229842 364116 229848
rect 364444 226982 364472 231676
rect 364812 230042 364840 231676
rect 364800 230036 364852 230042
rect 364800 229978 364852 229984
rect 364432 226976 364484 226982
rect 364432 226918 364484 226924
rect 365180 225554 365208 231676
rect 365548 226710 365576 231676
rect 365916 227390 365944 231676
rect 366284 229770 366312 231676
rect 366272 229764 366324 229770
rect 366272 229706 366324 229712
rect 365904 227384 365956 227390
rect 365904 227326 365956 227332
rect 365536 226704 365588 226710
rect 365536 226646 365588 226652
rect 365168 225548 365220 225554
rect 365168 225490 365220 225496
rect 363696 225480 363748 225486
rect 363696 225422 363748 225428
rect 366560 225350 366588 231676
rect 366928 229838 366956 231676
rect 366916 229832 366968 229838
rect 366916 229774 366968 229780
rect 366548 225344 366600 225350
rect 366548 225286 366600 225292
rect 365720 225276 365772 225282
rect 365720 225218 365772 225224
rect 363236 223576 363288 223582
rect 363236 223518 363288 223524
rect 363248 217410 363276 223518
rect 364984 223168 365036 223174
rect 364984 223110 365036 223116
rect 364340 223032 364392 223038
rect 364340 222974 364392 222980
rect 364352 217410 364380 222974
rect 364996 217410 365024 223110
rect 365732 221134 365760 225218
rect 365812 223372 365864 223378
rect 365812 223314 365864 223320
rect 365720 221128 365772 221134
rect 365720 221070 365772 221076
rect 365824 217410 365852 223314
rect 366640 221536 366692 221542
rect 366640 221478 366692 221484
rect 366652 217410 366680 221478
rect 367296 221202 367324 231676
rect 367468 222896 367520 222902
rect 367468 222838 367520 222844
rect 367284 221196 367336 221202
rect 367284 221138 367336 221144
rect 367480 217410 367508 222838
rect 367664 220182 367692 231676
rect 368032 225282 368060 231676
rect 368400 226778 368428 231676
rect 368768 227254 368796 231676
rect 369136 229566 369164 231676
rect 369124 229560 369176 229566
rect 369124 229502 369176 229508
rect 368756 227248 368808 227254
rect 368756 227190 368808 227196
rect 368388 226772 368440 226778
rect 368388 226714 368440 226720
rect 368020 225276 368072 225282
rect 368020 225218 368072 225224
rect 368572 225208 368624 225214
rect 368572 225150 368624 225156
rect 368296 223304 368348 223310
rect 368296 223246 368348 223252
rect 367652 220176 367704 220182
rect 367652 220118 367704 220124
rect 368308 217410 368336 223246
rect 368584 222902 368612 225150
rect 369412 224369 369440 231676
rect 369780 225214 369808 231676
rect 369768 225208 369820 225214
rect 369768 225150 369820 225156
rect 369398 224360 369454 224369
rect 369398 224295 369454 224304
rect 369124 223236 369176 223242
rect 369124 223178 369176 223184
rect 368572 222896 368624 222902
rect 368572 222838 368624 222844
rect 369136 217410 369164 223178
rect 370044 222964 370096 222970
rect 370044 222906 370096 222912
rect 370056 217410 370084 222906
rect 370148 220114 370176 231676
rect 370516 229634 370544 231676
rect 370504 229628 370556 229634
rect 370504 229570 370556 229576
rect 370884 224505 370912 231676
rect 371252 229498 371280 231676
rect 371240 229492 371292 229498
rect 371240 229434 371292 229440
rect 371620 227458 371648 231676
rect 371608 227452 371660 227458
rect 371608 227394 371660 227400
rect 370870 224496 370926 224505
rect 370870 224431 370926 224440
rect 371700 223100 371752 223106
rect 371700 223042 371752 223048
rect 370872 222828 370924 222834
rect 370872 222770 370924 222776
rect 370136 220108 370188 220114
rect 370136 220050 370188 220056
rect 370884 217410 370912 222770
rect 371712 217410 371740 223042
rect 371988 221270 372016 231676
rect 372068 227044 372120 227050
rect 372068 226986 372120 226992
rect 372080 223038 372108 226986
rect 372264 224777 372292 231676
rect 372632 229702 372660 231676
rect 372620 229696 372672 229702
rect 372620 229638 372672 229644
rect 373000 227050 373028 231676
rect 373368 229430 373396 231676
rect 373356 229424 373408 229430
rect 373356 229366 373408 229372
rect 372988 227044 373040 227050
rect 372988 226986 373040 226992
rect 372250 224768 372306 224777
rect 372250 224703 372306 224712
rect 373736 224641 373764 231676
rect 374000 228540 374052 228546
rect 374000 228482 374052 228488
rect 373722 224632 373778 224641
rect 373722 224567 373778 224576
rect 372068 223032 372120 223038
rect 372068 222974 372120 222980
rect 374012 222766 374040 228482
rect 374104 226506 374132 231676
rect 374472 227526 374500 231676
rect 374840 229362 374868 231676
rect 374828 229356 374880 229362
rect 374828 229298 374880 229304
rect 374460 227520 374512 227526
rect 374460 227462 374512 227468
rect 374092 226500 374144 226506
rect 374092 226442 374144 226448
rect 375116 223553 375144 231676
rect 375288 228608 375340 228614
rect 375288 228550 375340 228556
rect 375102 223544 375158 223553
rect 375102 223479 375158 223488
rect 372620 222760 372672 222766
rect 372620 222702 372672 222708
rect 374000 222760 374052 222766
rect 374000 222702 374052 222708
rect 371976 221264 372028 221270
rect 371976 221206 372028 221212
rect 372632 217410 372660 222702
rect 375300 222426 375328 228550
rect 375484 228546 375512 231676
rect 375472 228540 375524 228546
rect 375472 228482 375524 228488
rect 375380 222624 375432 222630
rect 375380 222566 375432 222572
rect 374184 222420 374236 222426
rect 374184 222362 374236 222368
rect 375288 222420 375340 222426
rect 375288 222362 375340 222368
rect 373356 221672 373408 221678
rect 373356 221614 373408 221620
rect 373368 217410 373396 221614
rect 374196 217410 374224 222362
rect 375392 217410 375420 222566
rect 375852 222057 375880 231676
rect 376220 229294 376248 231676
rect 376208 229288 376260 229294
rect 376208 229230 376260 229236
rect 376588 228682 376616 231676
rect 376576 228676 376628 228682
rect 376576 228618 376628 228624
rect 376852 228472 376904 228478
rect 376852 228414 376904 228420
rect 375932 228404 375984 228410
rect 375932 228346 375984 228352
rect 375838 222048 375894 222057
rect 375838 221983 375894 221992
rect 356532 217382 356868 217410
rect 357360 217382 357696 217410
rect 358280 217382 358616 217410
rect 359108 217382 359444 217410
rect 359936 217382 360272 217410
rect 360764 217382 361100 217410
rect 361776 217382 361928 217410
rect 362420 217382 362756 217410
rect 363248 217382 363584 217410
rect 364352 217382 364504 217410
rect 364996 217382 365332 217410
rect 365824 217382 366160 217410
rect 366652 217382 366988 217410
rect 367480 217382 367816 217410
rect 368308 217382 368644 217410
rect 369136 217382 369472 217410
rect 370056 217382 370392 217410
rect 370884 217382 371220 217410
rect 371712 217382 372048 217410
rect 372632 217382 372876 217410
rect 373368 217382 373704 217410
rect 374196 217382 374532 217410
rect 375360 217382 375420 217410
rect 375944 217410 375972 228346
rect 376760 222488 376812 222494
rect 376760 222430 376812 222436
rect 376772 217410 376800 222430
rect 376864 221066 376892 228414
rect 376956 227089 376984 231676
rect 377036 229084 377088 229090
rect 377036 229026 377088 229032
rect 376942 227080 376998 227089
rect 376942 227015 376998 227024
rect 377048 222494 377076 229026
rect 377324 227225 377352 231676
rect 377310 227216 377366 227225
rect 377310 227151 377366 227160
rect 377588 222692 377640 222698
rect 377588 222634 377640 222640
rect 377036 222488 377088 222494
rect 377036 222430 377088 222436
rect 376852 221060 376904 221066
rect 376852 221002 376904 221008
rect 377600 217410 377628 222634
rect 377692 221338 377720 231676
rect 377968 228614 377996 231676
rect 377956 228608 378008 228614
rect 377956 228550 378008 228556
rect 378140 227588 378192 227594
rect 378140 227530 378192 227536
rect 378152 223990 378180 227530
rect 378140 223984 378192 223990
rect 378140 223926 378192 223932
rect 378336 223417 378364 231676
rect 378508 228948 378560 228954
rect 378508 228890 378560 228896
rect 378322 223408 378378 223417
rect 378322 223343 378378 223352
rect 378520 222562 378548 228890
rect 378704 223281 378732 231676
rect 378690 223272 378746 223281
rect 378690 223207 378746 223216
rect 378416 222556 378468 222562
rect 378416 222498 378468 222504
rect 378508 222556 378560 222562
rect 378508 222498 378560 222504
rect 377680 221332 377732 221338
rect 377680 221274 377732 221280
rect 378428 217410 378456 222498
rect 379072 221406 379100 231676
rect 379440 228478 379468 231676
rect 379428 228472 379480 228478
rect 379428 228414 379480 228420
rect 379244 228268 379296 228274
rect 379244 228210 379296 228216
rect 379060 221400 379112 221406
rect 379060 221342 379112 221348
rect 379256 217410 379284 228210
rect 379808 227497 379836 231676
rect 379794 227488 379850 227497
rect 379794 227423 379850 227432
rect 380176 227361 380204 231676
rect 380162 227352 380218 227361
rect 380162 227287 380218 227296
rect 380072 221740 380124 221746
rect 380072 221682 380124 221688
rect 380084 217410 380112 221682
rect 380544 221542 380572 231676
rect 380532 221536 380584 221542
rect 380532 221478 380584 221484
rect 380820 221474 380848 231676
rect 380900 229016 380952 229022
rect 380900 228958 380952 228964
rect 380912 223922 380940 228958
rect 380900 223916 380952 223922
rect 380900 223858 380952 223864
rect 381188 223145 381216 231676
rect 381174 223136 381230 223145
rect 381174 223071 381230 223080
rect 381556 222873 381584 231676
rect 381542 222864 381598 222873
rect 381542 222799 381598 222808
rect 381082 222728 381138 222737
rect 381082 222663 381138 222672
rect 380808 221468 380860 221474
rect 380808 221410 380860 221416
rect 381096 217410 381124 222663
rect 381820 222352 381872 222358
rect 381820 222294 381872 222300
rect 381832 217410 381860 222294
rect 381924 222154 381952 231676
rect 382292 228410 382320 231676
rect 382660 228857 382688 231676
rect 382646 228848 382702 228857
rect 382646 228783 382702 228792
rect 382280 228404 382332 228410
rect 382280 228346 382332 228352
rect 382004 228336 382056 228342
rect 382004 228278 382056 228284
rect 381912 222148 381964 222154
rect 381912 222090 381964 222096
rect 382016 221610 382044 228278
rect 383028 227594 383056 231676
rect 383016 227588 383068 227594
rect 383016 227530 383068 227536
rect 383396 221746 383424 231676
rect 383672 223009 383700 231676
rect 383752 228880 383804 228886
rect 383752 228822 383804 228828
rect 383764 224058 383792 228822
rect 383752 224052 383804 224058
rect 383752 223994 383804 224000
rect 383658 223000 383714 223009
rect 383658 222935 383714 222944
rect 383658 222456 383714 222465
rect 383658 222391 383714 222400
rect 383384 221740 383436 221746
rect 383384 221682 383436 221688
rect 382004 221604 382056 221610
rect 382004 221546 382056 221552
rect 382648 221060 382700 221066
rect 382648 221002 382700 221008
rect 382660 217410 382688 221002
rect 383672 217410 383700 222391
rect 384040 221678 384068 231676
rect 384408 228342 384436 231676
rect 384776 228993 384804 231676
rect 384762 228984 384818 228993
rect 384762 228919 384818 228928
rect 384396 228336 384448 228342
rect 384396 228278 384448 228284
rect 385144 227662 385172 231676
rect 385132 227656 385184 227662
rect 385132 227598 385184 227604
rect 384302 222592 384358 222601
rect 384302 222527 384358 222536
rect 384028 221672 384080 221678
rect 384028 221614 384080 221620
rect 384316 217410 384344 222527
rect 385132 222284 385184 222290
rect 385132 222226 385184 222232
rect 385144 217410 385172 222226
rect 385512 221814 385540 231676
rect 385880 222737 385908 231676
rect 385960 228132 386012 228138
rect 385960 228074 386012 228080
rect 385866 222728 385922 222737
rect 385866 222663 385922 222672
rect 385500 221808 385552 221814
rect 385500 221750 385552 221756
rect 385972 217410 386000 228074
rect 386248 221882 386276 231676
rect 386524 228274 386552 231676
rect 386892 228721 386920 231676
rect 387260 228886 387288 231676
rect 387248 228880 387300 228886
rect 387248 228822 387300 228828
rect 386878 228712 386934 228721
rect 386878 228647 386934 228656
rect 386512 228268 386564 228274
rect 386512 228210 386564 228216
rect 387628 221950 387656 231676
rect 387996 222601 388024 231676
rect 388364 229022 388392 231676
rect 388352 229016 388404 229022
rect 388352 228958 388404 228964
rect 387982 222592 388038 222601
rect 387982 222527 388038 222536
rect 387706 222320 387762 222329
rect 387706 222255 387762 222264
rect 387616 221944 387668 221950
rect 387616 221886 387668 221892
rect 386236 221876 386288 221882
rect 386236 221818 386288 221824
rect 386786 221640 386842 221649
rect 386786 221575 386842 221584
rect 386800 217410 386828 221575
rect 387720 217410 387748 222255
rect 388732 222018 388760 231676
rect 389008 231662 389114 231690
rect 389008 222465 389036 231662
rect 389088 228744 389140 228750
rect 389088 228686 389140 228692
rect 388994 222456 389050 222465
rect 388994 222391 389050 222400
rect 388720 222012 388772 222018
rect 388720 221954 388772 221960
rect 388534 221776 388590 221785
rect 388534 221711 388590 221720
rect 388548 217410 388576 221711
rect 389100 221066 389128 228686
rect 389376 226137 389404 231676
rect 389744 228954 389772 231676
rect 389732 228948 389784 228954
rect 389732 228890 389784 228896
rect 390112 228585 390140 231676
rect 390098 228576 390154 228585
rect 390098 228511 390154 228520
rect 389362 226128 389418 226137
rect 389362 226063 389418 226072
rect 390480 226001 390508 231676
rect 390466 225992 390522 226001
rect 390466 225927 390522 225936
rect 390848 222358 390876 231676
rect 391020 222760 391072 222766
rect 391020 222702 391072 222708
rect 390836 222352 390888 222358
rect 390836 222294 390888 222300
rect 390190 222184 390246 222193
rect 390190 222119 390246 222128
rect 389364 221604 389416 221610
rect 389364 221546 389416 221552
rect 389088 221060 389140 221066
rect 389088 221002 389140 221008
rect 389376 217410 389404 221546
rect 390204 217410 390232 222119
rect 391032 217410 391060 222702
rect 391216 222329 391244 231676
rect 391584 225865 391612 231676
rect 391966 231662 392164 231690
rect 392136 229022 392164 231662
rect 392124 229016 392176 229022
rect 392124 228958 392176 228964
rect 391756 228812 391808 228818
rect 391756 228754 391808 228760
rect 391570 225856 391626 225865
rect 391570 225791 391626 225800
rect 391768 222698 391796 228754
rect 392228 228449 392256 231676
rect 392214 228440 392270 228449
rect 392214 228375 392270 228384
rect 391848 228200 391900 228206
rect 391848 228142 391900 228148
rect 391756 222692 391808 222698
rect 391756 222634 391808 222640
rect 391202 222320 391258 222329
rect 391860 222290 391888 228142
rect 391940 228064 391992 228070
rect 391940 228006 391992 228012
rect 391202 222255 391258 222264
rect 391848 222284 391900 222290
rect 391848 222226 391900 222232
rect 391952 217410 391980 228006
rect 392596 225729 392624 231676
rect 392978 231662 393268 231690
rect 392952 227928 393004 227934
rect 392952 227870 393004 227876
rect 392582 225720 392638 225729
rect 392582 225655 392638 225664
rect 392964 223582 392992 227870
rect 392952 223576 393004 223582
rect 392952 223518 393004 223524
rect 392676 222556 392728 222562
rect 392676 222498 392728 222504
rect 392688 217410 392716 222498
rect 393240 222086 393268 231662
rect 393332 222193 393360 231676
rect 393700 229226 393728 231676
rect 393688 229220 393740 229226
rect 393688 229162 393740 229168
rect 394068 228818 394096 231676
rect 394056 228812 394108 228818
rect 394056 228754 394108 228760
rect 394436 228313 394464 231676
rect 394422 228304 394478 228313
rect 394422 228239 394478 228248
rect 394804 225593 394832 231676
rect 394790 225584 394846 225593
rect 394790 225519 394846 225528
rect 394700 222420 394752 222426
rect 394700 222362 394752 222368
rect 393596 222216 393648 222222
rect 393318 222184 393374 222193
rect 393596 222158 393648 222164
rect 393318 222119 393374 222128
rect 393228 222080 393280 222086
rect 393228 222022 393280 222028
rect 393608 217410 393636 222158
rect 394712 217410 394740 222362
rect 395080 220862 395108 231676
rect 395252 223576 395304 223582
rect 395252 223518 395304 223524
rect 395068 220856 395120 220862
rect 395068 220798 395120 220804
rect 395264 217410 395292 223518
rect 395448 220930 395476 231676
rect 395816 226642 395844 231676
rect 396184 228750 396212 231676
rect 396172 228744 396224 228750
rect 396172 228686 396224 228692
rect 396552 228177 396580 231676
rect 396920 229158 396948 231676
rect 396908 229152 396960 229158
rect 396908 229094 396960 229100
rect 396538 228168 396594 228177
rect 396538 228103 396594 228112
rect 396540 227996 396592 228002
rect 396540 227938 396592 227944
rect 395804 226636 395856 226642
rect 395804 226578 395856 226584
rect 396552 222970 396580 227938
rect 397288 223446 397316 231676
rect 397368 229084 397420 229090
rect 397368 229026 397420 229032
rect 397380 226273 397408 229026
rect 397366 226264 397422 226273
rect 397366 226199 397422 226208
rect 397276 223440 397328 223446
rect 397276 223382 397328 223388
rect 396540 222964 396592 222970
rect 396540 222906 396592 222912
rect 396906 221912 396962 221921
rect 396906 221847 396962 221856
rect 396080 221060 396132 221066
rect 396080 221002 396132 221008
rect 395436 220924 395488 220930
rect 395436 220866 395488 220872
rect 396092 217410 396120 221002
rect 396920 217410 396948 221847
rect 397656 221066 397684 231676
rect 397932 225457 397960 231676
rect 397918 225448 397974 225457
rect 397918 225383 397974 225392
rect 398300 223378 398328 231676
rect 398668 228041 398696 231676
rect 398654 228032 398710 228041
rect 398654 227967 398710 227976
rect 398288 223372 398340 223378
rect 398288 223314 398340 223320
rect 399036 223310 399064 231676
rect 399024 223304 399076 223310
rect 399024 223246 399076 223252
rect 399404 223174 399432 231676
rect 399772 227905 399800 231676
rect 399758 227896 399814 227905
rect 399758 227831 399814 227840
rect 400140 223242 400168 231676
rect 400508 228206 400536 231676
rect 400496 228200 400548 228206
rect 400496 228142 400548 228148
rect 400404 224120 400456 224126
rect 400404 224062 400456 224068
rect 400128 223236 400180 223242
rect 400128 223178 400180 223184
rect 399392 223168 399444 223174
rect 399392 223110 399444 223116
rect 397736 223032 397788 223038
rect 397736 222974 397788 222980
rect 397644 221060 397696 221066
rect 397644 221002 397696 221008
rect 397748 217410 397776 222974
rect 398564 222896 398616 222902
rect 398564 222838 398616 222844
rect 398576 217410 398604 222838
rect 399484 222488 399536 222494
rect 399484 222430 399536 222436
rect 399496 217410 399524 222430
rect 400416 217410 400444 224062
rect 400784 223106 400812 231676
rect 401152 225321 401180 231676
rect 401534 231662 401824 231690
rect 401508 229084 401560 229090
rect 401508 229026 401560 229032
rect 401520 228886 401548 229026
rect 401508 228880 401560 228886
rect 401508 228822 401560 228828
rect 401138 225312 401194 225321
rect 401138 225247 401194 225256
rect 401508 224664 401560 224670
rect 401508 224606 401560 224612
rect 401520 223990 401548 224606
rect 401508 223984 401560 223990
rect 401508 223926 401560 223932
rect 400772 223100 400824 223106
rect 400772 223042 400824 223048
rect 401796 223038 401824 231662
rect 401784 223032 401836 223038
rect 401784 222974 401836 222980
rect 401888 222834 401916 231676
rect 401968 222964 402020 222970
rect 401968 222906 402020 222912
rect 401876 222828 401928 222834
rect 401876 222770 401928 222776
rect 401140 222284 401192 222290
rect 401140 222226 401192 222232
rect 401152 217410 401180 222226
rect 401416 222148 401468 222154
rect 401416 222090 401468 222096
rect 401428 221610 401456 222090
rect 401416 221604 401468 221610
rect 401416 221546 401468 221552
rect 401980 217410 402008 222906
rect 402256 222902 402284 231676
rect 402624 226574 402652 231676
rect 402992 228070 403020 231676
rect 403360 228818 403388 231676
rect 403348 228812 403400 228818
rect 403348 228754 403400 228760
rect 403636 228138 403664 231676
rect 403624 228132 403676 228138
rect 403624 228074 403676 228080
rect 402980 228064 403032 228070
rect 402980 228006 403032 228012
rect 403624 227860 403676 227866
rect 403624 227802 403676 227808
rect 402980 227792 403032 227798
rect 402980 227734 403032 227740
rect 402612 226568 402664 226574
rect 402612 226510 402664 226516
rect 402992 223582 403020 227734
rect 402980 223576 403032 223582
rect 402980 223518 403032 223524
rect 402244 222896 402296 222902
rect 402244 222838 402296 222844
rect 402980 222692 403032 222698
rect 402980 222634 403032 222640
rect 402992 217410 403020 222634
rect 403636 217410 403664 227802
rect 404004 227769 404032 231676
rect 403990 227760 404046 227769
rect 403990 227695 404046 227704
rect 404372 226438 404400 231676
rect 404544 226840 404596 226846
rect 404544 226782 404596 226788
rect 404360 226432 404412 226438
rect 404360 226374 404412 226380
rect 404556 224058 404584 226782
rect 404452 224052 404504 224058
rect 404452 223994 404504 224000
rect 404544 224052 404596 224058
rect 404544 223994 404596 224000
rect 404464 217410 404492 223994
rect 404740 222766 404768 231676
rect 404728 222760 404780 222766
rect 404728 222702 404780 222708
rect 405108 222630 405136 231676
rect 405476 225185 405504 231676
rect 405858 231662 406148 231690
rect 406226 231662 406424 231690
rect 405832 226704 405884 226710
rect 405832 226646 405884 226652
rect 405740 226500 405792 226506
rect 405740 226442 405792 226448
rect 405462 225176 405518 225185
rect 405462 225111 405518 225120
rect 405752 224602 405780 226442
rect 405648 224596 405700 224602
rect 405648 224538 405700 224544
rect 405740 224596 405792 224602
rect 405740 224538 405792 224544
rect 405660 224482 405688 224538
rect 405660 224454 405780 224482
rect 405096 222624 405148 222630
rect 405096 222566 405148 222572
rect 405752 217410 405780 224454
rect 405844 224126 405872 226646
rect 405832 224120 405884 224126
rect 405832 224062 405884 224068
rect 406120 222698 406148 231662
rect 406200 223576 406252 223582
rect 406200 223518 406252 223524
rect 406108 222692 406160 222698
rect 406108 222634 406160 222640
rect 375944 217382 376280 217410
rect 376772 217382 377108 217410
rect 377600 217382 377936 217410
rect 378428 217382 378764 217410
rect 379256 217382 379592 217410
rect 380084 217382 380420 217410
rect 381096 217382 381248 217410
rect 381832 217382 382168 217410
rect 382660 217382 382996 217410
rect 383672 217382 383824 217410
rect 384316 217382 384652 217410
rect 385144 217382 385480 217410
rect 385972 217382 386308 217410
rect 386800 217382 387136 217410
rect 387720 217382 388056 217410
rect 388548 217382 388884 217410
rect 389376 217382 389712 217410
rect 390204 217382 390540 217410
rect 391032 217382 391368 217410
rect 391952 217382 392196 217410
rect 392688 217382 393024 217410
rect 393608 217382 393944 217410
rect 394712 217382 394772 217410
rect 395264 217382 395600 217410
rect 396092 217382 396428 217410
rect 396920 217382 397256 217410
rect 397748 217382 398084 217410
rect 398576 217382 398912 217410
rect 399496 217382 399832 217410
rect 400416 217382 400660 217410
rect 401152 217382 401488 217410
rect 401980 217382 402316 217410
rect 402992 217382 403144 217410
rect 403636 217382 403972 217410
rect 404464 217382 404800 217410
rect 405720 217382 405780 217410
rect 406212 217410 406240 223518
rect 406396 222562 406424 231662
rect 406488 225049 406516 231676
rect 406856 228002 406884 231676
rect 406844 227996 406896 228002
rect 406844 227938 406896 227944
rect 407224 227798 407252 231676
rect 407212 227792 407264 227798
rect 407212 227734 407264 227740
rect 406474 225040 406530 225049
rect 406474 224975 406530 224984
rect 406568 223440 406620 223446
rect 406568 223382 406620 223388
rect 406580 223242 406608 223382
rect 406476 223236 406528 223242
rect 406476 223178 406528 223184
rect 406568 223236 406620 223242
rect 406568 223178 406620 223184
rect 406488 223038 406516 223178
rect 406476 223032 406528 223038
rect 406476 222974 406528 222980
rect 406384 222556 406436 222562
rect 406384 222498 406436 222504
rect 407592 222426 407620 231676
rect 407856 223848 407908 223854
rect 407856 223790 407908 223796
rect 407580 222420 407632 222426
rect 407580 222362 407632 222368
rect 407028 221128 407080 221134
rect 407028 221070 407080 221076
rect 407040 217410 407068 221070
rect 407868 217410 407896 223790
rect 407960 222494 407988 231676
rect 407948 222488 408000 222494
rect 407948 222430 408000 222436
rect 408328 222358 408356 231676
rect 408500 227316 408552 227322
rect 408500 227258 408552 227264
rect 408512 223650 408540 227258
rect 408696 226710 408724 231676
rect 409064 227934 409092 231676
rect 409052 227928 409104 227934
rect 409052 227870 409104 227876
rect 409340 227866 409368 231676
rect 409328 227860 409380 227866
rect 409328 227802 409380 227808
rect 409708 226846 409736 231676
rect 409696 226840 409748 226846
rect 409696 226782 409748 226788
rect 408776 226772 408828 226778
rect 408776 226714 408828 226720
rect 408684 226704 408736 226710
rect 408684 226646 408736 226652
rect 408788 224194 408816 226714
rect 408684 224188 408736 224194
rect 408684 224130 408736 224136
rect 408776 224188 408828 224194
rect 408776 224130 408828 224136
rect 408500 223644 408552 223650
rect 408500 223586 408552 223592
rect 408316 222352 408368 222358
rect 408316 222294 408368 222300
rect 408696 217410 408724 224130
rect 410076 222290 410104 231676
rect 410340 227724 410392 227730
rect 410340 227666 410392 227672
rect 410064 222284 410116 222290
rect 410064 222226 410116 222232
rect 409512 219292 409564 219298
rect 409512 219234 409564 219240
rect 409524 217410 409552 219234
rect 410352 217410 410380 227666
rect 410444 222222 410472 231676
rect 410812 224913 410840 231676
rect 411180 227633 411208 231676
rect 411548 227730 411576 231676
rect 414020 231192 414072 231198
rect 414020 231134 414072 231140
rect 411536 227724 411588 227730
rect 411536 227666 411588 227672
rect 411166 227624 411222 227633
rect 411166 227559 411222 227568
rect 413192 227180 413244 227186
rect 413192 227122 413244 227128
rect 410798 224904 410854 224913
rect 410798 224839 410854 224848
rect 413204 224262 413232 227122
rect 412088 224256 412140 224262
rect 412088 224198 412140 224204
rect 413192 224256 413244 224262
rect 413192 224198 413244 224204
rect 411260 223848 411312 223854
rect 411260 223790 411312 223796
rect 410432 222216 410484 222222
rect 410432 222158 410484 222164
rect 411272 217410 411300 223790
rect 412100 217410 412128 224198
rect 412916 220788 412968 220794
rect 412916 220730 412968 220736
rect 412928 217410 412956 220730
rect 414032 217410 414060 231134
rect 417148 231056 417200 231062
rect 417148 230998 417200 231004
rect 416780 228812 416832 228818
rect 416780 228754 416832 228760
rect 416872 228812 416924 228818
rect 416872 228754 416924 228760
rect 415308 227112 415360 227118
rect 415308 227054 415360 227060
rect 415320 224330 415348 227054
rect 416792 224942 416820 228754
rect 416884 228206 416912 228754
rect 416872 228200 416924 228206
rect 416872 228142 416924 228148
rect 416964 228200 417016 228206
rect 416964 228142 417016 228148
rect 416976 228070 417004 228142
rect 416964 228064 417016 228070
rect 416964 228006 417016 228012
rect 417056 228064 417108 228070
rect 417056 228006 417108 228012
rect 416872 226908 416924 226914
rect 416872 226850 416924 226856
rect 416688 224936 416740 224942
rect 416688 224878 416740 224884
rect 416780 224936 416832 224942
rect 416780 224878 416832 224884
rect 416700 224670 416728 224878
rect 416688 224664 416740 224670
rect 416688 224606 416740 224612
rect 416884 224466 416912 226850
rect 417068 226574 417096 228006
rect 417056 226568 417108 226574
rect 417056 226510 417108 226516
rect 415400 224460 415452 224466
rect 415400 224402 415452 224408
rect 416872 224460 416924 224466
rect 416872 224402 416924 224408
rect 414572 224324 414624 224330
rect 414572 224266 414624 224272
rect 415308 224324 415360 224330
rect 415308 224266 415360 224272
rect 414584 217410 414612 224266
rect 415412 217410 415440 224402
rect 416228 219360 416280 219366
rect 416228 219302 416280 219308
rect 416240 217410 416268 219302
rect 417160 217410 417188 230998
rect 418080 226334 418108 243063
rect 418158 240000 418214 240009
rect 418158 239935 418214 239944
rect 417896 226306 418108 226334
rect 406212 217382 406548 217410
rect 407040 217382 407376 217410
rect 407868 217382 408204 217410
rect 408696 217382 409032 217410
rect 409524 217382 409860 217410
rect 410352 217382 410688 217410
rect 411272 217382 411608 217410
rect 412100 217382 412436 217410
rect 412928 217382 413264 217410
rect 414032 217382 414092 217410
rect 414584 217382 414920 217410
rect 415412 217382 415748 217410
rect 416240 217382 416576 217410
rect 417160 217382 417496 217410
rect 63406 217288 63462 217297
rect 63406 217223 63462 217232
rect 417896 216850 417924 226306
rect 417976 224664 418028 224670
rect 417976 224606 418028 224612
rect 417988 217410 418016 224606
rect 418172 217870 418200 239935
rect 418434 236736 418490 236745
rect 418434 236671 418490 236680
rect 418160 217864 418212 217870
rect 418160 217806 418212 217812
rect 417988 217382 418324 217410
rect 418448 216986 418476 236671
rect 418526 233608 418582 233617
rect 418526 233543 418582 233552
rect 418540 217054 418568 233543
rect 437296 231124 437348 231130
rect 437296 231066 437348 231072
rect 420460 230920 420512 230926
rect 420460 230862 420512 230868
rect 418804 224392 418856 224398
rect 418804 224334 418856 224340
rect 418620 217864 418672 217870
rect 418620 217806 418672 217812
rect 418528 217048 418580 217054
rect 418528 216990 418580 216996
rect 418436 216980 418488 216986
rect 418436 216922 418488 216928
rect 418632 216918 418660 217806
rect 418816 217410 418844 224334
rect 419724 220652 419776 220658
rect 419724 220594 419776 220600
rect 419736 217410 419764 220594
rect 420472 217410 420500 230862
rect 427176 230852 427228 230858
rect 427176 230794 427228 230800
rect 425428 227384 425480 227390
rect 425428 227326 425480 227332
rect 422300 226976 422352 226982
rect 422300 226918 422352 226924
rect 422312 224670 422340 226918
rect 425060 226296 425112 226302
rect 425060 226238 425112 226244
rect 422300 224664 422352 224670
rect 422300 224606 422352 224612
rect 421288 224528 421340 224534
rect 421288 224470 421340 224476
rect 421300 217410 421328 224470
rect 422300 223984 422352 223990
rect 422300 223926 422352 223932
rect 422312 217410 422340 223926
rect 423864 223644 423916 223650
rect 423864 223586 423916 223592
rect 423036 220720 423088 220726
rect 423036 220662 423088 220668
rect 423048 217410 423076 220662
rect 423876 217410 423904 223586
rect 425072 217410 425100 226238
rect 425244 224800 425296 224806
rect 425244 224742 425296 224748
rect 425256 224534 425284 224742
rect 425440 224738 425468 227326
rect 425520 224800 425572 224806
rect 425520 224742 425572 224748
rect 425428 224732 425480 224738
rect 425428 224674 425480 224680
rect 425244 224528 425296 224534
rect 425244 224470 425296 224476
rect 418816 217382 419152 217410
rect 419736 217382 419980 217410
rect 420472 217382 420808 217410
rect 421300 217382 421636 217410
rect 422312 217382 422464 217410
rect 423048 217382 423384 217410
rect 423876 217382 424212 217410
rect 425040 217382 425100 217410
rect 425532 217410 425560 224742
rect 426348 220584 426400 220590
rect 426348 220526 426400 220532
rect 426360 217410 426388 220526
rect 427188 217410 427216 230794
rect 433892 230784 433944 230790
rect 433892 230726 433944 230732
rect 433156 227452 433208 227458
rect 433156 227394 433208 227400
rect 430396 227248 430448 227254
rect 430396 227190 430448 227196
rect 430408 226302 430436 227190
rect 430396 226296 430448 226302
rect 430396 226238 430448 226244
rect 433168 226234 433196 227394
rect 433248 227044 433300 227050
rect 433248 226986 433300 226992
rect 428924 226228 428976 226234
rect 428924 226170 428976 226176
rect 433156 226228 433208 226234
rect 433156 226170 433208 226176
rect 428004 224868 428056 224874
rect 428004 224810 428056 224816
rect 428016 217410 428044 224810
rect 428936 217410 428964 226170
rect 433260 226098 433288 226986
rect 431408 226092 431460 226098
rect 431408 226034 431460 226040
rect 433248 226092 433300 226098
rect 433248 226034 433300 226040
rect 429108 225888 429160 225894
rect 429108 225830 429160 225836
rect 429120 224806 429148 225830
rect 429108 224800 429160 224806
rect 429108 224742 429160 224748
rect 430580 224256 430632 224262
rect 430580 224198 430632 224204
rect 429752 220516 429804 220522
rect 429752 220458 429804 220464
rect 429764 217410 429792 220458
rect 430592 217410 430620 224198
rect 431420 217410 431448 226034
rect 432236 224528 432288 224534
rect 432236 224470 432288 224476
rect 432248 217410 432276 224470
rect 433340 220448 433392 220454
rect 433340 220390 433392 220396
rect 433352 217410 433380 220390
rect 433904 217410 433932 230726
rect 435732 227520 435784 227526
rect 435732 227462 435784 227468
rect 434812 226160 434864 226166
rect 434812 226102 434864 226108
rect 434628 225004 434680 225010
rect 434628 224946 434680 224952
rect 434640 224874 434668 224946
rect 434628 224868 434680 224874
rect 434628 224810 434680 224816
rect 434824 217410 434852 226102
rect 435744 225962 435772 227462
rect 435640 225956 435692 225962
rect 435640 225898 435692 225904
rect 435732 225956 435784 225962
rect 435732 225898 435784 225904
rect 435652 217410 435680 225898
rect 436468 220312 436520 220318
rect 436468 220254 436520 220260
rect 436480 217410 436508 220254
rect 437308 217410 437336 231066
rect 439780 230988 439832 230994
rect 439780 230930 439832 230936
rect 438768 226636 438820 226642
rect 438768 226578 438820 226584
rect 438780 225418 438808 226578
rect 439044 226024 439096 226030
rect 439044 225966 439096 225972
rect 438124 225412 438176 225418
rect 438124 225354 438176 225360
rect 438768 225412 438820 225418
rect 438768 225354 438820 225360
rect 438136 217410 438164 225354
rect 439056 217410 439084 225966
rect 439792 217410 439820 230930
rect 446588 230376 446640 230382
rect 446588 230318 446640 230324
rect 443184 230308 443236 230314
rect 443184 230250 443236 230256
rect 441620 226568 441672 226574
rect 441620 226510 441672 226516
rect 440332 225616 440384 225622
rect 440516 225616 440568 225622
rect 440384 225564 440516 225570
rect 440332 225558 440568 225564
rect 440344 225542 440556 225558
rect 441632 225146 441660 226510
rect 441620 225140 441672 225146
rect 441620 225082 441672 225088
rect 442356 225072 442408 225078
rect 442356 225014 442408 225020
rect 441620 224800 441672 224806
rect 441620 224742 441672 224748
rect 440700 220380 440752 220386
rect 440700 220322 440752 220328
rect 440712 217410 440740 220322
rect 441632 217410 441660 224742
rect 442368 217410 442396 225014
rect 443196 217410 443224 230250
rect 444380 226704 444432 226710
rect 444380 226646 444432 226652
rect 444392 225078 444420 226646
rect 444380 225072 444432 225078
rect 444380 225014 444432 225020
rect 444840 225004 444892 225010
rect 444840 224946 444892 224952
rect 444380 224324 444432 224330
rect 444380 224266 444432 224272
rect 444392 217410 444420 224266
rect 425532 217382 425868 217410
rect 426360 217382 426696 217410
rect 427188 217382 427524 217410
rect 428016 217382 428352 217410
rect 428936 217382 429272 217410
rect 429764 217382 430100 217410
rect 430592 217382 430928 217410
rect 431420 217382 431756 217410
rect 432248 217382 432584 217410
rect 433352 217382 433412 217410
rect 433904 217382 434240 217410
rect 434824 217382 435160 217410
rect 435652 217382 435988 217410
rect 436480 217382 436816 217410
rect 437308 217382 437644 217410
rect 438136 217382 438472 217410
rect 439056 217382 439300 217410
rect 439792 217382 440128 217410
rect 440712 217382 441048 217410
rect 441632 217382 441876 217410
rect 442368 217382 442704 217410
rect 443196 217382 443532 217410
rect 444360 217382 444420 217410
rect 444852 217410 444880 224946
rect 445668 224052 445720 224058
rect 445668 223994 445720 224000
rect 445680 217410 445708 223994
rect 446600 217410 446628 230318
rect 454132 230240 454184 230246
rect 454132 230182 454184 230188
rect 453304 230172 453356 230178
rect 453304 230114 453356 230120
rect 449900 230104 449952 230110
rect 449900 230046 449952 230052
rect 447140 226840 447192 226846
rect 447140 226782 447192 226788
rect 447152 225010 447180 226782
rect 448244 225888 448296 225894
rect 448244 225830 448296 225836
rect 447140 225004 447192 225010
rect 447140 224946 447192 224952
rect 447416 220244 447468 220250
rect 447416 220186 447468 220192
rect 447428 217410 447456 220186
rect 448256 217410 448284 225830
rect 449072 224868 449124 224874
rect 449072 224810 449124 224816
rect 449084 217410 449112 224810
rect 449912 217410 449940 230046
rect 452568 227588 452620 227594
rect 452568 227530 452620 227536
rect 452580 225826 452608 227530
rect 452568 225820 452620 225826
rect 452568 225762 452620 225768
rect 451556 225752 451608 225758
rect 451556 225694 451608 225700
rect 450728 224460 450780 224466
rect 450728 224402 450780 224408
rect 450740 217410 450768 224402
rect 451568 217410 451596 225694
rect 452660 225616 452712 225622
rect 452660 225558 452712 225564
rect 452672 217410 452700 225558
rect 453316 217410 453344 230114
rect 453856 227656 453908 227662
rect 453856 227598 453908 227604
rect 453868 225622 453896 227598
rect 453856 225616 453908 225622
rect 453856 225558 453908 225564
rect 454144 217410 454172 230182
rect 460020 230036 460072 230042
rect 460020 229978 460072 229984
rect 456616 229968 456668 229974
rect 456616 229910 456668 229916
rect 455788 229900 455840 229906
rect 455788 229842 455840 229848
rect 454960 225752 455012 225758
rect 454960 225694 455012 225700
rect 454972 217410 455000 225694
rect 455800 217410 455828 229842
rect 456628 217410 456656 229910
rect 458180 229084 458232 229090
rect 458180 229026 458232 229032
rect 458192 225486 458220 229026
rect 458456 225548 458508 225554
rect 458456 225490 458508 225496
rect 458180 225480 458232 225486
rect 458180 225422 458232 225428
rect 457444 224664 457496 224670
rect 457444 224606 457496 224612
rect 457456 217410 457484 224606
rect 458468 217410 458496 225490
rect 459192 224120 459244 224126
rect 459192 224062 459244 224068
rect 459204 217410 459232 224062
rect 460032 217410 460060 229978
rect 462504 229832 462556 229838
rect 462504 229774 462556 229780
rect 460940 228676 460992 228682
rect 460940 228618 460992 228624
rect 460952 225758 460980 228618
rect 460940 225752 460992 225758
rect 460940 225694 460992 225700
rect 461676 225684 461728 225690
rect 461676 225626 461728 225632
rect 460940 224732 460992 224738
rect 460940 224674 460992 224680
rect 460952 217410 460980 224674
rect 461688 217410 461716 225626
rect 462516 217410 462544 229774
rect 463700 229764 463752 229770
rect 463700 229706 463752 229712
rect 463712 217410 463740 229706
rect 476028 229696 476080 229702
rect 476028 229638 476080 229644
rect 473452 229628 473504 229634
rect 473452 229570 473504 229576
rect 470140 229560 470192 229566
rect 470140 229502 470192 229508
rect 467012 229016 467064 229022
rect 467012 228958 467064 228964
rect 464436 228948 464488 228954
rect 464436 228890 464488 228896
rect 464448 225554 464476 228890
rect 467024 225690 467052 228958
rect 469956 228880 470008 228886
rect 469956 228822 470008 228828
rect 467564 226296 467616 226302
rect 467564 226238 467616 226244
rect 467012 225684 467064 225690
rect 467012 225626 467064 225632
rect 464436 225548 464488 225554
rect 464436 225490 464488 225496
rect 465080 225344 465132 225350
rect 465080 225286 465132 225292
rect 464252 221196 464304 221202
rect 464252 221138 464304 221144
rect 444852 217382 445188 217410
rect 445680 217382 446016 217410
rect 446600 217382 446936 217410
rect 447428 217382 447764 217410
rect 448256 217382 448592 217410
rect 449084 217382 449420 217410
rect 449912 217382 450248 217410
rect 450740 217382 451076 217410
rect 451568 217382 451904 217410
rect 452672 217382 452824 217410
rect 453316 217382 453652 217410
rect 454144 217382 454480 217410
rect 454972 217382 455308 217410
rect 455800 217382 456136 217410
rect 456628 217382 456964 217410
rect 457456 217382 457792 217410
rect 458468 217382 458712 217410
rect 459204 217382 459540 217410
rect 460032 217382 460368 217410
rect 460952 217382 461196 217410
rect 461688 217382 462024 217410
rect 462516 217382 462852 217410
rect 463680 217382 463740 217410
rect 464264 217410 464292 221138
rect 465092 217410 465120 225286
rect 465908 224188 465960 224194
rect 465908 224130 465960 224136
rect 465920 217410 465948 224130
rect 466736 220176 466788 220182
rect 466736 220118 466788 220124
rect 466748 217410 466776 220118
rect 467576 217410 467604 226238
rect 469968 225350 469996 228822
rect 469956 225344 470008 225350
rect 469956 225286 470008 225292
rect 468392 225276 468444 225282
rect 468392 225218 468444 225224
rect 468404 217410 468432 225218
rect 469220 225208 469272 225214
rect 469220 225150 469272 225156
rect 469232 217410 469260 225150
rect 470152 217410 470180 229502
rect 472624 229492 472676 229498
rect 472624 229434 472676 229440
rect 471978 224360 472034 224369
rect 471978 224295 472034 224304
rect 470968 220108 471020 220114
rect 470968 220050 471020 220056
rect 470980 217410 471008 220050
rect 471992 217410 472020 224295
rect 472636 217410 472664 229434
rect 473268 228744 473320 228750
rect 473268 228686 473320 228692
rect 473280 225282 473308 228686
rect 473268 225276 473320 225282
rect 473268 225218 473320 225224
rect 473464 217410 473492 229570
rect 474740 228608 474792 228614
rect 474740 228550 474792 228556
rect 474280 226228 474332 226234
rect 474280 226170 474332 226176
rect 474292 217410 474320 226170
rect 474752 225894 474780 228550
rect 474740 225888 474792 225894
rect 474740 225830 474792 225836
rect 475106 224496 475162 224505
rect 475106 224431 475162 224440
rect 475120 217410 475148 224431
rect 476040 217410 476068 229638
rect 480352 229424 480404 229430
rect 480352 229366 480404 229372
rect 477500 228812 477552 228818
rect 477500 228754 477552 228760
rect 477512 225214 477540 228754
rect 480260 228540 480312 228546
rect 480260 228482 480312 228488
rect 477776 226092 477828 226098
rect 477776 226034 477828 226040
rect 477500 225208 477552 225214
rect 477500 225150 477552 225156
rect 476856 221264 476908 221270
rect 476856 221206 476908 221212
rect 476868 217410 476896 221206
rect 477788 217410 477816 226034
rect 478510 224768 478566 224777
rect 478510 224703 478566 224712
rect 478524 217410 478552 224703
rect 479340 224596 479392 224602
rect 479340 224538 479392 224544
rect 479352 217410 479380 224538
rect 480272 223650 480300 228482
rect 480260 223644 480312 223650
rect 480260 223586 480312 223592
rect 480364 217410 480392 229366
rect 483020 229356 483072 229362
rect 483020 229298 483072 229304
rect 480996 226024 481048 226030
rect 480996 225966 481048 225972
rect 481008 217410 481036 225966
rect 481914 224632 481970 224641
rect 481914 224567 481970 224576
rect 481928 217410 481956 224567
rect 483032 217410 483060 229298
rect 487160 229288 487212 229294
rect 487160 229230 487212 229236
rect 484400 223644 484452 223650
rect 484400 223586 484452 223592
rect 483846 223544 483902 223553
rect 483846 223479 483902 223488
rect 483860 217410 483888 223479
rect 484412 217410 484440 223586
rect 486330 222048 486386 222057
rect 486330 221983 486386 221992
rect 486344 217410 486372 221983
rect 487172 218074 487200 229230
rect 528376 229220 528428 229226
rect 528376 229162 528428 229168
rect 507398 228984 507454 228993
rect 507398 228919 507454 228928
rect 503810 228848 503866 228857
rect 503810 228783 503866 228792
rect 494520 228472 494572 228478
rect 494520 228414 494572 228420
rect 489734 227216 489790 227225
rect 489734 227151 489790 227160
rect 488906 227080 488962 227089
rect 488906 227015 488962 227024
rect 487804 225752 487856 225758
rect 487804 225694 487856 225700
rect 487160 218068 487212 218074
rect 487160 218010 487212 218016
rect 487172 217410 487200 218010
rect 487816 217410 487844 225694
rect 488920 217410 488948 227015
rect 489748 217546 489776 227151
rect 491300 225888 491352 225894
rect 491300 225830 491352 225836
rect 490288 221332 490340 221338
rect 490288 221274 490340 221280
rect 490300 218142 490328 221274
rect 490288 218136 490340 218142
rect 490288 218078 490340 218084
rect 489748 217518 489822 217546
rect 489794 217410 489822 217518
rect 490300 217410 490328 218078
rect 491312 217410 491340 225830
rect 494060 223508 494112 223514
rect 494060 223450 494112 223456
rect 491942 223408 491998 223417
rect 491942 223343 491998 223352
rect 491390 223272 491446 223281
rect 491390 223207 491446 223216
rect 491404 220969 491432 223207
rect 491390 220960 491446 220969
rect 491390 220895 491446 220904
rect 464264 217382 464600 217410
rect 465092 217382 465428 217410
rect 465920 217382 466256 217410
rect 466748 217382 467084 217410
rect 467576 217382 467912 217410
rect 468404 217382 468740 217410
rect 469232 217382 469568 217410
rect 470152 217382 470488 217410
rect 470980 217382 471316 217410
rect 471992 217382 472144 217410
rect 472636 217382 472972 217410
rect 473464 217382 473800 217410
rect 474292 217382 474628 217410
rect 475120 217382 475456 217410
rect 476040 217382 476376 217410
rect 476868 217382 477204 217410
rect 477788 217382 478032 217410
rect 478524 217382 478860 217410
rect 479352 217382 479688 217410
rect 480364 217382 480516 217410
rect 481008 217382 481344 217410
rect 481928 217382 482264 217410
rect 483032 217382 483092 217410
rect 483860 217382 484256 217410
rect 484412 217382 484748 217410
rect 486344 217382 486740 217410
rect 487172 217382 487232 217410
rect 487816 217382 488152 217410
rect 488920 217382 489316 217410
rect 489794 217396 489868 217410
rect 489808 217382 489868 217396
rect 490300 217382 490636 217410
rect 491312 217382 491464 217410
rect 418620 216912 418672 216918
rect 418620 216854 418672 216860
rect 417884 216844 417936 216850
rect 417884 216786 417936 216792
rect 59360 216708 59412 216714
rect 59360 216650 59412 216656
rect 62948 216708 63000 216714
rect 62948 216650 63000 216656
rect 59268 216640 59320 216646
rect 59268 216582 59320 216588
rect 484228 216442 484256 217382
rect 486712 216442 486740 217382
rect 489288 217122 489316 217382
rect 489276 217116 489328 217122
rect 489276 217058 489328 217064
rect 489840 216458 489868 217382
rect 491956 216458 491984 223343
rect 494072 221406 494100 223450
rect 494060 221400 494112 221406
rect 494060 221342 494112 221348
rect 493046 220960 493102 220969
rect 493046 220895 493102 220904
rect 493060 217410 493088 220895
rect 494072 217410 494100 221342
rect 493060 217382 493120 217410
rect 494040 217382 494100 217410
rect 494532 217410 494560 228414
rect 501236 228404 501288 228410
rect 501236 228346 501288 228352
rect 495346 227488 495402 227497
rect 495346 227423 495402 227432
rect 495360 221241 495388 227423
rect 496174 227352 496230 227361
rect 496174 227287 496230 227296
rect 495346 221232 495402 221241
rect 495346 221167 495402 221176
rect 495360 217410 495388 221167
rect 496188 217410 496216 227287
rect 499488 223440 499540 223446
rect 499488 223382 499540 223388
rect 498658 223136 498714 223145
rect 498658 223071 498714 223080
rect 497372 221536 497424 221542
rect 497372 221478 497424 221484
rect 497384 217410 497412 221478
rect 497832 221468 497884 221474
rect 497832 221410 497884 221416
rect 494532 217382 494868 217410
rect 495360 217382 495696 217410
rect 496188 217382 496676 217410
rect 497352 217382 497412 217410
rect 497844 217410 497872 221410
rect 497844 217382 498180 217410
rect 492588 216504 492640 216510
rect 489808 216442 490144 216458
rect 491956 216452 492588 216458
rect 491956 216446 492640 216452
rect 484216 216436 484268 216442
rect 484216 216378 484268 216384
rect 486700 216436 486752 216442
rect 489808 216436 490156 216442
rect 489808 216430 490104 216436
rect 486700 216378 486752 216384
rect 491956 216430 492628 216446
rect 496648 216442 496676 217382
rect 498672 216594 498700 223071
rect 499500 221542 499528 223382
rect 500222 222864 500278 222873
rect 500222 222799 500278 222808
rect 499488 221536 499540 221542
rect 499488 221478 499540 221484
rect 500236 221105 500264 222799
rect 500408 221604 500460 221610
rect 500408 221546 500460 221552
rect 500222 221096 500278 221105
rect 500222 221031 500278 221040
rect 500236 217410 500264 221031
rect 499928 217382 500264 217410
rect 500132 217116 500184 217122
rect 500132 217058 500184 217064
rect 498672 216578 499344 216594
rect 498672 216572 499356 216578
rect 498672 216566 499304 216572
rect 499304 216514 499356 216520
rect 500144 216442 500172 217058
rect 500420 216458 500448 221546
rect 501248 217410 501276 228346
rect 503168 225820 503220 225826
rect 503168 225762 503220 225768
rect 502708 221604 502760 221610
rect 502708 221546 502760 221552
rect 502720 217410 502748 221546
rect 503180 221270 503208 225762
rect 503824 223582 503852 228783
rect 506296 228336 506348 228342
rect 506296 228278 506348 228284
rect 503812 223576 503864 223582
rect 503812 223518 503864 223524
rect 503720 221740 503772 221746
rect 503720 221682 503772 221688
rect 503168 221264 503220 221270
rect 503168 221206 503220 221212
rect 501248 217382 501584 217410
rect 502412 217382 502748 217410
rect 503180 217410 503208 221206
rect 503732 217410 503760 221682
rect 503824 221610 503852 223518
rect 504822 223000 504878 223009
rect 504822 222935 504878 222944
rect 503812 221604 503864 221610
rect 503812 221546 503864 221552
rect 504836 217546 504864 222935
rect 505744 221672 505796 221678
rect 505744 221614 505796 221620
rect 505756 217546 505784 221614
rect 504836 217518 504910 217546
rect 505756 217518 505830 217546
rect 503180 217382 503240 217410
rect 503732 217382 504068 217410
rect 504882 216594 504910 217518
rect 505802 217410 505830 217518
rect 506308 217410 506336 228278
rect 507412 221377 507440 228919
rect 512182 228712 512238 228721
rect 512182 228647 512238 228656
rect 511356 228268 511408 228274
rect 511356 228210 511408 228216
rect 507952 225616 508004 225622
rect 507952 225558 508004 225564
rect 507964 221406 507992 225558
rect 509606 222728 509662 222737
rect 509606 222663 509662 222672
rect 508780 221808 508832 221814
rect 508780 221750 508832 221756
rect 507952 221400 508004 221406
rect 507398 221368 507454 221377
rect 507952 221342 508004 221348
rect 507398 221303 507454 221312
rect 507412 217410 507440 221303
rect 507964 217410 507992 221342
rect 508792 217410 508820 221750
rect 505802 217396 505876 217410
rect 505816 217382 505876 217396
rect 506308 217382 506644 217410
rect 507412 217382 507472 217410
rect 507964 217382 508300 217410
rect 508792 217382 509128 217410
rect 504882 216580 505048 216594
rect 504896 216566 505048 216580
rect 501052 216504 501104 216510
rect 500420 216452 501052 216458
rect 500420 216446 501104 216452
rect 496636 216436 496688 216442
rect 490104 216378 490156 216384
rect 496636 216378 496688 216384
rect 500132 216436 500184 216442
rect 500420 216430 501092 216446
rect 505020 216442 505048 216566
rect 505848 216458 505876 217382
rect 509620 216866 509648 222663
rect 510620 221876 510672 221882
rect 510620 221818 510672 221824
rect 510632 217138 510660 221818
rect 511368 217410 511396 228210
rect 512196 220998 512224 228647
rect 518990 228576 519046 228585
rect 518990 228511 519046 228520
rect 513470 226264 513526 226273
rect 513470 226199 513526 226208
rect 513380 225480 513432 225486
rect 513380 225422 513432 225428
rect 513392 221610 513420 225422
rect 513380 221604 513432 221610
rect 513380 221546 513432 221552
rect 512184 220992 512236 220998
rect 512184 220934 512236 220940
rect 512196 217410 512224 220934
rect 513392 217410 513420 221546
rect 513484 218210 513512 226199
rect 518714 226128 518770 226137
rect 518714 226063 518770 226072
rect 514666 222592 514722 222601
rect 514666 222527 514722 222536
rect 513840 221944 513892 221950
rect 513840 221886 513892 221892
rect 513472 218204 513524 218210
rect 513472 218146 513524 218152
rect 511368 217382 511704 217410
rect 512196 217382 512532 217410
rect 513360 217382 513420 217410
rect 513852 217410 513880 221886
rect 513852 217382 514188 217410
rect 511080 217184 511132 217190
rect 510632 217132 511080 217138
rect 510632 217126 511132 217132
rect 514680 217138 514708 222527
rect 517058 222456 517114 222465
rect 517058 222391 517114 222400
rect 516416 222012 516468 222018
rect 516416 221954 516468 221960
rect 515772 218204 515824 218210
rect 515772 218146 515824 218152
rect 515784 217410 515812 218146
rect 516428 217410 516456 221954
rect 517072 221134 517100 222391
rect 517060 221128 517112 221134
rect 517060 221070 517112 221076
rect 517612 221128 517664 221134
rect 517612 221070 517664 221076
rect 517624 217410 517652 221070
rect 518728 218278 518756 226063
rect 518900 225548 518952 225554
rect 518900 225490 518952 225496
rect 518716 218272 518768 218278
rect 518716 218214 518768 218220
rect 518728 217410 518756 218214
rect 515784 217382 515844 217410
rect 516428 217382 516672 217410
rect 517592 217382 517652 217410
rect 518420 217382 518756 217410
rect 518912 217410 518940 225490
rect 519004 221338 519032 228511
rect 525062 228440 525118 228449
rect 525062 228375 525118 228384
rect 520830 225992 520886 226001
rect 520830 225927 520886 225936
rect 518992 221332 519044 221338
rect 518992 221274 519044 221280
rect 520004 221332 520056 221338
rect 520004 221274 520056 221280
rect 520016 221202 520044 221274
rect 520004 221196 520056 221202
rect 520004 221138 520056 221144
rect 520016 217410 520044 221138
rect 520844 218346 520872 225927
rect 523406 225856 523462 225865
rect 523406 225791 523462 225800
rect 522210 222320 522266 222329
rect 522210 222255 522266 222264
rect 521660 222148 521712 222154
rect 521660 222090 521712 222096
rect 520832 218340 520884 218346
rect 520832 218282 520884 218288
rect 520844 217410 520872 218282
rect 521672 217410 521700 222090
rect 518912 217382 519248 217410
rect 520016 217382 520076 217410
rect 520844 217382 520904 217410
rect 521672 217382 521732 217410
rect 510632 217110 511120 217126
rect 514680 217122 515352 217138
rect 514680 217116 515364 217122
rect 514680 217110 515312 217116
rect 515312 217058 515364 217064
rect 516048 217116 516100 217122
rect 516048 217058 516100 217064
rect 509620 216852 509956 216866
rect 509620 216838 509970 216852
rect 506112 216572 506164 216578
rect 506112 216514 506164 216520
rect 506124 216458 506152 216514
rect 505008 216436 505060 216442
rect 500132 216378 500184 216384
rect 505816 216430 506152 216458
rect 509942 216418 509970 216838
rect 516060 216442 516088 217058
rect 522224 216458 522252 222255
rect 523420 218414 523448 225791
rect 523960 225684 524012 225690
rect 523960 225626 524012 225632
rect 523408 218408 523460 218414
rect 523408 218350 523460 218356
rect 523420 217410 523448 218350
rect 523972 217410 524000 225626
rect 525076 221338 525104 228375
rect 525798 225720 525854 225729
rect 525798 225655 525854 225664
rect 525064 221332 525116 221338
rect 525064 221274 525116 221280
rect 525076 217410 525104 221274
rect 525812 218482 525840 225655
rect 527270 222184 527326 222193
rect 527270 222119 527326 222128
rect 526444 222080 526496 222086
rect 526444 222022 526496 222028
rect 525800 218476 525852 218482
rect 525800 218418 525852 218424
rect 525812 217410 525840 218418
rect 526456 217410 526484 222022
rect 527284 217410 527312 222119
rect 528388 221814 528416 229162
rect 536656 229152 536708 229158
rect 536656 229094 536708 229100
rect 530122 228304 530178 228313
rect 530122 228239 530178 228248
rect 529020 225344 529072 225350
rect 529020 225286 529072 225292
rect 528376 221808 528428 221814
rect 528376 221750 528428 221756
rect 528388 217410 528416 221750
rect 529032 217410 529060 225286
rect 530136 221474 530164 228239
rect 534906 228168 534962 228177
rect 534906 228103 534962 228112
rect 530674 225584 530730 225593
rect 530674 225519 530730 225528
rect 530688 221950 530716 225519
rect 532700 225412 532752 225418
rect 532700 225354 532752 225360
rect 532712 222018 532740 225354
rect 533988 225276 534040 225282
rect 533988 225218 534040 225224
rect 532700 222012 532752 222018
rect 532700 221954 532752 221960
rect 533436 222012 533488 222018
rect 533436 221954 533488 221960
rect 530676 221944 530728 221950
rect 530676 221886 530728 221892
rect 530124 221468 530176 221474
rect 530124 221410 530176 221416
rect 530136 217410 530164 221410
rect 530688 217410 530716 221886
rect 532700 220924 532752 220930
rect 532700 220866 532752 220872
rect 531504 220856 531556 220862
rect 531504 220798 531556 220804
rect 531516 217410 531544 220798
rect 532712 217410 532740 220866
rect 533448 217410 533476 221954
rect 534000 217410 534028 225218
rect 534920 221542 534948 228103
rect 536288 223304 536340 223310
rect 536288 223246 536340 223252
rect 536380 223304 536432 223310
rect 536380 223246 536432 223252
rect 536300 222154 536328 223246
rect 536288 222148 536340 222154
rect 536288 222090 536340 222096
rect 534908 221536 534960 221542
rect 534908 221478 534960 221484
rect 534920 217410 534948 221478
rect 536392 217410 536420 223246
rect 536668 223242 536696 229094
rect 550272 228200 550324 228206
rect 550272 228142 550324 228148
rect 549260 228064 549312 228070
rect 538310 228032 538366 228041
rect 549260 228006 549312 228012
rect 538310 227967 538366 227976
rect 536564 223236 536616 223242
rect 536564 223178 536616 223184
rect 536656 223236 536708 223242
rect 536656 223178 536708 223184
rect 523420 217382 523480 217410
rect 523972 217382 524308 217410
rect 525076 217382 525136 217410
rect 525812 217382 525964 217410
rect 526456 217382 526792 217410
rect 527284 217382 527772 217410
rect 528388 217382 528448 217410
rect 529032 217382 529368 217410
rect 530136 217382 530196 217410
rect 530688 217382 531024 217410
rect 531516 217382 531852 217410
rect 532680 217382 532832 217410
rect 533448 217382 533508 217410
rect 534000 217382 534336 217410
rect 534920 217382 535256 217410
rect 536084 217382 536420 217410
rect 536576 217410 536604 223178
rect 538324 221678 538352 227967
rect 542726 227896 542782 227905
rect 542726 227831 542782 227840
rect 538862 225448 538918 225457
rect 538862 225383 538918 225392
rect 538876 222086 538904 225383
rect 539048 223372 539100 223378
rect 539048 223314 539100 223320
rect 538864 222080 538916 222086
rect 538864 222022 538916 222028
rect 538312 221672 538364 221678
rect 538312 221614 538364 221620
rect 537392 221060 537444 221066
rect 537392 221002 537444 221008
rect 536576 217382 536912 217410
rect 523040 217184 523092 217190
rect 523040 217126 523092 217132
rect 523052 216510 523080 217126
rect 527744 216510 527772 217382
rect 532804 217122 532832 217382
rect 532792 217116 532844 217122
rect 532792 217058 532844 217064
rect 537404 216594 537432 221002
rect 538876 217410 538904 222022
rect 538568 217382 538904 217410
rect 539060 217410 539088 223314
rect 541624 223168 541676 223174
rect 541624 223110 541676 223116
rect 541440 222148 541492 222154
rect 541440 222090 541492 222096
rect 540152 221672 540204 221678
rect 540152 221614 540204 221620
rect 540164 217410 540192 221614
rect 541452 220930 541480 222090
rect 541440 220924 541492 220930
rect 541440 220866 541492 220872
rect 541452 217410 541480 220866
rect 539060 217382 539396 217410
rect 540164 217382 540224 217410
rect 541144 217382 541480 217410
rect 541636 217410 541664 223110
rect 542740 221746 542768 227831
rect 545762 225312 545818 225321
rect 545762 225247 545818 225256
rect 544108 225208 544160 225214
rect 544108 225150 544160 225156
rect 543556 223032 543608 223038
rect 543556 222974 543608 222980
rect 542728 221740 542780 221746
rect 542728 221682 542780 221688
rect 542740 217410 542768 221682
rect 543568 220862 543596 222974
rect 543556 220856 543608 220862
rect 543556 220798 543608 220804
rect 543568 217410 543596 220798
rect 544120 217410 544148 225150
rect 545776 223106 545804 225247
rect 545120 223100 545172 223106
rect 545120 223042 545172 223048
rect 545764 223100 545816 223106
rect 545764 223042 545816 223048
rect 545132 217410 545160 223042
rect 545776 217410 545804 223042
rect 546684 222964 546736 222970
rect 546684 222906 546736 222912
rect 546696 217410 546724 222906
rect 548340 222896 548392 222902
rect 548340 222838 548392 222844
rect 547512 222828 547564 222834
rect 547512 222770 547564 222776
rect 547524 221882 547552 222770
rect 547512 221876 547564 221882
rect 547512 221818 547564 221824
rect 547524 217410 547552 221818
rect 548352 217410 548380 222838
rect 549272 217410 549300 228006
rect 549352 224936 549404 224942
rect 549352 224878 549404 224884
rect 549364 222902 549392 224878
rect 549352 222896 549404 222902
rect 549352 222838 549404 222844
rect 550284 217410 550312 228142
rect 552020 228132 552072 228138
rect 552020 228074 552072 228080
rect 551100 222896 551152 222902
rect 551100 222838 551152 222844
rect 551112 217410 551140 222838
rect 552032 217410 552060 228074
rect 559288 227996 559340 228002
rect 559288 227938 559340 227944
rect 552570 227760 552626 227769
rect 552570 227695 552626 227704
rect 552584 222086 552612 227695
rect 556066 225176 556122 225185
rect 554320 225140 554372 225146
rect 556066 225111 556122 225120
rect 554320 225082 554372 225088
rect 553768 222828 553820 222834
rect 553768 222770 553820 222776
rect 552572 222080 552624 222086
rect 552572 222022 552624 222028
rect 553216 222080 553268 222086
rect 553216 222022 553268 222028
rect 553228 217410 553256 222022
rect 553780 217410 553808 222770
rect 554332 222766 554360 225082
rect 554228 222760 554280 222766
rect 554228 222702 554280 222708
rect 554320 222760 554372 222766
rect 554320 222702 554372 222708
rect 541636 217382 541972 217410
rect 542740 217382 542800 217410
rect 543568 217382 543628 217410
rect 544120 217382 544456 217410
rect 545132 217382 545436 217410
rect 545776 217382 546112 217410
rect 546696 217382 547032 217410
rect 547524 217382 547860 217410
rect 548352 217382 548688 217410
rect 549272 217382 549516 217410
rect 550284 217382 550680 217410
rect 551112 217382 551172 217410
rect 552000 217382 552060 217410
rect 552920 217382 553256 217410
rect 553748 217382 553808 217410
rect 554240 217410 554268 222702
rect 556080 222630 556108 225111
rect 559102 225040 559158 225049
rect 559102 224975 559158 224984
rect 556712 222692 556764 222698
rect 556712 222634 556764 222640
rect 555056 222624 555108 222630
rect 555056 222566 555108 222572
rect 556068 222624 556120 222630
rect 556068 222566 556120 222572
rect 554240 217382 554576 217410
rect 545408 217190 545436 217382
rect 550652 217258 550680 217382
rect 555068 217274 555096 222566
rect 556080 217410 556108 222566
rect 556724 217410 556752 222634
rect 559116 222562 559144 224975
rect 558184 222556 558236 222562
rect 558184 222498 558236 222504
rect 559104 222556 559156 222562
rect 559104 222498 559156 222504
rect 558196 221066 558224 222498
rect 558184 221060 558236 221066
rect 558184 221002 558236 221008
rect 558196 217410 558224 221002
rect 559116 217410 559144 222498
rect 556080 217382 556232 217410
rect 556724 217382 557060 217410
rect 557888 217382 558224 217410
rect 558808 217382 559144 217410
rect 559300 217410 559328 227938
rect 560392 227792 560444 227798
rect 560392 227734 560444 227740
rect 560404 217410 560432 227734
rect 563704 225072 563756 225078
rect 563704 225014 563756 225020
rect 563716 222494 563744 225014
rect 561772 222488 561824 222494
rect 561772 222430 561824 222436
rect 563704 222488 563756 222494
rect 563704 222430 563756 222436
rect 561588 222420 561640 222426
rect 561588 222362 561640 222368
rect 560760 217456 560812 217462
rect 559300 217382 559636 217410
rect 560404 217404 560760 217410
rect 561600 217410 561628 222362
rect 560404 217398 560812 217404
rect 560404 217382 560800 217398
rect 561292 217382 561628 217410
rect 561784 217410 561812 222430
rect 562968 222352 563020 222358
rect 562968 222294 563020 222300
rect 562980 217410 563008 222294
rect 561784 217382 562120 217410
rect 562948 217382 563008 217410
rect 563716 217410 563744 222430
rect 564360 221785 564388 248406
rect 564532 245676 564584 245682
rect 564532 245618 564584 245624
rect 564440 227928 564492 227934
rect 564440 227870 564492 227876
rect 564346 221776 564402 221785
rect 564346 221711 564402 221720
rect 564452 217410 564480 227870
rect 564544 221513 564572 245618
rect 565452 227860 565504 227866
rect 565452 227802 565504 227808
rect 564530 221504 564586 221513
rect 564530 221439 564586 221448
rect 565464 217410 565492 227802
rect 566004 225004 566056 225010
rect 566004 224946 566056 224952
rect 566016 222970 566044 224946
rect 566004 222964 566056 222970
rect 566004 222906 566056 222912
rect 566016 217410 566044 222906
rect 566832 222284 566884 222290
rect 566832 222226 566884 222232
rect 566844 217410 566872 222226
rect 567120 221649 567148 251194
rect 648632 231334 648660 277578
rect 648724 269142 648752 278038
rect 654140 277568 654192 277574
rect 654140 277510 654192 277516
rect 648712 269136 648764 269142
rect 648712 269078 648764 269084
rect 648632 231306 650380 231334
rect 570236 227724 570288 227730
rect 570236 227666 570288 227672
rect 569314 227624 569370 227633
rect 569314 227559 569370 227568
rect 568578 224904 568634 224913
rect 568578 224839 568634 224848
rect 568592 222698 568620 224839
rect 568580 222692 568632 222698
rect 568580 222634 568632 222640
rect 567660 222216 567712 222222
rect 567660 222158 567712 222164
rect 567106 221640 567162 221649
rect 567106 221575 567162 221584
rect 567672 217410 567700 222158
rect 567982 217524 568034 217530
rect 567982 217466 568034 217472
rect 567994 217410 568022 217466
rect 563716 217382 563776 217410
rect 564452 217382 564696 217410
rect 565464 217394 565768 217410
rect 565464 217388 565780 217394
rect 565464 217382 565728 217388
rect 566016 217382 566352 217410
rect 566844 217382 567180 217410
rect 567672 217396 568022 217410
rect 568592 217410 568620 222634
rect 569328 217410 569356 227559
rect 570248 222290 570276 227666
rect 623412 223576 623464 223582
rect 623412 223518 623464 223524
rect 607588 223508 607640 223514
rect 607588 223450 607640 223456
rect 570236 222284 570288 222290
rect 570236 222226 570288 222232
rect 570880 222284 570932 222290
rect 570880 222226 570932 222232
rect 570892 217410 570920 222226
rect 574374 221640 574430 221649
rect 574374 221575 574430 221584
rect 573546 221504 573602 221513
rect 573546 221439 573602 221448
rect 567672 217382 568008 217396
rect 568592 217382 568836 217410
rect 569328 217382 569664 217410
rect 570584 217382 570920 217410
rect 573560 217410 573588 221439
rect 574388 217410 574416 221575
rect 575202 221504 575258 221513
rect 575202 221439 575258 221448
rect 575216 217410 575244 221439
rect 607128 218136 607180 218142
rect 607128 218078 607180 218084
rect 606668 218068 606720 218074
rect 606668 218010 606720 218016
rect 573560 217382 573896 217410
rect 574388 217382 574724 217410
rect 575216 217382 575552 217410
rect 565728 217330 565780 217336
rect 555700 217320 555752 217326
rect 555068 217268 555700 217274
rect 555068 217262 555752 217268
rect 550640 217252 550692 217258
rect 555068 217246 555740 217262
rect 550640 217194 550692 217200
rect 545396 217184 545448 217190
rect 545396 217126 545448 217132
rect 537404 216578 538076 216594
rect 537404 216572 538088 216578
rect 537404 216566 538036 216572
rect 538036 216514 538088 216520
rect 523040 216504 523092 216510
rect 522224 216442 522896 216458
rect 523040 216446 523092 216452
rect 527732 216504 527784 216510
rect 527732 216446 527784 216452
rect 516048 216436 516100 216442
rect 509942 216404 509978 216418
rect 505008 216378 505060 216384
rect 509932 216352 509938 216404
rect 509990 216352 509996 216404
rect 522224 216436 522908 216442
rect 522224 216430 522856 216436
rect 516048 216378 516100 216384
rect 522856 216378 522908 216384
rect 582286 216200 582342 216209
rect 582286 216135 582342 216144
rect 582300 215354 582328 216135
rect 582288 215348 582340 215354
rect 582288 215290 582340 215296
rect 600044 215348 600096 215354
rect 600044 215290 600096 215296
rect 582286 214704 582342 214713
rect 582286 214639 582342 214648
rect 580262 213208 580318 213217
rect 580262 213143 580318 213152
rect 580276 212566 580304 213143
rect 582300 212634 582328 214639
rect 582288 212628 582340 212634
rect 582288 212570 582340 212576
rect 599952 212628 600004 212634
rect 599952 212570 600004 212576
rect 580264 212560 580316 212566
rect 580264 212502 580316 212508
rect 599860 212560 599912 212566
rect 599860 212502 599912 212508
rect 580078 211712 580134 211721
rect 580078 211647 580134 211656
rect 580092 209846 580120 211647
rect 582286 210216 582342 210225
rect 582286 210151 582342 210160
rect 582300 209914 582328 210151
rect 582288 209908 582340 209914
rect 582288 209850 582340 209856
rect 580080 209840 580132 209846
rect 580080 209782 580132 209788
rect 581458 208720 581514 208729
rect 581458 208655 581514 208664
rect 581472 207058 581500 208655
rect 599872 207505 599900 212502
rect 599964 208593 599992 212570
rect 600056 209545 600084 215290
rect 606680 210202 606708 218010
rect 607140 210202 607168 218078
rect 607600 210202 607628 223450
rect 608048 223440 608100 223446
rect 608048 223382 608100 223388
rect 608060 210202 608088 223382
rect 615040 223236 615092 223242
rect 615040 223178 615092 223184
rect 614580 222012 614632 222018
rect 614580 221954 614632 221960
rect 614028 221944 614080 221950
rect 614028 221886 614080 221892
rect 613568 221808 613620 221814
rect 613568 221750 613620 221756
rect 610808 221604 610860 221610
rect 610808 221546 610860 221552
rect 609888 221400 609940 221406
rect 609888 221342 609940 221348
rect 608968 221264 609020 221270
rect 608968 221206 609020 221212
rect 608508 216232 608560 216238
rect 608508 216174 608560 216180
rect 608520 210202 608548 216174
rect 608980 210202 609008 221206
rect 609428 216368 609480 216374
rect 609428 216310 609480 216316
rect 609440 210202 609468 216310
rect 609900 210202 609928 221342
rect 610348 216436 610400 216442
rect 610348 216378 610400 216384
rect 610360 210202 610388 216378
rect 610820 210202 610848 221546
rect 613108 218476 613160 218482
rect 613108 218418 613160 218424
rect 612648 218408 612700 218414
rect 612648 218350 612700 218356
rect 612188 218340 612240 218346
rect 612188 218282 612240 218288
rect 611728 218272 611780 218278
rect 611728 218214 611780 218220
rect 611268 218204 611320 218210
rect 611268 218146 611320 218152
rect 611280 210202 611308 218146
rect 611740 210202 611768 218214
rect 612200 210202 612228 218282
rect 612660 210202 612688 218350
rect 613120 210202 613148 218418
rect 613580 210202 613608 221750
rect 614040 210202 614068 221886
rect 614592 210202 614620 221954
rect 615052 210202 615080 223178
rect 616880 223100 616932 223106
rect 616880 223042 616932 223048
rect 615500 222148 615552 222154
rect 615500 222090 615552 222096
rect 615512 210202 615540 222090
rect 615960 220924 616012 220930
rect 615960 220866 616012 220872
rect 615972 210202 616000 220866
rect 616420 220856 616472 220862
rect 616420 220798 616472 220804
rect 616432 210202 616460 220798
rect 616892 210202 616920 223042
rect 617340 223032 617392 223038
rect 617340 222974 617392 222980
rect 617352 210202 617380 222974
rect 620560 222964 620612 222970
rect 620560 222906 620612 222912
rect 617800 222896 617852 222902
rect 617800 222838 617852 222844
rect 617812 210202 617840 222838
rect 618260 222760 618312 222766
rect 618260 222702 618312 222708
rect 618272 210202 618300 222702
rect 618720 222624 618772 222630
rect 618720 222566 618772 222572
rect 618732 210202 618760 222566
rect 619180 222556 619232 222562
rect 619180 222498 619232 222504
rect 619192 210202 619220 222498
rect 620100 222488 620152 222494
rect 620100 222430 620152 222436
rect 619640 222420 619692 222426
rect 619640 222362 619692 222368
rect 619652 210202 619680 222362
rect 620112 210202 620140 222430
rect 620572 210202 620600 222906
rect 621020 222692 621072 222698
rect 621020 222634 621072 222640
rect 621032 210202 621060 222634
rect 622490 221232 622546 221241
rect 622490 221167 622546 221176
rect 622032 215892 622084 215898
rect 622032 215834 622084 215840
rect 621480 215824 621532 215830
rect 621480 215766 621532 215772
rect 621492 210202 621520 215766
rect 622044 210202 622072 215834
rect 622504 210202 622532 221167
rect 622952 215960 623004 215966
rect 622952 215902 623004 215908
rect 622964 210202 622992 215902
rect 623424 210202 623452 223518
rect 634544 222352 634596 222358
rect 634544 222294 634596 222300
rect 632704 222080 632756 222086
rect 632704 222022 632756 222028
rect 631784 221876 631836 221882
rect 631784 221818 631836 221824
rect 630864 221740 630916 221746
rect 630864 221682 630916 221688
rect 630404 221672 630456 221678
rect 630404 221614 630456 221620
rect 629484 221536 629536 221542
rect 629484 221478 629536 221484
rect 628472 221468 628524 221474
rect 628472 221410 628524 221416
rect 624330 221368 624386 221377
rect 624330 221303 624386 221312
rect 627552 221332 627604 221338
rect 623872 216028 623924 216034
rect 623872 215970 623924 215976
rect 623884 210202 623912 215970
rect 624344 210202 624372 221303
rect 627552 221274 627604 221280
rect 626632 221196 626684 221202
rect 626632 221138 626684 221144
rect 626172 221128 626224 221134
rect 626172 221070 626224 221076
rect 625252 220992 625304 220998
rect 625252 220934 625304 220940
rect 624792 216096 624844 216102
rect 624792 216038 624844 216044
rect 624804 210202 624832 216038
rect 625264 210202 625292 220934
rect 625712 216164 625764 216170
rect 625712 216106 625764 216112
rect 625724 210202 625752 216106
rect 626184 210202 626212 221070
rect 626644 210202 626672 221138
rect 627092 216300 627144 216306
rect 627092 216242 627144 216248
rect 627104 210202 627132 216242
rect 627564 210202 627592 221274
rect 628012 216504 628064 216510
rect 628012 216446 628064 216452
rect 628024 210202 628052 216446
rect 628484 210202 628512 221410
rect 628932 217116 628984 217122
rect 628932 217058 628984 217064
rect 628944 210202 628972 217058
rect 629496 210202 629524 221478
rect 629944 216572 629996 216578
rect 629944 216514 629996 216520
rect 629956 210202 629984 216514
rect 630416 210202 630444 221614
rect 630876 210202 630904 221682
rect 631324 217184 631376 217190
rect 631324 217126 631376 217132
rect 631336 210202 631364 217126
rect 631796 210202 631824 221818
rect 632244 217252 632296 217258
rect 632244 217194 632296 217200
rect 632256 210202 632284 217194
rect 632716 210202 632744 222022
rect 633624 221060 633676 221066
rect 633624 221002 633676 221008
rect 633164 217320 633216 217326
rect 633164 217262 633216 217268
rect 633176 210202 633204 217262
rect 633636 210202 633664 221002
rect 634084 217456 634136 217462
rect 634084 217398 634136 217404
rect 634096 210202 634124 217398
rect 634556 210202 634584 222294
rect 635924 222284 635976 222290
rect 635924 222226 635976 222232
rect 635464 217524 635516 217530
rect 635464 217466 635516 217472
rect 635004 217388 635056 217394
rect 635004 217330 635056 217336
rect 635016 210202 635044 217330
rect 635476 210202 635504 217466
rect 635936 210202 635964 222226
rect 637854 221096 637910 221105
rect 637854 221031 637910 221040
rect 636934 220960 636990 220969
rect 636934 220895 636990 220904
rect 636384 215688 636436 215694
rect 636384 215630 636436 215636
rect 636396 210202 636424 215630
rect 636948 210202 636976 220895
rect 637396 215756 637448 215762
rect 637396 215698 637448 215704
rect 637408 210202 637436 215698
rect 637868 210202 637896 221031
rect 650352 220346 650380 231306
rect 649552 220318 650380 220346
rect 639696 217048 639748 217054
rect 639696 216990 639748 216996
rect 638316 215620 638368 215626
rect 638316 215562 638368 215568
rect 638328 210202 638356 215562
rect 638776 215552 638828 215558
rect 638776 215494 638828 215500
rect 638788 210202 638816 215494
rect 639708 210202 639736 216990
rect 640616 216980 640668 216986
rect 640616 216922 640668 216928
rect 640156 216912 640208 216918
rect 640156 216854 640208 216860
rect 640168 210202 640196 216854
rect 640628 210202 640656 216922
rect 641076 216844 641128 216850
rect 641076 216786 641128 216792
rect 641088 210202 641116 216786
rect 648528 216776 648580 216782
rect 648528 216718 648580 216724
rect 643204 210310 643508 210338
rect 643204 210202 643232 210310
rect 606648 210174 606708 210202
rect 607108 210174 607168 210202
rect 607568 210174 607628 210202
rect 608028 210174 608088 210202
rect 608488 210174 608548 210202
rect 608948 210174 609008 210202
rect 609408 210174 609468 210202
rect 609868 210174 609928 210202
rect 610328 210174 610388 210202
rect 610788 210174 610848 210202
rect 611248 210174 611308 210202
rect 611708 210174 611768 210202
rect 612168 210174 612228 210202
rect 612628 210174 612688 210202
rect 613088 210174 613148 210202
rect 613548 210174 613608 210202
rect 614008 210174 614068 210202
rect 614560 210174 614620 210202
rect 615020 210174 615080 210202
rect 615480 210174 615540 210202
rect 615940 210174 616000 210202
rect 616400 210174 616460 210202
rect 616860 210174 616920 210202
rect 617320 210174 617380 210202
rect 617780 210174 617840 210202
rect 618240 210174 618300 210202
rect 618700 210174 618760 210202
rect 619160 210174 619220 210202
rect 619620 210174 619680 210202
rect 620080 210174 620140 210202
rect 620540 210174 620600 210202
rect 621000 210174 621060 210202
rect 621460 210174 621520 210202
rect 622012 210174 622072 210202
rect 622472 210174 622532 210202
rect 622932 210174 622992 210202
rect 623392 210174 623452 210202
rect 623852 210174 623912 210202
rect 624312 210174 624372 210202
rect 624772 210174 624832 210202
rect 625232 210174 625292 210202
rect 625692 210174 625752 210202
rect 626152 210174 626212 210202
rect 626612 210174 626672 210202
rect 627072 210174 627132 210202
rect 627532 210174 627592 210202
rect 627992 210174 628052 210202
rect 628452 210174 628512 210202
rect 628912 210174 628972 210202
rect 629464 210174 629524 210202
rect 629924 210174 629984 210202
rect 630384 210174 630444 210202
rect 630844 210174 630904 210202
rect 631304 210174 631364 210202
rect 631764 210174 631824 210202
rect 632224 210174 632284 210202
rect 632684 210174 632744 210202
rect 633144 210174 633204 210202
rect 633604 210174 633664 210202
rect 634064 210174 634124 210202
rect 634524 210174 634584 210202
rect 634984 210174 635044 210202
rect 635444 210174 635504 210202
rect 635904 210174 635964 210202
rect 636364 210174 636424 210202
rect 636916 210174 636976 210202
rect 637376 210174 637436 210202
rect 637836 210174 637896 210202
rect 638296 210174 638356 210202
rect 638756 210174 638816 210202
rect 639676 210174 639736 210202
rect 640136 210174 640196 210202
rect 640596 210174 640656 210202
rect 641056 210174 641116 210202
rect 642896 210174 643232 210202
rect 643480 210066 643508 210310
rect 646056 210310 646360 210338
rect 646056 210202 646084 210310
rect 645748 210174 646084 210202
rect 646332 210066 646360 210310
rect 648540 210202 648568 216718
rect 648816 210310 649120 210338
rect 648816 210202 648844 210310
rect 648508 210174 648844 210202
rect 649092 210066 649120 210310
rect 649552 210066 649580 220318
rect 651288 220040 651340 220046
rect 651288 219982 651340 219988
rect 650196 210310 650500 210338
rect 650196 210066 650224 210310
rect 643480 210038 643816 210066
rect 646332 210038 646668 210066
rect 649092 210038 649428 210066
rect 649552 210038 650224 210066
rect 650472 210066 650500 210310
rect 651300 210202 651328 219982
rect 652758 217288 652814 217297
rect 652758 217223 652814 217232
rect 651668 210310 651972 210338
rect 651668 210202 651696 210310
rect 651268 210174 651696 210202
rect 651944 210066 651972 210310
rect 652772 210202 652800 217223
rect 653048 210310 653352 210338
rect 653048 210202 653076 210310
rect 652740 210174 653076 210202
rect 653324 210066 653352 210310
rect 654152 210202 654180 277510
rect 655440 220862 655468 292703
rect 655518 291544 655574 291553
rect 655518 291479 655574 291488
rect 655532 221066 655560 291479
rect 655624 245614 655652 293927
rect 655702 290456 655758 290465
rect 655702 290391 655758 290400
rect 655612 245608 655664 245614
rect 655612 245550 655664 245556
rect 655716 221202 655744 290391
rect 655808 267782 655836 296239
rect 655978 295352 656034 295361
rect 655978 295287 656034 295296
rect 655992 267986 656020 295287
rect 656176 268122 656204 297463
rect 667020 289128 667072 289134
rect 667020 289070 667072 289076
rect 656806 287328 656862 287337
rect 656806 287263 656808 287272
rect 656860 287263 656862 287272
rect 666836 287292 666888 287298
rect 656808 287234 656860 287240
rect 666836 287234 666888 287240
rect 666744 284708 666796 284714
rect 666744 284650 666796 284656
rect 666652 278792 666704 278798
rect 666652 278734 666704 278740
rect 666560 277432 666612 277438
rect 666560 277374 666612 277380
rect 656164 268116 656216 268122
rect 656164 268058 656216 268064
rect 655980 267980 656032 267986
rect 655980 267922 656032 267928
rect 655796 267776 655848 267782
rect 655796 267718 655848 267724
rect 656900 230716 656952 230722
rect 656900 230658 656952 230664
rect 656912 226334 656940 230658
rect 659752 230648 659804 230654
rect 659752 230590 659804 230596
rect 659660 230580 659712 230586
rect 659660 230522 659712 230528
rect 656912 226306 657952 226334
rect 655704 221196 655756 221202
rect 655704 221138 655756 221144
rect 655520 221060 655572 221066
rect 655520 221002 655572 221008
rect 655428 220856 655480 220862
rect 655428 220798 655480 220804
rect 655520 219972 655572 219978
rect 655520 219914 655572 219920
rect 654428 210310 654732 210338
rect 654428 210202 654456 210310
rect 654120 210174 654456 210202
rect 654704 210066 654732 210310
rect 655532 210202 655560 219914
rect 656900 219768 656952 219774
rect 656900 219710 656952 219716
rect 655808 210310 656112 210338
rect 655808 210202 655836 210310
rect 655500 210174 655836 210202
rect 656084 210066 656112 210310
rect 656912 210202 656940 219710
rect 657188 210310 657492 210338
rect 657188 210202 657216 210310
rect 656880 210174 657216 210202
rect 657464 210066 657492 210310
rect 657924 210066 657952 226306
rect 659672 210338 659700 230522
rect 659764 226334 659792 230590
rect 662788 230512 662840 230518
rect 662788 230454 662840 230460
rect 659764 226306 660804 226334
rect 658568 210310 658872 210338
rect 659672 210310 659792 210338
rect 658568 210066 658596 210310
rect 650472 210038 650808 210066
rect 651944 210038 652280 210066
rect 653324 210038 653660 210066
rect 654704 210038 655040 210066
rect 656084 210038 656420 210066
rect 657464 210038 657800 210066
rect 657924 210038 658596 210066
rect 658844 210066 658872 210310
rect 659764 210202 659792 210310
rect 660040 210310 660344 210338
rect 660040 210202 660068 210310
rect 659732 210174 660068 210202
rect 660316 210066 660344 210310
rect 660776 210066 660804 226306
rect 662512 219496 662564 219502
rect 662512 219438 662564 219444
rect 661420 210310 661724 210338
rect 661420 210066 661448 210310
rect 658844 210038 659272 210066
rect 660316 210038 660652 210066
rect 660776 210038 661448 210066
rect 661696 210066 661724 210310
rect 662524 210202 662552 219438
rect 662492 210174 662552 210202
rect 662800 210118 662828 230454
rect 664352 219904 664404 219910
rect 664352 219846 664404 219852
rect 663892 219836 663944 219842
rect 663892 219778 663944 219784
rect 662972 219700 663024 219706
rect 662972 219642 663024 219648
rect 662984 210202 663012 219642
rect 663432 216708 663484 216714
rect 663432 216650 663484 216656
rect 663444 210202 663472 216650
rect 663904 210202 663932 219778
rect 664364 210202 664392 219846
rect 665732 217592 665784 217598
rect 665732 217534 665784 217540
rect 665272 215416 665324 215422
rect 665272 215358 665324 215364
rect 665284 210202 665312 215358
rect 665744 210202 665772 217534
rect 666572 216578 666600 277374
rect 666560 216572 666612 216578
rect 666560 216514 666612 216520
rect 666192 215484 666244 215490
rect 666192 215426 666244 215432
rect 666204 210202 666232 215426
rect 662952 210174 663012 210202
rect 663412 210174 663472 210202
rect 663872 210174 663932 210202
rect 664332 210174 664392 210202
rect 665252 210174 665312 210202
rect 665712 210174 665772 210202
rect 666172 210174 666232 210202
rect 662788 210112 662840 210118
rect 661696 210038 662032 210066
rect 662788 210054 662840 210060
rect 664444 210112 664496 210118
rect 664496 210060 664792 210066
rect 664444 210054 664792 210060
rect 664456 210038 664792 210054
rect 601148 209908 601200 209914
rect 601148 209850 601200 209856
rect 600780 209840 600832 209846
rect 600780 209782 600832 209788
rect 600042 209536 600098 209545
rect 600042 209471 600098 209480
rect 599950 208584 600006 208593
rect 599950 208519 600006 208528
rect 599858 207496 599914 207505
rect 599858 207431 599914 207440
rect 582288 207120 582340 207126
rect 582286 207088 582288 207097
rect 599676 207120 599728 207126
rect 582340 207088 582342 207097
rect 581460 207052 581512 207058
rect 599676 207062 599728 207068
rect 582286 207023 582342 207032
rect 581460 206994 581512 207000
rect 582286 205592 582342 205601
rect 582286 205527 582342 205536
rect 582300 204338 582328 205527
rect 582288 204332 582340 204338
rect 582288 204274 582340 204280
rect 580722 204096 580778 204105
rect 580722 204031 580778 204040
rect 580736 201550 580764 204031
rect 599688 203425 599716 207062
rect 600792 206553 600820 209782
rect 600778 206544 600834 206553
rect 600778 206479 600834 206488
rect 601160 205465 601188 209850
rect 641812 209840 641864 209846
rect 641516 209788 641812 209794
rect 641516 209782 641864 209788
rect 642088 209840 642140 209846
rect 644664 209840 644716 209846
rect 642140 209788 642436 209794
rect 642088 209782 642436 209788
rect 641516 209766 641852 209782
rect 642100 209766 642436 209782
rect 644368 209788 644664 209794
rect 644368 209782 644716 209788
rect 644940 209840 644992 209846
rect 647424 209840 647476 209846
rect 644992 209788 645288 209794
rect 644940 209782 645288 209788
rect 644368 209766 644704 209782
rect 644952 209766 645288 209782
rect 647128 209788 647424 209794
rect 647128 209782 647476 209788
rect 647700 209840 647752 209846
rect 647752 209788 648048 209794
rect 647700 209782 648048 209788
rect 647128 209766 647464 209782
rect 647712 209766 648048 209782
rect 666558 209264 666614 209273
rect 666558 209199 666614 209208
rect 601608 207052 601660 207058
rect 601608 206994 601660 207000
rect 601146 205456 601202 205465
rect 601146 205391 601202 205400
rect 601620 204513 601648 206994
rect 666572 205873 666600 209199
rect 666558 205864 666614 205873
rect 666558 205799 666614 205808
rect 601606 204504 601662 204513
rect 601606 204439 601662 204448
rect 599952 204332 600004 204338
rect 599952 204274 600004 204280
rect 599674 203416 599730 203425
rect 599674 203351 599730 203360
rect 581090 202600 581146 202609
rect 581090 202535 581146 202544
rect 581104 201618 581132 202535
rect 599964 202473 599992 204274
rect 666558 204232 666614 204241
rect 666558 204167 666614 204176
rect 599950 202464 600006 202473
rect 599950 202399 600006 202408
rect 581092 201612 581144 201618
rect 581092 201554 581144 201560
rect 599952 201612 600004 201618
rect 599952 201554 600004 201560
rect 580724 201544 580776 201550
rect 580724 201486 580776 201492
rect 598940 201544 598992 201550
rect 598940 201486 598992 201492
rect 598952 201385 598980 201486
rect 598938 201376 598994 201385
rect 598938 201311 598994 201320
rect 581090 201104 581146 201113
rect 581090 201039 581146 201048
rect 581104 200122 581132 201039
rect 599964 200433 599992 201554
rect 666572 200841 666600 204167
rect 666558 200832 666614 200841
rect 666558 200767 666614 200776
rect 599950 200424 600006 200433
rect 599950 200359 600006 200368
rect 581092 200116 581144 200122
rect 581092 200058 581144 200064
rect 599952 200116 600004 200122
rect 599952 200058 600004 200064
rect 582286 199608 582342 199617
rect 582286 199543 582342 199552
rect 582300 198762 582328 199543
rect 599964 199345 599992 200058
rect 599950 199336 600006 199345
rect 599950 199271 600006 199280
rect 666558 199064 666614 199073
rect 666558 198999 666614 199008
rect 582288 198756 582340 198762
rect 582288 198698 582340 198704
rect 599952 198756 600004 198762
rect 599952 198698 600004 198704
rect 599964 198393 599992 198698
rect 599950 198384 600006 198393
rect 599950 198319 600006 198328
rect 582286 197976 582342 197985
rect 582286 197911 582342 197920
rect 582300 197402 582328 197911
rect 582288 197396 582340 197402
rect 582288 197338 582340 197344
rect 599400 197396 599452 197402
rect 599400 197338 599452 197344
rect 580724 197328 580776 197334
rect 580724 197270 580776 197276
rect 580736 196489 580764 197270
rect 580722 196480 580778 196489
rect 580722 196415 580778 196424
rect 599412 196353 599440 197338
rect 599952 197328 600004 197334
rect 599950 197296 599952 197305
rect 600004 197296 600006 197305
rect 599950 197231 600006 197240
rect 599398 196344 599454 196353
rect 599398 196279 599454 196288
rect 666572 195673 666600 198999
rect 666558 195664 666614 195673
rect 666558 195599 666614 195608
rect 599858 195256 599914 195265
rect 599858 195191 599914 195200
rect 582286 194984 582342 194993
rect 582286 194919 582342 194928
rect 582196 194676 582248 194682
rect 582196 194618 582248 194624
rect 582208 193497 582236 194618
rect 582300 194614 582328 194919
rect 599872 194614 599900 195191
rect 599952 194676 600004 194682
rect 599952 194618 600004 194624
rect 582288 194608 582340 194614
rect 582288 194550 582340 194556
rect 599860 194608 599912 194614
rect 599860 194550 599912 194556
rect 599964 194313 599992 194618
rect 599950 194304 600006 194313
rect 599950 194239 600006 194248
rect 582194 193488 582250 193497
rect 582194 193423 582250 193432
rect 599490 193216 599546 193225
rect 599490 193151 599546 193160
rect 582286 191992 582342 192001
rect 582286 191927 582342 191936
rect 582300 191894 582328 191927
rect 599504 191894 599532 193151
rect 599950 192264 600006 192273
rect 599950 192199 600006 192208
rect 582288 191888 582340 191894
rect 582288 191830 582340 191836
rect 599492 191888 599544 191894
rect 599492 191830 599544 191836
rect 599964 191826 599992 192199
rect 581276 191820 581328 191826
rect 581276 191762 581328 191768
rect 599952 191820 600004 191826
rect 599952 191762 600004 191768
rect 581288 190505 581316 191762
rect 599950 191176 600006 191185
rect 599950 191111 600006 191120
rect 581274 190496 581330 190505
rect 579712 190460 579764 190466
rect 599964 190466 599992 191111
rect 581274 190431 581330 190440
rect 599952 190460 600004 190466
rect 579712 190402 579764 190408
rect 599952 190402 600004 190408
rect 579724 188873 579752 190402
rect 601514 190224 601570 190233
rect 601514 190159 601570 190168
rect 579710 188864 579766 188873
rect 579710 188799 579766 188808
rect 599122 188184 599178 188193
rect 599122 188119 599178 188128
rect 582288 187672 582340 187678
rect 582288 187614 582340 187620
rect 579896 187604 579948 187610
rect 579896 187546 579948 187552
rect 579908 185881 579936 187546
rect 582300 187377 582328 187614
rect 582286 187368 582342 187377
rect 582286 187303 582342 187312
rect 579894 185872 579950 185881
rect 579894 185807 579950 185816
rect 580264 184884 580316 184890
rect 580264 184826 580316 184832
rect 580276 182889 580304 184826
rect 599136 184822 599164 188119
rect 601528 187678 601556 190159
rect 601606 189136 601662 189145
rect 601606 189071 601662 189080
rect 601516 187672 601568 187678
rect 601516 187614 601568 187620
rect 601620 187610 601648 189071
rect 666558 189000 666614 189009
rect 666558 188935 666614 188944
rect 601608 187604 601660 187610
rect 601608 187546 601660 187552
rect 599950 187096 600006 187105
rect 599950 187031 600006 187040
rect 599858 185056 599914 185065
rect 599858 184991 599914 185000
rect 580908 184816 580960 184822
rect 580908 184758 580960 184764
rect 599124 184816 599176 184822
rect 599124 184758 599176 184764
rect 580920 184385 580948 184758
rect 580906 184376 580962 184385
rect 580906 184311 580962 184320
rect 598938 183016 598994 183025
rect 598938 182951 598994 182960
rect 580262 182880 580318 182889
rect 580262 182815 580318 182824
rect 580632 182164 580684 182170
rect 580632 182106 580684 182112
rect 580540 182096 580592 182102
rect 580540 182038 580592 182044
rect 580552 179761 580580 182038
rect 580644 181393 580672 182106
rect 580630 181384 580686 181393
rect 580630 181319 580686 181328
rect 580538 179752 580594 179761
rect 580538 179687 580594 179696
rect 598952 179382 598980 182951
rect 599872 182102 599900 184991
rect 599964 184890 599992 187031
rect 600042 186144 600098 186153
rect 600042 186079 600098 186088
rect 599952 184884 600004 184890
rect 599952 184826 600004 184832
rect 599950 184104 600006 184113
rect 599950 184039 600006 184048
rect 599860 182096 599912 182102
rect 599860 182038 599912 182044
rect 599858 180024 599914 180033
rect 599858 179959 599914 179968
rect 580724 179376 580776 179382
rect 580724 179318 580776 179324
rect 598940 179376 598992 179382
rect 598940 179318 598992 179324
rect 580736 176769 580764 179318
rect 581092 179308 581144 179314
rect 581092 179250 581144 179256
rect 581104 178265 581132 179250
rect 599674 178936 599730 178945
rect 599674 178871 599730 178880
rect 581090 178256 581146 178265
rect 581090 178191 581146 178200
rect 580722 176760 580778 176769
rect 580722 176695 580778 176704
rect 581092 176724 581144 176730
rect 581092 176666 581144 176672
rect 579712 173868 579764 173874
rect 579712 173810 579764 173816
rect 579724 172281 579752 173810
rect 579710 172272 579766 172281
rect 579710 172207 579766 172216
rect 579896 171148 579948 171154
rect 579896 171090 579948 171096
rect 579804 168496 579856 168502
rect 579804 168438 579856 168444
rect 579816 158545 579844 168438
rect 579908 161537 579936 171090
rect 580540 171012 580592 171018
rect 580540 170954 580592 170960
rect 580552 170649 580580 170954
rect 580538 170640 580594 170649
rect 580538 170575 580594 170584
rect 580448 168564 580500 168570
rect 580448 168506 580500 168512
rect 580264 168428 580316 168434
rect 580264 168370 580316 168376
rect 580172 168360 580224 168366
rect 580172 168302 580224 168308
rect 580184 166161 580212 168302
rect 580170 166152 580226 166161
rect 580170 166087 580226 166096
rect 580080 162988 580132 162994
rect 580080 162930 580132 162936
rect 579894 161528 579950 161537
rect 579894 161463 579950 161472
rect 579802 158536 579858 158545
rect 579802 158471 579858 158480
rect 580092 149433 580120 162930
rect 580276 155553 580304 168370
rect 580460 157049 580488 168506
rect 581104 167657 581132 176666
rect 581460 176656 581512 176662
rect 581460 176598 581512 176604
rect 581472 175273 581500 176598
rect 581458 175264 581514 175273
rect 581458 175199 581514 175208
rect 581644 173936 581696 173942
rect 581644 173878 581696 173884
rect 581090 167648 581146 167657
rect 581090 167583 581146 167592
rect 581276 165640 581328 165646
rect 581276 165582 581328 165588
rect 581184 162920 581236 162926
rect 581184 162862 581236 162868
rect 581092 157548 581144 157554
rect 581092 157490 581144 157496
rect 580908 157480 580960 157486
rect 580908 157422 580960 157428
rect 580632 157412 580684 157418
rect 580632 157354 580684 157360
rect 580446 157040 580502 157049
rect 580446 156975 580502 156984
rect 580262 155544 580318 155553
rect 580262 155479 580318 155488
rect 580540 154624 580592 154630
rect 580540 154566 580592 154572
rect 580078 149424 580134 149433
rect 580078 149359 580134 149368
rect 580552 138825 580580 154566
rect 580644 143313 580672 157354
rect 580724 154692 580776 154698
rect 580724 154634 580776 154640
rect 580630 143304 580686 143313
rect 580630 143239 580686 143248
rect 580538 138816 580594 138825
rect 580538 138751 580594 138760
rect 579712 138100 579764 138106
rect 579712 138042 579764 138048
rect 579724 112985 579752 138042
rect 579896 138032 579948 138038
rect 579896 137974 579948 137980
rect 579710 112976 579766 112985
rect 579710 112911 579766 112920
rect 579908 111489 579936 137974
rect 580736 135833 580764 154634
rect 580816 151836 580868 151842
rect 580816 151778 580868 151784
rect 580722 135824 580778 135833
rect 580722 135759 580778 135768
rect 580080 135380 580132 135386
rect 580080 135322 580132 135328
rect 579988 132524 580040 132530
rect 579988 132466 580040 132472
rect 579894 111480 579950 111489
rect 579894 111415 579950 111424
rect 580000 105369 580028 132466
rect 580092 108497 580120 135322
rect 580172 135312 580224 135318
rect 580172 135254 580224 135260
rect 580078 108488 580134 108497
rect 580078 108423 580134 108432
rect 580184 106865 580212 135254
rect 580828 132705 580856 151778
rect 580920 137329 580948 157422
rect 581104 141817 581132 157490
rect 581196 147937 581224 162862
rect 581288 154057 581316 165582
rect 581656 164665 581684 173878
rect 582288 173800 582340 173806
rect 582286 173768 582288 173777
rect 582340 173768 582342 173777
rect 582286 173703 582342 173712
rect 599490 172816 599546 172825
rect 599490 172751 599546 172760
rect 582104 171216 582156 171222
rect 582104 171158 582156 171164
rect 582012 171080 582064 171086
rect 582012 171022 582064 171028
rect 582024 169153 582052 171022
rect 582010 169144 582066 169153
rect 582010 169079 582066 169088
rect 582116 168374 582144 171158
rect 599504 171154 599532 172751
rect 599492 171148 599544 171154
rect 599492 171090 599544 171096
rect 599688 171018 599716 178871
rect 599766 177984 599822 177993
rect 599766 177919 599822 177928
rect 599780 171086 599808 177919
rect 599872 173874 599900 179959
rect 599964 179314 599992 184039
rect 600056 182170 600084 186079
rect 666572 185609 666600 188935
rect 666558 185600 666614 185609
rect 666558 185535 666614 185544
rect 666558 183832 666614 183841
rect 666558 183767 666614 183776
rect 600044 182164 600096 182170
rect 600044 182106 600096 182112
rect 600042 182064 600098 182073
rect 600042 181999 600098 182008
rect 599952 179308 600004 179314
rect 599952 179250 600004 179256
rect 599950 176896 600006 176905
rect 599950 176831 600006 176840
rect 599964 176730 599992 176831
rect 599952 176724 600004 176730
rect 599952 176666 600004 176672
rect 600056 176662 600084 181999
rect 600134 180976 600190 180985
rect 600134 180911 600190 180920
rect 600044 176656 600096 176662
rect 600044 176598 600096 176604
rect 599950 174856 600006 174865
rect 599950 174791 600006 174800
rect 599964 173942 599992 174791
rect 599952 173936 600004 173942
rect 599952 173878 600004 173884
rect 599860 173868 599912 173874
rect 599860 173810 599912 173816
rect 600148 173806 600176 180911
rect 666572 180441 666600 183767
rect 666558 180432 666614 180441
rect 666558 180367 666614 180376
rect 600410 175944 600466 175953
rect 600410 175879 600466 175888
rect 600136 173800 600188 173806
rect 600136 173742 600188 173748
rect 599950 171864 600006 171873
rect 599950 171799 600006 171808
rect 599964 171222 599992 171799
rect 599952 171216 600004 171222
rect 599952 171158 600004 171164
rect 599768 171080 599820 171086
rect 599768 171022 599820 171028
rect 599676 171012 599728 171018
rect 599676 170954 599728 170960
rect 599858 170776 599914 170785
rect 599858 170711 599914 170720
rect 599490 168736 599546 168745
rect 599490 168671 599546 168680
rect 599504 168434 599532 168671
rect 599872 168502 599900 170711
rect 599950 169824 600006 169833
rect 599950 169759 600006 169768
rect 599964 168570 599992 169759
rect 599952 168564 600004 168570
rect 599952 168506 600004 168512
rect 599860 168496 599912 168502
rect 599860 168438 599912 168444
rect 582024 168346 582144 168374
rect 599492 168428 599544 168434
rect 599492 168370 599544 168376
rect 600424 168366 600452 175879
rect 601330 173904 601386 173913
rect 601330 173839 601386 173848
rect 600412 168360 600464 168366
rect 581828 165572 581880 165578
rect 581828 165514 581880 165520
rect 581642 164656 581698 164665
rect 581642 164591 581698 164600
rect 581840 163169 581868 165514
rect 581826 163160 581882 163169
rect 581826 163095 581882 163104
rect 581644 160200 581696 160206
rect 581644 160142 581696 160148
rect 581274 154048 581330 154057
rect 581274 153983 581330 153992
rect 581552 149184 581604 149190
rect 581552 149126 581604 149132
rect 581368 149116 581420 149122
rect 581368 149058 581420 149064
rect 581182 147928 581238 147937
rect 581182 147863 581238 147872
rect 581276 143608 581328 143614
rect 581276 143550 581328 143556
rect 581090 141808 581146 141817
rect 581090 141743 581146 141752
rect 581000 140888 581052 140894
rect 581000 140830 581052 140836
rect 580906 137320 580962 137329
rect 580906 137255 580962 137264
rect 580814 132696 580870 132705
rect 580814 132631 580870 132640
rect 580908 132660 580960 132666
rect 580908 132602 580960 132608
rect 580264 132592 580316 132598
rect 580264 132534 580316 132540
rect 580170 106856 580226 106865
rect 580170 106791 580226 106800
rect 579986 105360 580042 105369
rect 579986 105295 580042 105304
rect 580276 103873 580304 132534
rect 580356 129940 580408 129946
rect 580356 129882 580408 129888
rect 580262 103864 580318 103873
rect 580262 103799 580318 103808
rect 580368 100881 580396 129882
rect 580632 129872 580684 129878
rect 580632 129814 580684 129820
rect 580448 129804 580500 129810
rect 580448 129746 580500 129752
rect 580354 100872 580410 100881
rect 580354 100807 580410 100816
rect 580460 97753 580488 129746
rect 580540 127016 580592 127022
rect 580540 126958 580592 126964
rect 580446 97744 580502 97753
rect 580446 97679 580502 97688
rect 575664 95260 575716 95266
rect 575664 95202 575716 95208
rect 84824 52686 85160 52714
rect 150328 52686 150388 52714
rect 215832 52686 216168 52714
rect 281336 52686 281488 52714
rect 52276 47116 52328 47122
rect 52276 47058 52328 47064
rect 85132 45762 85160 52686
rect 145380 52488 145432 52494
rect 145380 52430 145432 52436
rect 145392 50810 145420 52430
rect 145084 50782 145420 50810
rect 150360 48346 150388 52686
rect 198648 52488 198700 52494
rect 198648 52430 198700 52436
rect 198660 51066 198688 52430
rect 213828 51128 213880 51134
rect 213828 51070 213880 51076
rect 198648 51060 198700 51066
rect 198648 51002 198700 51008
rect 207020 51060 207072 51066
rect 207020 51002 207072 51008
rect 150348 48340 150400 48346
rect 150348 48282 150400 48288
rect 150360 47122 150388 48282
rect 150348 47116 150400 47122
rect 150348 47058 150400 47064
rect 141804 46702 142370 46730
rect 85120 45756 85172 45762
rect 85120 45698 85172 45704
rect 52184 42764 52236 42770
rect 52184 42706 52236 42712
rect 141804 40202 141832 46702
rect 194416 44124 194468 44130
rect 194416 44066 194468 44072
rect 194428 42106 194456 44066
rect 194074 42078 194456 42106
rect 187606 41848 187662 41857
rect 187358 41806 187606 41834
rect 187606 41783 187662 41792
rect 141758 40174 141832 40202
rect 141758 39984 141786 40174
rect 207032 17490 207060 51002
rect 212448 45552 212500 45558
rect 212448 45494 212500 45500
rect 212460 41313 212488 45494
rect 209778 41304 209834 41313
rect 209778 41239 209834 41248
rect 212446 41304 212502 41313
rect 212446 41239 212502 41248
rect 209792 17490 209820 41239
rect 213840 24818 213868 51070
rect 216140 48249 216168 52686
rect 281460 48346 281488 52686
rect 346504 52686 346900 52714
rect 412344 52686 412680 52714
rect 477848 52686 478184 52714
rect 346504 51134 346532 52686
rect 346872 52426 346900 52686
rect 346860 52420 346912 52426
rect 346860 52362 346912 52368
rect 346492 51128 346544 51134
rect 346492 51070 346544 51076
rect 412652 48414 412680 52686
rect 478156 48482 478184 52686
rect 543016 52686 543352 52714
rect 478144 48476 478196 48482
rect 478144 48418 478196 48424
rect 526168 48476 526220 48482
rect 526168 48418 526220 48424
rect 412640 48408 412692 48414
rect 412640 48350 412692 48356
rect 506388 48408 506440 48414
rect 506388 48350 506440 48356
rect 218060 48340 218112 48346
rect 218060 48282 218112 48288
rect 281448 48340 281500 48346
rect 281448 48282 281500 48288
rect 502248 48340 502300 48346
rect 502248 48282 502300 48288
rect 216126 48240 216182 48249
rect 216126 48175 216182 48184
rect 218072 46918 218100 48282
rect 218060 46912 218112 46918
rect 218060 46854 218112 46860
rect 215300 42764 215352 42770
rect 215300 42706 215352 42712
rect 213184 24812 213236 24818
rect 213184 24754 213236 24760
rect 213828 24812 213880 24818
rect 213828 24754 213880 24760
rect 213196 17490 213224 24754
rect 207032 17462 207184 17490
rect 209792 17462 210036 17490
rect 212888 17462 213224 17490
rect 215312 17490 215340 42706
rect 218072 33134 218100 46854
rect 460664 46028 460716 46034
rect 460664 45970 460716 45976
rect 367100 45960 367152 45966
rect 367100 45902 367152 45908
rect 311900 45892 311952 45898
rect 311900 45834 311952 45840
rect 230940 45824 230992 45830
rect 230940 45766 230992 45772
rect 230388 45688 230440 45694
rect 230388 45630 230440 45636
rect 226248 43172 226300 43178
rect 226248 43114 226300 43120
rect 223488 43104 223540 43110
rect 223488 43046 223540 43052
rect 218072 33106 218192 33134
rect 218164 17490 218192 33106
rect 223500 22574 223528 43046
rect 226260 23050 226288 43114
rect 224592 23044 224644 23050
rect 224592 22986 224644 22992
rect 226248 23044 226300 23050
rect 226248 22986 226300 22992
rect 221740 22568 221792 22574
rect 221740 22510 221792 22516
rect 223488 22568 223540 22574
rect 223488 22510 223540 22516
rect 221752 17490 221780 22510
rect 224604 17490 224632 22986
rect 215312 17462 215740 17490
rect 218164 17462 218592 17490
rect 221444 17462 221780 17490
rect 224296 17462 224632 17490
rect 230400 10713 230428 45630
rect 230480 43512 230532 43518
rect 230480 43454 230532 43460
rect 230386 10704 230442 10713
rect 230386 10639 230442 10648
rect 230492 7721 230520 43454
rect 230664 43444 230716 43450
rect 230664 43386 230716 43392
rect 230572 43308 230624 43314
rect 230572 43250 230624 43256
rect 230584 9217 230612 43250
rect 230676 13705 230704 43386
rect 230848 43376 230900 43382
rect 230848 43318 230900 43324
rect 230756 43240 230808 43246
rect 230756 43182 230808 43188
rect 230768 15201 230796 43182
rect 230754 15192 230810 15201
rect 230754 15127 230810 15136
rect 230662 13696 230718 13705
rect 230662 13631 230718 13640
rect 230860 12209 230888 43318
rect 230952 16697 230980 45766
rect 233148 45620 233200 45626
rect 233148 45562 233200 45568
rect 230938 16688 230994 16697
rect 230938 16623 230994 16632
rect 230846 12200 230902 12209
rect 230846 12135 230902 12144
rect 230570 9208 230626 9217
rect 230570 9143 230626 9152
rect 230478 7712 230534 7721
rect 230478 7647 230534 7656
rect 233160 6526 233188 45562
rect 311912 43858 311940 45834
rect 367112 43926 367140 45902
rect 365168 43920 365220 43926
rect 365168 43862 365220 43868
rect 367100 43920 367152 43926
rect 367100 43862 367152 43868
rect 310428 43852 310480 43858
rect 310428 43794 310480 43800
rect 311900 43852 311952 43858
rect 311900 43794 311952 43800
rect 307298 43208 307354 43217
rect 307298 43143 307354 43152
rect 307312 42106 307340 43143
rect 310440 42106 310468 43794
rect 365180 42106 365208 43862
rect 416594 43480 416650 43489
rect 416594 43415 416650 43424
rect 415398 43344 415454 43353
rect 415398 43279 415454 43288
rect 415412 42636 415440 43279
rect 307004 42078 307340 42106
rect 310132 42078 310468 42106
rect 364918 42078 365208 42106
rect 416608 42092 416636 43415
rect 460676 42106 460704 45970
rect 475568 45756 475620 45762
rect 475568 45698 475620 45704
rect 470138 43616 470194 43625
rect 470138 43551 470194 43560
rect 470152 42650 470180 43551
rect 470152 42622 470198 42650
rect 475476 42628 475528 42634
rect 475476 42570 475528 42576
rect 460368 42078 460704 42106
rect 405582 41954 405872 41970
rect 405582 41948 405884 41954
rect 405582 41942 405832 41948
rect 405832 41890 405884 41896
rect 426348 41948 426400 41954
rect 426348 41890 426400 41896
rect 361946 41848 362002 41857
rect 361790 41806 361946 41834
rect 419998 41848 420054 41857
rect 419750 41806 419998 41834
rect 361946 41783 362002 41792
rect 419998 41783 420054 41792
rect 426360 41478 426388 41890
rect 427910 41848 427966 41857
rect 471702 41848 471758 41857
rect 471408 41806 471702 41834
rect 427910 41783 427966 41792
rect 471702 41783 471758 41792
rect 426348 41472 426400 41478
rect 426348 41414 426400 41420
rect 427924 41177 427952 41783
rect 427910 41168 427966 41177
rect 427910 41103 427966 41112
rect 475488 41041 475516 42570
rect 475474 41032 475530 41041
rect 475474 40967 475530 40976
rect 475580 38622 475608 45698
rect 502260 41290 502288 48282
rect 506400 41410 506428 48350
rect 521750 42120 521806 42129
rect 521806 42078 521870 42106
rect 526180 42092 526208 48418
rect 543016 42770 543044 52686
rect 571800 48408 571852 48414
rect 571800 48350 571852 48356
rect 549260 48340 549312 48346
rect 549260 48282 549312 48288
rect 529664 42764 529716 42770
rect 529664 42706 529716 42712
rect 543004 42764 543056 42770
rect 543004 42706 543056 42712
rect 529676 42106 529704 42706
rect 529322 42078 529704 42106
rect 521750 42055 521806 42064
rect 513932 42016 513984 42022
rect 520372 42016 520424 42022
rect 513932 41958 513984 41964
rect 513286 41848 513342 41857
rect 513286 41783 513342 41792
rect 513300 41410 513328 41783
rect 506388 41404 506440 41410
rect 506388 41346 506440 41352
rect 513288 41404 513340 41410
rect 513288 41346 513340 41352
rect 502260 41262 502380 41290
rect 475568 38616 475620 38622
rect 475568 38558 475620 38564
rect 502352 38554 502380 41262
rect 513944 38554 513972 41958
rect 514864 41954 515154 41970
rect 520424 41964 520674 41970
rect 520372 41958 520674 41964
rect 514024 41948 514076 41954
rect 514024 41890 514076 41896
rect 514852 41948 515154 41954
rect 514904 41942 515154 41948
rect 520384 41942 520674 41958
rect 514852 41890 514904 41896
rect 514036 38622 514064 41890
rect 518530 41848 518586 41857
rect 518586 41806 518830 41834
rect 518530 41783 518586 41792
rect 530400 41404 530452 41410
rect 530400 41346 530452 41352
rect 530308 41336 530360 41342
rect 530306 41304 530308 41313
rect 530360 41304 530362 41313
rect 530306 41239 530362 41248
rect 530412 41177 530440 41346
rect 530398 41168 530454 41177
rect 530398 41103 530454 41112
rect 549272 41041 549300 48282
rect 568580 47252 568632 47258
rect 568580 47194 568632 47200
rect 568592 41449 568620 47194
rect 568578 41440 568634 41449
rect 568578 41375 568634 41384
rect 571812 41342 571840 48350
rect 575676 43217 575704 95202
rect 580552 94761 580580 126958
rect 580644 99385 580672 129814
rect 580724 127084 580776 127090
rect 580724 127026 580776 127032
rect 580630 99376 580686 99385
rect 580630 99311 580686 99320
rect 580736 96257 580764 127026
rect 580816 124228 580868 124234
rect 580816 124170 580868 124176
rect 580722 96248 580778 96257
rect 580722 96183 580778 96192
rect 580538 94752 580594 94761
rect 580538 94687 580594 94696
rect 580828 91769 580856 124170
rect 580920 102377 580948 132602
rect 581012 117609 581040 140830
rect 581184 140820 581236 140826
rect 581184 140762 581236 140768
rect 581092 138168 581144 138174
rect 581092 138110 581144 138116
rect 580998 117600 581054 117609
rect 580998 117535 581054 117544
rect 581000 110492 581052 110498
rect 581000 110434 581052 110440
rect 580906 102368 580962 102377
rect 580906 102303 580962 102312
rect 580908 99408 580960 99414
rect 580908 99350 580960 99356
rect 580814 91760 580870 91769
rect 580814 91695 580870 91704
rect 580724 84244 580776 84250
rect 580724 84186 580776 84192
rect 579620 82680 579672 82686
rect 579618 82648 579620 82657
rect 579672 82648 579674 82657
rect 579618 82583 579674 82592
rect 575848 78668 575900 78674
rect 575848 78610 575900 78616
rect 575756 74996 575808 75002
rect 575756 74938 575808 74944
rect 575768 47258 575796 74938
rect 575756 47252 575808 47258
rect 575756 47194 575808 47200
rect 575860 43625 575888 78610
rect 580736 68921 580764 84186
rect 580816 84176 580868 84182
rect 580816 84118 580868 84124
rect 580722 68912 580778 68921
rect 580722 68847 580778 68856
rect 579620 66224 579672 66230
rect 579620 66166 579672 66172
rect 579632 65929 579660 66166
rect 579618 65920 579674 65929
rect 579618 65855 579674 65864
rect 580828 62937 580856 84118
rect 580814 62928 580870 62937
rect 580814 62863 580870 62872
rect 580920 53825 580948 99350
rect 581012 70417 581040 110434
rect 581104 109993 581132 138110
rect 581196 114481 581224 140762
rect 581288 120601 581316 143550
rect 581380 126721 581408 149058
rect 581460 146328 581512 146334
rect 581460 146270 581512 146276
rect 581366 126712 581422 126721
rect 581366 126647 581422 126656
rect 581472 123593 581500 146270
rect 581564 125089 581592 149126
rect 581656 144945 581684 160142
rect 581736 160132 581788 160138
rect 581736 160074 581788 160080
rect 581748 146441 581776 160074
rect 582024 160041 582052 168346
rect 600412 168302 600464 168308
rect 599490 167784 599546 167793
rect 599490 167719 599546 167728
rect 582288 165776 582340 165782
rect 582288 165718 582340 165724
rect 582196 165708 582248 165714
rect 582196 165650 582248 165656
rect 582104 160268 582156 160274
rect 582104 160210 582156 160216
rect 582010 160032 582066 160041
rect 582010 159967 582066 159976
rect 581828 151904 581880 151910
rect 581828 151846 581880 151852
rect 581734 146432 581790 146441
rect 581734 146367 581790 146376
rect 581642 144936 581698 144945
rect 581642 144871 581698 144880
rect 581736 143676 581788 143682
rect 581736 143618 581788 143624
rect 581644 140956 581696 140962
rect 581644 140898 581696 140904
rect 581550 125080 581606 125089
rect 581550 125015 581606 125024
rect 581458 123584 581514 123593
rect 581458 123519 581514 123528
rect 581274 120592 581330 120601
rect 581274 120527 581330 120536
rect 581460 118720 581512 118726
rect 581460 118662 581512 118668
rect 581276 116000 581328 116006
rect 581276 115942 581328 115948
rect 581182 114472 581238 114481
rect 581182 114407 581238 114416
rect 581090 109984 581146 109993
rect 581090 109919 581146 109928
rect 581184 107704 581236 107710
rect 581184 107646 581236 107652
rect 581092 104916 581144 104922
rect 581092 104858 581144 104864
rect 580998 70408 581054 70417
rect 580998 70343 581054 70352
rect 581104 64433 581132 104858
rect 581196 67425 581224 107646
rect 581288 79529 581316 115942
rect 581368 113212 581420 113218
rect 581368 113154 581420 113160
rect 581274 79520 581330 79529
rect 581274 79455 581330 79464
rect 581380 76537 581408 113154
rect 581472 81161 581500 118662
rect 581656 115977 581684 140898
rect 581748 119105 581776 143618
rect 581840 131209 581868 151846
rect 582012 149252 582064 149258
rect 582012 149194 582064 149200
rect 581920 143744 581972 143750
rect 581920 143686 581972 143692
rect 581826 131200 581882 131209
rect 581826 131135 581882 131144
rect 581828 124296 581880 124302
rect 581828 124238 581880 124244
rect 581734 119096 581790 119105
rect 581734 119031 581790 119040
rect 581736 116068 581788 116074
rect 581736 116010 581788 116016
rect 581642 115968 581698 115977
rect 581642 115903 581698 115912
rect 581644 113280 581696 113286
rect 581644 113222 581696 113228
rect 581552 110560 581604 110566
rect 581552 110502 581604 110508
rect 581458 81152 581514 81161
rect 581458 81087 581514 81096
rect 581366 76528 581422 76537
rect 581366 76463 581422 76472
rect 581564 72049 581592 110502
rect 581656 75041 581684 113222
rect 581748 78033 581776 116010
rect 581840 90273 581868 124238
rect 581932 122097 581960 143686
rect 582024 129713 582052 149194
rect 582116 140321 582144 160210
rect 582208 150929 582236 165650
rect 582300 152425 582328 165718
rect 599504 165646 599532 167719
rect 600042 166696 600098 166705
rect 600042 166631 600098 166640
rect 600056 165782 600084 166631
rect 600044 165776 600096 165782
rect 599950 165744 600006 165753
rect 600044 165718 600096 165724
rect 599950 165679 599952 165688
rect 600004 165679 600006 165688
rect 599952 165650 600004 165656
rect 599492 165640 599544 165646
rect 599492 165582 599544 165588
rect 601344 165578 601372 173839
rect 666558 173632 666614 173641
rect 666558 173567 666614 173576
rect 666572 170241 666600 173567
rect 666558 170232 666614 170241
rect 666664 170202 666692 278734
rect 666756 177970 666784 284650
rect 666848 216730 666876 287234
rect 667032 226334 667060 289070
rect 670240 287088 670292 287094
rect 670240 287030 670292 287036
rect 669964 283212 670016 283218
rect 669964 283154 670016 283160
rect 667032 226306 667152 226334
rect 666848 216702 667060 216730
rect 666836 216572 666888 216578
rect 666836 216514 666888 216520
rect 666848 178090 666876 216514
rect 666928 213308 666980 213314
rect 666928 213250 666980 213256
rect 666836 178084 666888 178090
rect 666836 178026 666888 178032
rect 666756 177942 666876 177970
rect 666744 177880 666796 177886
rect 666744 177822 666796 177828
rect 666558 170167 666614 170176
rect 666652 170196 666704 170202
rect 666652 170138 666704 170144
rect 666756 170082 666784 177822
rect 666572 170054 666784 170082
rect 601332 165572 601384 165578
rect 601332 165514 601384 165520
rect 600042 164656 600098 164665
rect 600042 164591 600098 164600
rect 599950 163704 600006 163713
rect 599950 163639 600006 163648
rect 599964 162926 599992 163639
rect 600056 162994 600084 164591
rect 600044 162988 600096 162994
rect 600044 162930 600096 162936
rect 599952 162920 600004 162926
rect 599952 162862 600004 162868
rect 600042 162616 600098 162625
rect 600042 162551 600098 162560
rect 599858 161664 599914 161673
rect 599858 161599 599914 161608
rect 599872 160206 599900 161599
rect 599950 160576 600006 160585
rect 599950 160511 600006 160520
rect 599964 160274 599992 160511
rect 599952 160268 600004 160274
rect 599952 160210 600004 160216
rect 599860 160200 599912 160206
rect 599860 160142 599912 160148
rect 600056 160138 600084 162551
rect 600044 160132 600096 160138
rect 600044 160074 600096 160080
rect 599858 159624 599914 159633
rect 599858 159559 599914 159568
rect 599872 157554 599900 159559
rect 600042 158536 600098 158545
rect 600042 158471 600098 158480
rect 599950 157584 600006 157593
rect 599860 157548 599912 157554
rect 599950 157519 600006 157528
rect 599860 157490 599912 157496
rect 599964 157486 599992 157519
rect 599952 157480 600004 157486
rect 599952 157422 600004 157428
rect 600056 157418 600084 158471
rect 600044 157412 600096 157418
rect 600044 157354 600096 157360
rect 599858 156496 599914 156505
rect 599858 156431 599914 156440
rect 599872 154630 599900 156431
rect 599950 155544 600006 155553
rect 599950 155479 600006 155488
rect 599964 154698 599992 155479
rect 599952 154692 600004 154698
rect 599952 154634 600004 154640
rect 599860 154624 599912 154630
rect 599860 154566 599912 154572
rect 599858 154456 599914 154465
rect 599858 154391 599914 154400
rect 582286 152416 582342 152425
rect 582286 152351 582342 152360
rect 599872 151978 599900 154391
rect 600042 153504 600098 153513
rect 600042 153439 600098 153448
rect 599950 152416 600006 152425
rect 599950 152351 600006 152360
rect 582288 151972 582340 151978
rect 582288 151914 582340 151920
rect 599860 151972 599912 151978
rect 599860 151914 599912 151920
rect 582194 150920 582250 150929
rect 582194 150855 582250 150864
rect 582196 146396 582248 146402
rect 582196 146338 582248 146344
rect 582102 140312 582158 140321
rect 582102 140247 582158 140256
rect 582010 129704 582066 129713
rect 582010 129639 582066 129648
rect 582208 128217 582236 146338
rect 582300 134201 582328 151914
rect 599964 151910 599992 152351
rect 599952 151904 600004 151910
rect 599952 151846 600004 151852
rect 600056 151842 600084 153439
rect 600044 151836 600096 151842
rect 600044 151778 600096 151784
rect 600042 151464 600098 151473
rect 600042 151399 600098 151408
rect 599858 150376 599914 150385
rect 599858 150311 599914 150320
rect 599872 149190 599900 150311
rect 599950 149424 600006 149433
rect 599950 149359 600006 149368
rect 599860 149184 599912 149190
rect 599860 149126 599912 149132
rect 599964 149122 599992 149359
rect 600056 149258 600084 151399
rect 600044 149252 600096 149258
rect 600044 149194 600096 149200
rect 599952 149116 600004 149122
rect 599952 149058 600004 149064
rect 599858 148336 599914 148345
rect 599858 148271 599914 148280
rect 599872 146402 599900 148271
rect 599950 147384 600006 147393
rect 599950 147319 600006 147328
rect 599860 146396 599912 146402
rect 599860 146338 599912 146344
rect 599964 146334 599992 147319
rect 599952 146328 600004 146334
rect 599858 146296 599914 146305
rect 599952 146270 600004 146276
rect 599858 146231 599914 146240
rect 599872 143750 599900 146231
rect 600042 145344 600098 145353
rect 600042 145279 600098 145288
rect 599950 144256 600006 144265
rect 599950 144191 600006 144200
rect 599860 143744 599912 143750
rect 599860 143686 599912 143692
rect 599964 143682 599992 144191
rect 599952 143676 600004 143682
rect 599952 143618 600004 143624
rect 600056 143614 600084 145279
rect 600044 143608 600096 143614
rect 600044 143550 600096 143556
rect 600042 143304 600098 143313
rect 600042 143239 600098 143248
rect 599950 142216 600006 142225
rect 599950 142151 600006 142160
rect 599858 141264 599914 141273
rect 599858 141199 599914 141208
rect 599872 140826 599900 141199
rect 599964 140962 599992 142151
rect 599952 140956 600004 140962
rect 599952 140898 600004 140904
rect 600056 140894 600084 143239
rect 600044 140888 600096 140894
rect 600044 140830 600096 140836
rect 599860 140820 599912 140826
rect 599860 140762 599912 140768
rect 600042 140176 600098 140185
rect 600042 140111 600098 140120
rect 599858 139224 599914 139233
rect 599858 139159 599914 139168
rect 599872 138038 599900 139159
rect 599952 138168 600004 138174
rect 599950 138136 599952 138145
rect 600004 138136 600006 138145
rect 600056 138106 600084 140111
rect 599950 138071 600006 138080
rect 600044 138100 600096 138106
rect 600044 138042 600096 138048
rect 599860 138032 599912 138038
rect 599860 137974 599912 137980
rect 599858 137184 599914 137193
rect 599858 137119 599914 137128
rect 599872 135386 599900 137119
rect 599950 136096 600006 136105
rect 599950 136031 600006 136040
rect 599860 135380 599912 135386
rect 599860 135322 599912 135328
rect 599964 135318 599992 136031
rect 599952 135312 600004 135318
rect 599952 135254 600004 135260
rect 600042 135144 600098 135153
rect 600042 135079 600098 135088
rect 582286 134192 582342 134201
rect 582286 134127 582342 134136
rect 599858 134056 599914 134065
rect 599858 133991 599914 134000
rect 599872 132598 599900 133991
rect 599950 133104 600006 133113
rect 599950 133039 600006 133048
rect 599964 132666 599992 133039
rect 599952 132660 600004 132666
rect 599952 132602 600004 132608
rect 599860 132592 599912 132598
rect 599860 132534 599912 132540
rect 600056 132530 600084 135079
rect 600044 132524 600096 132530
rect 600044 132466 600096 132472
rect 600042 132016 600098 132025
rect 600042 131951 600098 131960
rect 599858 131064 599914 131073
rect 599858 130999 599914 131008
rect 599872 129878 599900 130999
rect 599950 129976 600006 129985
rect 600056 129946 600084 131951
rect 599950 129911 600006 129920
rect 600044 129940 600096 129946
rect 599860 129872 599912 129878
rect 599860 129814 599912 129820
rect 599964 129810 599992 129911
rect 600044 129882 600096 129888
rect 599952 129804 600004 129810
rect 599952 129746 600004 129752
rect 599858 129024 599914 129033
rect 599858 128959 599914 128968
rect 582194 128208 582250 128217
rect 582194 128143 582250 128152
rect 599872 127090 599900 128959
rect 599950 127936 600006 127945
rect 599950 127871 600006 127880
rect 599860 127084 599912 127090
rect 599860 127026 599912 127032
rect 599964 127022 599992 127871
rect 599952 127016 600004 127022
rect 599858 126984 599914 126993
rect 599952 126958 600004 126964
rect 599858 126919 599914 126928
rect 599766 124944 599822 124953
rect 599766 124879 599822 124888
rect 582288 124364 582340 124370
rect 582288 124306 582340 124312
rect 581918 122088 581974 122097
rect 581918 122023 581974 122032
rect 582196 121644 582248 121650
rect 582196 121586 582248 121592
rect 582012 121576 582064 121582
rect 582012 121518 582064 121524
rect 581920 118788 581972 118794
rect 581920 118730 581972 118736
rect 581826 90264 581882 90273
rect 581826 90199 581882 90208
rect 581828 84448 581880 84454
rect 581828 84390 581880 84396
rect 581734 78024 581790 78033
rect 581734 77959 581790 77968
rect 581642 75032 581698 75041
rect 581642 74967 581698 74976
rect 581550 72040 581606 72049
rect 581550 71975 581606 71984
rect 581182 67416 581238 67425
rect 581182 67351 581238 67360
rect 581090 64424 581146 64433
rect 581090 64359 581146 64368
rect 581840 56817 581868 84390
rect 581932 84153 581960 118730
rect 582024 87145 582052 121518
rect 582104 121508 582156 121514
rect 582104 121450 582156 121456
rect 582116 88641 582144 121450
rect 582102 88632 582158 88641
rect 582102 88567 582158 88576
rect 582010 87136 582066 87145
rect 582010 87071 582066 87080
rect 582208 85649 582236 121586
rect 582300 93265 582328 124306
rect 599780 124302 599808 124879
rect 599872 124370 599900 126919
rect 599950 125896 600006 125905
rect 599950 125831 600006 125840
rect 599860 124364 599912 124370
rect 599860 124306 599912 124312
rect 599768 124296 599820 124302
rect 599768 124238 599820 124244
rect 599964 124234 599992 125831
rect 599952 124228 600004 124234
rect 599952 124170 600004 124176
rect 600042 123856 600098 123865
rect 600042 123791 600098 123800
rect 599858 122904 599914 122913
rect 599858 122839 599914 122848
rect 599872 121582 599900 122839
rect 599950 121816 600006 121825
rect 599950 121751 600006 121760
rect 599964 121650 599992 121751
rect 599952 121644 600004 121650
rect 599952 121586 600004 121592
rect 599860 121576 599912 121582
rect 599860 121518 599912 121524
rect 600056 121514 600084 123791
rect 600044 121508 600096 121514
rect 600044 121450 600096 121456
rect 600042 120864 600098 120873
rect 600042 120799 600098 120808
rect 599950 119776 600006 119785
rect 599950 119711 600006 119720
rect 599964 118862 599992 119711
rect 583668 118856 583720 118862
rect 599952 118856 600004 118862
rect 583668 118798 583720 118804
rect 599858 118824 599914 118833
rect 582286 93256 582342 93265
rect 582286 93191 582342 93200
rect 582194 85640 582250 85649
rect 582194 85575 582250 85584
rect 582196 84584 582248 84590
rect 582196 84526 582248 84532
rect 582012 84380 582064 84386
rect 582012 84322 582064 84328
rect 581918 84144 581974 84153
rect 581918 84079 581974 84088
rect 581826 56808 581882 56817
rect 581826 56743 581882 56752
rect 582024 55321 582052 84322
rect 582104 84312 582156 84318
rect 582104 84254 582156 84260
rect 582116 59809 582144 84254
rect 582208 61305 582236 84526
rect 582288 84516 582340 84522
rect 582288 84458 582340 84464
rect 582194 61296 582250 61305
rect 582194 61231 582250 61240
rect 582102 59800 582158 59809
rect 582102 59735 582158 59744
rect 582300 58313 582328 84458
rect 583680 82686 583708 118798
rect 599952 118798 600004 118804
rect 600056 118794 600084 120799
rect 599858 118759 599914 118768
rect 600044 118788 600096 118794
rect 599872 118726 599900 118759
rect 600044 118730 600096 118736
rect 599860 118720 599912 118726
rect 599860 118662 599912 118668
rect 600042 117736 600098 117745
rect 600042 117671 600098 117680
rect 599950 116784 600006 116793
rect 599950 116719 600006 116728
rect 599964 116074 599992 116719
rect 599952 116068 600004 116074
rect 599952 116010 600004 116016
rect 600056 116006 600084 117671
rect 600044 116000 600096 116006
rect 600044 115942 600096 115948
rect 599858 115696 599914 115705
rect 599858 115631 599914 115640
rect 599872 113218 599900 115631
rect 599950 114744 600006 114753
rect 599950 114679 600006 114688
rect 599964 113286 599992 114679
rect 599952 113280 600004 113286
rect 599952 113222 600004 113228
rect 599860 113212 599912 113218
rect 599860 113154 599912 113160
rect 599858 112704 599914 112713
rect 599858 112639 599914 112648
rect 599872 110566 599900 112639
rect 599950 111616 600006 111625
rect 599950 111551 600006 111560
rect 599860 110560 599912 110566
rect 599860 110502 599912 110508
rect 599964 110498 599992 111551
rect 600226 110664 600282 110673
rect 600226 110599 600282 110608
rect 599952 110492 600004 110498
rect 599952 110434 600004 110440
rect 599306 109576 599362 109585
rect 599306 109511 599362 109520
rect 599320 107710 599348 109511
rect 599308 107704 599360 107710
rect 599308 107646 599360 107652
rect 599950 107536 600006 107545
rect 599950 107471 600006 107480
rect 599964 104922 599992 107471
rect 599952 104916 600004 104922
rect 599952 104858 600004 104864
rect 599950 100464 600006 100473
rect 599950 100399 600006 100408
rect 599964 99414 599992 100399
rect 599952 99408 600004 99414
rect 599952 99350 600004 99356
rect 591948 95396 592000 95402
rect 591948 95338 592000 95344
rect 589188 95328 589240 95334
rect 589188 95270 589240 95276
rect 583760 84652 583812 84658
rect 583760 84594 583812 84600
rect 583668 82680 583720 82686
rect 583668 82622 583720 82628
rect 583668 73160 583720 73166
rect 583668 73102 583720 73108
rect 582286 58304 582342 58313
rect 582286 58239 582342 58248
rect 582010 55312 582066 55321
rect 582010 55247 582066 55256
rect 580906 53816 580962 53825
rect 580906 53751 580962 53760
rect 581644 53236 581696 53242
rect 581644 53178 581696 53184
rect 581656 48414 581684 53178
rect 581644 48408 581696 48414
rect 581644 48350 581696 48356
rect 583680 47122 583708 73102
rect 583772 66230 583800 84594
rect 589200 75002 589228 95270
rect 589188 74996 589240 75002
rect 589188 74938 589240 74944
rect 591960 72690 591988 95338
rect 600240 84250 600268 110599
rect 600318 108624 600374 108633
rect 600318 108559 600374 108568
rect 600332 84658 600360 108559
rect 600594 106584 600650 106593
rect 600594 106519 600650 106528
rect 600410 105496 600466 105505
rect 600410 105431 600466 105440
rect 600320 84652 600372 84658
rect 600320 84594 600372 84600
rect 600424 84590 600452 105431
rect 600502 102504 600558 102513
rect 600502 102439 600558 102448
rect 600412 84584 600464 84590
rect 600412 84526 600464 84532
rect 600516 84454 600544 102439
rect 600504 84448 600556 84454
rect 600504 84390 600556 84396
rect 600228 84244 600280 84250
rect 600228 84186 600280 84192
rect 600608 84182 600636 106519
rect 600870 104544 600926 104553
rect 600870 104479 600926 104488
rect 600686 103456 600742 103465
rect 600686 103391 600742 103400
rect 600700 84522 600728 103391
rect 600778 101416 600834 101425
rect 600778 101351 600834 101360
rect 600688 84516 600740 84522
rect 600688 84458 600740 84464
rect 600792 84386 600820 101351
rect 600780 84380 600832 84386
rect 600780 84322 600832 84328
rect 600884 84318 600912 104479
rect 606404 100014 606740 100042
rect 606404 95606 606432 100014
rect 607370 99770 607398 100028
rect 607324 99742 607398 99770
rect 607692 100014 608028 100042
rect 608152 100014 608672 100042
rect 608980 100014 609316 100042
rect 609960 100014 610204 100042
rect 604460 95600 604512 95606
rect 604460 95542 604512 95548
rect 606392 95600 606444 95606
rect 606392 95542 606444 95548
rect 600872 84312 600924 84318
rect 600872 84254 600924 84260
rect 600596 84176 600648 84182
rect 600596 84118 600648 84124
rect 596916 83156 596968 83162
rect 596916 83098 596968 83104
rect 596928 78674 596956 83098
rect 604472 82890 604500 95542
rect 607220 93900 607272 93906
rect 607220 93842 607272 93848
rect 607232 83162 607260 93842
rect 607220 83156 607272 83162
rect 607220 83098 607272 83104
rect 597468 82884 597520 82890
rect 597468 82826 597520 82832
rect 604460 82884 604512 82890
rect 604460 82826 604512 82832
rect 596916 78668 596968 78674
rect 596916 78610 596968 78616
rect 586428 72684 586480 72690
rect 586428 72626 586480 72632
rect 591948 72684 592000 72690
rect 591948 72626 592000 72632
rect 583760 66224 583812 66230
rect 583760 66166 583812 66172
rect 577964 47116 578016 47122
rect 577964 47058 578016 47064
rect 583668 47116 583720 47122
rect 583668 47058 583720 47064
rect 575846 43616 575902 43625
rect 575846 43551 575902 43560
rect 577976 43489 578004 47058
rect 577962 43480 578018 43489
rect 577962 43415 578018 43424
rect 586440 43353 586468 72626
rect 594708 66292 594760 66298
rect 594708 66234 594760 66240
rect 587900 62348 587952 62354
rect 587900 62290 587952 62296
rect 587912 53242 587940 62290
rect 587900 53236 587952 53242
rect 587900 53178 587952 53184
rect 594720 48346 594748 66234
rect 597480 62354 597508 82826
rect 600228 80164 600280 80170
rect 600228 80106 600280 80112
rect 600240 66298 600268 80106
rect 600228 66292 600280 66298
rect 600228 66234 600280 66240
rect 602988 66292 603040 66298
rect 602988 66234 603040 66240
rect 597468 62348 597520 62354
rect 597468 62290 597520 62296
rect 594708 48340 594760 48346
rect 594708 48282 594760 48288
rect 586426 43344 586482 43353
rect 586426 43279 586482 43288
rect 575662 43208 575718 43217
rect 575662 43143 575718 43152
rect 603000 41410 603028 66234
rect 607324 45966 607352 99742
rect 607496 95600 607548 95606
rect 607496 95542 607548 95548
rect 607312 45960 607364 45966
rect 607312 45902 607364 45908
rect 607508 41478 607536 95542
rect 607692 95266 607720 100014
rect 607680 95260 607732 95266
rect 607680 95202 607732 95208
rect 608152 91094 608180 100014
rect 608980 95606 609008 100014
rect 608968 95600 609020 95606
rect 608968 95542 609020 95548
rect 607600 91066 608180 91094
rect 607600 45898 607628 91066
rect 610176 73166 610204 100014
rect 610360 100014 610604 100042
rect 610728 100014 611248 100042
rect 611556 100014 611892 100042
rect 612200 100014 612536 100042
rect 612936 100014 613180 100042
rect 613304 100014 613916 100042
rect 614560 100014 614804 100042
rect 610256 95600 610308 95606
rect 610256 95542 610308 95548
rect 610164 73160 610216 73166
rect 610164 73102 610216 73108
rect 610268 46034 610296 95542
rect 610360 95402 610388 100014
rect 610348 95396 610400 95402
rect 610348 95338 610400 95344
rect 610728 91094 610756 100014
rect 611556 95606 611584 100014
rect 611544 95600 611596 95606
rect 611544 95542 611596 95548
rect 612200 95334 612228 100014
rect 612188 95328 612240 95334
rect 612188 95270 612240 95276
rect 612936 93906 612964 100014
rect 613304 94602 613332 100014
rect 614776 95810 614804 100014
rect 614868 100014 615204 100042
rect 615848 100014 616184 100042
rect 616492 100014 616828 100042
rect 617136 100014 617472 100042
rect 617780 100014 618116 100042
rect 618424 100014 618760 100042
rect 619068 100014 619404 100042
rect 619712 100014 620048 100042
rect 614764 95804 614816 95810
rect 614764 95746 614816 95752
rect 613028 94574 613332 94602
rect 612924 93900 612976 93906
rect 612924 93842 612976 93848
rect 613028 93786 613056 94574
rect 610360 91066 610756 91094
rect 612844 93758 613056 93786
rect 610360 66298 610388 91066
rect 612844 80170 612872 93758
rect 614868 93702 614896 100014
rect 616156 95742 616184 100014
rect 616144 95736 616196 95742
rect 616144 95678 616196 95684
rect 616800 94926 616828 100014
rect 617444 95402 617472 100014
rect 617432 95396 617484 95402
rect 617432 95338 617484 95344
rect 616788 94920 616840 94926
rect 616788 94862 616840 94868
rect 618088 94178 618116 100014
rect 618260 95600 618312 95606
rect 618260 95542 618312 95548
rect 618076 94172 618128 94178
rect 618076 94114 618128 94120
rect 613016 93696 613068 93702
rect 613016 93638 613068 93644
rect 614856 93696 614908 93702
rect 614856 93638 614908 93644
rect 612832 80164 612884 80170
rect 612832 80106 612884 80112
rect 610348 66292 610400 66298
rect 610348 66234 610400 66240
rect 610256 46028 610308 46034
rect 610256 45970 610308 45976
rect 607588 45892 607640 45898
rect 607588 45834 607640 45840
rect 613028 45830 613056 93638
rect 613016 45824 613068 45830
rect 613016 45766 613068 45772
rect 618272 43518 618300 95542
rect 618732 94790 618760 100014
rect 619376 95130 619404 100014
rect 620020 95470 620048 100014
rect 620112 100014 620448 100042
rect 621092 100014 621152 100042
rect 620112 95606 620140 100014
rect 620100 95600 620152 95606
rect 620100 95542 620152 95548
rect 620008 95464 620060 95470
rect 620008 95406 620060 95412
rect 619364 95124 619416 95130
rect 619364 95066 619416 95072
rect 618720 94784 618772 94790
rect 618720 94726 618772 94732
rect 618260 43512 618312 43518
rect 618260 43454 618312 43460
rect 621124 43314 621152 100014
rect 621400 100014 621736 100042
rect 622044 100014 622380 100042
rect 622688 100014 623024 100042
rect 623332 100014 623668 100042
rect 623792 100014 624312 100042
rect 624620 100014 624956 100042
rect 625600 100014 625936 100042
rect 626244 100014 626488 100042
rect 626980 100014 627316 100042
rect 627624 100014 627960 100042
rect 628268 100014 628328 100042
rect 621296 95668 621348 95674
rect 621296 95610 621348 95616
rect 621204 95532 621256 95538
rect 621204 95474 621256 95480
rect 621216 43382 621244 95474
rect 621204 43376 621256 43382
rect 621204 43318 621256 43324
rect 621112 43308 621164 43314
rect 621112 43250 621164 43256
rect 621308 43246 621336 95610
rect 621400 45694 621428 100014
rect 621480 95600 621532 95606
rect 621480 95542 621532 95548
rect 621388 45688 621440 45694
rect 621388 45630 621440 45636
rect 621492 43450 621520 95542
rect 622044 95538 622072 100014
rect 622492 95736 622544 95742
rect 622492 95678 622544 95684
rect 622032 95532 622084 95538
rect 622032 95474 622084 95480
rect 622124 95396 622176 95402
rect 622124 95338 622176 95344
rect 622136 83201 622164 95338
rect 622504 87961 622532 95678
rect 622688 95606 622716 100014
rect 623332 95674 623360 100014
rect 623320 95668 623372 95674
rect 623320 95610 623372 95616
rect 622676 95600 622728 95606
rect 622676 95542 622728 95548
rect 623412 95464 623464 95470
rect 623412 95406 623464 95412
rect 623228 94920 623280 94926
rect 623228 94862 623280 94868
rect 623136 94172 623188 94178
rect 623136 94114 623188 94120
rect 622490 87952 622546 87961
rect 622490 87887 622546 87896
rect 623148 84153 623176 94114
rect 623240 88913 623268 94862
rect 623320 94784 623372 94790
rect 623320 94726 623372 94732
rect 623226 88904 623282 88913
rect 623226 88839 623282 88848
rect 623332 85105 623360 94726
rect 623424 87009 623452 95406
rect 623504 95124 623556 95130
rect 623504 95066 623556 95072
rect 623410 87000 623466 87009
rect 623410 86935 623466 86944
rect 623516 86057 623544 95066
rect 623792 89729 623820 100014
rect 624620 91094 624648 100014
rect 625908 91633 625936 100014
rect 626460 92585 626488 100014
rect 627288 93537 627316 100014
rect 627932 94489 627960 100014
rect 628300 95985 628328 100014
rect 628760 100014 628912 100042
rect 629556 100014 629708 100042
rect 630200 100014 630628 100042
rect 630844 100014 631180 100042
rect 631488 100014 631824 100042
rect 632132 100014 632468 100042
rect 632776 100014 633112 100042
rect 633512 100014 633848 100042
rect 634156 100014 634492 100042
rect 634800 100014 635136 100042
rect 635444 100014 635780 100042
rect 636088 100014 636332 100042
rect 636732 100014 637068 100042
rect 637376 100014 637528 100042
rect 638020 100014 638356 100042
rect 638664 100014 638908 100042
rect 639308 100014 639644 100042
rect 639952 100014 640104 100042
rect 640688 100014 640932 100042
rect 641332 100014 641668 100042
rect 641976 100014 642312 100042
rect 642620 100014 642680 100042
rect 643264 100014 643600 100042
rect 643908 100014 644244 100042
rect 644552 100014 644796 100042
rect 628286 95976 628342 95985
rect 628286 95911 628342 95920
rect 628760 95826 628788 100014
rect 628728 95798 628788 95826
rect 629680 95826 629708 100014
rect 630600 95826 630628 100014
rect 631152 96082 631180 100014
rect 631140 96076 631192 96082
rect 631140 96018 631192 96024
rect 631796 95946 631824 100014
rect 632440 96082 632468 100014
rect 633084 96626 633112 100014
rect 633072 96620 633124 96626
rect 633072 96562 633124 96568
rect 633820 96558 633848 100014
rect 633808 96552 633860 96558
rect 633808 96494 633860 96500
rect 634464 96490 634492 100014
rect 634452 96484 634504 96490
rect 634452 96426 634504 96432
rect 635108 96082 635136 100014
rect 635280 96620 635332 96626
rect 635280 96562 635332 96568
rect 632106 96076 632158 96082
rect 632106 96018 632158 96024
rect 632428 96076 632480 96082
rect 632428 96018 632480 96024
rect 634406 96076 634458 96082
rect 634406 96018 634458 96024
rect 635096 96076 635148 96082
rect 635096 96018 635148 96024
rect 631784 95940 631836 95946
rect 631784 95882 631836 95888
rect 629680 95798 629832 95826
rect 630600 95798 631028 95826
rect 632118 95812 632146 96018
rect 632980 95940 633032 95946
rect 632980 95882 633032 95888
rect 632992 95826 633020 95882
rect 632992 95798 633328 95826
rect 634418 95812 634446 96018
rect 635292 95826 635320 96562
rect 635752 96422 635780 100014
rect 636304 96626 636332 100014
rect 636292 96620 636344 96626
rect 636292 96562 636344 96568
rect 637040 96558 637068 100014
rect 636384 96552 636436 96558
rect 636384 96494 636436 96500
rect 637028 96552 637080 96558
rect 637028 96494 637080 96500
rect 635740 96416 635792 96422
rect 635740 96358 635792 96364
rect 636396 95826 636424 96494
rect 635292 95798 635628 95826
rect 636396 95798 636732 95826
rect 637500 95742 637528 100014
rect 637580 96484 637632 96490
rect 637580 96426 637632 96432
rect 637592 95826 637620 96426
rect 637592 95798 637928 95826
rect 637488 95736 637540 95742
rect 637488 95678 637540 95684
rect 638328 95606 638356 100014
rect 638880 95878 638908 100014
rect 639006 96076 639058 96082
rect 639006 96018 639058 96024
rect 638868 95872 638920 95878
rect 638868 95814 638920 95820
rect 639018 95812 639046 96018
rect 639616 95810 639644 100014
rect 639880 96416 639932 96422
rect 639880 96358 639932 96364
rect 639892 95826 639920 96358
rect 640076 95946 640104 100014
rect 640064 95940 640116 95946
rect 640064 95882 640116 95888
rect 639604 95804 639656 95810
rect 639892 95798 640228 95826
rect 639604 95746 639656 95752
rect 640904 95742 640932 100014
rect 640984 96620 641036 96626
rect 640984 96562 641036 96568
rect 640996 95826 641024 96562
rect 640996 95798 641332 95826
rect 640524 95736 640576 95742
rect 640522 95704 640524 95713
rect 640892 95736 640944 95742
rect 640576 95704 640578 95713
rect 640892 95678 640944 95684
rect 641640 95674 641668 100014
rect 640522 95639 640578 95648
rect 641628 95668 641680 95674
rect 641628 95610 641680 95616
rect 642284 95606 642312 100014
rect 642364 96552 642416 96558
rect 642364 96494 642416 96500
rect 642376 95826 642404 96494
rect 642376 95798 642528 95826
rect 638316 95600 638368 95606
rect 638316 95542 638368 95548
rect 642272 95600 642324 95606
rect 642272 95542 642324 95548
rect 627918 94480 627974 94489
rect 627918 94415 627974 94424
rect 627274 93528 627330 93537
rect 627274 93463 627330 93472
rect 626446 92576 626502 92585
rect 626446 92511 626502 92520
rect 625894 91624 625950 91633
rect 625894 91559 625950 91568
rect 623976 91066 624648 91094
rect 623976 90681 624004 91066
rect 623962 90672 624018 90681
rect 623962 90607 624018 90616
rect 623778 89720 623834 89729
rect 623778 89655 623834 89664
rect 623502 86048 623558 86057
rect 623502 85983 623558 85992
rect 623318 85096 623374 85105
rect 623318 85031 623374 85040
rect 623134 84144 623190 84153
rect 623134 84079 623190 84088
rect 622122 83192 622178 83201
rect 622122 83127 622178 83136
rect 622306 82240 622362 82249
rect 622306 82175 622362 82184
rect 621480 43444 621532 43450
rect 621480 43386 621532 43392
rect 621296 43240 621348 43246
rect 621296 43182 621348 43188
rect 622320 43110 622348 82175
rect 622490 81424 622546 81433
rect 622490 81359 622546 81368
rect 622504 43178 622532 81359
rect 631856 80974 631916 81002
rect 639308 80974 639368 81002
rect 631888 51066 631916 80974
rect 631876 51060 631928 51066
rect 631876 51002 631928 51008
rect 639340 45558 639368 80974
rect 642652 46918 642680 100014
rect 642824 95668 642876 95674
rect 642824 95610 642876 95616
rect 642732 95532 642784 95538
rect 642732 95474 642784 95480
rect 642744 92721 642772 95474
rect 642730 92712 642786 92721
rect 642730 92647 642786 92656
rect 642640 46912 642692 46918
rect 642640 46854 642692 46860
rect 642836 45626 642864 95610
rect 642916 95600 642968 95606
rect 642916 95542 642968 95548
rect 642928 52426 642956 95542
rect 643468 95124 643520 95130
rect 643468 95066 643520 95072
rect 643480 85270 643508 95066
rect 643572 94246 643600 100014
rect 643560 94240 643612 94246
rect 643560 94182 643612 94188
rect 644216 94110 644244 100014
rect 644204 94104 644256 94110
rect 644204 94046 644256 94052
rect 644768 93906 644796 100014
rect 644860 100014 645196 100042
rect 645840 100014 646176 100042
rect 646484 100014 646820 100042
rect 647220 100014 647556 100042
rect 647864 100014 648108 100042
rect 644860 95130 644888 100014
rect 646044 95940 646096 95946
rect 646044 95882 646096 95888
rect 645860 95872 645912 95878
rect 645860 95814 645912 95820
rect 644848 95124 644900 95130
rect 644848 95066 644900 95072
rect 644756 93900 644808 93906
rect 644756 93842 644808 93848
rect 645872 89729 645900 95814
rect 645952 95736 646004 95742
rect 645952 95678 646004 95684
rect 645858 89720 645914 89729
rect 645858 89655 645914 89664
rect 643468 85264 643520 85270
rect 643468 85206 643520 85212
rect 645964 82249 645992 95678
rect 646056 95554 646084 95882
rect 646148 95878 646176 100014
rect 646136 95872 646188 95878
rect 646136 95814 646188 95820
rect 646056 95526 646176 95554
rect 646044 95464 646096 95470
rect 646044 95406 646096 95412
rect 646056 87145 646084 95406
rect 646042 87136 646098 87145
rect 646042 87071 646098 87080
rect 646148 84697 646176 95526
rect 646792 95470 646820 100014
rect 647528 96354 647556 100014
rect 647516 96348 647568 96354
rect 647516 96290 647568 96296
rect 646780 95464 646832 95470
rect 646780 95406 646832 95412
rect 646596 94784 646648 94790
rect 646596 94726 646648 94732
rect 646608 85202 646636 94726
rect 648080 94518 648108 100014
rect 648172 100014 648508 100042
rect 649152 100014 649396 100042
rect 648172 94790 648200 100014
rect 648620 95396 648672 95402
rect 648620 95338 648672 95344
rect 648160 94784 648212 94790
rect 648160 94726 648212 94732
rect 648068 94512 648120 94518
rect 648068 94454 648120 94460
rect 648632 85542 648660 95338
rect 648804 94988 648856 94994
rect 648804 94930 648856 94936
rect 648620 85536 648672 85542
rect 648620 85478 648672 85484
rect 648816 85338 648844 94930
rect 648896 94852 648948 94858
rect 648896 94794 648948 94800
rect 648908 85406 648936 94794
rect 649368 94042 649396 100014
rect 649460 100014 649796 100042
rect 650104 100014 650440 100042
rect 650748 100014 651084 100042
rect 651728 100014 652064 100042
rect 652372 100014 652708 100042
rect 653016 100014 653352 100042
rect 649460 94858 649488 100014
rect 650104 94994 650132 100014
rect 650748 95402 650776 100014
rect 652036 95810 652064 100014
rect 652024 95804 652076 95810
rect 652024 95746 652076 95752
rect 652680 95674 652708 100014
rect 652668 95668 652720 95674
rect 652668 95610 652720 95616
rect 651840 95600 651892 95606
rect 651840 95542 651892 95548
rect 650736 95396 650788 95402
rect 650736 95338 650788 95344
rect 650092 94988 650144 94994
rect 650092 94930 650144 94936
rect 649448 94852 649500 94858
rect 649448 94794 649500 94800
rect 649356 94036 649408 94042
rect 649356 93978 649408 93984
rect 651852 85474 651880 95542
rect 653324 94790 653352 100014
rect 653416 100014 653752 100042
rect 654396 100014 654732 100042
rect 655040 100014 655376 100042
rect 655684 100014 656020 100042
rect 656328 100014 656664 100042
rect 656972 100014 657308 100042
rect 653416 95606 653444 100014
rect 654704 96558 654732 100014
rect 654692 96552 654744 96558
rect 654692 96494 654744 96500
rect 653956 96348 654008 96354
rect 653956 96290 654008 96296
rect 653404 95600 653456 95606
rect 653404 95542 653456 95548
rect 653312 94784 653364 94790
rect 653312 94726 653364 94732
rect 653128 93900 653180 93906
rect 653128 93842 653180 93848
rect 653140 90681 653168 93842
rect 653968 92585 653996 96290
rect 654048 94104 654100 94110
rect 654048 94046 654100 94052
rect 653954 92576 654010 92585
rect 653954 92511 654010 92520
rect 654060 91497 654088 94046
rect 655348 93401 655376 100014
rect 655992 96626 656020 100014
rect 655980 96620 656032 96626
rect 655980 96562 656032 96568
rect 656636 94722 656664 100014
rect 656992 95600 657044 95606
rect 656992 95542 657044 95548
rect 656624 94716 656676 94722
rect 656624 94658 656676 94664
rect 656900 94580 656952 94586
rect 656900 94522 656952 94528
rect 656912 94042 656940 94522
rect 656900 94036 656952 94042
rect 656900 93978 656952 93984
rect 655334 93392 655390 93401
rect 655334 93327 655390 93336
rect 654046 91488 654102 91497
rect 654046 91423 654102 91432
rect 653126 90672 653182 90681
rect 653126 90607 653182 90616
rect 657004 90409 657032 95542
rect 657084 95260 657136 95266
rect 657084 95202 657136 95208
rect 656990 90400 657046 90409
rect 656990 90335 657046 90344
rect 657096 88874 657124 95202
rect 657280 94654 657308 100014
rect 657372 100014 657616 100042
rect 657924 100014 658260 100042
rect 658904 100014 659148 100042
rect 657372 94761 657400 100014
rect 657728 99816 657780 99822
rect 657728 99758 657780 99764
rect 657740 95132 657768 99758
rect 657924 95266 657952 100014
rect 659120 96558 659148 100014
rect 659212 100014 659548 100042
rect 660284 100014 660620 100042
rect 658280 96552 658332 96558
rect 658280 96494 658332 96500
rect 659108 96552 659160 96558
rect 659108 96494 659160 96500
rect 657912 95260 657964 95266
rect 657912 95202 657964 95208
rect 658292 95132 658320 96494
rect 659212 95606 659240 100014
rect 659568 96620 659620 96626
rect 659568 96562 659620 96568
rect 659200 95600 659252 95606
rect 659200 95542 659252 95548
rect 659580 95132 659608 96562
rect 660592 95538 660620 100014
rect 660914 99822 660942 100028
rect 661572 100014 661908 100042
rect 662216 100014 662276 100042
rect 662860 100014 663288 100042
rect 660902 99816 660954 99822
rect 660902 99758 660954 99764
rect 661880 96626 661908 100014
rect 661868 96620 661920 96626
rect 661868 96562 661920 96568
rect 661960 95804 662012 95810
rect 661960 95746 662012 95752
rect 660580 95532 660632 95538
rect 660580 95474 660632 95480
rect 661408 95532 661460 95538
rect 661408 95474 661460 95480
rect 661420 95132 661448 95474
rect 661972 95132 662000 95746
rect 662248 95577 662276 100014
rect 663064 96620 663116 96626
rect 663064 96562 663116 96568
rect 662512 96552 662564 96558
rect 662512 96494 662564 96500
rect 662234 95568 662290 95577
rect 662234 95503 662290 95512
rect 662524 95132 662552 96494
rect 663076 95132 663104 96562
rect 657358 94752 657414 94761
rect 657358 94687 657414 94696
rect 657268 94648 657320 94654
rect 657268 94590 657320 94596
rect 658568 94586 658858 94602
rect 658556 94580 658858 94586
rect 658608 94574 658858 94580
rect 658556 94522 658608 94528
rect 659844 94512 659896 94518
rect 660396 94512 660448 94518
rect 659896 94460 660146 94466
rect 659844 94454 660146 94460
rect 660448 94460 660698 94466
rect 660396 94454 660698 94460
rect 659856 94438 660146 94454
rect 660408 94438 660698 94454
rect 663260 93809 663288 100014
rect 663352 100014 663504 100042
rect 663246 93800 663302 93809
rect 663246 93735 663302 93744
rect 663352 93378 663380 100014
rect 663524 95872 663576 95878
rect 663524 95814 663576 95820
rect 663432 95396 663484 95402
rect 663432 95338 663484 95344
rect 663168 93350 663380 93378
rect 658016 88874 658306 88890
rect 657084 88868 657136 88874
rect 657084 88810 657136 88816
rect 658004 88868 658306 88874
rect 658056 88862 658306 88868
rect 658004 88810 658056 88816
rect 663168 88806 663196 93350
rect 663444 93129 663472 95338
rect 663430 93120 663486 93129
rect 663430 93055 663486 93064
rect 663536 92313 663564 95814
rect 663892 95668 663944 95674
rect 663892 95610 663944 95616
rect 663800 94784 663852 94790
rect 663800 94726 663852 94732
rect 663708 94716 663760 94722
rect 663708 94658 663760 94664
rect 663616 94648 663668 94654
rect 663616 94590 663668 94596
rect 663522 92304 663578 92313
rect 663522 92239 663578 92248
rect 663628 91474 663656 94590
rect 663444 91446 663656 91474
rect 663248 91112 663300 91118
rect 663248 91054 663300 91060
rect 659476 88800 659528 88806
rect 663156 88800 663208 88806
rect 662142 88768 662198 88777
rect 659528 88748 659594 88754
rect 659476 88742 659594 88748
rect 659488 88726 659594 88742
rect 661986 88726 662142 88754
rect 663156 88742 663208 88748
rect 662142 88703 662198 88712
rect 663260 88618 663288 91054
rect 663444 89593 663472 91446
rect 663720 91338 663748 94658
rect 663536 91310 663748 91338
rect 663536 91089 663564 91310
rect 663812 91094 663840 94726
rect 663904 91118 663932 95610
rect 665180 95192 665232 95198
rect 665180 95134 665232 95140
rect 663522 91080 663578 91089
rect 663522 91015 663578 91024
rect 663628 91066 663840 91094
rect 663892 91112 663944 91118
rect 663628 90409 663656 91066
rect 663892 91054 663944 91060
rect 663614 90400 663670 90409
rect 663614 90335 663670 90344
rect 663430 89584 663486 89593
rect 663430 89519 663486 89528
rect 662538 88590 663288 88618
rect 657188 85542 657216 88196
rect 657176 85536 657228 85542
rect 657176 85478 657228 85484
rect 651840 85468 651892 85474
rect 651840 85410 651892 85416
rect 648896 85400 648948 85406
rect 648896 85342 648948 85348
rect 657740 85338 657768 88196
rect 658844 85474 658872 88196
rect 658832 85468 658884 85474
rect 658832 85410 658884 85416
rect 648804 85332 648856 85338
rect 648804 85274 648856 85280
rect 657728 85332 657780 85338
rect 657728 85274 657780 85280
rect 660132 85270 660160 88196
rect 660684 85406 660712 88196
rect 660672 85400 660724 85406
rect 660672 85342 660724 85348
rect 660120 85264 660172 85270
rect 660120 85206 660172 85212
rect 661420 85202 661448 88196
rect 646596 85196 646648 85202
rect 646596 85138 646648 85144
rect 661408 85196 661460 85202
rect 661408 85138 661460 85144
rect 646134 84688 646190 84697
rect 646134 84623 646190 84632
rect 645950 82240 646006 82249
rect 645950 82175 646006 82184
rect 642916 52420 642968 52426
rect 642916 52362 642968 52368
rect 661130 47560 661186 47569
rect 661130 47495 661186 47504
rect 642824 45620 642876 45626
rect 642824 45562 642876 45568
rect 639328 45552 639380 45558
rect 639328 45494 639380 45500
rect 661144 44130 661172 47495
rect 665192 47433 665220 95134
rect 666572 48521 666600 170054
rect 666652 169992 666704 169998
rect 666652 169934 666704 169940
rect 666664 128058 666692 169934
rect 666742 168600 666798 168609
rect 666742 168535 666798 168544
rect 666756 165209 666784 168535
rect 666742 165200 666798 165209
rect 666742 165135 666798 165144
rect 666742 163568 666798 163577
rect 666742 163503 666798 163512
rect 666756 160177 666784 163503
rect 666848 161022 666876 177942
rect 666836 161016 666888 161022
rect 666836 160958 666888 160964
rect 666742 160168 666798 160177
rect 666742 160103 666798 160112
rect 666742 158400 666798 158409
rect 666742 158335 666798 158344
rect 666756 155009 666784 158335
rect 666742 155000 666798 155009
rect 666742 154935 666798 154944
rect 666742 153368 666798 153377
rect 666742 153303 666798 153312
rect 666756 149977 666784 153303
rect 666742 149968 666798 149977
rect 666742 149903 666798 149912
rect 666742 148200 666798 148209
rect 666742 148135 666798 148144
rect 666756 144945 666784 148135
rect 666742 144936 666798 144945
rect 666742 144871 666798 144880
rect 666742 143168 666798 143177
rect 666742 143103 666798 143112
rect 666756 139777 666784 143103
rect 666742 139768 666798 139777
rect 666742 139703 666798 139712
rect 666742 132968 666798 132977
rect 666742 132903 666798 132912
rect 666756 129577 666784 132903
rect 666742 129568 666798 129577
rect 666742 129503 666798 129512
rect 666664 128030 666784 128058
rect 666650 127936 666706 127945
rect 666650 127871 666706 127880
rect 666664 124545 666692 127871
rect 666650 124536 666706 124545
rect 666650 124471 666706 124480
rect 666650 122904 666706 122913
rect 666650 122839 666706 122848
rect 666664 119513 666692 122839
rect 666650 119504 666706 119513
rect 666650 119439 666706 119448
rect 666756 115938 666784 128030
rect 666744 115932 666796 115938
rect 666744 115874 666796 115880
rect 666940 107545 666968 213250
rect 667032 176866 667060 216702
rect 667124 206009 667152 226306
rect 667110 206000 667166 206009
rect 667110 205935 667166 205944
rect 667020 176860 667072 176866
rect 667020 176802 667072 176808
rect 669976 132666 670004 283154
rect 670056 281580 670108 281586
rect 670056 281522 670108 281528
rect 670068 132802 670096 281522
rect 670148 280424 670200 280430
rect 670148 280366 670200 280372
rect 670160 132938 670188 280366
rect 670252 177002 670280 287030
rect 670332 284980 670384 284986
rect 670332 284922 670384 284928
rect 670344 177138 670372 284922
rect 671632 278390 671660 311850
rect 671712 310276 671764 310282
rect 671712 310218 671764 310224
rect 671620 278384 671672 278390
rect 671620 278326 671672 278332
rect 671724 278322 671752 310218
rect 671804 309460 671856 309466
rect 671804 309402 671856 309408
rect 671712 278316 671764 278322
rect 671712 278258 671764 278264
rect 671816 278118 671844 309402
rect 671804 278112 671856 278118
rect 671804 278054 671856 278060
rect 671894 217152 671950 217161
rect 671894 217087 671950 217096
rect 670698 194032 670754 194041
rect 670698 193967 670754 193976
rect 670712 190641 670740 193967
rect 670698 190632 670754 190641
rect 670698 190567 670754 190576
rect 670698 178800 670754 178809
rect 670698 178735 670754 178744
rect 670332 177132 670384 177138
rect 670332 177074 670384 177080
rect 670240 176996 670292 177002
rect 670240 176938 670292 176944
rect 670712 175409 670740 178735
rect 670698 175400 670754 175409
rect 670698 175335 670754 175344
rect 670698 138136 670754 138145
rect 670698 138071 670754 138080
rect 670712 134745 670740 138071
rect 670698 134736 670754 134745
rect 670698 134671 670754 134680
rect 670148 132932 670200 132938
rect 670148 132874 670200 132880
rect 670056 132796 670108 132802
rect 670056 132738 670108 132744
rect 669964 132660 670016 132666
rect 669964 132602 670016 132608
rect 671908 130082 671936 217087
rect 672000 178809 672028 883186
rect 673380 739694 673408 894610
rect 675956 894402 675984 896679
rect 676034 896336 676090 896345
rect 676034 896271 676090 896280
rect 676048 894538 676076 896271
rect 676126 895248 676182 895257
rect 676126 895183 676182 895192
rect 676036 894532 676088 894538
rect 676036 894474 676088 894480
rect 676140 894470 676168 895183
rect 676128 894464 676180 894470
rect 676128 894406 676180 894412
rect 675944 894396 675996 894402
rect 675944 894338 675996 894344
rect 676034 893888 676090 893897
rect 676034 893823 676036 893832
rect 676088 893823 676090 893832
rect 676036 893794 676088 893800
rect 676034 893072 676090 893081
rect 676034 893007 676036 893016
rect 676088 893007 676090 893016
rect 676036 892978 676088 892984
rect 679622 892664 679678 892673
rect 679622 892599 679678 892608
rect 676034 892256 676090 892265
rect 676034 892191 676090 892200
rect 676048 891546 676076 892191
rect 679346 891848 679402 891857
rect 679346 891783 679402 891792
rect 674288 891540 674340 891546
rect 674288 891482 674340 891488
rect 676036 891540 676088 891546
rect 676036 891482 676088 891488
rect 673828 887868 673880 887874
rect 673828 887810 673880 887816
rect 673736 886100 673788 886106
rect 673736 886042 673788 886048
rect 673748 873662 673776 886042
rect 673736 873656 673788 873662
rect 673736 873598 673788 873604
rect 673840 872370 673868 887810
rect 673828 872364 673880 872370
rect 673828 872306 673880 872312
rect 674300 865774 674328 891482
rect 679162 891440 679218 891449
rect 679162 891375 679218 891384
rect 676034 891032 676090 891041
rect 676034 890967 676090 890976
rect 676048 890730 676076 890967
rect 674748 890724 674800 890730
rect 674748 890666 674800 890672
rect 676036 890724 676088 890730
rect 676036 890666 676088 890672
rect 674564 888820 674616 888826
rect 674564 888762 674616 888768
rect 674472 886032 674524 886038
rect 674472 885974 674524 885980
rect 674484 869990 674512 885974
rect 674472 869984 674524 869990
rect 674472 869926 674524 869932
rect 674576 867610 674604 888762
rect 674656 880252 674708 880258
rect 674656 880194 674708 880200
rect 674668 873798 674696 880194
rect 674656 873792 674708 873798
rect 674656 873734 674708 873740
rect 674656 873656 674708 873662
rect 674656 873598 674708 873604
rect 674668 868766 674696 873598
rect 674760 872506 674788 890666
rect 676034 890624 676090 890633
rect 676034 890559 676090 890568
rect 675942 888992 675998 889001
rect 675942 888927 675998 888936
rect 675956 888826 675984 888927
rect 675944 888820 675996 888826
rect 675944 888762 675996 888768
rect 676048 888758 676076 890559
rect 678978 890216 679034 890225
rect 678978 890151 679034 890160
rect 675024 888752 675076 888758
rect 675024 888694 675076 888700
rect 676036 888752 676088 888758
rect 676036 888694 676088 888700
rect 674840 883040 674892 883046
rect 674840 882982 674892 882988
rect 674852 877334 674880 882982
rect 674932 880456 674984 880462
rect 674932 880398 674984 880404
rect 674840 877328 674892 877334
rect 674840 877270 674892 877276
rect 674944 872658 674972 880398
rect 675036 872778 675064 888694
rect 676034 888584 676090 888593
rect 676034 888519 676090 888528
rect 676048 887874 676076 888519
rect 676036 887868 676088 887874
rect 676036 887810 676088 887816
rect 676034 887768 676090 887777
rect 676034 887703 676090 887712
rect 675942 887360 675998 887369
rect 675942 887295 675998 887304
rect 675956 886106 675984 887295
rect 675944 886100 675996 886106
rect 675944 886042 675996 886048
rect 676048 886038 676076 887703
rect 676036 886032 676088 886038
rect 676036 885974 676088 885980
rect 675392 883312 675444 883318
rect 675392 883254 675444 883260
rect 675300 883176 675352 883182
rect 675300 883118 675352 883124
rect 675208 880388 675260 880394
rect 675208 880330 675260 880336
rect 675116 880320 675168 880326
rect 675116 880262 675168 880268
rect 675128 873882 675156 880262
rect 675220 874934 675248 880330
rect 675312 877418 675340 883118
rect 675404 878084 675432 883254
rect 678992 883182 679020 890151
rect 679070 888176 679126 888185
rect 679070 888111 679126 888120
rect 678980 883176 679032 883182
rect 678980 883118 679032 883124
rect 675760 883108 675812 883114
rect 675760 883050 675812 883056
rect 675772 878422 675800 883050
rect 679084 880462 679112 888111
rect 679072 880456 679124 880462
rect 679072 880398 679124 880404
rect 679176 880394 679204 891375
rect 679254 889808 679310 889817
rect 679254 889743 679310 889752
rect 679164 880388 679216 880394
rect 679164 880330 679216 880336
rect 679268 880326 679296 889743
rect 679360 883114 679388 891783
rect 679438 889400 679494 889409
rect 679438 889335 679494 889344
rect 679348 883108 679400 883114
rect 679348 883050 679400 883056
rect 679256 880320 679308 880326
rect 679256 880262 679308 880268
rect 679452 880258 679480 889335
rect 679530 885048 679586 885057
rect 679530 884983 679586 884992
rect 679544 883250 679572 884983
rect 679532 883244 679584 883250
rect 679532 883186 679584 883192
rect 679636 883046 679664 892599
rect 679624 883040 679676 883046
rect 679624 882982 679676 882988
rect 679440 880252 679492 880258
rect 679440 880194 679492 880200
rect 675760 878416 675812 878422
rect 675760 878358 675812 878364
rect 675760 877804 675812 877810
rect 675760 877746 675812 877752
rect 675772 877540 675800 877746
rect 675312 877390 675432 877418
rect 675300 877328 675352 877334
rect 675300 877270 675352 877276
rect 675312 876262 675340 877270
rect 675404 876860 675432 877390
rect 675312 876234 675418 876262
rect 675220 874906 675524 874934
rect 675496 874412 675524 874906
rect 675128 873854 675340 873882
rect 675116 873792 675168 873798
rect 675116 873734 675168 873740
rect 675312 873746 675340 873854
rect 675404 873746 675432 873868
rect 675128 873202 675156 873734
rect 675312 873718 675432 873746
rect 675128 873174 675418 873202
rect 675024 872772 675076 872778
rect 675024 872714 675076 872720
rect 674944 872630 675156 872658
rect 675128 872590 675156 872630
rect 675024 872568 675076 872574
rect 675128 872562 675340 872590
rect 675024 872510 675076 872516
rect 675312 872522 675340 872562
rect 675404 872522 675432 872576
rect 674748 872500 674800 872506
rect 674748 872442 674800 872448
rect 674748 872364 674800 872370
rect 674748 872306 674800 872312
rect 674760 869446 674788 872306
rect 674748 869440 674800 869446
rect 674748 869382 674800 869388
rect 674656 868760 674708 868766
rect 674656 868702 674708 868708
rect 674564 867604 674616 867610
rect 674564 867546 674616 867552
rect 674288 865768 674340 865774
rect 674288 865710 674340 865716
rect 675036 863342 675064 872510
rect 675208 872500 675260 872506
rect 675312 872494 675432 872522
rect 675208 872442 675260 872448
rect 675116 872228 675168 872234
rect 675116 872170 675168 872176
rect 675128 867694 675156 872170
rect 675220 870074 675248 872442
rect 675220 870046 675418 870074
rect 675208 869984 675260 869990
rect 675208 869926 675260 869932
rect 675220 869530 675248 869926
rect 675220 869502 675418 869530
rect 675208 869440 675260 869446
rect 675208 869382 675260 869388
rect 675220 868889 675248 869382
rect 675220 868861 675418 868889
rect 675208 868760 675260 868766
rect 675208 868702 675260 868708
rect 675220 868238 675248 868702
rect 675220 868210 675418 868238
rect 675128 867666 675418 867694
rect 675116 867604 675168 867610
rect 675116 867546 675168 867552
rect 675128 867049 675156 867546
rect 675128 867021 675418 867049
rect 675128 865830 675418 865858
rect 675128 863870 675156 865830
rect 675208 865768 675260 865774
rect 675208 865710 675260 865716
rect 675220 865209 675248 865710
rect 675220 865181 675418 865209
rect 675116 863864 675168 863870
rect 675116 863806 675168 863812
rect 675312 863382 675432 863410
rect 675312 863342 675340 863382
rect 675036 863314 675340 863342
rect 675404 863328 675432 863382
rect 675392 792192 675444 792198
rect 675392 792134 675444 792140
rect 675404 788868 675432 792134
rect 675114 788352 675170 788361
rect 675170 788310 675418 788338
rect 675114 788287 675170 788296
rect 675128 787665 675418 787693
rect 675128 787273 675156 787665
rect 675114 787264 675170 787273
rect 675114 787199 675170 787208
rect 675128 787018 675418 787046
rect 675128 786729 675156 787018
rect 675114 786720 675170 786729
rect 675114 786655 675170 786664
rect 675128 785182 675418 785210
rect 675128 784786 675156 785182
rect 673736 784780 673788 784786
rect 673736 784722 673788 784728
rect 675116 784780 675168 784786
rect 675116 784722 675168 784728
rect 673644 780972 673696 780978
rect 673644 780914 673696 780920
rect 673552 744184 673604 744190
rect 673552 744126 673604 744132
rect 673564 739694 673592 744126
rect 673196 739666 673408 739694
rect 673472 739666 673592 739694
rect 673196 720374 673224 739666
rect 673472 732442 673500 739666
rect 673552 733916 673604 733922
rect 673552 733858 673604 733864
rect 673288 732414 673500 732442
rect 673288 727938 673316 732414
rect 673460 732352 673512 732358
rect 673460 732294 673512 732300
rect 673276 727932 673328 727938
rect 673276 727874 673328 727880
rect 673196 720346 673408 720374
rect 673380 714542 673408 720346
rect 673472 718758 673500 732294
rect 673564 718894 673592 733858
rect 673552 718888 673604 718894
rect 673552 718830 673604 718836
rect 673460 718752 673512 718758
rect 673460 718694 673512 718700
rect 673368 714536 673420 714542
rect 673368 714478 673420 714484
rect 673276 714060 673328 714066
rect 673276 714002 673328 714008
rect 672080 705152 672132 705158
rect 672080 705094 672132 705100
rect 671986 178800 672042 178809
rect 671986 178735 672042 178744
rect 672092 173641 672120 705094
rect 673288 669390 673316 714002
rect 673656 707878 673684 780914
rect 673748 711550 673776 784722
rect 674760 784638 675418 784666
rect 674656 783896 674708 783902
rect 674656 783838 674708 783844
rect 674564 780156 674616 780162
rect 674564 780098 674616 780104
rect 674288 779136 674340 779142
rect 674288 779078 674340 779084
rect 673828 778660 673880 778666
rect 673828 778602 673880 778608
rect 673840 745385 673868 778602
rect 673826 745376 673882 745385
rect 673826 745311 673882 745320
rect 673828 734188 673880 734194
rect 673828 734130 673880 734136
rect 673736 711544 673788 711550
rect 673736 711486 673788 711492
rect 673644 707872 673696 707878
rect 673644 707814 673696 707820
rect 673736 690192 673788 690198
rect 673736 690134 673788 690140
rect 673644 689172 673696 689178
rect 673644 689114 673696 689120
rect 673368 688628 673420 688634
rect 673368 688570 673420 688576
rect 673276 669384 673328 669390
rect 673276 669326 673328 669332
rect 672172 659728 672224 659734
rect 672172 659670 672224 659676
rect 672078 173632 672134 173641
rect 672078 173567 672134 173576
rect 672184 168609 672212 659670
rect 673276 644292 673328 644298
rect 673276 644234 673328 644240
rect 673288 637974 673316 644234
rect 673276 637968 673328 637974
rect 673276 637910 673328 637916
rect 673276 623824 673328 623830
rect 673276 623766 673328 623772
rect 672264 614644 672316 614650
rect 672264 614586 672316 614592
rect 672170 168600 672226 168609
rect 672170 168535 672226 168544
rect 671988 167068 672040 167074
rect 671988 167010 672040 167016
rect 671896 130076 671948 130082
rect 671896 130018 671948 130024
rect 672000 114345 672028 167010
rect 672276 163577 672304 614586
rect 673288 579086 673316 623766
rect 673380 616758 673408 688570
rect 673552 687880 673604 687886
rect 673552 687822 673604 687828
rect 673460 647760 673512 647766
rect 673460 647702 673512 647708
rect 673472 637158 673500 647702
rect 673460 637152 673512 637158
rect 673460 637094 673512 637100
rect 673564 620158 673592 687822
rect 673552 620152 673604 620158
rect 673552 620094 673604 620100
rect 673656 618118 673684 689114
rect 673748 680406 673776 690134
rect 673736 680400 673788 680406
rect 673736 680342 673788 680348
rect 673840 663134 673868 734130
rect 674300 708286 674328 779078
rect 674472 777368 674524 777374
rect 674472 777310 674524 777316
rect 674484 708898 674512 777310
rect 674576 745249 674604 780098
rect 674668 779618 674696 783838
rect 674656 779612 674708 779618
rect 674656 779554 674708 779560
rect 674760 773362 674788 784638
rect 675312 784094 675432 784122
rect 675312 783986 675340 784094
rect 674944 783958 675340 783986
rect 675404 783972 675432 784094
rect 674944 780722 674972 783958
rect 675220 783346 675418 783374
rect 675220 780978 675248 783346
rect 675208 780972 675260 780978
rect 675208 780914 675260 780920
rect 675312 780966 675432 780994
rect 675312 780858 675340 780966
rect 675220 780830 675340 780858
rect 675404 780844 675432 780966
rect 674944 780694 675064 780722
rect 675036 780094 675064 780694
rect 675024 780088 675076 780094
rect 675024 780030 675076 780036
rect 675220 779906 675248 780830
rect 675496 780162 675524 780300
rect 675484 780156 675536 780162
rect 675484 780098 675536 780104
rect 674944 779878 675248 779906
rect 674748 773356 674800 773362
rect 674748 773298 674800 773304
rect 674840 769684 674892 769690
rect 674840 769626 674892 769632
rect 674852 747974 674880 769626
rect 674668 747946 674880 747974
rect 674562 745240 674618 745249
rect 674562 745175 674618 745184
rect 674668 739694 674696 747946
rect 674668 739666 674788 739694
rect 674564 737316 674616 737322
rect 674564 737258 674616 737264
rect 674576 728142 674604 737258
rect 674656 735684 674708 735690
rect 674656 735626 674708 735632
rect 674668 728822 674696 735626
rect 674760 734913 674788 739666
rect 674840 736976 674892 736982
rect 674840 736918 674892 736924
rect 674746 734904 674802 734913
rect 674746 734839 674802 734848
rect 674748 734800 674800 734806
rect 674748 734742 674800 734748
rect 674760 730674 674788 734742
rect 674852 732086 674880 736918
rect 674840 732080 674892 732086
rect 674840 732022 674892 732028
rect 674760 730646 674880 730674
rect 674748 730516 674800 730522
rect 674748 730458 674800 730464
rect 674656 728816 674708 728822
rect 674656 728758 674708 728764
rect 674656 728680 674708 728686
rect 674656 728622 674708 728628
rect 674564 728136 674616 728142
rect 674564 728078 674616 728084
rect 674564 728000 674616 728006
rect 674564 727942 674616 727948
rect 674472 708892 674524 708898
rect 674472 708834 674524 708840
rect 674288 708280 674340 708286
rect 674288 708222 674340 708228
rect 674472 687336 674524 687342
rect 674472 687278 674524 687284
rect 674286 687168 674342 687177
rect 674286 687103 674342 687112
rect 674300 683942 674328 687103
rect 674288 683936 674340 683942
rect 674288 683878 674340 683884
rect 674288 680400 674340 680406
rect 674288 680342 674340 680348
rect 673828 663128 673880 663134
rect 673828 663070 673880 663076
rect 673736 649596 673788 649602
rect 673736 649538 673788 649544
rect 673748 644298 673776 649538
rect 673828 644632 673880 644638
rect 673828 644574 673880 644580
rect 673736 644292 673788 644298
rect 673736 644234 673788 644240
rect 673736 644156 673788 644162
rect 673736 644098 673788 644104
rect 673748 638110 673776 644098
rect 673736 638104 673788 638110
rect 673736 638046 673788 638052
rect 673736 637968 673788 637974
rect 673736 637910 673788 637916
rect 673644 618112 673696 618118
rect 673644 618054 673696 618060
rect 673368 616752 673420 616758
rect 673368 616694 673420 616700
rect 673644 603492 673696 603498
rect 673644 603434 673696 603440
rect 673552 600432 673604 600438
rect 673552 600374 673604 600380
rect 673460 598596 673512 598602
rect 673460 598538 673512 598544
rect 673472 583778 673500 598538
rect 673564 597310 673592 600374
rect 673552 597304 673604 597310
rect 673552 597246 673604 597252
rect 673552 597168 673604 597174
rect 673552 597110 673604 597116
rect 673460 583772 673512 583778
rect 673460 583714 673512 583720
rect 673564 583642 673592 597110
rect 673552 583636 673604 583642
rect 673552 583578 673604 583584
rect 673276 579080 673328 579086
rect 673276 579022 673328 579028
rect 673368 578468 673420 578474
rect 673368 578410 673420 578416
rect 672356 568608 672408 568614
rect 672356 568550 672408 568556
rect 672262 163568 672318 163577
rect 672262 163503 672318 163512
rect 672368 158409 672396 568550
rect 673092 554736 673144 554742
rect 673092 554678 673144 554684
rect 673104 548010 673132 554678
rect 673184 552220 673236 552226
rect 673184 552162 673236 552168
rect 673092 548004 673144 548010
rect 673092 547946 673144 547952
rect 673196 547670 673224 552162
rect 673276 549024 673328 549030
rect 673276 548966 673328 548972
rect 673184 547664 673236 547670
rect 673184 547606 673236 547612
rect 673288 544474 673316 548966
rect 673276 544468 673328 544474
rect 673276 544410 673328 544416
rect 673380 534138 673408 578410
rect 673460 568812 673512 568818
rect 673460 568754 673512 568760
rect 673472 554742 673500 568754
rect 673460 554736 673512 554742
rect 673460 554678 673512 554684
rect 673550 554704 673606 554713
rect 673550 554639 673606 554648
rect 673460 554600 673512 554606
rect 673460 554542 673512 554548
rect 673472 549030 673500 554542
rect 673460 549024 673512 549030
rect 673460 548966 673512 548972
rect 673460 548888 673512 548894
rect 673460 548830 673512 548836
rect 673368 534132 673420 534138
rect 673368 534074 673420 534080
rect 672448 524476 672500 524482
rect 672448 524418 672500 524424
rect 672354 158400 672410 158409
rect 672354 158335 672410 158344
rect 672460 153377 672488 524418
rect 673472 492590 673500 548830
rect 673460 492584 673512 492590
rect 673460 492526 673512 492532
rect 673564 483478 673592 554639
rect 673656 529854 673684 603434
rect 673748 576774 673776 637910
rect 673840 637294 673868 644574
rect 673828 637288 673880 637294
rect 673828 637230 673880 637236
rect 673828 637152 673880 637158
rect 673828 637094 673880 637100
rect 673736 576768 673788 576774
rect 673736 576710 673788 576716
rect 673840 572422 673868 637094
rect 674300 620974 674328 680342
rect 674288 620968 674340 620974
rect 674288 620910 674340 620916
rect 674484 618254 674512 687278
rect 674576 665990 674604 727942
rect 674668 718842 674696 728622
rect 674760 718978 674788 730458
rect 674852 727870 674880 730646
rect 674840 727864 674892 727870
rect 674840 727806 674892 727812
rect 674944 720374 674972 779878
rect 675024 779748 675076 779754
rect 675024 779690 675076 779696
rect 675036 773430 675064 779690
rect 675220 779674 675418 779702
rect 675116 779612 675168 779618
rect 675116 779554 675168 779560
rect 675128 778478 675156 779554
rect 675220 779142 675248 779674
rect 675208 779136 675260 779142
rect 675208 779078 675260 779084
rect 675312 779062 675432 779090
rect 675312 779022 675340 779062
rect 675220 778994 675340 779022
rect 675404 779008 675432 779062
rect 675220 778666 675248 778994
rect 675208 778660 675260 778666
rect 675208 778602 675260 778608
rect 675128 778450 675418 778478
rect 675404 777374 675432 777852
rect 675392 777368 675444 777374
rect 675392 777310 675444 777316
rect 675128 776614 675418 776642
rect 675128 775538 675156 776614
rect 675220 776002 675340 776030
rect 675116 775532 675168 775538
rect 675116 775474 675168 775480
rect 675024 773424 675076 773430
rect 675024 773366 675076 773372
rect 675220 737322 675248 776002
rect 675312 775962 675340 776002
rect 675404 775962 675432 776016
rect 675312 775934 675432 775962
rect 675404 773650 675432 774180
rect 675312 773622 675432 773650
rect 675312 769690 675340 773622
rect 675668 773424 675720 773430
rect 675668 773366 675720 773372
rect 675300 769684 675352 769690
rect 675300 769626 675352 769632
rect 675680 767294 675708 773366
rect 675760 773356 675812 773362
rect 675760 773298 675812 773304
rect 675312 767266 675708 767294
rect 675208 737316 675260 737322
rect 675208 737258 675260 737264
rect 675208 737044 675260 737050
rect 675208 736986 675260 736992
rect 675220 733666 675248 736986
rect 675312 733854 675340 767266
rect 675392 747992 675444 747998
rect 675392 747934 675444 747940
rect 675404 743852 675432 747934
rect 675772 744190 675800 773298
rect 675760 744184 675812 744190
rect 675760 744126 675812 744132
rect 675404 742937 675432 743308
rect 675390 742928 675446 742937
rect 675390 742863 675446 742872
rect 675404 742529 675432 742696
rect 675390 742520 675446 742529
rect 675390 742455 675446 742464
rect 675496 741713 675524 742016
rect 675482 741704 675538 741713
rect 675482 741639 675538 741648
rect 675404 739809 675432 740180
rect 675390 739800 675446 739809
rect 675390 739735 675446 739744
rect 675404 739129 675432 739636
rect 675390 739120 675446 739129
rect 675390 739055 675446 739064
rect 675404 738721 675432 739024
rect 675390 738712 675446 738721
rect 675390 738647 675446 738656
rect 675404 738041 675432 738344
rect 675390 738032 675446 738041
rect 675390 737967 675446 737976
rect 675404 735690 675432 735896
rect 675392 735684 675444 735690
rect 675392 735626 675444 735632
rect 675404 734806 675432 735319
rect 675392 734800 675444 734806
rect 675392 734742 675444 734748
rect 675404 734194 675432 734672
rect 675392 734188 675444 734194
rect 675392 734130 675444 734136
rect 675404 733922 675432 734031
rect 675392 733916 675444 733922
rect 675392 733858 675444 733864
rect 675300 733848 675352 733854
rect 675300 733790 675352 733796
rect 675220 733638 675432 733666
rect 675300 733508 675352 733514
rect 675404 733479 675432 733638
rect 675300 733450 675352 733456
rect 675206 733408 675262 733417
rect 675206 733343 675262 733352
rect 675220 728074 675248 733343
rect 675208 728068 675260 728074
rect 675208 728010 675260 728016
rect 675208 727932 675260 727938
rect 675208 727874 675260 727880
rect 675116 727864 675168 727870
rect 675116 727806 675168 727812
rect 674944 720346 675064 720374
rect 674760 718950 674880 718978
rect 674668 718814 674788 718842
rect 674656 718752 674708 718758
rect 674656 718694 674708 718700
rect 674564 665984 674616 665990
rect 674564 665926 674616 665932
rect 674668 664358 674696 718694
rect 674760 665106 674788 718814
rect 674852 709334 674880 718950
rect 675036 712162 675064 720346
rect 675024 712156 675076 712162
rect 675024 712098 675076 712104
rect 675128 709334 675156 727806
rect 675220 714950 675248 727874
rect 675312 718978 675340 733450
rect 675404 732358 675432 732836
rect 675392 732352 675444 732358
rect 675392 732294 675444 732300
rect 675392 732080 675444 732086
rect 675392 732022 675444 732028
rect 675404 731612 675432 732022
rect 675404 730522 675432 731000
rect 675392 730516 675444 730522
rect 675392 730458 675444 730464
rect 675404 728686 675432 729164
rect 675392 728680 675444 728686
rect 675392 728622 675444 728628
rect 676128 728136 676180 728142
rect 676128 728078 676180 728084
rect 675312 718950 675708 718978
rect 675576 718888 675628 718894
rect 675576 718830 675628 718836
rect 675208 714944 675260 714950
rect 675208 714886 675260 714892
rect 674852 709306 675064 709334
rect 675128 709306 675524 709334
rect 675036 701054 675064 709306
rect 675392 703860 675444 703866
rect 675392 703802 675444 703808
rect 674944 701026 675064 701054
rect 674944 684162 674972 701026
rect 675404 698875 675432 703802
rect 675496 699417 675524 709306
rect 675482 699408 675538 699417
rect 675482 699343 675538 699352
rect 675588 699281 675616 718830
rect 675680 708801 675708 718950
rect 675758 716544 675814 716553
rect 675758 716479 675814 716488
rect 675772 715154 675800 716479
rect 675850 716136 675906 716145
rect 675850 716071 675906 716080
rect 675760 715148 675812 715154
rect 675760 715090 675812 715096
rect 675864 715018 675892 716071
rect 675942 715728 675998 715737
rect 675942 715663 675998 715672
rect 675956 715290 675984 715663
rect 676036 715420 676088 715426
rect 676036 715362 676088 715368
rect 676048 715329 676076 715362
rect 676034 715320 676090 715329
rect 675944 715284 675996 715290
rect 676034 715255 676090 715264
rect 675944 715226 675996 715232
rect 675852 715012 675904 715018
rect 675852 714954 675904 714960
rect 675760 714944 675812 714950
rect 675760 714886 675812 714892
rect 676034 714912 676090 714921
rect 675772 709209 675800 714886
rect 676034 714847 676036 714856
rect 676088 714847 676090 714856
rect 676036 714818 676088 714824
rect 676036 714536 676088 714542
rect 676034 714504 676036 714513
rect 676088 714504 676090 714513
rect 676034 714439 676090 714448
rect 676034 714096 676090 714105
rect 676034 714031 676036 714040
rect 676088 714031 676090 714040
rect 676036 714002 676088 714008
rect 676034 713688 676090 713697
rect 676034 713623 676090 713632
rect 675850 713280 675906 713289
rect 675850 713215 675906 713224
rect 675864 712230 675892 713215
rect 675942 712872 675998 712881
rect 675942 712807 675998 712816
rect 675956 712366 675984 712807
rect 676048 712570 676076 713623
rect 676036 712564 676088 712570
rect 676036 712506 676088 712512
rect 676034 712464 676090 712473
rect 676034 712399 676090 712408
rect 675944 712360 675996 712366
rect 675944 712302 675996 712308
rect 676048 712298 676076 712399
rect 676036 712292 676088 712298
rect 676036 712234 676088 712240
rect 675852 712224 675904 712230
rect 675852 712166 675904 712172
rect 675944 712156 675996 712162
rect 675944 712098 675996 712104
rect 675956 710433 675984 712098
rect 676034 711648 676090 711657
rect 676140 711634 676168 728078
rect 678980 728068 679032 728074
rect 678980 728010 679032 728016
rect 676090 711606 676168 711634
rect 676034 711583 676090 711592
rect 676036 711544 676088 711550
rect 676036 711486 676088 711492
rect 676048 710841 676076 711486
rect 676034 710832 676090 710841
rect 676034 710767 676090 710776
rect 675942 710424 675998 710433
rect 675942 710359 675998 710368
rect 678992 710025 679020 728010
rect 703694 717196 703722 717332
rect 704154 717196 704182 717332
rect 704614 717196 704642 717332
rect 705074 717196 705102 717332
rect 705534 717196 705562 717332
rect 705994 717196 706022 717332
rect 706454 717196 706482 717332
rect 706914 717196 706942 717332
rect 707374 717196 707402 717332
rect 707834 717196 707862 717332
rect 708294 717196 708322 717332
rect 708754 717196 708782 717332
rect 709214 717196 709242 717332
rect 678978 710016 679034 710025
rect 678978 709951 679034 709960
rect 675758 709200 675814 709209
rect 675758 709135 675814 709144
rect 676036 708892 676088 708898
rect 676036 708834 676088 708840
rect 675666 708792 675722 708801
rect 675666 708727 675722 708736
rect 676048 708393 676076 708834
rect 676034 708384 676090 708393
rect 676034 708319 676090 708328
rect 676036 708280 676088 708286
rect 676036 708222 676088 708228
rect 676048 707985 676076 708222
rect 676034 707976 676090 707985
rect 676034 707911 676090 707920
rect 676036 707872 676088 707878
rect 676036 707814 676088 707820
rect 676048 707577 676076 707814
rect 676034 707568 676090 707577
rect 676034 707503 676090 707512
rect 676034 706344 676090 706353
rect 676034 706279 676090 706288
rect 676048 705158 676076 706279
rect 676036 705152 676088 705158
rect 676034 705120 676036 705129
rect 676088 705120 676090 705129
rect 676034 705055 676090 705064
rect 676048 705029 676076 705055
rect 675574 699272 675630 699281
rect 675574 699207 675630 699216
rect 675128 698329 675418 698337
rect 675114 698320 675418 698329
rect 675170 698309 675418 698320
rect 675114 698255 675170 698264
rect 675772 697241 675800 697680
rect 675758 697232 675814 697241
rect 675758 697167 675814 697176
rect 675128 697021 675418 697049
rect 675128 695609 675156 697021
rect 675114 695600 675170 695609
rect 675114 695535 675170 695544
rect 675128 695181 675418 695209
rect 675128 694793 675156 695181
rect 675114 694784 675170 694793
rect 675114 694719 675170 694728
rect 675312 694742 675432 694770
rect 675114 694648 675170 694657
rect 675312 694634 675340 694742
rect 675170 694606 675340 694634
rect 675404 694620 675432 694742
rect 675114 694583 675170 694592
rect 675128 693994 675418 694022
rect 675128 687886 675156 693994
rect 675772 693025 675800 693328
rect 675758 693016 675814 693025
rect 675758 692951 675814 692960
rect 675208 692912 675260 692918
rect 675208 692854 675260 692860
rect 675220 688770 675248 692854
rect 675312 690866 675418 690894
rect 675312 690198 675340 690866
rect 675300 690192 675352 690198
rect 675772 690169 675800 690336
rect 675300 690134 675352 690140
rect 675758 690160 675814 690169
rect 675758 690095 675814 690104
rect 675300 690056 675352 690062
rect 675300 689998 675352 690004
rect 675208 688764 675260 688770
rect 675208 688706 675260 688712
rect 675312 688650 675340 689998
rect 675496 689178 675524 689656
rect 675484 689172 675536 689178
rect 675484 689114 675536 689120
rect 675220 688622 675340 688650
rect 675404 688634 675432 689044
rect 675484 688764 675536 688770
rect 675484 688706 675536 688712
rect 675392 688628 675444 688634
rect 675116 687880 675168 687886
rect 675116 687822 675168 687828
rect 675220 686678 675248 688622
rect 675392 688570 675444 688576
rect 675496 688500 675524 688706
rect 675404 687342 675432 687820
rect 675392 687336 675444 687342
rect 675392 687278 675444 687284
rect 675220 686650 675340 686678
rect 675312 686610 675340 686650
rect 675404 686610 675432 686664
rect 675312 686582 675432 686610
rect 675128 685970 675418 685998
rect 675128 684282 675156 685970
rect 675206 685808 675262 685817
rect 675206 685743 675262 685752
rect 675220 684282 675248 685743
rect 675116 684276 675168 684282
rect 675116 684218 675168 684224
rect 675208 684276 675260 684282
rect 675208 684218 675260 684224
rect 674944 684134 675340 684162
rect 675024 684072 675076 684078
rect 674944 684020 675024 684026
rect 674944 684014 675076 684020
rect 674944 683998 675064 684014
rect 674748 665100 674800 665106
rect 674748 665042 674800 665048
rect 674656 664352 674708 664358
rect 674656 664294 674708 664300
rect 674656 648984 674708 648990
rect 674656 648926 674708 648932
rect 674564 648916 674616 648922
rect 674564 648858 674616 648864
rect 674576 638246 674604 648858
rect 674668 642258 674696 648926
rect 674748 645244 674800 645250
rect 674748 645186 674800 645192
rect 674656 642252 674708 642258
rect 674656 642194 674708 642200
rect 674656 642116 674708 642122
rect 674656 642058 674708 642064
rect 674564 638240 674616 638246
rect 674564 638182 674616 638188
rect 674564 638104 674616 638110
rect 674564 638046 674616 638052
rect 674472 618248 674524 618254
rect 674472 618190 674524 618196
rect 674288 609000 674340 609006
rect 674288 608942 674340 608948
rect 674300 599962 674328 608942
rect 674472 605124 674524 605130
rect 674472 605066 674524 605072
rect 674484 600438 674512 605066
rect 674472 600432 674524 600438
rect 674472 600374 674524 600380
rect 674472 600296 674524 600302
rect 674472 600238 674524 600244
rect 674288 599956 674340 599962
rect 674288 599898 674340 599904
rect 674288 599820 674340 599826
rect 674288 599762 674340 599768
rect 673828 572416 673880 572422
rect 673828 572358 673880 572364
rect 674300 571577 674328 599762
rect 674484 589286 674512 600238
rect 674472 589280 674524 589286
rect 674472 589222 674524 589228
rect 674472 583772 674524 583778
rect 674472 583714 674524 583720
rect 674286 571568 674342 571577
rect 674286 571503 674342 571512
rect 673828 564460 673880 564466
rect 673828 564402 673880 564408
rect 673736 553852 673788 553858
rect 673736 553794 673788 553800
rect 673748 544610 673776 553794
rect 673840 552226 673868 564402
rect 674288 558272 674340 558278
rect 674288 558214 674340 558220
rect 673828 552220 673880 552226
rect 673828 552162 673880 552168
rect 673828 552084 673880 552090
rect 673828 552026 673880 552032
rect 673840 545290 673868 552026
rect 673828 545284 673880 545290
rect 673828 545226 673880 545232
rect 674300 545154 674328 558214
rect 673828 545148 673880 545154
rect 673828 545090 673880 545096
rect 674288 545148 674340 545154
rect 674288 545090 674340 545096
rect 673736 544604 673788 544610
rect 673736 544546 673788 544552
rect 673736 544468 673788 544474
rect 673736 544410 673788 544416
rect 673644 529848 673696 529854
rect 673644 529790 673696 529796
rect 673552 483472 673604 483478
rect 673552 483414 673604 483420
rect 673748 482934 673776 544410
rect 673840 485654 673868 545090
rect 674288 544604 674340 544610
rect 674288 544546 674340 544552
rect 673828 485648 673880 485654
rect 673828 485590 673880 485596
rect 674300 483002 674328 544546
rect 674484 527134 674512 583714
rect 674576 572830 674604 638046
rect 674668 637378 674696 642058
rect 674760 637838 674788 645186
rect 674748 637832 674800 637838
rect 674748 637774 674800 637780
rect 674668 637350 674788 637378
rect 674656 637288 674708 637294
rect 674656 637230 674708 637236
rect 674668 610201 674696 637230
rect 674654 610192 674710 610201
rect 674654 610127 674710 610136
rect 674656 599956 674708 599962
rect 674656 599898 674708 599904
rect 674668 595474 674696 599898
rect 674656 595468 674708 595474
rect 674656 595410 674708 595416
rect 674656 595332 674708 595338
rect 674656 595274 674708 595280
rect 674668 583778 674696 595274
rect 674656 583772 674708 583778
rect 674656 583714 674708 583720
rect 674656 583636 674708 583642
rect 674656 583578 674708 583584
rect 674564 572824 674616 572830
rect 674564 572766 674616 572772
rect 674564 558068 674616 558074
rect 674564 558010 674616 558016
rect 674576 552090 674604 558010
rect 674564 552084 674616 552090
rect 674564 552026 674616 552032
rect 674564 551948 674616 551954
rect 674564 551890 674616 551896
rect 674472 527128 674524 527134
rect 674472 527070 674524 527076
rect 674576 485722 674604 551890
rect 674668 529922 674696 583578
rect 674760 573714 674788 637350
rect 674944 623762 674972 683998
rect 675024 683936 675076 683942
rect 675024 683878 675076 683884
rect 675208 683936 675260 683942
rect 675208 683878 675260 683884
rect 675036 665174 675064 683878
rect 675116 683664 675168 683670
rect 675116 683606 675168 683612
rect 675024 665168 675076 665174
rect 675024 665110 675076 665116
rect 675128 648990 675156 683606
rect 675220 667894 675248 683878
rect 675312 678978 675340 684134
rect 675404 683670 675432 684148
rect 675392 683664 675444 683670
rect 675392 683606 675444 683612
rect 675300 678972 675352 678978
rect 675300 678914 675352 678920
rect 679072 678972 679124 678978
rect 679072 678914 679124 678920
rect 676126 677968 676182 677977
rect 676126 677903 676182 677912
rect 676140 676481 676168 677903
rect 676126 676472 676182 676481
rect 676126 676407 676182 676416
rect 676218 671120 676274 671129
rect 676218 671055 676274 671064
rect 676034 670984 676090 670993
rect 676232 670954 676260 671055
rect 676034 670919 676090 670928
rect 676220 670948 676272 670954
rect 676048 670818 676076 670919
rect 676220 670890 676272 670896
rect 676036 670812 676088 670818
rect 676036 670754 676088 670760
rect 678978 670304 679034 670313
rect 678978 670239 679034 670248
rect 676126 669896 676182 669905
rect 676126 669831 676182 669840
rect 676036 669384 676088 669390
rect 676034 669352 676036 669361
rect 676088 669352 676090 669361
rect 676034 669287 676090 669296
rect 676140 668234 676168 669831
rect 676310 669488 676366 669497
rect 676310 669423 676366 669432
rect 676218 668264 676274 668273
rect 676128 668228 676180 668234
rect 676218 668199 676274 668208
rect 676128 668170 676180 668176
rect 676232 668166 676260 668199
rect 676220 668160 676272 668166
rect 675298 668128 675354 668137
rect 676220 668102 676272 668108
rect 675298 668063 675354 668072
rect 675208 667888 675260 667894
rect 675208 667830 675260 667836
rect 675116 648984 675168 648990
rect 675116 648926 675168 648932
rect 675312 648922 675340 668063
rect 676324 668030 676352 669423
rect 678992 668098 679020 670239
rect 678980 668092 679032 668098
rect 678980 668034 679032 668040
rect 676312 668024 676364 668030
rect 676312 667966 676364 667972
rect 676036 667888 676088 667894
rect 676036 667830 676088 667836
rect 676048 666097 676076 667830
rect 678978 667448 679034 667457
rect 678978 667383 679034 667392
rect 676218 667040 676274 667049
rect 676218 666975 676274 666984
rect 676034 666088 676090 666097
rect 676034 666023 676090 666032
rect 676036 665984 676088 665990
rect 676036 665926 676088 665932
rect 676048 665281 676076 665926
rect 676232 665310 676260 666975
rect 676220 665304 676272 665310
rect 676034 665272 676090 665281
rect 676220 665246 676272 665252
rect 678992 665242 679020 667383
rect 679084 666641 679112 678914
rect 679162 678872 679218 678881
rect 679162 678807 679218 678816
rect 679176 667049 679204 678807
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 679162 667040 679218 667049
rect 679162 666975 679218 666984
rect 679070 666632 679126 666641
rect 679070 666567 679126 666576
rect 676034 665207 676090 665216
rect 678980 665236 679032 665242
rect 678980 665178 679032 665184
rect 676036 665168 676088 665174
rect 676036 665110 676088 665116
rect 676048 664465 676076 665110
rect 676128 665100 676180 665106
rect 676128 665042 676180 665048
rect 676140 665009 676168 665042
rect 676126 665000 676182 665009
rect 676126 664935 676182 664944
rect 676034 664456 676090 664465
rect 676034 664391 676090 664400
rect 676036 664352 676088 664358
rect 676036 664294 676088 664300
rect 676048 663241 676076 664294
rect 676034 663232 676090 663241
rect 676034 663167 676090 663176
rect 676036 663128 676088 663134
rect 676036 663070 676088 663076
rect 676048 662833 676076 663070
rect 676034 662824 676090 662833
rect 676034 662759 676090 662768
rect 678978 660920 679034 660929
rect 678978 660855 679034 660864
rect 678992 660113 679020 660855
rect 678978 660104 679034 660113
rect 678978 660039 679034 660048
rect 678992 659734 679020 660039
rect 678980 659728 679032 659734
rect 678980 659670 679032 659676
rect 675392 656940 675444 656946
rect 675392 656882 675444 656888
rect 675404 653684 675432 656882
rect 675404 652905 675432 653140
rect 675390 652896 675446 652905
rect 675390 652831 675446 652840
rect 675496 652225 675524 652460
rect 675482 652216 675538 652225
rect 675482 652151 675538 652160
rect 675404 651681 675432 651848
rect 675390 651672 675446 651681
rect 675390 651607 675446 651616
rect 675404 649602 675432 650012
rect 675392 649596 675444 649602
rect 675392 649538 675444 649544
rect 675404 649233 675432 649468
rect 675390 649224 675446 649233
rect 675390 649159 675446 649168
rect 675300 648916 675352 648922
rect 675300 648858 675352 648864
rect 675036 648774 675418 648802
rect 675036 640370 675064 648774
rect 675116 648644 675168 648650
rect 675116 648586 675168 648592
rect 675128 643550 675156 648586
rect 675404 647766 675432 648176
rect 675392 647760 675444 647766
rect 675392 647702 675444 647708
rect 675208 645924 675260 645930
rect 675208 645866 675260 645872
rect 675220 643770 675248 645866
rect 675404 645250 675432 645660
rect 675392 645244 675444 645250
rect 675392 645186 675444 645192
rect 675404 644638 675432 645116
rect 675392 644632 675444 644638
rect 675392 644574 675444 644580
rect 675404 644162 675432 644475
rect 675392 644156 675444 644162
rect 675392 644098 675444 644104
rect 675220 643742 675340 643770
rect 675116 643544 675168 643550
rect 675116 643486 675168 643492
rect 675208 643408 675260 643414
rect 675208 643350 675260 643356
rect 675116 642252 675168 642258
rect 675116 642194 675168 642200
rect 675128 640830 675156 642194
rect 675116 640824 675168 640830
rect 675116 640766 675168 640772
rect 675036 640342 675156 640370
rect 675024 640280 675076 640286
rect 675024 640222 675076 640228
rect 674932 623756 674984 623762
rect 674932 623698 674984 623704
rect 674932 599004 674984 599010
rect 674932 598946 674984 598952
rect 674944 589422 674972 598946
rect 674932 589416 674984 589422
rect 674932 589358 674984 589364
rect 674932 589280 674984 589286
rect 674932 589222 674984 589228
rect 674748 573708 674800 573714
rect 674748 573650 674800 573656
rect 674748 555280 674800 555286
rect 674748 555222 674800 555228
rect 674760 545306 674788 555222
rect 674760 545278 674880 545306
rect 674748 545148 674800 545154
rect 674748 545090 674800 545096
rect 674656 529916 674708 529922
rect 674656 529858 674708 529864
rect 674760 493406 674788 545090
rect 674852 544814 674880 545278
rect 674840 544808 674892 544814
rect 674840 544750 674892 544756
rect 674840 542156 674892 542162
rect 674840 542098 674892 542104
rect 674748 493400 674800 493406
rect 674748 493342 674800 493348
rect 674852 485790 674880 542098
rect 674944 532846 674972 589222
rect 675036 576842 675064 640222
rect 675128 638602 675156 640342
rect 675220 638722 675248 643350
rect 675312 641458 675340 643742
rect 675496 643618 675524 643824
rect 675484 643612 675536 643618
rect 675484 643554 675536 643560
rect 675392 643544 675444 643550
rect 675392 643486 675444 643492
rect 675404 643280 675432 643486
rect 675404 642122 675432 642635
rect 675392 642116 675444 642122
rect 675392 642058 675444 642064
rect 675312 641430 675418 641458
rect 675300 640756 675352 640762
rect 675300 640698 675352 640704
rect 675312 638874 675340 640698
rect 675404 640286 675432 640795
rect 675392 640280 675444 640286
rect 675392 640222 675444 640228
rect 675312 638846 675432 638874
rect 675208 638716 675260 638722
rect 675208 638658 675260 638664
rect 675128 638574 675340 638602
rect 675208 638512 675260 638518
rect 675208 638454 675260 638460
rect 675116 638444 675168 638450
rect 675116 638386 675168 638392
rect 675024 576836 675076 576842
rect 675024 576778 675076 576784
rect 675128 576094 675156 638386
rect 675220 637922 675248 638454
rect 675312 638194 675340 638574
rect 675404 638489 675432 638846
rect 675390 638480 675446 638489
rect 675496 638450 675524 638928
rect 675390 638415 675446 638424
rect 675484 638444 675536 638450
rect 675484 638386 675536 638392
rect 675760 638240 675812 638246
rect 675666 638208 675722 638217
rect 675312 638166 675616 638194
rect 675220 637894 675340 637922
rect 675208 637832 675260 637838
rect 675208 637774 675260 637780
rect 675220 605130 675248 637774
rect 675312 610065 675340 637894
rect 675298 610056 675354 610065
rect 675298 609991 675354 610000
rect 675588 609006 675616 638166
rect 675760 638182 675812 638188
rect 675666 638143 675722 638152
rect 675680 637566 675708 638143
rect 675668 637560 675720 637566
rect 675668 637502 675720 637508
rect 675772 623506 675800 638182
rect 679072 637560 679124 637566
rect 679072 637502 679124 637508
rect 678978 626104 679034 626113
rect 678978 626039 679034 626048
rect 676310 625696 676366 625705
rect 676310 625631 676366 625640
rect 676034 625560 676090 625569
rect 676034 625495 676090 625504
rect 675942 623928 675998 623937
rect 676048 623898 676076 625495
rect 676218 624880 676274 624889
rect 676218 624815 676274 624824
rect 676126 624472 676182 624481
rect 676126 624407 676182 624416
rect 676140 623966 676168 624407
rect 676232 624102 676260 624815
rect 676220 624096 676272 624102
rect 676220 624038 676272 624044
rect 676324 624034 676352 625631
rect 678992 624170 679020 626039
rect 678980 624164 679032 624170
rect 678980 624106 679032 624112
rect 676312 624028 676364 624034
rect 676312 623970 676364 623976
rect 676128 623960 676180 623966
rect 676128 623902 676180 623908
rect 675942 623863 675998 623872
rect 676036 623892 676088 623898
rect 675956 623830 675984 623863
rect 676036 623834 676088 623840
rect 675944 623824 675996 623830
rect 675944 623766 675996 623772
rect 676036 623756 676088 623762
rect 676036 623698 676088 623704
rect 675942 623520 675998 623529
rect 675772 623478 675942 623506
rect 675942 623455 675998 623464
rect 675956 623454 675984 623455
rect 676048 621489 676076 623698
rect 676126 622840 676182 622849
rect 676126 622775 676182 622784
rect 676034 621480 676090 621489
rect 676034 621415 676090 621424
rect 676140 621178 676168 622775
rect 676310 622432 676366 622441
rect 676310 622367 676366 622376
rect 676218 622024 676274 622033
rect 676218 621959 676274 621968
rect 676128 621172 676180 621178
rect 676128 621114 676180 621120
rect 676232 621110 676260 621959
rect 676220 621104 676272 621110
rect 676220 621046 676272 621052
rect 676324 621042 676352 622367
rect 676312 621036 676364 621042
rect 676312 620978 676364 620984
rect 676036 620968 676088 620974
rect 676036 620910 676088 620916
rect 676048 620265 676076 620910
rect 676034 620256 676090 620265
rect 676034 620191 676090 620200
rect 676036 620152 676088 620158
rect 676036 620094 676088 620100
rect 676048 618633 676076 620094
rect 679084 619993 679112 637502
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 679070 619984 679126 619993
rect 679070 619919 679126 619928
rect 676034 618624 676090 618633
rect 676034 618559 676090 618568
rect 676036 618248 676088 618254
rect 676034 618216 676036 618225
rect 676088 618216 676090 618225
rect 676034 618151 676090 618160
rect 676036 618112 676088 618118
rect 676036 618054 676088 618060
rect 676048 617817 676076 618054
rect 676034 617808 676090 617817
rect 676034 617743 676090 617752
rect 676220 616752 676272 616758
rect 676218 616720 676220 616729
rect 676272 616720 676274 616729
rect 676218 616655 676274 616664
rect 679070 615904 679126 615913
rect 679070 615839 679126 615848
rect 679084 615097 679112 615839
rect 679070 615088 679126 615097
rect 679070 615023 679126 615032
rect 679084 614650 679112 615023
rect 679072 614644 679124 614650
rect 679072 614586 679124 614592
rect 675668 612876 675720 612882
rect 675668 612818 675720 612824
rect 675576 609000 675628 609006
rect 675576 608942 675628 608948
rect 675680 608668 675708 612818
rect 675298 608152 675354 608161
rect 675354 608110 675418 608138
rect 675298 608087 675354 608096
rect 675312 607465 675418 607493
rect 675312 607345 675340 607465
rect 675298 607336 675354 607345
rect 675298 607271 675354 607280
rect 675312 606818 675418 606846
rect 675312 605169 675340 606818
rect 675298 605160 675354 605169
rect 675208 605124 675260 605130
rect 675298 605095 675354 605104
rect 675208 605066 675260 605072
rect 675206 605024 675262 605033
rect 675262 604982 675418 605010
rect 675206 604959 675262 604968
rect 675206 604480 675262 604489
rect 675262 604438 675418 604466
rect 675206 604415 675262 604424
rect 675496 603498 675524 603772
rect 675484 603492 675536 603498
rect 675484 603434 675536 603440
rect 675220 603146 675418 603174
rect 675220 601905 675248 603146
rect 675206 601896 675262 601905
rect 675206 601831 675262 601840
rect 675208 601792 675260 601798
rect 675208 601734 675260 601740
rect 675220 598942 675248 601734
rect 675300 601724 675352 601730
rect 675300 601666 675352 601672
rect 675208 598936 675260 598942
rect 675208 598878 675260 598884
rect 675312 598874 675340 601666
rect 675496 600302 675524 600644
rect 675484 600296 675536 600302
rect 675484 600238 675536 600244
rect 675496 599826 675524 600100
rect 675484 599820 675536 599826
rect 675484 599762 675536 599768
rect 675404 599010 675432 599488
rect 675392 599004 675444 599010
rect 675392 598946 675444 598952
rect 675300 598868 675352 598874
rect 675300 598810 675352 598816
rect 675392 598732 675444 598738
rect 675392 598674 675444 598680
rect 675300 598664 675352 598670
rect 675300 598606 675352 598612
rect 675208 597304 675260 597310
rect 675208 597246 675260 597252
rect 675220 596306 675248 597246
rect 675312 596442 675340 598606
rect 675404 598264 675432 598674
rect 675496 598602 675524 598808
rect 675484 598596 675536 598602
rect 675484 598538 675536 598544
rect 675404 597174 675432 597652
rect 675392 597168 675444 597174
rect 675392 597110 675444 597116
rect 675312 596414 675418 596442
rect 675220 596278 675340 596306
rect 675208 595468 675260 595474
rect 675208 595410 675260 595416
rect 675220 593230 675248 595410
rect 675312 593570 675340 596278
rect 675404 595338 675432 595816
rect 675392 595332 675444 595338
rect 675392 595274 675444 595280
rect 675300 593564 675352 593570
rect 675300 593506 675352 593512
rect 675404 593450 675432 593980
rect 675312 593422 675432 593450
rect 675208 593224 675260 593230
rect 675208 593166 675260 593172
rect 675312 593178 675340 593422
rect 675576 593224 675628 593230
rect 675312 593150 675432 593178
rect 675576 593166 675628 593172
rect 675300 589416 675352 589422
rect 675300 589358 675352 589364
rect 675208 583772 675260 583778
rect 675208 583714 675260 583720
rect 675116 576088 675168 576094
rect 675116 576030 675168 576036
rect 675220 574094 675248 583714
rect 675128 574066 675248 574094
rect 675128 559722 675156 574066
rect 675312 564466 675340 589358
rect 675404 568818 675432 593150
rect 675588 573345 675616 593166
rect 678980 592804 679032 592810
rect 678980 592746 679032 592752
rect 676126 580952 676182 580961
rect 676126 580887 676182 580896
rect 676140 579970 676168 580887
rect 676310 580544 676366 580553
rect 676310 580479 676366 580488
rect 676218 580136 676274 580145
rect 676218 580071 676220 580080
rect 676272 580071 676274 580080
rect 676220 580042 676272 580048
rect 676128 579964 676180 579970
rect 676128 579906 676180 579912
rect 676324 579834 676352 580479
rect 676312 579828 676364 579834
rect 676312 579770 676364 579776
rect 676218 579728 676274 579737
rect 676218 579663 676220 579672
rect 676272 579663 676274 579672
rect 676220 579634 676272 579640
rect 676036 579080 676088 579086
rect 676034 579048 676036 579057
rect 676088 579048 676090 579057
rect 676034 578983 676090 578992
rect 676218 578504 676274 578513
rect 676218 578439 676220 578448
rect 676272 578439 676274 578448
rect 676220 578410 676272 578416
rect 676126 578096 676182 578105
rect 676126 578031 676182 578040
rect 676140 576910 676168 578031
rect 676218 577280 676274 577289
rect 676218 577215 676274 577224
rect 676232 576978 676260 577215
rect 676220 576972 676272 576978
rect 676220 576914 676272 576920
rect 676128 576904 676180 576910
rect 676128 576846 676180 576852
rect 676036 576836 676088 576842
rect 676036 576778 676088 576784
rect 675944 576768 675996 576774
rect 675944 576710 675996 576716
rect 675956 575385 675984 576710
rect 676048 576201 676076 576778
rect 676034 576192 676090 576201
rect 676034 576127 676090 576136
rect 676036 576088 676088 576094
rect 676036 576030 676088 576036
rect 675942 575376 675998 575385
rect 675942 575311 675998 575320
rect 676048 574569 676076 576030
rect 678992 575249 679020 592746
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 678978 575240 679034 575249
rect 678978 575175 679034 575184
rect 676034 574560 676090 574569
rect 676034 574495 676090 574504
rect 676036 573708 676088 573714
rect 676036 573650 676088 573656
rect 675574 573336 675630 573345
rect 675574 573271 675630 573280
rect 676048 572937 676076 573650
rect 676034 572928 676090 572937
rect 676034 572863 676090 572872
rect 676036 572824 676088 572830
rect 676036 572766 676088 572772
rect 676048 572529 676076 572766
rect 676034 572520 676090 572529
rect 676034 572455 676090 572464
rect 676036 572416 676088 572422
rect 676036 572358 676088 572364
rect 676048 572121 676076 572358
rect 676034 572112 676090 572121
rect 676034 572047 676090 572056
rect 678978 570752 679034 570761
rect 678978 570687 679034 570696
rect 678992 569945 679020 570687
rect 678978 569936 679034 569945
rect 678978 569871 679034 569880
rect 675392 568812 675444 568818
rect 675392 568754 675444 568760
rect 675392 568676 675444 568682
rect 675392 568618 675444 568624
rect 675300 564460 675352 564466
rect 675300 564402 675352 564408
rect 675404 563448 675432 568618
rect 678992 568614 679020 569871
rect 678980 568608 679032 568614
rect 678980 568550 679032 568556
rect 675496 562737 675524 562904
rect 675482 562728 675538 562737
rect 675482 562663 675538 562672
rect 675298 562320 675354 562329
rect 675354 562278 675418 562306
rect 675298 562255 675354 562264
rect 675496 561241 675524 561612
rect 675482 561232 675538 561241
rect 675482 561167 675538 561176
rect 675128 559694 675248 559722
rect 675024 559564 675076 559570
rect 675024 559506 675076 559512
rect 675036 545154 675064 559506
rect 675116 557592 675168 557598
rect 675116 557534 675168 557540
rect 675128 553518 675156 557534
rect 675116 553512 675168 553518
rect 675116 553454 675168 553460
rect 675116 553376 675168 553382
rect 675116 553318 675168 553324
rect 675024 545148 675076 545154
rect 675024 545090 675076 545096
rect 675128 544898 675156 553318
rect 675036 544870 675156 544898
rect 674932 532840 674984 532846
rect 674932 532782 674984 532788
rect 674840 485784 674892 485790
rect 674840 485726 674892 485732
rect 674564 485716 674616 485722
rect 674564 485658 674616 485664
rect 675036 485518 675064 544870
rect 675116 544808 675168 544814
rect 675116 544750 675168 544756
rect 675128 486033 675156 544750
rect 675220 532778 675248 559694
rect 675496 559570 675524 559776
rect 675484 559564 675536 559570
rect 675484 559506 675536 559512
rect 675312 559218 675418 559246
rect 675312 558074 675340 559218
rect 675404 558278 675432 558620
rect 675392 558272 675444 558278
rect 675392 558214 675444 558220
rect 675300 558068 675352 558074
rect 675300 558010 675352 558016
rect 675312 557926 675418 557954
rect 675312 554985 675340 557926
rect 675404 555286 675432 555492
rect 675392 555280 675444 555286
rect 675392 555222 675444 555228
rect 675298 554976 675354 554985
rect 675298 554911 675354 554920
rect 675300 554804 675352 554810
rect 675300 554746 675352 554752
rect 675312 551253 675340 554746
rect 675404 554606 675432 554919
rect 675392 554600 675444 554606
rect 675392 554542 675444 554548
rect 675496 553790 675524 554268
rect 675576 553852 675628 553858
rect 675576 553794 675628 553800
rect 675484 553784 675536 553790
rect 675484 553726 675536 553732
rect 675588 553656 675616 553794
rect 675392 553512 675444 553518
rect 675392 553454 675444 553460
rect 675404 553079 675432 553454
rect 675404 551954 675432 552432
rect 675392 551948 675444 551954
rect 675392 551890 675444 551896
rect 675312 551225 675418 551253
rect 675312 550582 675418 550610
rect 675312 548894 675340 550582
rect 675300 548888 675352 548894
rect 675300 548830 675352 548836
rect 675312 548746 675418 548774
rect 675312 542162 675340 548746
rect 675392 548004 675444 548010
rect 675392 547946 675444 547952
rect 675404 543726 675432 547946
rect 677600 547664 677652 547670
rect 677600 547606 677652 547612
rect 677506 546544 677562 546553
rect 677506 546479 677562 546488
rect 675576 545284 675628 545290
rect 675576 545226 675628 545232
rect 675392 543720 675444 543726
rect 675392 543662 675444 543668
rect 675300 542156 675352 542162
rect 675300 542098 675352 542104
rect 675208 532772 675260 532778
rect 675208 532714 675260 532720
rect 675484 492584 675536 492590
rect 675484 492526 675536 492532
rect 675392 492380 675444 492386
rect 675392 492322 675444 492328
rect 675404 489297 675432 492322
rect 675390 489288 675446 489297
rect 675390 489223 675446 489232
rect 675404 489216 675432 489223
rect 675496 487257 675524 492526
rect 675482 487248 675538 487257
rect 675482 487183 675538 487192
rect 675114 486024 675170 486033
rect 675114 485959 675170 485968
rect 675024 485512 675076 485518
rect 675024 485454 675076 485460
rect 675588 484809 675616 545226
rect 675942 543348 675998 543357
rect 675942 543283 675998 543292
rect 675956 539625 675984 543283
rect 675942 539616 675998 539625
rect 675942 539551 675998 539560
rect 676218 535936 676274 535945
rect 676218 535871 676274 535880
rect 676036 535764 676088 535770
rect 676034 535732 676036 535741
rect 676088 535732 676090 535741
rect 676034 535667 676090 535676
rect 676232 535634 676260 535871
rect 676220 535628 676272 535634
rect 676220 535570 676272 535576
rect 675850 534508 675906 534517
rect 675850 534443 675906 534452
rect 675760 529848 675812 529854
rect 675760 529790 675812 529796
rect 675772 528397 675800 529790
rect 675758 528388 675814 528397
rect 675758 528323 675814 528332
rect 675864 496814 675892 534443
rect 676036 534132 676088 534138
rect 676034 534100 676036 534109
rect 676088 534100 676090 534109
rect 676034 534035 676090 534044
rect 677414 533488 677470 533497
rect 677414 533423 677470 533432
rect 676034 532808 676090 532817
rect 676034 532743 676090 532752
rect 676220 532772 676272 532778
rect 675942 532060 675998 532069
rect 675942 531995 675998 532004
rect 675772 496786 675892 496814
rect 675772 491609 675800 496786
rect 675852 493400 675904 493406
rect 675852 493342 675904 493348
rect 675758 491600 675814 491609
rect 675758 491535 675814 491544
rect 675758 491464 675814 491473
rect 675758 491399 675814 491408
rect 675666 491328 675722 491337
rect 675666 491263 675722 491272
rect 675680 487665 675708 491263
rect 675666 487656 675722 487665
rect 675666 487591 675722 487600
rect 675772 486849 675800 491399
rect 675758 486840 675814 486849
rect 675758 486775 675814 486784
rect 675864 486441 675892 493342
rect 675956 492266 675984 531995
rect 676048 531661 676076 532743
rect 676220 532714 676272 532720
rect 676126 532672 676182 532681
rect 676126 532607 676182 532616
rect 676034 531652 676090 531661
rect 676034 531587 676090 531596
rect 676036 529916 676088 529922
rect 676036 529858 676088 529864
rect 676048 527989 676076 529858
rect 676034 527980 676090 527989
rect 676034 527915 676090 527924
rect 676036 527128 676088 527134
rect 676036 527070 676088 527076
rect 676048 526357 676076 527070
rect 676034 526348 676090 526357
rect 676034 526283 676090 526292
rect 676140 516134 676168 532607
rect 676232 531457 676260 532714
rect 676218 531448 676274 531457
rect 676218 531383 676274 531392
rect 676048 516106 676168 516134
rect 676048 492386 676076 516106
rect 676036 492380 676088 492386
rect 676036 492322 676088 492328
rect 675956 492238 676168 492266
rect 675942 492144 675998 492153
rect 675942 492079 675998 492088
rect 675956 491434 675984 492079
rect 676034 491736 676090 491745
rect 676034 491671 676036 491680
rect 676088 491671 676090 491680
rect 676036 491642 676088 491648
rect 676036 491564 676088 491570
rect 676036 491506 676088 491512
rect 675944 491428 675996 491434
rect 675944 491370 675996 491376
rect 676048 491337 676076 491506
rect 676034 491328 676090 491337
rect 676034 491263 676090 491272
rect 676140 491178 676168 492238
rect 677428 491298 677456 533423
rect 677520 527377 677548 546479
rect 677612 527785 677640 547606
rect 679440 543720 679492 543726
rect 679162 543688 679218 543697
rect 679440 543662 679492 543668
rect 679162 543623 679218 543632
rect 678978 535120 679034 535129
rect 678978 535055 679034 535064
rect 678992 532914 679020 535055
rect 679070 533080 679126 533089
rect 679070 533015 679126 533024
rect 678980 532908 679032 532914
rect 678980 532850 679032 532856
rect 678980 532772 679032 532778
rect 678980 532714 679032 532720
rect 678992 530233 679020 532714
rect 679084 530641 679112 533015
rect 679070 530632 679126 530641
rect 679070 530567 679126 530576
rect 678978 530224 679034 530233
rect 678978 530159 679034 530168
rect 679176 529009 679204 543623
rect 679346 543552 679402 543561
rect 679346 543487 679402 543496
rect 679254 533896 679310 533905
rect 679254 533831 679310 533840
rect 679268 531049 679296 533831
rect 679254 531040 679310 531049
rect 679254 530975 679310 530984
rect 679360 529417 679388 543487
rect 679452 529825 679480 543662
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 679438 529816 679494 529825
rect 679438 529751 679494 529760
rect 679346 529408 679402 529417
rect 679346 529343 679402 529352
rect 679162 529000 679218 529009
rect 679162 528935 679218 528944
rect 677598 527776 677654 527785
rect 677598 527711 677654 527720
rect 677506 527368 677562 527377
rect 677506 527303 677562 527312
rect 678978 525736 679034 525745
rect 678978 525671 679034 525680
rect 678992 524929 679020 525671
rect 678978 524920 679034 524929
rect 678978 524855 679034 524864
rect 678992 524482 679020 524855
rect 678980 524476 679032 524482
rect 678980 524418 679032 524424
rect 703694 492796 703722 492932
rect 704154 492796 704182 492932
rect 704614 492796 704642 492932
rect 705074 492796 705102 492932
rect 705534 492796 705562 492932
rect 705994 492796 706022 492932
rect 706454 492796 706482 492932
rect 706914 492796 706942 492932
rect 707374 492796 707402 492932
rect 707834 492796 707862 492932
rect 708294 492796 708322 492932
rect 708754 492796 708782 492932
rect 709214 492796 709242 492932
rect 676220 491292 676272 491298
rect 676220 491234 676272 491240
rect 677416 491292 677468 491298
rect 677416 491234 677468 491240
rect 675956 491150 676168 491178
rect 675956 488481 675984 491150
rect 676034 490104 676090 490113
rect 676232 490090 676260 491234
rect 679438 490512 679494 490521
rect 679438 490447 679494 490456
rect 676090 490062 676260 490090
rect 676034 490039 676090 490048
rect 676034 489696 676090 489705
rect 676090 489654 676260 489682
rect 676034 489631 676090 489640
rect 676232 488578 676260 489654
rect 676220 488572 676272 488578
rect 676220 488514 676272 488520
rect 677488 488572 677540 488578
rect 677488 488514 677540 488520
rect 675942 488472 675998 488481
rect 675942 488407 675998 488416
rect 675956 488388 675984 488407
rect 675850 486432 675906 486441
rect 675850 486367 675906 486376
rect 676036 485784 676088 485790
rect 676036 485726 676088 485732
rect 675944 485716 675996 485722
rect 675944 485658 675996 485664
rect 675852 485648 675904 485654
rect 675852 485590 675904 485596
rect 675574 484800 675630 484809
rect 675574 484735 675630 484744
rect 675864 484401 675892 485590
rect 675850 484392 675906 484401
rect 675850 484327 675906 484336
rect 675956 483993 675984 485658
rect 676048 485625 676076 485726
rect 676034 485616 676090 485625
rect 676034 485551 676090 485560
rect 676036 485512 676088 485518
rect 676036 485454 676088 485460
rect 675942 483984 675998 483993
rect 675942 483919 675998 483928
rect 676048 483585 676076 485454
rect 676034 483576 676090 483585
rect 676034 483511 676090 483520
rect 676036 483472 676088 483478
rect 676036 483414 676088 483420
rect 676048 483177 676076 483414
rect 676034 483168 676090 483177
rect 676034 483103 676090 483112
rect 674288 482996 674340 483002
rect 674288 482938 674340 482944
rect 676036 482996 676088 483002
rect 676036 482938 676088 482944
rect 673736 482928 673788 482934
rect 673736 482870 673788 482876
rect 675944 482928 675996 482934
rect 675944 482870 675996 482876
rect 675956 482769 675984 482870
rect 675942 482760 675998 482769
rect 675942 482695 675998 482704
rect 676048 482361 676076 482938
rect 676034 482352 676090 482361
rect 676034 482287 676090 482296
rect 676034 481944 676090 481953
rect 676034 481879 676090 481888
rect 676048 480758 676076 481879
rect 672540 480752 672592 480758
rect 676036 480752 676088 480758
rect 672540 480694 672592 480700
rect 676034 480720 676036 480729
rect 676088 480720 676090 480729
rect 672446 153368 672502 153377
rect 672446 153303 672502 153312
rect 672552 148209 672580 480694
rect 676034 480655 676090 480664
rect 676048 480629 676076 480655
rect 676128 475448 676180 475454
rect 676128 475390 676180 475396
rect 676036 475260 676088 475266
rect 676036 475202 676088 475208
rect 675944 475068 675996 475074
rect 675944 475010 675996 475016
rect 675850 403064 675906 403073
rect 675850 402999 675852 403008
rect 675904 402999 675906 403008
rect 675852 402970 675904 402976
rect 675956 402665 675984 475010
rect 675942 402656 675998 402665
rect 675942 402591 675998 402600
rect 675298 401432 675354 401441
rect 675298 401367 675354 401376
rect 674472 398268 674524 398274
rect 674472 398210 674524 398216
rect 673736 397588 673788 397594
rect 673736 397530 673788 397536
rect 673460 395412 673512 395418
rect 673460 395354 673512 395360
rect 672816 392080 672868 392086
rect 672816 392022 672868 392028
rect 672632 256828 672684 256834
rect 672632 256770 672684 256776
rect 672538 148200 672594 148209
rect 672538 148135 672594 148144
rect 672172 131708 672224 131714
rect 672172 131650 672224 131656
rect 672080 130076 672132 130082
rect 672080 130018 672132 130024
rect 671986 114336 672042 114345
rect 671986 114271 672042 114280
rect 666926 107536 666982 107545
rect 666926 107471 666982 107480
rect 672092 100881 672120 130018
rect 672184 104145 672212 131650
rect 672264 130892 672316 130898
rect 672264 130834 672316 130840
rect 672276 105913 672304 130834
rect 672356 129464 672408 129470
rect 672356 129406 672408 129412
rect 672262 105904 672318 105913
rect 672262 105839 672318 105848
rect 672170 104136 672226 104145
rect 672170 104071 672226 104080
rect 672368 102513 672396 129406
rect 672644 127945 672672 256770
rect 672724 212084 672776 212090
rect 672724 212026 672776 212032
rect 672630 127936 672686 127945
rect 672630 127871 672686 127880
rect 672736 122913 672764 212026
rect 672828 143177 672856 392022
rect 673368 386028 673420 386034
rect 673368 385970 673420 385976
rect 673380 384742 673408 385970
rect 673368 384736 673420 384742
rect 673368 384678 673420 384684
rect 673472 375766 673500 395354
rect 673552 394936 673604 394942
rect 673552 394878 673604 394884
rect 673564 377466 673592 394878
rect 673644 394188 673696 394194
rect 673644 394130 673696 394136
rect 673656 384826 673684 394130
rect 673748 385014 673776 397530
rect 674288 397044 674340 397050
rect 674288 396986 674340 396992
rect 673828 392012 673880 392018
rect 673828 391954 673880 391960
rect 673736 385008 673788 385014
rect 673736 384950 673788 384956
rect 673656 384798 673776 384826
rect 673644 384736 673696 384742
rect 673644 384678 673696 384684
rect 673656 378826 673684 384678
rect 673644 378820 673696 378826
rect 673644 378762 673696 378768
rect 673748 378214 673776 384798
rect 673736 378208 673788 378214
rect 673736 378150 673788 378156
rect 673552 377460 673604 377466
rect 673552 377402 673604 377408
rect 673840 376990 673868 391954
rect 674300 381206 674328 396986
rect 674484 384810 674512 398210
rect 674564 397656 674616 397662
rect 674564 397598 674616 397604
rect 674576 386034 674604 397598
rect 674656 397520 674708 397526
rect 674656 397462 674708 397468
rect 674564 386028 674616 386034
rect 674564 385970 674616 385976
rect 674564 385892 674616 385898
rect 674564 385834 674616 385840
rect 674472 384804 674524 384810
rect 674472 384746 674524 384752
rect 674288 381200 674340 381206
rect 674288 381142 674340 381148
rect 673828 376984 673880 376990
rect 673828 376926 673880 376932
rect 673460 375760 673512 375766
rect 673460 375702 673512 375708
rect 674576 372570 674604 385834
rect 674668 383178 674696 397462
rect 674840 395004 674892 395010
rect 674840 394946 674892 394952
rect 674656 383172 674708 383178
rect 674656 383114 674708 383120
rect 674852 381954 674880 394946
rect 675024 394868 675076 394874
rect 675024 394810 675076 394816
rect 675036 382498 675064 394810
rect 675116 394800 675168 394806
rect 675116 394742 675168 394748
rect 675024 382492 675076 382498
rect 675024 382434 675076 382440
rect 674840 381948 674892 381954
rect 674840 381890 674892 381896
rect 675128 381342 675156 394742
rect 675208 394732 675260 394738
rect 675208 394674 675260 394680
rect 675220 385626 675248 394674
rect 675208 385620 675260 385626
rect 675208 385562 675260 385568
rect 675208 385008 675260 385014
rect 675208 384950 675260 384956
rect 675116 381336 675168 381342
rect 675116 381278 675168 381284
rect 675116 381200 675168 381206
rect 675116 381142 675168 381148
rect 675024 373516 675076 373522
rect 675024 373458 675076 373464
rect 674564 372564 674616 372570
rect 674564 372506 674616 372512
rect 675036 361574 675064 373458
rect 675128 371566 675156 381142
rect 675220 373266 675248 384950
rect 675312 373522 675340 401367
rect 676048 401033 676076 475202
rect 676034 401024 676090 401033
rect 676034 400959 676090 400968
rect 676048 400944 676076 400959
rect 676034 400214 676090 400217
rect 676140 400214 676168 475390
rect 676310 403744 676366 403753
rect 676310 403679 676366 403688
rect 676218 403336 676274 403345
rect 676218 403271 676274 403280
rect 676232 403170 676260 403271
rect 676220 403164 676272 403170
rect 676220 403106 676272 403112
rect 676324 403102 676352 403679
rect 676312 403096 676364 403102
rect 676312 403038 676364 403044
rect 677500 402121 677528 488514
rect 679162 488064 679218 488073
rect 679162 487999 679218 488008
rect 679176 475454 679204 487999
rect 679166 475448 679218 475454
rect 679166 475390 679218 475396
rect 679452 475074 679480 490447
rect 679622 488880 679678 488889
rect 679622 488815 679678 488824
rect 679636 475266 679664 488815
rect 679624 475260 679676 475266
rect 679624 475202 679676 475208
rect 679440 475068 679492 475074
rect 679440 475010 679492 475016
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 677486 402112 677542 402121
rect 677486 402047 677542 402056
rect 676034 400208 676168 400214
rect 676090 400186 676168 400208
rect 676034 400143 676090 400152
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 675758 398576 675814 398585
rect 675758 398511 675814 398520
rect 675772 386646 675800 398511
rect 676048 398274 676076 399327
rect 676126 398848 676182 398857
rect 676126 398783 676182 398792
rect 676036 398268 676088 398274
rect 676036 398210 676088 398216
rect 676034 398168 676090 398177
rect 676034 398103 676090 398112
rect 675942 397760 675998 397769
rect 675942 397695 675998 397704
rect 675956 397662 675984 397695
rect 675944 397656 675996 397662
rect 675944 397598 675996 397604
rect 676048 397526 676076 398103
rect 676140 397594 676168 398783
rect 676128 397588 676180 397594
rect 676128 397530 676180 397536
rect 676036 397520 676088 397526
rect 676036 397462 676088 397468
rect 676034 397352 676090 397361
rect 676034 397287 676090 397296
rect 676048 397050 676076 397287
rect 676036 397044 676088 397050
rect 676036 396986 676088 396992
rect 676034 396944 676090 396953
rect 676034 396879 676090 396888
rect 675942 396128 675998 396137
rect 675942 396063 675998 396072
rect 675850 395720 675906 395729
rect 675850 395655 675906 395664
rect 675864 395418 675892 395655
rect 675852 395412 675904 395418
rect 675852 395354 675904 395360
rect 675850 395312 675906 395321
rect 675850 395247 675906 395256
rect 675864 394942 675892 395247
rect 675956 395010 675984 396063
rect 675944 395004 675996 395010
rect 675944 394946 675996 394952
rect 675852 394936 675904 394942
rect 675852 394878 675904 394884
rect 675942 394904 675998 394913
rect 675942 394839 675998 394848
rect 675956 394806 675984 394839
rect 675944 394800 675996 394806
rect 675944 394742 675996 394748
rect 676048 394738 676076 396879
rect 676126 396400 676182 396409
rect 676126 396335 676182 396344
rect 676140 394874 676168 396335
rect 676128 394868 676180 394874
rect 676128 394810 676180 394816
rect 676036 394732 676088 394738
rect 676036 394674 676088 394680
rect 676034 394496 676090 394505
rect 676034 394431 676090 394440
rect 676048 394194 676076 394431
rect 676036 394188 676088 394194
rect 676036 394130 676088 394136
rect 676034 394088 676090 394097
rect 676034 394023 676090 394032
rect 676048 392018 676076 394023
rect 678978 393544 679034 393553
rect 678978 393479 679034 393488
rect 678992 392737 679020 393479
rect 678978 392728 679034 392737
rect 678978 392663 679034 392672
rect 678992 392086 679020 392663
rect 678980 392080 679032 392086
rect 678980 392022 679032 392028
rect 676036 392012 676088 392018
rect 676036 391954 676088 391960
rect 675760 386640 675812 386646
rect 675760 386582 675812 386588
rect 675404 386034 675432 386275
rect 675392 386028 675444 386034
rect 675392 385970 675444 385976
rect 675760 386028 675812 386034
rect 675760 385970 675812 385976
rect 675772 385696 675800 385970
rect 675392 385620 675444 385626
rect 675392 385562 675444 385568
rect 675404 385084 675432 385562
rect 675392 384804 675444 384810
rect 675392 384746 675444 384752
rect 675404 384435 675432 384746
rect 675392 383172 675444 383178
rect 675392 383114 675444 383120
rect 675404 382568 675432 383114
rect 675392 382492 675444 382498
rect 675392 382434 675444 382440
rect 675404 382024 675432 382434
rect 675392 381948 675444 381954
rect 675392 381890 675444 381896
rect 675404 381412 675432 381890
rect 675392 381336 675444 381342
rect 675392 381278 675444 381284
rect 675404 380732 675432 381278
rect 675392 378820 675444 378826
rect 675392 378762 675444 378768
rect 675404 378284 675432 378762
rect 675484 378208 675536 378214
rect 675484 378150 675536 378156
rect 675496 377740 675524 378150
rect 675392 377460 675444 377466
rect 675392 377402 675444 377408
rect 675404 377060 675432 377402
rect 675484 376984 675536 376990
rect 675484 376926 675536 376932
rect 675496 376448 675524 376926
rect 675392 375760 675444 375766
rect 675392 375702 675444 375708
rect 675404 375224 675432 375702
rect 675300 373516 675352 373522
rect 675300 373458 675352 373464
rect 675404 373266 675432 373388
rect 675220 373238 675432 373266
rect 675220 371606 675432 371634
rect 675220 371566 675248 371606
rect 675128 371538 675248 371566
rect 675404 371552 675432 371606
rect 675036 361546 675800 361574
rect 675666 357096 675722 357105
rect 673092 357060 673144 357066
rect 675666 357031 675668 357040
rect 673092 357002 673144 357008
rect 675720 357031 675722 357040
rect 675668 357002 675720 357008
rect 672908 347268 672960 347274
rect 672908 347210 672960 347216
rect 672814 143168 672870 143177
rect 672814 143103 672870 143112
rect 672920 138465 672948 347210
rect 673104 312458 673132 357002
rect 675772 356697 675800 361546
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 675850 358728 675906 358737
rect 675850 358663 675906 358672
rect 675758 356688 675814 356697
rect 675758 356623 675814 356632
rect 675864 356250 675892 358663
rect 675942 358320 675998 358329
rect 675942 358255 675998 358264
rect 675956 356522 675984 358255
rect 676034 357912 676090 357921
rect 676034 357847 676090 357856
rect 675944 356516 675996 356522
rect 675944 356458 675996 356464
rect 676048 356386 676076 357847
rect 676036 356380 676088 356386
rect 676036 356322 676088 356328
rect 676034 356280 676090 356289
rect 675852 356244 675904 356250
rect 676034 356215 676090 356224
rect 675852 356186 675904 356192
rect 676048 356182 676076 356215
rect 673368 356176 673420 356182
rect 673368 356118 673420 356124
rect 676036 356176 676088 356182
rect 676036 356118 676088 356124
rect 673184 355428 673236 355434
rect 673184 355370 673236 355376
rect 673092 312452 673144 312458
rect 673092 312394 673144 312400
rect 673104 312392 673132 312394
rect 673196 310690 673224 355370
rect 673276 354612 673328 354618
rect 673276 354554 673328 354560
rect 673184 310684 673236 310690
rect 673184 310626 673236 310632
rect 673196 310624 673224 310626
rect 673288 309874 673316 354554
rect 673380 311710 673408 356118
rect 676034 355464 676090 355473
rect 676034 355399 676036 355408
rect 676088 355399 676090 355408
rect 676036 355370 676088 355376
rect 676034 354648 676090 354657
rect 676034 354583 676036 354592
rect 676088 354583 676090 354592
rect 676036 354554 676088 354560
rect 676034 354240 676090 354249
rect 676034 354175 676090 354184
rect 675390 353832 675446 353841
rect 675390 353767 675446 353776
rect 674656 353524 674708 353530
rect 674656 353466 674708 353472
rect 673736 351076 673788 351082
rect 673736 351018 673788 351024
rect 673552 350872 673604 350878
rect 673552 350814 673604 350820
rect 673460 350736 673512 350742
rect 673460 350678 673512 350684
rect 673472 331158 673500 350678
rect 673460 331152 673512 331158
rect 673460 331094 673512 331100
rect 673564 326942 673592 350814
rect 673644 347948 673696 347954
rect 673644 347890 673696 347896
rect 673656 331770 673684 347890
rect 673748 335442 673776 351018
rect 674564 350668 674616 350674
rect 674564 350610 674616 350616
rect 674288 349852 674340 349858
rect 674288 349794 674340 349800
rect 674300 341834 674328 349794
rect 674472 347880 674524 347886
rect 674472 347822 674524 347828
rect 673828 341828 673880 341834
rect 673828 341770 673880 341776
rect 674288 341828 674340 341834
rect 674288 341770 674340 341776
rect 673736 335436 673788 335442
rect 673736 335378 673788 335384
rect 673840 332450 673868 341770
rect 674484 341698 674512 347822
rect 674288 341692 674340 341698
rect 674288 341634 674340 341640
rect 674472 341692 674524 341698
rect 674472 341634 674524 341640
rect 674300 335510 674328 341634
rect 674576 341578 674604 350610
rect 674484 341550 674604 341578
rect 674484 336734 674512 341550
rect 674564 341420 674616 341426
rect 674564 341362 674616 341368
rect 674472 336728 674524 336734
rect 674472 336670 674524 336676
rect 674288 335504 674340 335510
rect 674288 335446 674340 335452
rect 673828 332444 673880 332450
rect 673828 332386 673880 332392
rect 673644 331764 673696 331770
rect 673644 331706 673696 331712
rect 674576 328778 674604 341362
rect 674668 339590 674696 353466
rect 675116 353320 675168 353326
rect 675116 353262 675168 353268
rect 674840 351484 674892 351490
rect 674840 351426 674892 351432
rect 674656 339584 674708 339590
rect 674656 339526 674708 339532
rect 674852 337958 674880 351426
rect 675024 347812 675076 347818
rect 675024 347754 675076 347760
rect 675036 340814 675064 347754
rect 675128 340882 675156 353262
rect 675298 351792 675354 351801
rect 675298 351727 675354 351736
rect 675208 350600 675260 350606
rect 675208 350542 675260 350548
rect 675116 340876 675168 340882
rect 675116 340818 675168 340824
rect 675024 340808 675076 340814
rect 675024 340750 675076 340756
rect 675024 340672 675076 340678
rect 675024 340614 675076 340620
rect 674840 337952 674892 337958
rect 674840 337894 674892 337900
rect 675036 335374 675064 340614
rect 675116 340468 675168 340474
rect 675116 340410 675168 340416
rect 675128 335594 675156 340410
rect 675220 336857 675248 350542
rect 675312 339878 675340 351727
rect 675404 341426 675432 353767
rect 676048 353530 676076 354175
rect 676036 353524 676088 353530
rect 676036 353466 676088 353472
rect 676034 353424 676090 353433
rect 676034 353359 676090 353368
rect 676048 353326 676076 353359
rect 676036 353320 676088 353326
rect 676036 353262 676088 353268
rect 676034 353016 676090 353025
rect 676034 352951 676090 352960
rect 675942 352608 675998 352617
rect 675942 352543 675998 352552
rect 675850 352200 675906 352209
rect 675850 352135 675906 352144
rect 675864 350878 675892 352135
rect 675956 351082 675984 352543
rect 676048 351490 676076 352951
rect 676036 351484 676088 351490
rect 676036 351426 676088 351432
rect 676034 351384 676090 351393
rect 676034 351319 676090 351328
rect 675944 351076 675996 351082
rect 675944 351018 675996 351024
rect 675942 350976 675998 350985
rect 675942 350911 675998 350920
rect 675852 350872 675904 350878
rect 675852 350814 675904 350820
rect 675852 350736 675904 350742
rect 675852 350678 675904 350684
rect 675864 350577 675892 350678
rect 675956 350674 675984 350911
rect 675944 350668 675996 350674
rect 675944 350610 675996 350616
rect 676048 350606 676076 351319
rect 676036 350600 676088 350606
rect 675850 350568 675906 350577
rect 676036 350542 676088 350548
rect 675850 350503 675906 350512
rect 676034 350160 676090 350169
rect 676034 350095 676090 350104
rect 676048 349858 676076 350095
rect 676036 349852 676088 349858
rect 676036 349794 676088 349800
rect 676034 349752 676090 349761
rect 676034 349687 676090 349696
rect 675942 349344 675998 349353
rect 675942 349279 675998 349288
rect 675850 348936 675906 348945
rect 675850 348871 675906 348880
rect 675864 347954 675892 348871
rect 675852 347948 675904 347954
rect 675852 347890 675904 347896
rect 675956 347886 675984 349279
rect 675944 347880 675996 347886
rect 675944 347822 675996 347828
rect 676048 347818 676076 349687
rect 676036 347812 676088 347818
rect 676036 347754 676088 347760
rect 676034 347304 676090 347313
rect 676034 347239 676036 347248
rect 676088 347239 676090 347248
rect 676036 347210 676088 347216
rect 675392 341420 675444 341426
rect 675392 341362 675444 341368
rect 675404 340678 675432 341088
rect 675484 340808 675536 340814
rect 675484 340750 675536 340756
rect 675392 340672 675444 340678
rect 675392 340614 675444 340620
rect 675496 340544 675524 340750
rect 675312 339850 675418 339878
rect 675484 339584 675536 339590
rect 675484 339526 675536 339532
rect 675496 339252 675524 339526
rect 675484 337952 675536 337958
rect 675484 337894 675536 337900
rect 675496 337416 675524 337894
rect 675220 336829 675418 336857
rect 675208 336728 675260 336734
rect 675208 336670 675260 336676
rect 675220 336206 675248 336670
rect 675220 336178 675418 336206
rect 675128 335566 675340 335594
rect 675116 335504 675168 335510
rect 675116 335446 675168 335452
rect 675312 335458 675340 335566
rect 675404 335458 675432 335580
rect 675024 335368 675076 335374
rect 675024 335310 675076 335316
rect 675128 332534 675156 335446
rect 675208 335436 675260 335442
rect 675312 335430 675432 335458
rect 675208 335378 675260 335384
rect 675220 333078 675248 335378
rect 675220 333050 675418 333078
rect 675128 332506 675418 332534
rect 675116 332444 675168 332450
rect 675116 332386 675168 332392
rect 675128 331889 675156 332386
rect 675128 331861 675418 331889
rect 675116 331764 675168 331770
rect 675116 331706 675168 331712
rect 675128 331242 675156 331706
rect 675128 331214 675418 331242
rect 675116 331152 675168 331158
rect 675116 331094 675168 331100
rect 675128 330049 675156 331094
rect 675128 330021 675418 330049
rect 674564 328772 674616 328778
rect 674564 328714 674616 328720
rect 675392 328772 675444 328778
rect 675392 328714 675444 328720
rect 675404 328168 675432 328714
rect 673552 326936 673604 326942
rect 673552 326878 673604 326884
rect 675392 326936 675444 326942
rect 675392 326878 675444 326884
rect 675404 326332 675432 326878
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676310 313576 676366 313585
rect 676310 313511 676366 313520
rect 676126 313168 676182 313177
rect 676126 313103 676182 313112
rect 676034 312488 676090 312497
rect 676034 312423 676036 312432
rect 676088 312423 676090 312432
rect 676036 312394 676088 312400
rect 676140 311982 676168 313103
rect 676218 312760 676274 312769
rect 676218 312695 676274 312704
rect 676232 312186 676260 312695
rect 676220 312180 676272 312186
rect 676220 312122 676272 312128
rect 676324 312050 676352 313511
rect 676312 312044 676364 312050
rect 676312 311986 676364 311992
rect 676128 311976 676180 311982
rect 676128 311918 676180 311924
rect 676218 311944 676274 311953
rect 676218 311879 676220 311888
rect 676272 311879 676274 311888
rect 676220 311850 676272 311856
rect 673368 311704 673420 311710
rect 676036 311704 676088 311710
rect 673368 311646 673420 311652
rect 676034 311672 676036 311681
rect 676088 311672 676090 311681
rect 676034 311607 676090 311616
rect 676218 311128 676274 311137
rect 673368 311092 673420 311098
rect 676218 311063 676220 311072
rect 673368 311034 673420 311040
rect 676272 311063 676274 311072
rect 676220 311034 676272 311040
rect 673276 309868 673328 309874
rect 673276 309810 673328 309816
rect 673000 300892 673052 300898
rect 673000 300834 673052 300840
rect 672906 138456 672962 138465
rect 672906 138391 672962 138400
rect 673012 132977 673040 300834
rect 673380 266694 673408 311034
rect 676218 310720 676274 310729
rect 676218 310655 676220 310664
rect 676272 310655 676274 310664
rect 676220 310626 676272 310632
rect 676218 310312 676274 310321
rect 676218 310247 676220 310256
rect 676272 310247 676274 310256
rect 676220 310218 676272 310224
rect 676218 309904 676274 309913
rect 676218 309839 676220 309848
rect 676272 309839 676274 309848
rect 676220 309810 676272 309816
rect 676218 309496 676274 309505
rect 676218 309431 676220 309440
rect 676272 309431 676274 309440
rect 676220 309402 676272 309408
rect 676034 309224 676090 309233
rect 674656 309188 674708 309194
rect 676034 309159 676036 309168
rect 674656 309130 674708 309136
rect 676088 309159 676090 309168
rect 676036 309130 676088 309136
rect 673460 308100 673512 308106
rect 673460 308042 673512 308048
rect 673472 286822 673500 308042
rect 674472 306876 674524 306882
rect 674472 306818 674524 306824
rect 673552 306400 673604 306406
rect 673552 306342 673604 306348
rect 673564 288658 673592 306342
rect 673644 305108 673696 305114
rect 673644 305050 673696 305056
rect 673552 288652 673604 288658
rect 673552 288594 673604 288600
rect 673460 286816 673512 286822
rect 673460 286758 673512 286764
rect 673656 286754 673684 305050
rect 673828 304360 673880 304366
rect 673828 304302 673880 304308
rect 673736 303748 673788 303754
rect 673736 303690 673788 303696
rect 673644 286748 673696 286754
rect 673644 286690 673696 286696
rect 673460 286680 673512 286686
rect 673460 286622 673512 286628
rect 673472 282878 673500 286622
rect 673748 286618 673776 303690
rect 673840 287434 673868 304302
rect 674288 303952 674340 303958
rect 674288 303894 674340 303900
rect 674300 290494 674328 303894
rect 674484 294166 674512 306818
rect 674564 306468 674616 306474
rect 674564 306410 674616 306416
rect 674576 295254 674604 306410
rect 674668 295458 674696 309130
rect 676034 308816 676090 308825
rect 676034 308751 676090 308760
rect 675298 308408 675354 308417
rect 675298 308343 675354 308352
rect 675208 306060 675260 306066
rect 675208 306002 675260 306008
rect 675024 304836 675076 304842
rect 675024 304778 675076 304784
rect 674840 304224 674892 304230
rect 674840 304166 674892 304172
rect 674656 295452 674708 295458
rect 674656 295394 674708 295400
rect 674564 295248 674616 295254
rect 674564 295190 674616 295196
rect 674472 294160 674524 294166
rect 674472 294102 674524 294108
rect 674564 293956 674616 293962
rect 674564 293898 674616 293904
rect 674288 290488 674340 290494
rect 674288 290430 674340 290436
rect 673828 287428 673880 287434
rect 673828 287370 673880 287376
rect 674576 286686 674604 293898
rect 674852 291310 674880 304166
rect 674840 291304 674892 291310
rect 674840 291246 674892 291252
rect 675036 291190 675064 304778
rect 675116 298308 675168 298314
rect 675116 298250 675168 298256
rect 675128 293962 675156 298250
rect 675116 293956 675168 293962
rect 675116 293898 675168 293904
rect 675220 291870 675248 306002
rect 675312 295542 675340 308343
rect 676048 308106 676076 308751
rect 676036 308100 676088 308106
rect 676036 308042 676088 308048
rect 676034 308000 676090 308009
rect 676034 307935 676090 307944
rect 675390 307184 675446 307193
rect 675390 307119 675446 307128
rect 675404 298314 675432 307119
rect 676048 306882 676076 307935
rect 676126 307456 676182 307465
rect 676126 307391 676182 307400
rect 676036 306876 676088 306882
rect 676036 306818 676088 306824
rect 676034 306776 676090 306785
rect 676034 306711 676090 306720
rect 676048 306474 676076 306711
rect 676036 306468 676088 306474
rect 676036 306410 676088 306416
rect 676140 306406 676168 307391
rect 676128 306400 676180 306406
rect 676034 306368 676090 306377
rect 676128 306342 676180 306348
rect 676034 306303 676090 306312
rect 676048 306066 676076 306303
rect 676036 306060 676088 306066
rect 676036 306002 676088 306008
rect 676034 305960 676090 305969
rect 676034 305895 676090 305904
rect 676048 304842 676076 305895
rect 676126 305416 676182 305425
rect 676126 305351 676182 305360
rect 676140 305114 676168 305351
rect 676128 305108 676180 305114
rect 676128 305050 676180 305056
rect 676126 305008 676182 305017
rect 676126 304943 676182 304952
rect 676036 304836 676088 304842
rect 676036 304778 676088 304784
rect 676034 304736 676090 304745
rect 676034 304671 676090 304680
rect 676048 304230 676076 304671
rect 676140 304366 676168 304943
rect 676128 304360 676180 304366
rect 676128 304302 676180 304308
rect 676036 304224 676088 304230
rect 676036 304166 676088 304172
rect 676126 304192 676182 304201
rect 676126 304127 676182 304136
rect 676140 303958 676168 304127
rect 676128 303952 676180 303958
rect 676034 303920 676090 303929
rect 676128 303894 676180 303900
rect 676034 303855 676090 303864
rect 676048 303754 676076 303855
rect 676036 303748 676088 303754
rect 676036 303690 676088 303696
rect 678978 303376 679034 303385
rect 678978 303311 679034 303320
rect 678992 302569 679020 303311
rect 678978 302560 679034 302569
rect 678978 302495 679034 302504
rect 678992 300898 679020 302495
rect 678980 300892 679032 300898
rect 678980 300834 679032 300840
rect 675392 298308 675444 298314
rect 675392 298250 675444 298256
rect 675392 298172 675444 298178
rect 675392 298114 675444 298120
rect 675404 296072 675432 298114
rect 675312 295514 675418 295542
rect 675300 295452 675352 295458
rect 675300 295394 675352 295400
rect 675312 294250 675340 295394
rect 675392 295248 675444 295254
rect 675392 295190 675444 295196
rect 675404 294879 675432 295190
rect 675312 294222 675418 294250
rect 675300 294160 675352 294166
rect 675300 294102 675352 294108
rect 675312 292414 675340 294102
rect 675312 292386 675418 292414
rect 675220 291842 675418 291870
rect 675312 291230 675432 291258
rect 675312 291190 675340 291230
rect 675036 291162 675340 291190
rect 675404 291176 675432 291230
rect 675116 291100 675168 291106
rect 675116 291042 675168 291048
rect 675128 290578 675156 291042
rect 675128 290550 675418 290578
rect 675116 290488 675168 290494
rect 675116 290430 675168 290436
rect 675128 287518 675156 290430
rect 675392 288652 675444 288658
rect 675392 288594 675444 288600
rect 675404 288048 675432 288594
rect 675128 287490 675418 287518
rect 675116 287428 675168 287434
rect 675116 287370 675168 287376
rect 675128 286906 675156 287370
rect 675128 286878 675340 286906
rect 675116 286816 675168 286822
rect 675116 286758 675168 286764
rect 675312 286770 675340 286878
rect 675404 286770 675432 286892
rect 674564 286680 674616 286686
rect 674564 286622 674616 286628
rect 673736 286612 673788 286618
rect 673736 286554 673788 286560
rect 675128 283234 675156 286758
rect 675208 286748 675260 286754
rect 675312 286742 675432 286770
rect 675208 286690 675260 286696
rect 675220 285070 675248 286690
rect 675392 286612 675444 286618
rect 675392 286554 675444 286560
rect 675404 286212 675432 286554
rect 675220 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675128 283206 675340 283234
rect 675312 283098 675340 283206
rect 675404 283098 675432 283220
rect 675312 283070 675432 283098
rect 673460 282872 673512 282878
rect 673460 282814 673512 282820
rect 675116 282872 675168 282878
rect 675116 282814 675168 282820
rect 675128 281369 675156 282814
rect 675128 281341 675418 281369
rect 678980 278384 679032 278390
rect 678980 278326 679032 278332
rect 676126 268560 676182 268569
rect 676126 268495 676182 268504
rect 676036 267980 676088 267986
rect 676036 267922 676088 267928
rect 676048 267889 676076 267922
rect 676034 267880 676090 267889
rect 676034 267815 676090 267824
rect 676140 267782 676168 268495
rect 676218 268152 676274 268161
rect 676218 268087 676220 268096
rect 676272 268087 676274 268096
rect 676220 268058 676272 268064
rect 676128 267776 676180 267782
rect 678992 267753 679020 278326
rect 679072 278316 679124 278322
rect 679072 278258 679124 278264
rect 676128 267718 676180 267724
rect 678978 267744 679034 267753
rect 678978 267679 679034 267688
rect 675680 267073 675708 267082
rect 675666 267064 675722 267073
rect 675666 266999 675722 267008
rect 673368 266688 673420 266694
rect 673368 266630 673420 266636
rect 675208 265600 675260 265606
rect 675208 265542 675260 265548
rect 675220 264974 675248 265542
rect 675680 264974 675708 266999
rect 676036 266688 676088 266694
rect 676034 266656 676036 266665
rect 676088 266656 676090 266665
rect 676034 266591 676090 266600
rect 676034 266248 676090 266257
rect 676034 266183 676090 266192
rect 676048 265606 676076 266183
rect 679084 266121 679112 278258
rect 679164 278112 679216 278118
rect 679164 278054 679216 278060
rect 679070 266112 679126 266121
rect 679070 266047 679126 266056
rect 676036 265600 676088 265606
rect 676036 265542 676088 265548
rect 675772 265441 675800 265454
rect 675758 265432 675814 265441
rect 675758 265367 675814 265376
rect 675128 264946 675248 264974
rect 675312 264946 675708 264974
rect 673828 263084 673880 263090
rect 673828 263026 673880 263032
rect 673460 262540 673512 262546
rect 673460 262482 673512 262488
rect 673472 252770 673500 262482
rect 673552 262336 673604 262342
rect 673552 262278 673604 262284
rect 673380 252742 673500 252770
rect 673564 252754 673592 262278
rect 673644 260228 673696 260234
rect 673644 260170 673696 260176
rect 673552 252748 673604 252754
rect 673380 249558 673408 252742
rect 673552 252690 673604 252696
rect 673656 252634 673684 260170
rect 673736 259752 673788 259758
rect 673736 259694 673788 259700
rect 673472 252606 673684 252634
rect 673368 249552 673420 249558
rect 673368 249494 673420 249500
rect 673472 241126 673500 252606
rect 673552 252544 673604 252550
rect 673748 252498 673776 259694
rect 673552 252486 673604 252492
rect 673564 243642 673592 252486
rect 673656 252470 673776 252498
rect 673552 243636 673604 243642
rect 673552 243578 673604 243584
rect 673656 242214 673684 252470
rect 673736 252340 673788 252346
rect 673736 252282 673788 252288
rect 673748 242962 673776 252282
rect 673840 249626 673868 263026
rect 674472 262268 674524 262274
rect 674472 262210 674524 262216
rect 674288 259004 674340 259010
rect 674288 258946 674340 258952
rect 674300 252346 674328 258946
rect 674288 252340 674340 252346
rect 674288 252282 674340 252288
rect 674288 252204 674340 252210
rect 674288 252146 674340 252152
rect 673828 249620 673880 249626
rect 673828 249562 673880 249568
rect 674300 245478 674328 252146
rect 674484 249694 674512 262210
rect 674932 261860 674984 261866
rect 674932 261802 674984 261808
rect 674748 259684 674800 259690
rect 674748 259626 674800 259632
rect 674656 259616 674708 259622
rect 674656 259558 674708 259564
rect 674564 256760 674616 256766
rect 674564 256702 674616 256708
rect 674576 252210 674604 256702
rect 674564 252204 674616 252210
rect 674564 252146 674616 252152
rect 674668 252090 674696 259558
rect 674576 252062 674696 252090
rect 674472 249688 674524 249694
rect 674472 249630 674524 249636
rect 674472 249552 674524 249558
rect 674472 249494 674524 249500
rect 674288 245472 674340 245478
rect 674288 245414 674340 245420
rect 673736 242956 673788 242962
rect 673736 242898 673788 242904
rect 673644 242208 673696 242214
rect 673644 242150 673696 242156
rect 673460 241120 673512 241126
rect 673460 241062 673512 241068
rect 674484 239970 674512 249494
rect 674576 246566 674604 252062
rect 674656 251932 674708 251938
rect 674656 251874 674708 251880
rect 674564 246560 674616 246566
rect 674564 246502 674616 246508
rect 674668 246090 674696 251874
rect 674760 251818 674788 259626
rect 674840 259548 674892 259554
rect 674840 259490 674892 259496
rect 674852 251938 674880 259490
rect 674840 251932 674892 251938
rect 674840 251874 674892 251880
rect 674760 251790 674880 251818
rect 674748 251252 674800 251258
rect 674748 251194 674800 251200
rect 674656 246084 674708 246090
rect 674656 246026 674708 246032
rect 674472 239964 674524 239970
rect 674472 239906 674524 239912
rect 674760 235550 674788 251194
rect 674852 247314 674880 251790
rect 674840 247308 674892 247314
rect 674840 247250 674892 247256
rect 674944 247042 674972 261802
rect 675024 259480 675076 259486
rect 675024 259422 675076 259428
rect 675036 250238 675064 259422
rect 675024 250232 675076 250238
rect 675024 250174 675076 250180
rect 675024 249824 675076 249830
rect 675024 249766 675076 249772
rect 674932 247036 674984 247042
rect 674932 246978 674984 246984
rect 675036 246922 675064 249766
rect 674944 246894 675064 246922
rect 674944 235618 674972 246894
rect 675128 237374 675156 264946
rect 675312 251258 675340 264946
rect 675666 260536 675722 260545
rect 675666 260471 675722 260480
rect 675680 260234 675708 260471
rect 675668 260228 675720 260234
rect 675668 260170 675720 260176
rect 675666 260128 675722 260137
rect 675666 260063 675722 260072
rect 675680 259758 675708 260063
rect 675668 259752 675720 259758
rect 675668 259694 675720 259700
rect 675772 256694 675800 265367
rect 679176 265305 679204 278054
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 679162 265296 679218 265305
rect 679162 265231 679218 265240
rect 676034 264208 676090 264217
rect 676034 264143 676090 264152
rect 675850 263392 675906 263401
rect 675850 263327 675906 263336
rect 675680 256666 675800 256694
rect 675680 251394 675708 256666
rect 675864 253586 675892 263327
rect 676048 263090 676076 264143
rect 676126 263664 676182 263673
rect 676126 263599 676182 263608
rect 676036 263084 676088 263090
rect 676036 263026 676088 263032
rect 676034 262984 676090 262993
rect 676034 262919 676090 262928
rect 676048 262274 676076 262919
rect 676140 262546 676168 263599
rect 676128 262540 676180 262546
rect 676128 262482 676180 262488
rect 676126 262440 676182 262449
rect 676126 262375 676182 262384
rect 676140 262342 676168 262375
rect 676128 262336 676180 262342
rect 676128 262278 676180 262284
rect 676036 262268 676088 262274
rect 676036 262210 676088 262216
rect 676034 262168 676090 262177
rect 676034 262103 676090 262112
rect 676048 261866 676076 262103
rect 676036 261860 676088 261866
rect 676036 261802 676088 261808
rect 676034 261760 676090 261769
rect 676034 261695 676090 261704
rect 675942 260944 675998 260953
rect 675942 260879 675998 260888
rect 675956 259622 675984 260879
rect 675944 259616 675996 259622
rect 675944 259558 675996 259564
rect 676048 259486 676076 261695
rect 676126 261216 676182 261225
rect 676126 261151 676182 261160
rect 676140 259690 676168 261151
rect 676128 259684 676180 259690
rect 676128 259626 676180 259632
rect 676126 259584 676182 259593
rect 676126 259519 676128 259528
rect 676180 259519 676182 259528
rect 676128 259490 676180 259496
rect 676036 259480 676088 259486
rect 676036 259422 676088 259428
rect 676034 259312 676090 259321
rect 676034 259247 676090 259256
rect 676048 259010 676076 259247
rect 676036 259004 676088 259010
rect 676036 258946 676088 258952
rect 676034 258904 676090 258913
rect 676034 258839 676090 258848
rect 676048 256766 676076 258839
rect 678978 258360 679034 258369
rect 678978 258295 679034 258304
rect 678992 257553 679020 258295
rect 678978 257544 679034 257553
rect 678978 257479 679034 257488
rect 678992 256834 679020 257479
rect 678980 256828 679032 256834
rect 678980 256770 679032 256776
rect 676036 256760 676088 256766
rect 676036 256702 676088 256708
rect 675772 253558 675892 253586
rect 675772 251394 675800 253558
rect 675668 251388 675720 251394
rect 675668 251330 675720 251336
rect 675760 251388 675812 251394
rect 675760 251330 675812 251336
rect 675300 251252 675352 251258
rect 675300 251194 675352 251200
rect 675312 251110 675432 251138
rect 675312 251070 675340 251110
rect 675220 251042 675340 251070
rect 675404 251056 675432 251110
rect 675220 247194 675248 251042
rect 675300 250980 675352 250986
rect 675300 250922 675352 250928
rect 675312 249830 675340 250922
rect 675760 250776 675812 250782
rect 675760 250718 675812 250724
rect 675772 250512 675800 250718
rect 675484 250232 675536 250238
rect 675484 250174 675536 250180
rect 675496 249900 675524 250174
rect 675300 249824 675352 249830
rect 675300 249766 675352 249772
rect 675300 249688 675352 249694
rect 675300 249630 675352 249636
rect 675312 247398 675340 249630
rect 675392 249620 675444 249626
rect 675392 249562 675444 249568
rect 675404 249220 675432 249562
rect 675312 247370 675418 247398
rect 675392 247308 675444 247314
rect 675392 247250 675444 247256
rect 675220 247166 675340 247194
rect 675208 247036 675260 247042
rect 675208 246978 675260 246984
rect 675036 237346 675156 237374
rect 674932 235612 674984 235618
rect 674932 235554 674984 235560
rect 674748 235544 674800 235550
rect 674748 235486 674800 235492
rect 675036 221513 675064 237346
rect 675220 236382 675248 246978
rect 675312 245614 675340 247166
rect 675404 246840 675432 247250
rect 675392 246560 675444 246566
rect 675392 246502 675444 246508
rect 675404 246199 675432 246502
rect 675392 246084 675444 246090
rect 675392 246026 675444 246032
rect 675300 245608 675352 245614
rect 675300 245550 675352 245556
rect 675404 245548 675432 246026
rect 675300 245472 675352 245478
rect 675300 245414 675352 245420
rect 675312 241245 675340 245414
rect 675392 243636 675444 243642
rect 675392 243578 675444 243584
rect 675404 243071 675432 243578
rect 675392 242956 675444 242962
rect 675392 242898 675444 242904
rect 675404 242519 675432 242898
rect 675392 242208 675444 242214
rect 675392 242150 675444 242156
rect 675404 241876 675432 242150
rect 675312 241217 675418 241245
rect 675300 241120 675352 241126
rect 675300 241062 675352 241068
rect 675312 240054 675340 241062
rect 675312 240026 675418 240054
rect 675300 239964 675352 239970
rect 675300 239906 675352 239912
rect 675312 238218 675340 239906
rect 675312 238190 675418 238218
rect 675220 236354 675418 236382
rect 675760 235612 675812 235618
rect 675760 235554 675812 235560
rect 675668 235544 675720 235550
rect 675668 235486 675720 235492
rect 675680 222329 675708 235486
rect 675666 222320 675722 222329
rect 675666 222255 675722 222264
rect 675588 221921 675616 221942
rect 675574 221912 675630 221921
rect 675312 221870 675574 221898
rect 675022 221504 675078 221513
rect 675022 221439 675078 221448
rect 674472 218340 674524 218346
rect 674472 218282 674524 218288
rect 673090 216880 673146 216889
rect 673090 216815 673146 216824
rect 672998 132968 673054 132977
rect 672998 132903 673054 132912
rect 673104 129470 673132 216815
rect 673274 216608 673330 216617
rect 673274 216543 673330 216552
rect 673288 131714 673316 216543
rect 674288 216300 674340 216306
rect 674288 216242 674340 216248
rect 673552 215552 673604 215558
rect 673552 215494 673604 215500
rect 673460 212628 673512 212634
rect 673460 212570 673512 212576
rect 673472 207330 673500 212570
rect 673460 207324 673512 207330
rect 673460 207266 673512 207272
rect 673564 207210 673592 215494
rect 673736 215484 673788 215490
rect 673736 215426 673788 215432
rect 673644 214668 673696 214674
rect 673644 214610 673696 214616
rect 673380 207182 673592 207210
rect 673380 204270 673408 207182
rect 673552 207120 673604 207126
rect 673552 207062 673604 207068
rect 673460 207052 673512 207058
rect 673460 206994 673512 207000
rect 673368 204264 673420 204270
rect 673368 204206 673420 204212
rect 673472 197606 673500 206994
rect 673460 197600 673512 197606
rect 673460 197542 673512 197548
rect 673564 191690 673592 207062
rect 673656 197198 673684 214610
rect 673748 201550 673776 215426
rect 673828 212560 673880 212566
rect 673828 212502 673880 212508
rect 673736 201544 673788 201550
rect 673736 201486 673788 201492
rect 673840 200734 673868 212502
rect 673828 200728 673880 200734
rect 673828 200670 673880 200676
rect 674300 198422 674328 216242
rect 674484 204406 674512 218282
rect 674748 218068 674800 218074
rect 674748 218010 674800 218016
rect 674656 216708 674708 216714
rect 674656 216650 674708 216656
rect 674564 215416 674616 215422
rect 674564 215358 674616 215364
rect 674472 204400 674524 204406
rect 674472 204342 674524 204348
rect 674472 204264 674524 204270
rect 674472 204206 674524 204212
rect 674288 198416 674340 198422
rect 674288 198358 674340 198364
rect 673644 197192 673696 197198
rect 673644 197134 673696 197140
rect 674484 195362 674512 204206
rect 674576 201890 674604 215358
rect 674668 202774 674696 216650
rect 674760 205630 674788 218010
rect 674932 215892 674984 215898
rect 674932 215834 674984 215840
rect 674840 215348 674892 215354
rect 674840 215290 674892 215296
rect 674748 205624 674800 205630
rect 674748 205566 674800 205572
rect 674748 205488 674800 205494
rect 674748 205430 674800 205436
rect 674656 202768 674708 202774
rect 674656 202710 674708 202716
rect 674564 201884 674616 201890
rect 674564 201826 674616 201832
rect 674760 196450 674788 205430
rect 674852 205018 674880 215290
rect 674944 207126 674972 215834
rect 674932 207120 674984 207126
rect 674932 207062 674984 207068
rect 674932 206372 674984 206378
rect 674932 206314 674984 206320
rect 674840 205012 674892 205018
rect 674840 204954 674892 204960
rect 674838 204912 674894 204921
rect 674838 204847 674894 204856
rect 674748 196444 674800 196450
rect 674748 196386 674800 196392
rect 674472 195356 674524 195362
rect 674472 195298 674524 195304
rect 674852 192794 674880 204847
rect 674944 192914 674972 206314
rect 675024 206304 675076 206310
rect 675024 206246 675076 206252
rect 675036 196586 675064 206246
rect 675208 206236 675260 206242
rect 675208 206178 675260 206184
rect 675024 196580 675076 196586
rect 675024 196522 675076 196528
rect 675024 196444 675076 196450
rect 675024 196386 675076 196392
rect 674932 192908 674984 192914
rect 674932 192850 674984 192856
rect 674760 192766 674880 192794
rect 673552 191684 673604 191690
rect 673552 191626 673604 191632
rect 673368 176044 673420 176050
rect 673368 175986 673420 175992
rect 673276 131708 673328 131714
rect 673276 131650 673328 131656
rect 673380 131510 673408 175986
rect 674760 175574 674788 192766
rect 674930 176896 674986 176905
rect 674930 176831 674986 176840
rect 674748 175568 674800 175574
rect 674748 175510 674800 175516
rect 674944 175114 674972 176831
rect 675036 176390 675064 196386
rect 675220 193474 675248 206178
rect 675312 193594 675340 221870
rect 675574 221847 675630 221856
rect 675390 221096 675446 221105
rect 675390 221031 675446 221040
rect 675404 206378 675432 221031
rect 675772 220697 675800 235554
rect 703694 224196 703722 224332
rect 704154 224196 704182 224332
rect 704614 224196 704642 224332
rect 705074 224196 705102 224332
rect 705534 224196 705562 224332
rect 705994 224196 706022 224332
rect 706454 224196 706482 224332
rect 706914 224196 706942 224332
rect 707374 224196 707402 224332
rect 707834 224196 707862 224332
rect 708294 224196 708322 224332
rect 708754 224196 708782 224332
rect 709214 224196 709242 224332
rect 675850 223544 675906 223553
rect 675850 223479 675906 223488
rect 675864 221066 675892 223479
rect 675942 223136 675998 223145
rect 675942 223071 675998 223080
rect 675852 221060 675904 221066
rect 675852 221002 675904 221008
rect 675956 220862 675984 223071
rect 676034 222728 676090 222737
rect 676034 222663 676090 222672
rect 676048 221202 676076 222663
rect 676036 221196 676088 221202
rect 676036 221138 676088 221144
rect 675944 220856 675996 220862
rect 675944 220798 675996 220804
rect 675758 220688 675814 220697
rect 675758 220623 675814 220632
rect 675942 220280 675998 220289
rect 675942 220215 675998 220224
rect 675576 219632 675628 219638
rect 675576 219574 675628 219580
rect 675482 218648 675538 218657
rect 675482 218583 675538 218592
rect 675392 206372 675444 206378
rect 675392 206314 675444 206320
rect 675496 206242 675524 218583
rect 675588 206281 675616 219574
rect 675956 219570 675984 220215
rect 676036 219632 676088 219638
rect 676036 219574 676088 219580
rect 675668 219564 675720 219570
rect 675668 219506 675720 219512
rect 675944 219564 675996 219570
rect 675944 219506 675996 219512
rect 675574 206272 675630 206281
rect 675484 206236 675536 206242
rect 675680 206242 675708 219506
rect 676048 219473 676076 219574
rect 676034 219464 676090 219473
rect 676034 219399 676090 219408
rect 676034 219056 676090 219065
rect 676034 218991 676090 219000
rect 676048 218346 676076 218991
rect 676036 218340 676088 218346
rect 676036 218282 676088 218288
rect 676034 218240 676090 218249
rect 676034 218175 676090 218184
rect 676048 218074 676076 218175
rect 676036 218068 676088 218074
rect 676036 218010 676088 218016
rect 676034 217832 676090 217841
rect 676034 217767 676090 217776
rect 675942 217424 675998 217433
rect 675942 217359 675998 217368
rect 675850 217016 675906 217025
rect 675850 216951 675906 216960
rect 675864 215898 675892 216951
rect 675956 216306 675984 217359
rect 676048 216714 676076 217767
rect 676036 216708 676088 216714
rect 676036 216650 676088 216656
rect 676034 216608 676090 216617
rect 676034 216543 676090 216552
rect 675944 216300 675996 216306
rect 675944 216242 675996 216248
rect 675942 216200 675998 216209
rect 675942 216135 675998 216144
rect 675852 215892 675904 215898
rect 675852 215834 675904 215840
rect 675850 215792 675906 215801
rect 675850 215727 675906 215736
rect 675760 215552 675812 215558
rect 675760 215494 675812 215500
rect 675772 215393 675800 215494
rect 675864 215490 675892 215727
rect 675852 215484 675904 215490
rect 675852 215426 675904 215432
rect 675956 215422 675984 216135
rect 675944 215416 675996 215422
rect 675758 215384 675814 215393
rect 675944 215358 675996 215364
rect 676048 215354 676076 216543
rect 675758 215319 675814 215328
rect 676036 215348 676088 215354
rect 676036 215290 676088 215296
rect 676034 214976 676090 214985
rect 676034 214911 676090 214920
rect 676048 214674 676076 214911
rect 676036 214668 676088 214674
rect 676036 214610 676088 214616
rect 676034 214568 676090 214577
rect 676034 214503 676090 214512
rect 675942 214160 675998 214169
rect 675942 214095 675998 214104
rect 675758 213752 675814 213761
rect 675758 213687 675814 213696
rect 675772 206310 675800 213687
rect 675956 212634 675984 214095
rect 675944 212628 675996 212634
rect 675944 212570 675996 212576
rect 676048 212566 676076 214503
rect 676036 212560 676088 212566
rect 676036 212502 676088 212508
rect 676034 212120 676090 212129
rect 676034 212055 676036 212064
rect 676088 212055 676090 212064
rect 676036 212026 676088 212032
rect 675760 206304 675812 206310
rect 675760 206246 675812 206252
rect 675574 206207 675630 206216
rect 675668 206236 675720 206242
rect 675484 206178 675536 206184
rect 675668 206178 675720 206184
rect 675390 206000 675446 206009
rect 675390 205935 675446 205944
rect 675404 205875 675432 205935
rect 675392 205624 675444 205630
rect 675392 205566 675444 205572
rect 675404 205323 675432 205566
rect 675392 205012 675444 205018
rect 675392 204954 675444 204960
rect 675404 204680 675432 204954
rect 675392 204400 675444 204406
rect 675392 204342 675444 204348
rect 675404 204035 675432 204342
rect 675392 202768 675444 202774
rect 675392 202710 675444 202716
rect 675404 202195 675432 202710
rect 675392 201884 675444 201890
rect 675392 201826 675444 201832
rect 675404 201620 675432 201826
rect 675392 201544 675444 201550
rect 675392 201486 675444 201492
rect 675404 201008 675432 201486
rect 675392 200728 675444 200734
rect 675392 200670 675444 200676
rect 675404 200328 675432 200670
rect 675392 198416 675444 198422
rect 675392 198358 675444 198364
rect 675404 197880 675432 198358
rect 675484 197600 675536 197606
rect 675484 197542 675536 197548
rect 675496 197336 675524 197542
rect 675392 197192 675444 197198
rect 675392 197134 675444 197140
rect 675404 196656 675432 197134
rect 675392 196580 675444 196586
rect 675392 196522 675444 196528
rect 675404 196044 675432 196522
rect 675392 195356 675444 195362
rect 675392 195298 675444 195304
rect 675404 194820 675432 195298
rect 675300 193588 675352 193594
rect 675300 193530 675352 193536
rect 675220 193446 675432 193474
rect 675300 193384 675352 193390
rect 675300 193326 675352 193332
rect 675208 192908 675260 192914
rect 675208 192850 675260 192856
rect 675220 176662 675248 192850
rect 675312 177313 675340 193326
rect 675404 192984 675432 193446
rect 675392 191684 675444 191690
rect 675392 191626 675444 191632
rect 675404 191148 675432 191626
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 675850 178528 675906 178537
rect 675850 178463 675906 178472
rect 675298 177304 675354 177313
rect 675298 177239 675354 177248
rect 675864 176866 675892 178463
rect 675942 178120 675998 178129
rect 675942 178055 675998 178064
rect 675956 177002 675984 178055
rect 676034 177712 676090 177721
rect 676034 177647 676090 177656
rect 676048 177138 676076 177647
rect 676036 177132 676088 177138
rect 676036 177074 676088 177080
rect 675944 176996 675996 177002
rect 675944 176938 675996 176944
rect 675852 176860 675904 176866
rect 675852 176802 675904 176808
rect 675208 176656 675260 176662
rect 675208 176598 675260 176604
rect 676036 176656 676088 176662
rect 676036 176598 676088 176604
rect 676048 176497 676076 176598
rect 676034 176488 676090 176497
rect 676034 176423 676090 176432
rect 675024 176384 675076 176390
rect 675024 176326 675076 176332
rect 676036 176384 676088 176390
rect 676036 176326 676088 176332
rect 675942 176080 675998 176089
rect 675942 176015 675944 176024
rect 675996 176015 675998 176024
rect 675944 175986 675996 175992
rect 676048 175681 676076 176326
rect 676034 175672 676090 175681
rect 676034 175607 676090 175616
rect 676036 175568 676088 175574
rect 676036 175510 676088 175516
rect 675390 175264 675446 175273
rect 675364 175222 675390 175250
rect 675390 175199 675446 175208
rect 674944 175086 675248 175114
rect 674748 173936 674800 173942
rect 674748 173878 674800 173884
rect 673552 172916 673604 172922
rect 673552 172858 673604 172864
rect 673460 164892 673512 164898
rect 673460 164834 673512 164840
rect 673472 150414 673500 164834
rect 673460 150408 673512 150414
rect 673460 150350 673512 150356
rect 673564 148578 673592 172858
rect 674288 172100 674340 172106
rect 674288 172042 674340 172048
rect 673736 170060 673788 170066
rect 673736 170002 673788 170008
rect 673644 169244 673696 169250
rect 673644 169186 673696 169192
rect 673656 152250 673684 169186
rect 673748 164898 673776 170002
rect 673828 168564 673880 168570
rect 673828 168506 673880 168512
rect 673736 164892 673788 164898
rect 673736 164834 673788 164840
rect 673840 164778 673868 168506
rect 673748 164750 673868 164778
rect 673644 152244 673696 152250
rect 673644 152186 673696 152192
rect 673748 151570 673776 164750
rect 674300 164626 674328 172042
rect 674564 171216 674616 171222
rect 674564 171158 674616 171164
rect 674472 168632 674524 168638
rect 674472 168574 674524 168580
rect 673828 164620 673880 164626
rect 673828 164562 673880 164568
rect 674288 164620 674340 164626
rect 674288 164562 674340 164568
rect 673840 153406 673868 164562
rect 674484 164490 674512 168574
rect 674288 164484 674340 164490
rect 674288 164426 674340 164432
rect 674472 164484 674524 164490
rect 674472 164426 674524 164432
rect 674300 155854 674328 164426
rect 674472 164348 674524 164354
rect 674472 164290 674524 164296
rect 674484 156942 674512 164290
rect 674472 156936 674524 156942
rect 674472 156878 674524 156884
rect 674288 155848 674340 155854
rect 674288 155790 674340 155796
rect 673828 153400 673880 153406
rect 673828 153342 673880 153348
rect 673736 151564 673788 151570
rect 673736 151506 673788 151512
rect 673552 148572 673604 148578
rect 673552 148514 673604 148520
rect 674576 146742 674604 171158
rect 674656 171148 674708 171154
rect 674656 171090 674708 171096
rect 674668 164354 674696 171090
rect 674656 164348 674708 164354
rect 674656 164290 674708 164296
rect 674656 164212 674708 164218
rect 674656 164154 674708 164160
rect 674668 158098 674696 164154
rect 674760 159390 674788 173878
rect 674840 171284 674892 171290
rect 674840 171226 674892 171232
rect 674748 159384 674800 159390
rect 674748 159326 674800 159332
rect 674656 158092 674708 158098
rect 674656 158034 674708 158040
rect 674852 157758 674880 171226
rect 674932 169652 674984 169658
rect 674932 169594 674984 169600
rect 674944 164218 674972 169594
rect 675024 168972 675076 168978
rect 675024 168914 675076 168920
rect 674932 164212 674984 164218
rect 674932 164154 674984 164160
rect 675036 164098 675064 168914
rect 675116 164484 675168 164490
rect 675116 164426 675168 164432
rect 674944 164070 675064 164098
rect 674840 157752 674892 157758
rect 674840 157694 674892 157700
rect 674944 155922 674972 164070
rect 675024 164008 675076 164014
rect 675024 163950 675076 163956
rect 675036 160206 675064 163950
rect 675024 160200 675076 160206
rect 675024 160142 675076 160148
rect 675024 160064 675076 160070
rect 675024 160006 675076 160012
rect 674932 155916 674984 155922
rect 674932 155858 674984 155864
rect 674564 146736 674616 146742
rect 674564 146678 674616 146684
rect 675036 140774 675064 160006
rect 675128 150482 675156 164426
rect 675116 150476 675168 150482
rect 675116 150418 675168 150424
rect 675036 140746 675156 140774
rect 673368 131504 673420 131510
rect 673368 131446 673420 131452
rect 675128 129734 675156 140746
rect 675220 132462 675248 175086
rect 675404 164490 675432 175199
rect 676048 174865 676076 175510
rect 676034 174856 676090 174865
rect 676034 174791 676090 174800
rect 675758 174448 675814 174457
rect 675758 174383 675814 174392
rect 675574 173224 675630 173233
rect 675574 173159 675630 173168
rect 675392 164484 675444 164490
rect 675392 164426 675444 164432
rect 675588 164370 675616 173159
rect 675666 171592 675722 171601
rect 675666 171527 675722 171536
rect 675312 164342 675616 164370
rect 675312 160290 675340 164342
rect 675680 164014 675708 171527
rect 675668 164008 675720 164014
rect 675668 163950 675720 163956
rect 675772 161226 675800 174383
rect 676034 174040 676090 174049
rect 676034 173975 676090 173984
rect 676048 173942 676076 173975
rect 676036 173936 676088 173942
rect 676036 173878 676088 173884
rect 676034 173632 676090 173641
rect 676034 173567 676090 173576
rect 676048 172922 676076 173567
rect 676036 172916 676088 172922
rect 676036 172858 676088 172864
rect 676034 172816 676090 172825
rect 676034 172751 676090 172760
rect 675942 172408 675998 172417
rect 675942 172343 675998 172352
rect 675956 172106 675984 172343
rect 675944 172100 675996 172106
rect 675944 172042 675996 172048
rect 675942 172000 675998 172009
rect 675942 171935 675998 171944
rect 675956 171222 675984 171935
rect 676048 171290 676076 172751
rect 676036 171284 676088 171290
rect 676036 171226 676088 171232
rect 675944 171216 675996 171222
rect 675944 171158 675996 171164
rect 676034 171184 676090 171193
rect 676034 171119 676036 171128
rect 676088 171119 676090 171128
rect 676036 171090 676088 171096
rect 676034 170776 676090 170785
rect 676034 170711 676090 170720
rect 675942 170368 675998 170377
rect 675942 170303 675998 170312
rect 675956 170066 675984 170303
rect 675944 170060 675996 170066
rect 675944 170002 675996 170008
rect 675942 169960 675998 169969
rect 675942 169895 675998 169904
rect 675956 169250 675984 169895
rect 676048 169658 676076 170711
rect 676036 169652 676088 169658
rect 676036 169594 676088 169600
rect 676034 169552 676090 169561
rect 676034 169487 676090 169496
rect 675944 169244 675996 169250
rect 675944 169186 675996 169192
rect 675942 169144 675998 169153
rect 675942 169079 675998 169088
rect 675956 168638 675984 169079
rect 676048 168978 676076 169487
rect 676036 168972 676088 168978
rect 676036 168914 676088 168920
rect 676034 168736 676090 168745
rect 676034 168671 676090 168680
rect 675944 168632 675996 168638
rect 675944 168574 675996 168580
rect 676048 168570 676076 168671
rect 676036 168564 676088 168570
rect 676036 168506 676088 168512
rect 676034 167104 676090 167113
rect 676034 167039 676036 167048
rect 676088 167039 676090 167048
rect 676036 167010 676088 167016
rect 675760 161220 675812 161226
rect 675760 161162 675812 161168
rect 675392 161016 675444 161022
rect 675392 160958 675444 160964
rect 675404 160888 675432 160958
rect 675404 160290 675432 160344
rect 675312 160262 675432 160290
rect 675300 160200 675352 160206
rect 675300 160142 675352 160148
rect 675312 159678 675340 160142
rect 675312 159650 675418 159678
rect 675484 159384 675536 159390
rect 675484 159326 675536 159332
rect 675496 159052 675524 159326
rect 675300 158092 675352 158098
rect 675300 158034 675352 158040
rect 675312 156006 675340 158034
rect 675484 157752 675536 157758
rect 675484 157694 675536 157700
rect 675496 157216 675524 157694
rect 675392 156936 675444 156942
rect 675392 156878 675444 156884
rect 675404 156643 675432 156878
rect 675312 155978 675418 156006
rect 675484 155916 675536 155922
rect 675484 155858 675536 155864
rect 675300 155848 675352 155854
rect 675300 155790 675352 155796
rect 675312 152334 675340 155790
rect 675496 155380 675524 155858
rect 675392 153400 675444 153406
rect 675392 153342 675444 153348
rect 675404 152864 675432 153342
rect 675312 152306 675418 152334
rect 675300 152244 675352 152250
rect 675300 152186 675352 152192
rect 675312 151689 675340 152186
rect 675312 151661 675418 151689
rect 675300 151564 675352 151570
rect 675300 151506 675352 151512
rect 675312 151042 675340 151506
rect 675312 151014 675418 151042
rect 675300 150476 675352 150482
rect 675300 150418 675352 150424
rect 675208 132456 675260 132462
rect 675208 132398 675260 132404
rect 675312 130529 675340 150418
rect 675392 150408 675444 150414
rect 675392 150350 675444 150356
rect 675404 149835 675432 150350
rect 675392 148572 675444 148578
rect 675392 148514 675444 148520
rect 675404 147968 675432 148514
rect 675392 146736 675444 146742
rect 675392 146678 675444 146684
rect 675404 146132 675432 146678
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 676126 133104 676182 133113
rect 676126 133039 676182 133048
rect 676034 132968 676090 132977
rect 676034 132903 676090 132912
rect 676048 132666 676076 132903
rect 676140 132802 676168 133039
rect 676220 132932 676272 132938
rect 676220 132874 676272 132880
rect 676128 132796 676180 132802
rect 676128 132738 676180 132744
rect 676232 132705 676260 132874
rect 676218 132696 676274 132705
rect 676036 132660 676088 132666
rect 676218 132631 676274 132640
rect 676036 132602 676088 132608
rect 676036 132456 676088 132462
rect 676036 132398 676088 132404
rect 676048 132161 676076 132398
rect 676034 132152 676090 132161
rect 676034 132087 676090 132096
rect 676034 131744 676090 131753
rect 676034 131679 676036 131688
rect 676088 131679 676090 131688
rect 676036 131650 676088 131656
rect 676220 131504 676272 131510
rect 676218 131472 676220 131481
rect 676272 131472 676274 131481
rect 676218 131407 676274 131416
rect 676034 130928 676090 130937
rect 676034 130863 676036 130872
rect 676088 130863 676090 130872
rect 676036 130834 676088 130840
rect 675298 130520 675354 130529
rect 675298 130455 675354 130464
rect 676034 130112 676090 130121
rect 676034 130047 676036 130056
rect 676088 130047 676090 130056
rect 676036 130018 676088 130024
rect 675128 129713 675800 129734
rect 675128 129706 675814 129713
rect 675758 129704 675814 129706
rect 675758 129639 675814 129648
rect 673092 129464 673144 129470
rect 676220 129464 676272 129470
rect 673092 129406 673144 129412
rect 676218 129432 676220 129441
rect 676272 129432 676274 129441
rect 676218 129367 676274 129376
rect 676034 128888 676090 128897
rect 676034 128823 676090 128832
rect 675942 128480 675998 128489
rect 675942 128415 675998 128424
rect 675574 128072 675630 128081
rect 675574 128007 675630 128016
rect 674748 127764 674800 127770
rect 674748 127706 674800 127712
rect 673552 127356 673604 127362
rect 673552 127298 673604 127304
rect 672722 122904 672778 122913
rect 672722 122839 672778 122848
rect 672448 121644 672500 121650
rect 672448 121586 672500 121592
rect 672460 109313 672488 121586
rect 672446 109304 672502 109313
rect 672446 109239 672502 109248
rect 673564 104582 673592 127298
rect 673828 127084 673880 127090
rect 673828 127026 673880 127032
rect 673644 124908 673696 124914
rect 673644 124850 673696 124856
rect 673656 106350 673684 124850
rect 673736 124500 673788 124506
rect 673736 124442 673788 124448
rect 673748 110090 673776 124442
rect 673736 110084 673788 110090
rect 673736 110026 673788 110032
rect 673840 108254 673868 127026
rect 674656 126540 674708 126546
rect 674656 126482 674708 126488
rect 674288 121576 674340 121582
rect 674288 121518 674340 121524
rect 673828 108248 673880 108254
rect 673828 108190 673880 108196
rect 674300 106418 674328 121518
rect 674472 121508 674524 121514
rect 674472 121450 674524 121456
rect 674668 121454 674696 126482
rect 674484 107574 674512 121450
rect 674576 121426 674696 121454
rect 674576 110514 674604 121426
rect 674760 121378 674788 127706
rect 674840 127016 674892 127022
rect 674840 126958 674892 126964
rect 674748 121372 674800 121378
rect 674748 121314 674800 121320
rect 674748 121168 674800 121174
rect 674748 121110 674800 121116
rect 674760 114374 674788 121110
rect 674748 114368 674800 114374
rect 674748 114310 674800 114316
rect 674852 113762 674880 126958
rect 675298 126032 675354 126041
rect 675298 125967 675354 125976
rect 675206 125624 675262 125633
rect 675206 125559 675262 125568
rect 674932 124296 674984 124302
rect 674932 124238 674984 124244
rect 674944 121446 674972 124238
rect 675024 124228 675076 124234
rect 675024 124170 675076 124176
rect 674932 121440 674984 121446
rect 674932 121382 674984 121388
rect 674932 121168 674984 121174
rect 674932 121110 674984 121116
rect 674840 113756 674892 113762
rect 674840 113698 674892 113704
rect 674576 110486 674788 110514
rect 674472 107568 674524 107574
rect 674472 107510 674524 107516
rect 674288 106412 674340 106418
rect 674288 106354 674340 106360
rect 673644 106344 673696 106350
rect 673644 106286 673696 106292
rect 673552 104576 673604 104582
rect 673552 104518 673604 104524
rect 672354 102504 672410 102513
rect 672354 102439 672410 102448
rect 674760 102134 674788 110486
rect 674944 110174 674972 121110
rect 675036 115054 675064 124170
rect 675220 121454 675248 125559
rect 675128 121426 675248 121454
rect 675024 115048 675076 115054
rect 675024 114990 675076 114996
rect 675128 110786 675156 121426
rect 675312 118402 675340 125967
rect 675220 118374 675340 118402
rect 675220 111466 675248 118374
rect 675588 118266 675616 128007
rect 675956 127362 675984 128415
rect 676048 127770 676076 128823
rect 676036 127764 676088 127770
rect 676036 127706 676088 127712
rect 676034 127664 676090 127673
rect 676034 127599 676090 127608
rect 675944 127356 675996 127362
rect 675944 127298 675996 127304
rect 675942 127256 675998 127265
rect 675942 127191 675998 127200
rect 675956 127090 675984 127191
rect 675944 127084 675996 127090
rect 675944 127026 675996 127032
rect 676048 127022 676076 127599
rect 676036 127016 676088 127022
rect 676036 126958 676088 126964
rect 676034 126848 676090 126857
rect 676034 126783 676090 126792
rect 676048 126546 676076 126783
rect 676036 126540 676088 126546
rect 676036 126482 676088 126488
rect 676034 126440 676090 126449
rect 676034 126375 676090 126384
rect 675942 125216 675998 125225
rect 675942 125151 675998 125160
rect 675956 124914 675984 125151
rect 675944 124908 675996 124914
rect 675944 124850 675996 124856
rect 675942 124808 675998 124817
rect 675942 124743 675998 124752
rect 675956 124506 675984 124743
rect 675944 124500 675996 124506
rect 675944 124442 675996 124448
rect 675942 124400 675998 124409
rect 675942 124335 675998 124344
rect 675956 124302 675984 124335
rect 675944 124296 675996 124302
rect 675944 124238 675996 124244
rect 676048 124234 676076 126375
rect 676036 124228 676088 124234
rect 676036 124170 676088 124176
rect 676034 123992 676090 124001
rect 676034 123927 676090 123936
rect 675942 123584 675998 123593
rect 675942 123519 675998 123528
rect 675956 121582 675984 123519
rect 675944 121576 675996 121582
rect 675944 121518 675996 121524
rect 676048 121514 676076 123927
rect 676218 121680 676274 121689
rect 676218 121615 676220 121624
rect 676272 121615 676274 121624
rect 676220 121586 676272 121592
rect 676036 121508 676088 121514
rect 676036 121450 676088 121456
rect 675312 118238 675616 118266
rect 675312 115138 675340 118238
rect 675392 115932 675444 115938
rect 675392 115874 675444 115880
rect 675404 115668 675432 115874
rect 675312 115110 675418 115138
rect 675300 115048 675352 115054
rect 675300 114990 675352 114996
rect 675312 114493 675340 114990
rect 675312 114465 675418 114493
rect 675300 114368 675352 114374
rect 675300 114310 675352 114316
rect 675312 113846 675340 114310
rect 675312 113818 675418 113846
rect 675300 113756 675352 113762
rect 675300 113698 675352 113704
rect 675312 112010 675340 113698
rect 675312 111982 675418 112010
rect 675220 111438 675418 111466
rect 675312 110894 675432 110922
rect 675312 110786 675340 110894
rect 675128 110758 675340 110786
rect 675404 110772 675432 110894
rect 674944 110146 675418 110174
rect 675116 110084 675168 110090
rect 675116 110026 675168 110032
rect 675128 106502 675156 110026
rect 675392 108248 675444 108254
rect 675392 108190 675444 108196
rect 675404 107644 675432 108190
rect 675392 107568 675444 107574
rect 675392 107510 675444 107516
rect 675404 107100 675432 107510
rect 675128 106474 675418 106502
rect 675392 106412 675444 106418
rect 675392 106354 675444 106360
rect 675116 106344 675168 106350
rect 675116 106286 675168 106292
rect 675128 104666 675156 106286
rect 675404 105808 675432 106354
rect 675128 104638 675340 104666
rect 675116 104576 675168 104582
rect 675116 104518 675168 104524
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675128 102830 675156 104518
rect 675312 104502 675432 104530
rect 675128 102802 675340 102830
rect 675312 102762 675340 102802
rect 675404 102762 675432 102816
rect 675312 102734 675432 102762
rect 674760 102106 674880 102134
rect 674852 100994 674880 102106
rect 674852 100966 675340 100994
rect 672078 100872 672134 100881
rect 675312 100858 675340 100966
rect 675404 100858 675432 100980
rect 675312 100830 675432 100858
rect 672078 100807 672134 100816
rect 666558 48512 666614 48521
rect 666558 48447 666614 48456
rect 665178 47424 665234 47433
rect 665178 47359 665234 47368
rect 661132 44124 661184 44130
rect 661132 44066 661184 44072
rect 622492 43172 622544 43178
rect 622492 43114 622544 43120
rect 622308 43104 622360 43110
rect 622308 43046 622360 43052
rect 607496 41472 607548 41478
rect 607496 41414 607548 41420
rect 602988 41404 603040 41410
rect 602988 41346 603040 41352
rect 571800 41336 571852 41342
rect 571800 41278 571852 41284
rect 549258 41032 549314 41041
rect 549258 40967 549314 40976
rect 514024 38616 514076 38622
rect 514024 38558 514076 38564
rect 502340 38548 502392 38554
rect 502340 38490 502392 38496
rect 513932 38548 513984 38554
rect 513932 38490 513984 38496
rect 229376 6520 229428 6526
rect 229376 6462 229428 6468
rect 233148 6520 233200 6526
rect 233148 6462 233200 6468
rect 229388 6225 229416 6462
rect 229374 6216 229430 6225
rect 229374 6151 229430 6160
<< via2 >>
rect 483570 1004692 483626 1004728
rect 483570 1004672 483572 1004692
rect 483572 1004672 483624 1004692
rect 483624 1004672 483626 1004692
rect 676034 897096 676090 897152
rect 675942 896688 675998 896744
rect 675850 894668 675906 894704
rect 675850 894648 675852 894668
rect 675852 894648 675904 894668
rect 675904 894648 675906 894668
rect 655518 867584 655574 867640
rect 655426 866496 655482 866552
rect 655702 868808 655758 868864
rect 655610 865272 655666 865328
rect 655794 863776 655850 863832
rect 656806 862552 656862 862608
rect 41786 817692 41842 817728
rect 41786 817672 41788 817692
rect 41788 817672 41840 817692
rect 41840 817672 41842 817692
rect 41786 817284 41842 817320
rect 41786 817264 41788 817284
rect 41788 817264 41840 817284
rect 41840 817264 41842 817284
rect 41786 816856 41842 816912
rect 44594 816070 44654 816130
rect 43626 815224 43682 815280
rect 41786 814544 41842 814600
rect 43442 813184 43498 813240
rect 42706 812776 42762 812832
rect 42246 811144 42302 811200
rect 41970 809104 42026 809160
rect 41878 808696 41934 808752
rect 41786 808308 41842 808344
rect 41786 808288 41788 808308
rect 41788 808288 41840 808308
rect 41840 808288 41842 808308
rect 41786 807472 41842 807528
rect 41786 806248 41842 806304
rect 42614 809512 42670 809568
rect 42338 806248 42394 806304
rect 43074 812368 43130 812424
rect 42798 811960 42854 812016
rect 42890 811552 42946 811608
rect 41878 794960 41934 795016
rect 41510 774732 41512 774752
rect 41512 774732 41564 774752
rect 41564 774732 41566 774752
rect 41510 774696 41566 774732
rect 41510 773900 41566 773936
rect 41510 773880 41512 773900
rect 41512 773880 41564 773900
rect 41564 773880 41566 773900
rect 41510 773492 41566 773528
rect 41510 773472 41512 773492
rect 41512 773472 41564 773492
rect 41564 773472 41566 773492
rect 43718 810736 43774 810792
rect 43810 810328 43866 810384
rect 43902 809920 43958 809976
rect 44686 814408 44746 814468
rect 44594 773254 44654 773314
rect 44594 772870 44654 772930
rect 43626 772384 43682 772440
rect 43718 771976 43774 772032
rect 42338 769528 42394 769584
rect 38290 767760 38346 767816
rect 38198 767352 38254 767408
rect 41510 764904 41566 764960
rect 38566 764496 38622 764552
rect 41602 764088 41658 764144
rect 41602 762884 41658 762920
rect 41602 762864 41604 762884
rect 41604 762864 41656 762884
rect 41656 762864 41658 762884
rect 43626 769120 43682 769176
rect 43074 768712 43130 768768
rect 42706 768304 42762 768360
rect 42430 765448 42486 765504
rect 43166 766264 43222 766320
rect 43258 765856 43314 765912
rect 44086 769936 44142 769992
rect 43902 767080 43958 767136
rect 43810 766672 43866 766728
rect 44306 731040 44362 731096
rect 44128 730632 44184 730688
rect 43902 730224 43958 730280
rect 41510 729408 41566 729464
rect 44778 813616 44838 813676
rect 44686 771618 44746 771678
rect 44686 771208 44746 771268
rect 44594 730054 44654 730114
rect 44594 729670 44654 729730
rect 44306 729136 44362 729192
rect 44138 729000 44194 729056
rect 43718 728864 43774 728920
rect 43902 728864 43958 728920
rect 43166 726824 43222 726880
rect 41786 724784 41842 724840
rect 41418 723288 41474 723344
rect 41510 720840 41566 720896
rect 41510 719616 41566 719672
rect 42246 723152 42302 723208
rect 42706 722744 42762 722800
rect 42338 721928 42394 721984
rect 43350 726416 43406 726472
rect 43258 722336 43314 722392
rect 43442 723968 43498 724024
rect 43626 721520 43682 721576
rect 41510 688356 41566 688392
rect 41510 688336 41512 688356
rect 41512 688336 41564 688356
rect 41564 688336 41566 688356
rect 41786 687676 41842 687712
rect 41786 687656 41788 687676
rect 41788 687656 41840 687676
rect 41840 687656 41842 687676
rect 41786 687268 41842 687304
rect 41786 687248 41788 687268
rect 41788 687248 41840 687268
rect 41840 687248 41842 687268
rect 43810 726008 43866 726064
rect 43994 725600 44050 725656
rect 43902 725192 43958 725248
rect 44086 724376 44142 724432
rect 59266 814544 59322 814600
rect 58254 790880 58310 790936
rect 58530 789284 58532 789304
rect 58532 789284 58584 789304
rect 58584 789284 58586 789304
rect 58530 789248 58586 789284
rect 58070 788432 58126 788488
rect 59266 787344 59322 787400
rect 58530 786120 58586 786176
rect 58438 784896 58494 784952
rect 44778 770828 44838 770888
rect 44778 770416 44838 770476
rect 44686 728418 44746 728478
rect 44686 728008 44746 728068
rect 44594 686854 44654 686914
rect 44594 686470 44654 686530
rect 43718 686024 43774 686080
rect 43074 685616 43130 685672
rect 42246 683168 42302 683224
rect 41878 681944 41934 682000
rect 41694 681400 41750 681456
rect 41786 678680 41842 678736
rect 41786 678272 41842 678328
rect 5446 676232 5502 676288
rect 5538 676096 5594 676152
rect 30562 675960 30618 676016
rect 42062 680312 42118 680368
rect 42062 670656 42118 670712
rect 42338 681128 42394 681184
rect 42430 679496 42486 679552
rect 43258 683576 43314 683632
rect 43534 682760 43590 682816
rect 43442 682352 43498 682408
rect 43258 665080 43314 665136
rect 43718 680720 43774 680776
rect 43626 679904 43682 679960
rect 41786 644884 41842 644940
rect 41510 644680 41566 644736
rect 41786 644088 41842 644124
rect 41786 644068 41788 644088
rect 41788 644068 41840 644088
rect 41840 644068 41842 644088
rect 44778 727628 44838 727688
rect 44778 727216 44838 727276
rect 44686 685218 44746 685278
rect 44686 684808 44746 684868
rect 44594 643654 44654 643714
rect 44594 643270 44654 643330
rect 43994 643048 44050 643104
rect 43902 642232 43958 642288
rect 43074 640328 43130 640384
rect 42338 639784 42394 639840
rect 42246 638152 42302 638208
rect 30194 637744 30250 637800
rect 30102 637336 30158 637392
rect 38474 634888 38530 634944
rect 24766 632576 24822 632632
rect 30102 632576 30158 632632
rect 41510 634480 41566 634536
rect 41510 633276 41566 633312
rect 41510 633256 41512 633276
rect 41512 633256 41564 633276
rect 41564 633256 41566 633276
rect 42706 636928 42762 636984
rect 42430 627408 42486 627464
rect 43166 638968 43222 639024
rect 43626 638560 43682 638616
rect 43258 636520 43314 636576
rect 42338 620880 42394 620936
rect 43074 622104 43130 622160
rect 43442 636112 43498 636168
rect 43350 635296 43406 635352
rect 43718 635704 43774 635760
rect 43626 627000 43682 627056
rect 41786 601724 41842 601760
rect 41786 601704 41788 601724
rect 41788 601704 41840 601724
rect 41840 601704 41842 601724
rect 44086 639376 44142 639432
rect 41510 601432 41566 601488
rect 43902 601432 43958 601488
rect 42706 601024 42762 601080
rect 41510 599800 41566 599856
rect 43074 600616 43130 600672
rect 42706 599120 42762 599176
rect 44778 684428 44838 684488
rect 44778 684016 44838 684076
rect 44686 642018 44746 642078
rect 44686 641608 44746 641668
rect 44594 600454 44654 600514
rect 44594 600070 44654 600130
rect 43902 599256 43958 599312
rect 43074 598984 43130 599040
rect 43166 596808 43222 596864
rect 41786 595176 41842 595232
rect 38566 593272 38622 593328
rect 41510 591232 41566 591288
rect 41510 590008 41566 590064
rect 42430 594768 42486 594824
rect 43718 596400 43774 596456
rect 43350 595584 43406 595640
rect 43442 594360 43498 594416
rect 43166 591912 43222 591968
rect 43074 585248 43130 585304
rect 43074 581304 43130 581360
rect 43350 583752 43406 583808
rect 43534 593952 43590 594008
rect 43626 592320 43682 592376
rect 43534 583752 43590 583808
rect 43810 593136 43866 593192
rect 44086 597216 44142 597272
rect 43994 595992 44050 596048
rect 44086 592728 44142 592784
rect 41510 558764 41512 558784
rect 41512 558764 41564 558784
rect 41564 558764 41566 558784
rect 41510 558728 41566 558764
rect 41510 558320 41566 558376
rect 41510 557540 41512 557560
rect 41512 557540 41564 557560
rect 41564 557540 41566 557560
rect 41510 557504 41566 557540
rect 44778 641228 44838 641288
rect 44778 640816 44838 640876
rect 44686 598818 44746 598878
rect 44686 598408 44746 598468
rect 44594 557254 44654 557314
rect 44594 556870 44654 556930
rect 43902 556416 43958 556472
rect 38106 555464 38162 555520
rect 43350 553560 43406 553616
rect 41786 551928 41842 551984
rect 41602 549752 41658 549808
rect 41418 549344 41474 549400
rect 38106 546352 38162 546408
rect 41510 548936 41566 548992
rect 41510 548528 41566 548584
rect 41510 548120 41566 548176
rect 41510 546916 41566 546952
rect 41510 546896 41512 546916
rect 41512 546896 41564 546916
rect 41564 546896 41566 546916
rect 43166 550296 43222 550352
rect 42246 535744 42302 535800
rect 42154 532752 42210 532808
rect 43350 538736 43406 538792
rect 43074 533024 43130 533080
rect 42430 532752 42486 532808
rect 42338 530168 42394 530224
rect 43166 530712 43222 530768
rect 42430 455912 42486 455968
rect 42430 450744 42486 450800
rect 42430 445848 42486 445904
rect 42430 440680 42486 440736
rect 41786 430908 41842 430944
rect 41786 430888 41788 430908
rect 41788 430888 41840 430908
rect 41840 430888 41842 430908
rect 41786 430480 41842 430536
rect 30102 428032 30158 428088
rect 42062 430072 42118 430128
rect 44778 598028 44838 598088
rect 44778 597616 44838 597676
rect 44686 555618 44746 555678
rect 44686 555208 44746 555268
rect 44594 429654 44654 429714
rect 44594 429270 44654 429330
rect 43718 428440 43774 428496
rect 42054 428256 42110 428312
rect 41786 427816 41842 427872
rect 30010 427624 30066 427680
rect 43442 426400 43498 426456
rect 42338 425992 42394 426048
rect 42246 424360 42302 424416
rect 41878 422728 41934 422784
rect 41786 420688 41842 420744
rect 41786 419484 41842 419520
rect 41786 419464 41788 419484
rect 41788 419464 41840 419484
rect 41840 419464 41842 419484
rect 41970 422320 42026 422376
rect 42706 425584 42762 425640
rect 43350 421504 43406 421560
rect 43258 421096 43314 421152
rect 43534 425176 43590 425232
rect 43626 424768 43682 424824
rect 41786 387640 41842 387696
rect 41510 387504 41566 387560
rect 41510 386708 41566 386744
rect 41510 386688 41512 386708
rect 41512 386688 41564 386708
rect 41564 386688 41566 386708
rect 43902 423952 43958 424008
rect 43810 423544 43866 423600
rect 43994 423136 44050 423192
rect 44086 421912 44142 421968
rect 44778 554828 44838 554888
rect 44778 554416 44838 554476
rect 44686 428024 44746 428084
rect 44686 427608 44746 427668
rect 44594 386454 44654 386514
rect 44594 386070 44654 386130
rect 43718 385600 43774 385656
rect 43534 385192 43590 385248
rect 43442 383152 43498 383208
rect 42706 382744 42762 382800
rect 38198 380976 38254 381032
rect 41970 379888 42026 379944
rect 41602 378528 41658 378584
rect 41418 378120 41474 378176
rect 41510 377712 41566 377768
rect 41786 377440 41842 377496
rect 41786 376236 41842 376272
rect 41786 376216 41788 376236
rect 41788 376216 41840 376236
rect 41840 376216 41842 376236
rect 43074 381928 43130 381984
rect 43258 381520 43314 381576
rect 43166 379480 43222 379536
rect 43718 382336 43774 382392
rect 43442 379072 43498 379128
rect 43718 380704 43774 380760
rect 43902 380296 43958 380352
rect 41510 344276 41566 344312
rect 41510 344256 41512 344276
rect 41512 344256 41564 344276
rect 41564 344256 41566 344276
rect 41510 343868 41566 343904
rect 41510 343848 41512 343868
rect 41512 343848 41564 343868
rect 41564 343848 41566 343868
rect 41510 343460 41566 343496
rect 41510 343440 41512 343460
rect 41512 343440 41564 343460
rect 41564 343440 41566 343460
rect 44778 427228 44838 427288
rect 44778 426816 44838 426876
rect 44686 384818 44746 384878
rect 44686 384408 44746 384468
rect 44594 343254 44654 343314
rect 44594 342870 44654 342930
rect 41510 342624 41566 342680
rect 43350 342080 43406 342136
rect 32862 339768 32918 339824
rect 33046 339768 33102 339824
rect 43166 338408 43222 338464
rect 41786 338000 41842 338056
rect 41510 336912 41566 336968
rect 41418 336504 41474 336560
rect 41602 334056 41658 334112
rect 41602 332852 41658 332888
rect 41602 332832 41604 332852
rect 41604 332832 41656 332852
rect 41656 332832 41658 332852
rect 32862 329704 32918 329760
rect 42338 336368 42394 336424
rect 42706 335552 42762 335608
rect 43258 335960 43314 336016
rect 41970 315560 42026 315616
rect 42154 313792 42210 313848
rect 41786 313112 41842 313168
rect 41786 312296 41842 312352
rect 41786 301316 41788 301336
rect 41788 301316 41840 301336
rect 41840 301316 41842 301336
rect 41786 301280 41842 301316
rect 43626 335144 43682 335200
rect 43442 334736 43498 334792
rect 41878 300872 41934 300928
rect 42706 300464 42762 300520
rect 41786 299240 41842 299296
rect 44778 384028 44838 384088
rect 44778 383616 44838 383676
rect 44686 341618 44746 341678
rect 44686 341208 44746 341268
rect 44594 300054 44654 300114
rect 44594 299670 44654 299730
rect 43074 298832 43130 298888
rect 42706 298152 42762 298208
rect 41878 294752 41934 294808
rect 30010 292712 30066 292768
rect 41786 291916 41842 291952
rect 41786 291896 41788 291916
rect 41788 291896 41840 291916
rect 41840 291896 41842 291916
rect 41786 291488 41842 291544
rect 42430 293936 42486 293992
rect 43626 296384 43682 296440
rect 43258 295976 43314 296032
rect 43166 293120 43222 293176
rect 41786 270408 41842 270464
rect 43534 295160 43590 295216
rect 43718 295568 43774 295624
rect 41786 258068 41788 258088
rect 41788 258068 41840 258088
rect 41840 258068 41842 258088
rect 41786 258032 41842 258068
rect 41510 257932 41512 257952
rect 41512 257932 41564 257952
rect 41564 257932 41566 257952
rect 41510 257896 41566 257932
rect 41510 257524 41512 257544
rect 41512 257524 41564 257544
rect 41564 257524 41566 257544
rect 41510 257488 41566 257524
rect 43902 294344 43958 294400
rect 43994 293528 44050 293584
rect 44086 292304 44142 292360
rect 44778 340828 44838 340888
rect 44778 340416 44838 340476
rect 44686 298418 44746 298478
rect 44686 298008 44746 298068
rect 44594 256854 44654 256914
rect 44594 256470 44654 256530
rect 43718 255992 43774 256048
rect 42246 255584 42302 255640
rect 30102 251368 30158 251424
rect 38106 248920 38162 248976
rect 38198 248512 38254 248568
rect 41510 248104 41566 248160
rect 41418 247716 41474 247752
rect 41418 247696 41420 247716
rect 41420 247696 41472 247716
rect 41472 247696 41474 247716
rect 41418 247288 41474 247344
rect 41510 246472 41566 246528
rect 42338 253544 42394 253600
rect 43810 253136 43866 253192
rect 43258 252320 43314 252376
rect 42706 249872 42762 249928
rect 41786 225936 41842 225992
rect 30102 204040 30158 204096
rect 41694 215056 41750 215112
rect 41510 214648 41566 214704
rect 41418 214240 41474 214296
rect 43074 249464 43130 249520
rect 43534 251912 43590 251968
rect 43626 251096 43682 251152
rect 43718 250688 43774 250744
rect 43994 250280 44050 250336
rect 44778 297628 44838 297688
rect 44778 297216 44838 297276
rect 44686 255218 44746 255278
rect 44686 254808 44746 254868
rect 44592 213654 44648 213710
rect 42338 212880 42394 212936
rect 41510 212608 41566 212664
rect 44778 254428 44838 254488
rect 44778 254016 44838 254076
rect 44688 212020 44744 212076
rect 58438 747632 58494 747688
rect 59266 746408 59322 746464
rect 58438 744912 58494 744968
rect 58530 744096 58586 744152
rect 57978 742348 58034 742384
rect 57978 742328 57980 742348
rect 57980 742328 58032 742348
rect 58032 742328 58034 742348
rect 58438 741784 58494 741840
rect 59634 729136 59690 729192
rect 59266 729000 59322 729056
rect 59450 728864 59506 728920
rect 50986 290672 51042 290728
rect 48594 289856 48650 289912
rect 47298 217086 47358 217146
rect 47390 216820 47450 216880
rect 47298 211620 47358 211680
rect 44778 211210 44834 211266
rect 47482 216544 47542 216604
rect 47482 213248 47542 213308
rect 47390 210806 47450 210866
rect 37830 210160 37886 210216
rect 31666 203632 31722 203688
rect 8206 202408 8262 202464
rect 30102 202408 30158 202464
rect 38014 209752 38070 209808
rect 37922 206896 37978 206952
rect 38290 209344 38346 209400
rect 38198 208936 38254 208992
rect 38106 208528 38162 208584
rect 38566 208120 38622 208176
rect 38382 207712 38438 207768
rect 38474 207304 38530 207360
rect 38382 204856 38438 204912
rect 38290 204448 38346 204504
rect 42706 206760 42762 206816
rect 42338 205128 42394 205184
rect 37830 198736 37886 198792
rect 43258 206352 43314 206408
rect 43074 205536 43130 205592
rect 43442 205944 43498 206000
rect 48226 204720 48282 204776
rect 41878 184184 41934 184240
rect 41786 183368 41842 183424
rect 41786 182688 41842 182744
rect 58530 702072 58586 702128
rect 59358 704384 59414 704440
rect 59266 703296 59322 703352
rect 59450 700848 59506 700904
rect 59634 699624 59690 699680
rect 59174 698128 59230 698184
rect 60646 661136 60702 661192
rect 58530 659504 58586 659560
rect 58438 658824 58494 658880
rect 58622 657600 58678 657656
rect 58990 656512 59046 656568
rect 58438 655288 58494 655344
rect 58162 617752 58218 617808
rect 58530 616800 58586 616856
rect 58530 615476 58532 615496
rect 58532 615476 58584 615496
rect 58584 615476 58586 615496
rect 58530 615440 58586 615476
rect 58162 614488 58218 614544
rect 57978 612584 58034 612640
rect 57978 612076 57980 612096
rect 57980 612076 58032 612096
rect 58032 612076 58034 612096
rect 57978 612040 58034 612076
rect 59266 599120 59322 599176
rect 58530 574776 58586 574832
rect 58714 570016 58770 570072
rect 59450 598984 59506 599040
rect 59358 573552 59414 573608
rect 60646 572328 60702 572384
rect 59450 571240 59506 571296
rect 59266 568520 59322 568576
rect 59450 531664 59506 531720
rect 59266 530576 59322 530632
rect 58530 529352 58586 529408
rect 58346 528128 58402 528184
rect 60646 527076 60648 527096
rect 60648 527076 60700 527096
rect 60700 527076 60702 527096
rect 60646 527040 60702 527076
rect 59358 525816 59414 525872
rect 59266 428032 59322 428088
rect 58162 404096 58218 404152
rect 58162 402908 58164 402928
rect 58164 402908 58216 402928
rect 58216 402908 58218 402928
rect 58162 402872 58218 402908
rect 58898 400696 58954 400752
rect 58162 399336 58218 399392
rect 59450 427896 59506 427952
rect 59266 400016 59322 400072
rect 59450 398248 59506 398304
rect 58162 360848 58218 360904
rect 58346 359760 58402 359816
rect 58622 357448 58678 357504
rect 58530 357312 58586 357368
rect 58070 355988 58072 356008
rect 58072 355988 58124 356008
rect 58124 355988 58126 356008
rect 58070 355952 58126 355988
rect 59358 355000 59414 355056
rect 58438 317328 58494 317384
rect 58162 316512 58218 316568
rect 58346 314744 58402 314800
rect 58162 312976 58218 313032
rect 58530 314064 58586 314120
rect 58530 311788 58532 311808
rect 58532 311788 58584 311808
rect 58584 311788 58586 311808
rect 58530 311752 58586 311788
rect 58438 298152 58494 298208
rect 58346 293936 58402 293992
rect 58530 295432 58586 295488
rect 59450 292712 59506 292768
rect 58438 292440 58494 292496
rect 57886 291488 57942 291544
rect 58530 289756 58532 289776
rect 58532 289756 58584 289776
rect 58584 289756 58586 289776
rect 58530 289720 58586 289756
rect 57978 287952 58034 288008
rect 58530 287136 58586 287192
rect 56046 227568 56102 227624
rect 54390 222128 54446 222184
rect 57978 285640 58034 285696
rect 58530 284416 58586 284472
rect 57978 283192 58034 283248
rect 59266 282104 59322 282160
rect 57610 227704 57666 227760
rect 56874 224848 56930 224904
rect 58622 224984 58678 225040
rect 59174 222264 59230 222320
rect 59358 279656 59414 279712
rect 61842 291080 61898 291136
rect 59542 280880 59598 280936
rect 61106 222400 61162 222456
rect 655426 778368 655482 778424
rect 654966 773472 655022 773528
rect 655150 730224 655206 730280
rect 655610 777008 655666 777064
rect 655518 775512 655574 775568
rect 655518 731448 655574 731504
rect 655426 687248 655482 687304
rect 654230 685752 654286 685808
rect 654138 684392 654194 684448
rect 654414 639376 654470 639432
rect 655794 775920 655850 775976
rect 655702 734304 655758 734360
rect 655610 689424 655666 689480
rect 655518 643184 655574 643240
rect 655426 595312 655482 595368
rect 656530 774696 656586 774752
rect 655886 732672 655942 732728
rect 655794 688200 655850 688256
rect 655702 640192 655758 640248
rect 655978 731312 656034 731368
rect 656070 728592 656126 728648
rect 655978 686976 656034 687032
rect 655978 641824 656034 641880
rect 655886 597760 655942 597816
rect 655702 596536 655758 596592
rect 655610 593000 655666 593056
rect 655610 553288 655666 553344
rect 655426 552064 655482 552120
rect 654230 549208 654286 549264
rect 654138 548528 654194 548584
rect 655518 550976 655574 551032
rect 655794 595448 655850 595504
rect 656162 640600 656218 640656
rect 656438 638152 656494 638208
rect 656806 594224 656862 594280
rect 655978 550840 656034 550896
rect 655702 374448 655758 374504
rect 655518 373224 655574 373280
rect 655426 372136 655482 372192
rect 654506 370912 654562 370968
rect 655518 329840 655574 329896
rect 655610 328208 655666 328264
rect 655426 327392 655482 327448
rect 655978 325624 656034 325680
rect 655518 303320 655574 303376
rect 655702 302096 655758 302152
rect 655426 300736 655482 300792
rect 655058 298696 655114 298752
rect 656162 297472 656218 297528
rect 655794 296248 655850 296304
rect 655610 293936 655666 293992
rect 655426 292712 655482 292768
rect 654138 289176 654194 289232
rect 654138 287952 654194 288008
rect 655242 285640 655298 285696
rect 654506 284708 654562 284744
rect 654506 284688 654508 284708
rect 654508 284688 654560 284708
rect 654560 284688 654562 284708
rect 654230 283600 654286 283656
rect 655242 282104 655298 282160
rect 654138 280880 654194 280936
rect 654874 279656 654930 279712
rect 63406 275984 63462 276040
rect 62670 227840 62726 227896
rect 63314 225120 63370 225176
rect 70582 271904 70638 271960
rect 69386 271768 69442 271824
rect 71778 269048 71834 269104
rect 80058 272312 80114 272368
rect 81254 272040 81310 272096
rect 83646 272176 83702 272232
rect 85946 269728 86002 269784
rect 84750 269592 84806 269648
rect 78862 269456 78918 269512
rect 88338 272584 88394 272640
rect 90730 272448 90786 272504
rect 93030 269864 93086 269920
rect 96618 272856 96674 272912
rect 99010 272720 99066 272776
rect 101310 270136 101366 270192
rect 100114 270000 100170 270056
rect 103702 272992 103758 273048
rect 106094 273128 106150 273184
rect 107198 270272 107254 270328
rect 111982 271632 112038 271688
rect 110786 271360 110842 271416
rect 115478 271496 115534 271552
rect 77666 269320 77722 269376
rect 76470 269184 76526 269240
rect 117870 271224 117926 271280
rect 120262 270408 120318 270464
rect 122562 271088 122618 271144
rect 128542 268912 128598 268968
rect 146206 268776 146262 268832
rect 150990 268640 151046 268696
rect 158074 268504 158130 268560
rect 159270 268368 159326 268424
rect 194138 271904 194194 271960
rect 193678 271768 193734 271824
rect 194598 269048 194654 269104
rect 196898 272312 196954 272368
rect 196806 269320 196862 269376
rect 196346 269184 196402 269240
rect 195978 268232 196034 268288
rect 198094 272040 198150 272096
rect 197726 269456 197782 269512
rect 199106 272176 199162 272232
rect 199014 269592 199070 269648
rect 199934 269728 199990 269784
rect 201222 272584 201278 272640
rect 201682 272448 201738 272504
rect 202142 268232 202198 268288
rect 203062 269864 203118 269920
rect 204350 272856 204406 272912
rect 204810 272720 204866 272776
rect 205270 270136 205326 270192
rect 205730 270000 205786 270056
rect 207478 273128 207534 273184
rect 207018 272992 207074 273048
rect 208398 270272 208454 270328
rect 209226 271632 209282 271688
rect 209686 271360 209742 271416
rect 210606 271496 210662 271552
rect 212354 271224 212410 271280
rect 213274 271088 213330 271144
rect 212814 270408 212870 270464
rect 216402 268912 216458 268968
rect 221738 268776 221794 268832
rect 223946 268640 224002 268696
rect 226614 268504 226670 268560
rect 227534 268368 227590 268424
rect 353022 271088 353078 271144
rect 352194 268368 352250 268424
rect 353942 268504 353998 268560
rect 355322 271224 355378 271280
rect 354862 268640 354918 268696
rect 357530 268912 357586 268968
rect 356610 268776 356666 268832
rect 357990 271360 358046 271416
rect 358910 271496 358966 271552
rect 361026 271632 361082 271688
rect 362866 270408 362922 270464
rect 362038 270272 362094 270328
rect 364062 273128 364118 273184
rect 365534 270136 365590 270192
rect 365994 268232 366050 268288
rect 366914 272992 366970 273048
rect 368662 272856 368718 272912
rect 369674 272720 369730 272776
rect 370042 270000 370098 270056
rect 370870 269864 370926 269920
rect 372618 272584 372674 272640
rect 372434 272448 372490 272504
rect 372066 268232 372122 268288
rect 376666 269728 376722 269784
rect 380714 272312 380770 272368
rect 382002 269592 382058 269648
rect 386970 267144 387026 267200
rect 389638 267008 389694 267064
rect 390466 266872 390522 266928
rect 391386 269456 391442 269512
rect 391846 266736 391902 266792
rect 393594 274216 393650 274272
rect 393134 266600 393190 266656
rect 395434 272176 395490 272232
rect 394514 266464 394570 266520
rect 396262 275712 396318 275768
rect 395802 274352 395858 274408
rect 397366 275848 397422 275904
rect 398930 275576 398986 275632
rect 398470 275440 398526 275496
rect 397642 267416 397698 267472
rect 399850 275168 399906 275224
rect 401138 275304 401194 275360
rect 401966 275032 402022 275088
rect 402518 274896 402574 274952
rect 405186 274760 405242 274816
rect 403438 269320 403494 269376
rect 402978 267552 403034 267608
rect 404726 272040 404782 272096
rect 408314 274624 408370 274680
rect 407854 274488 407910 274544
rect 406106 269184 406162 269240
rect 405646 267688 405702 267744
rect 406934 267280 406990 267336
rect 410522 271904 410578 271960
rect 410062 271768 410118 271824
rect 410982 269048 411038 269104
rect 441802 267688 441858 267744
rect 455970 267552 456026 267608
rect 472530 267416 472586 267472
rect 485042 267280 485098 267336
rect 491390 271088 491446 271144
rect 494886 268504 494942 268560
rect 490194 268368 490250 268424
rect 498474 271224 498530 271280
rect 497278 268640 497334 268696
rect 501970 268776 502026 268832
rect 507950 271496 508006 271552
rect 505558 271360 505614 271416
rect 504362 268912 504418 268968
rect 512642 271632 512698 271688
rect 516230 270272 516286 270328
rect 522118 273128 522174 273184
rect 518530 270408 518586 270464
rect 529202 272992 529258 273048
rect 525614 270136 525670 270192
rect 533894 272856 533950 272912
rect 536286 272720 536342 272776
rect 537482 270000 537538 270056
rect 540978 272584 541034 272640
rect 543370 272448 543426 272504
rect 539874 269864 539930 269920
rect 555238 269728 555294 269784
rect 565818 272312 565874 272368
rect 569406 269592 569462 269648
rect 582378 267144 582434 267200
rect 589462 267008 589518 267064
rect 594246 269456 594302 269512
rect 591854 266872 591910 266928
rect 595350 266736 595406 266792
rect 600134 274216 600190 274272
rect 598938 266600 598994 266656
rect 607218 275712 607274 275768
rect 606022 274352 606078 274408
rect 604826 272176 604882 272232
rect 609610 275848 609666 275904
rect 614302 275576 614358 275632
rect 613106 275440 613162 275496
rect 616694 275168 616750 275224
rect 620190 275304 620246 275360
rect 621386 275032 621442 275088
rect 623778 274896 623834 274952
rect 630862 274760 630918 274816
rect 629666 272040 629722 272096
rect 626078 269320 626134 269376
rect 639142 274624 639198 274680
rect 637946 274488 638002 274544
rect 633254 269184 633310 269240
rect 645030 271904 645086 271960
rect 643834 271768 643890 271824
rect 646226 269048 646282 269104
rect 602434 266464 602490 266520
rect 184938 258576 184994 258632
rect 416778 252728 416834 252784
rect 416778 249464 416834 249520
rect 184938 247968 184994 248024
rect 416778 246336 416834 246392
rect 418066 243072 418122 243128
rect 184938 237396 184940 237416
rect 184940 237396 184992 237416
rect 184992 237396 184994 237416
rect 184938 237360 184994 237396
rect 84658 228928 84714 228984
rect 82726 228520 82782 228576
rect 77942 228384 77998 228440
rect 76286 228248 76342 228304
rect 71226 228112 71282 228168
rect 64510 227976 64566 228032
rect 66166 222672 66222 222728
rect 67822 222536 67878 222592
rect 70398 225256 70454 225312
rect 72882 222944 72938 223000
rect 74446 222808 74502 222864
rect 77114 225392 77170 225448
rect 80426 225528 80482 225584
rect 79598 223080 79654 223136
rect 83830 225664 83886 225720
rect 88062 228792 88118 228848
rect 86314 228656 86370 228712
rect 93030 227432 93086 227488
rect 94778 227296 94834 227352
rect 101494 227160 101550 227216
rect 99838 227024 99894 227080
rect 98918 225936 98974 225992
rect 96434 223216 96490 223272
rect 98090 223352 98146 223408
rect 106554 226888 106610 226944
rect 103978 226072 104034 226128
rect 102046 225800 102102 225856
rect 103150 223488 103206 223544
rect 104806 221992 104862 222048
rect 113086 226752 113142 226808
rect 109038 226208 109094 226264
rect 109866 221856 109922 221912
rect 112442 224712 112498 224768
rect 111614 221720 111670 221776
rect 115754 224576 115810 224632
rect 117502 224440 117558 224496
rect 118330 221312 118386 221368
rect 120814 224304 120870 224360
rect 119986 221584 120042 221640
rect 121366 221448 121422 221504
rect 160098 224168 160154 224224
rect 172426 224032 172482 224088
rect 194782 227704 194838 227760
rect 194414 227568 194470 227624
rect 194046 224984 194102 225040
rect 193678 224848 193734 224904
rect 193310 222128 193366 222184
rect 195794 222264 195850 222320
rect 197634 227976 197690 228032
rect 197266 227840 197322 227896
rect 196530 225120 196586 225176
rect 196162 222400 196218 222456
rect 198646 222672 198702 222728
rect 200486 228112 200542 228168
rect 199382 225256 199438 225312
rect 199014 222536 199070 222592
rect 201682 226480 201738 226536
rect 201498 222944 201554 223000
rect 203338 228384 203394 228440
rect 202970 228248 203026 228304
rect 202234 225392 202290 225448
rect 201866 222808 201922 222864
rect 203706 225528 203762 225584
rect 204350 223080 204406 223136
rect 205086 225664 205142 225720
rect 206190 228928 206246 228984
rect 205822 228520 205878 228576
rect 207018 228928 207074 228984
rect 207570 228792 207626 228848
rect 207202 228656 207258 228712
rect 206558 224032 206614 224088
rect 208674 226480 208730 226536
rect 207938 224168 207994 224224
rect 210054 227432 210110 227488
rect 210790 228928 210846 228984
rect 210790 227568 210846 227624
rect 210422 227296 210478 227352
rect 211158 225936 211214 225992
rect 211526 223216 211582 223272
rect 212354 227704 212410 227760
rect 211894 223352 211950 223408
rect 213274 227160 213330 227216
rect 212906 227024 212962 227080
rect 213642 226072 213698 226128
rect 212538 225800 212594 225856
rect 214378 223488 214434 223544
rect 215758 226888 215814 226944
rect 215390 226208 215446 226264
rect 214746 221992 214802 222048
rect 216862 224712 216918 224768
rect 217230 221856 217286 221912
rect 217598 227840 217654 227896
rect 217322 221720 217378 221776
rect 219254 228112 219310 228168
rect 218610 226752 218666 226808
rect 218242 224576 218298 224632
rect 219346 224440 219402 224496
rect 220726 227976 220782 228032
rect 220450 221312 220506 221368
rect 220818 224304 220874 224360
rect 221462 221584 221518 221640
rect 221830 221448 221886 221504
rect 225970 228248 226026 228304
rect 236734 228384 236790 228440
rect 237010 228520 237066 228576
rect 245658 228792 245714 228848
rect 259182 227024 259238 227080
rect 259642 228520 259698 228576
rect 260378 227704 260434 227760
rect 260010 227568 260066 227624
rect 261390 228792 261446 228848
rect 261758 227024 261814 227080
rect 262494 228384 262550 228440
rect 263230 228112 263286 228168
rect 262862 227840 262918 227896
rect 264242 227976 264298 228032
rect 266082 228248 266138 228304
rect 330942 222672 330998 222728
rect 332322 222536 332378 222592
rect 333058 222400 333114 222456
rect 333794 222264 333850 222320
rect 334530 221584 334586 221640
rect 335910 222128 335966 222184
rect 335818 221720 335874 221776
rect 338762 221856 338818 221912
rect 369398 224304 369454 224360
rect 370870 224440 370926 224496
rect 372250 224712 372306 224768
rect 373722 224576 373778 224632
rect 375102 223488 375158 223544
rect 375838 221992 375894 222048
rect 376942 227024 376998 227080
rect 377310 227160 377366 227216
rect 378322 223352 378378 223408
rect 378690 223216 378746 223272
rect 379794 227432 379850 227488
rect 380162 227296 380218 227352
rect 381174 223080 381230 223136
rect 381542 222808 381598 222864
rect 381082 222672 381138 222728
rect 382646 228792 382702 228848
rect 383658 222944 383714 223000
rect 383658 222400 383714 222456
rect 384762 228928 384818 228984
rect 384302 222536 384358 222592
rect 385866 222672 385922 222728
rect 386878 228656 386934 228712
rect 387982 222536 388038 222592
rect 387706 222264 387762 222320
rect 386786 221584 386842 221640
rect 388994 222400 389050 222456
rect 388534 221720 388590 221776
rect 390098 228520 390154 228576
rect 389362 226072 389418 226128
rect 390466 225936 390522 225992
rect 390190 222128 390246 222184
rect 391570 225800 391626 225856
rect 392214 228384 392270 228440
rect 391202 222264 391258 222320
rect 392582 225664 392638 225720
rect 394422 228248 394478 228304
rect 394790 225528 394846 225584
rect 393318 222128 393374 222184
rect 396538 228112 396594 228168
rect 397366 226208 397422 226264
rect 396906 221856 396962 221912
rect 397918 225392 397974 225448
rect 398654 227976 398710 228032
rect 399758 227840 399814 227896
rect 401138 225256 401194 225312
rect 403990 227704 404046 227760
rect 405462 225120 405518 225176
rect 406474 224984 406530 225040
rect 411166 227568 411222 227624
rect 410798 224848 410854 224904
rect 418158 239944 418214 240000
rect 63406 217232 63462 217288
rect 418434 236680 418490 236736
rect 418526 233552 418582 233608
rect 471978 224304 472034 224360
rect 475106 224440 475162 224496
rect 478510 224712 478566 224768
rect 481914 224576 481970 224632
rect 483846 223488 483902 223544
rect 486330 221992 486386 222048
rect 507398 228928 507454 228984
rect 503810 228792 503866 228848
rect 489734 227160 489790 227216
rect 488906 227024 488962 227080
rect 491942 223352 491998 223408
rect 491390 223216 491446 223272
rect 491390 220904 491446 220960
rect 493046 220904 493102 220960
rect 495346 227432 495402 227488
rect 496174 227296 496230 227352
rect 495346 221176 495402 221232
rect 498658 223080 498714 223136
rect 500222 222808 500278 222864
rect 500222 221040 500278 221096
rect 504822 222944 504878 223000
rect 512182 228656 512238 228712
rect 509606 222672 509662 222728
rect 507398 221312 507454 221368
rect 518990 228520 519046 228576
rect 513470 226208 513526 226264
rect 518714 226072 518770 226128
rect 514666 222536 514722 222592
rect 517058 222400 517114 222456
rect 525062 228384 525118 228440
rect 520830 225936 520886 225992
rect 523406 225800 523462 225856
rect 522210 222264 522266 222320
rect 525798 225664 525854 225720
rect 527270 222128 527326 222184
rect 530122 228248 530178 228304
rect 534906 228112 534962 228168
rect 530674 225528 530730 225584
rect 538310 227976 538366 228032
rect 542726 227840 542782 227896
rect 538862 225392 538918 225448
rect 545762 225256 545818 225312
rect 552570 227704 552626 227760
rect 556066 225120 556122 225176
rect 559102 224984 559158 225040
rect 564346 221720 564402 221776
rect 564530 221448 564586 221504
rect 569314 227568 569370 227624
rect 568578 224848 568634 224904
rect 567106 221584 567162 221640
rect 574374 221584 574430 221640
rect 573546 221448 573602 221504
rect 575202 221448 575258 221504
rect 582286 216144 582342 216200
rect 582286 214648 582342 214704
rect 580262 213152 580318 213208
rect 580078 211656 580134 211712
rect 582286 210160 582342 210216
rect 581458 208664 581514 208720
rect 622490 221176 622546 221232
rect 624330 221312 624386 221368
rect 637854 221040 637910 221096
rect 636934 220904 636990 220960
rect 652758 217232 652814 217288
rect 655518 291488 655574 291544
rect 655702 290400 655758 290456
rect 655978 295296 656034 295352
rect 656806 287292 656862 287328
rect 656806 287272 656808 287292
rect 656808 287272 656860 287292
rect 656860 287272 656862 287292
rect 600042 209480 600098 209536
rect 599950 208528 600006 208584
rect 599858 207440 599914 207496
rect 582286 207068 582288 207088
rect 582288 207068 582340 207088
rect 582340 207068 582342 207088
rect 582286 207032 582342 207068
rect 582286 205536 582342 205592
rect 580722 204040 580778 204096
rect 600778 206488 600834 206544
rect 666558 209208 666614 209264
rect 601146 205400 601202 205456
rect 666558 205808 666614 205864
rect 601606 204448 601662 204504
rect 599674 203360 599730 203416
rect 581090 202544 581146 202600
rect 666558 204176 666614 204232
rect 599950 202408 600006 202464
rect 598938 201320 598994 201376
rect 581090 201048 581146 201104
rect 666558 200776 666614 200832
rect 599950 200368 600006 200424
rect 582286 199552 582342 199608
rect 599950 199280 600006 199336
rect 666558 199008 666614 199064
rect 599950 198328 600006 198384
rect 582286 197920 582342 197976
rect 580722 196424 580778 196480
rect 599950 197276 599952 197296
rect 599952 197276 600004 197296
rect 600004 197276 600006 197296
rect 599950 197240 600006 197276
rect 599398 196288 599454 196344
rect 666558 195608 666614 195664
rect 599858 195200 599914 195256
rect 582286 194928 582342 194984
rect 599950 194248 600006 194304
rect 582194 193432 582250 193488
rect 599490 193160 599546 193216
rect 582286 191936 582342 191992
rect 599950 192208 600006 192264
rect 599950 191120 600006 191176
rect 581274 190440 581330 190496
rect 601514 190168 601570 190224
rect 579710 188808 579766 188864
rect 599122 188128 599178 188184
rect 582286 187312 582342 187368
rect 579894 185816 579950 185872
rect 601606 189080 601662 189136
rect 666558 188944 666614 189000
rect 599950 187040 600006 187096
rect 599858 185000 599914 185056
rect 580906 184320 580962 184376
rect 598938 182960 598994 183016
rect 580262 182824 580318 182880
rect 580630 181328 580686 181384
rect 580538 179696 580594 179752
rect 600042 186088 600098 186144
rect 599950 184048 600006 184104
rect 599858 179968 599914 180024
rect 599674 178880 599730 178936
rect 581090 178200 581146 178256
rect 580722 176704 580778 176760
rect 579710 172216 579766 172272
rect 580538 170584 580594 170640
rect 580170 166096 580226 166152
rect 579894 161472 579950 161528
rect 579802 158480 579858 158536
rect 581458 175208 581514 175264
rect 581090 167592 581146 167648
rect 580446 156984 580502 157040
rect 580262 155488 580318 155544
rect 580078 149368 580134 149424
rect 580630 143248 580686 143304
rect 580538 138760 580594 138816
rect 579710 112920 579766 112976
rect 580722 135768 580778 135824
rect 579894 111424 579950 111480
rect 580078 108432 580134 108488
rect 582286 173748 582288 173768
rect 582288 173748 582340 173768
rect 582340 173748 582342 173768
rect 582286 173712 582342 173748
rect 599490 172760 599546 172816
rect 582010 169088 582066 169144
rect 599766 177928 599822 177984
rect 666558 185544 666614 185600
rect 666558 183776 666614 183832
rect 600042 182008 600098 182064
rect 599950 176840 600006 176896
rect 600134 180920 600190 180976
rect 599950 174800 600006 174856
rect 666558 180376 666614 180432
rect 600410 175888 600466 175944
rect 599950 171808 600006 171864
rect 599858 170720 599914 170776
rect 599490 168680 599546 168736
rect 599950 169768 600006 169824
rect 601330 173848 601386 173904
rect 581642 164600 581698 164656
rect 581826 163104 581882 163160
rect 581274 153992 581330 154048
rect 581182 147872 581238 147928
rect 581090 141752 581146 141808
rect 580906 137264 580962 137320
rect 580814 132640 580870 132696
rect 580170 106800 580226 106856
rect 579986 105304 580042 105360
rect 580262 103808 580318 103864
rect 580354 100816 580410 100872
rect 580446 97688 580502 97744
rect 187606 41792 187662 41848
rect 209778 41248 209834 41304
rect 212446 41248 212502 41304
rect 216126 48184 216182 48240
rect 230386 10648 230442 10704
rect 230754 15136 230810 15192
rect 230662 13640 230718 13696
rect 230938 16632 230994 16688
rect 230846 12144 230902 12200
rect 230570 9152 230626 9208
rect 230478 7656 230534 7712
rect 307298 43152 307354 43208
rect 416594 43424 416650 43480
rect 415398 43288 415454 43344
rect 470138 43560 470194 43616
rect 361946 41792 362002 41848
rect 419998 41792 420054 41848
rect 427910 41792 427966 41848
rect 471702 41792 471758 41848
rect 427910 41112 427966 41168
rect 475474 40976 475530 41032
rect 521750 42064 521806 42120
rect 513286 41792 513342 41848
rect 518530 41792 518586 41848
rect 530306 41284 530308 41304
rect 530308 41284 530360 41304
rect 530360 41284 530362 41304
rect 530306 41248 530362 41284
rect 530398 41112 530454 41168
rect 568578 41384 568634 41440
rect 580630 99320 580686 99376
rect 580722 96192 580778 96248
rect 580538 94696 580594 94752
rect 580998 117544 581054 117600
rect 580906 102312 580962 102368
rect 580814 91704 580870 91760
rect 579618 82628 579620 82648
rect 579620 82628 579672 82648
rect 579672 82628 579674 82648
rect 579618 82592 579674 82628
rect 580722 68856 580778 68912
rect 579618 65864 579674 65920
rect 580814 62872 580870 62928
rect 581366 126656 581422 126712
rect 599490 167728 599546 167784
rect 582010 159976 582066 160032
rect 581734 146376 581790 146432
rect 581642 144880 581698 144936
rect 581550 125024 581606 125080
rect 581458 123528 581514 123584
rect 581274 120536 581330 120592
rect 581182 114416 581238 114472
rect 581090 109928 581146 109984
rect 580998 70352 581054 70408
rect 581274 79464 581330 79520
rect 581826 131144 581882 131200
rect 581734 119040 581790 119096
rect 581642 115912 581698 115968
rect 581458 81096 581514 81152
rect 581366 76472 581422 76528
rect 600042 166640 600098 166696
rect 599950 165708 600006 165744
rect 599950 165688 599952 165708
rect 599952 165688 600004 165708
rect 600004 165688 600006 165708
rect 666558 173576 666614 173632
rect 666558 170176 666614 170232
rect 600042 164600 600098 164656
rect 599950 163648 600006 163704
rect 600042 162560 600098 162616
rect 599858 161608 599914 161664
rect 599950 160520 600006 160576
rect 599858 159568 599914 159624
rect 600042 158480 600098 158536
rect 599950 157528 600006 157584
rect 599858 156440 599914 156496
rect 599950 155488 600006 155544
rect 599858 154400 599914 154456
rect 582286 152360 582342 152416
rect 600042 153448 600098 153504
rect 599950 152360 600006 152416
rect 582194 150864 582250 150920
rect 582102 140256 582158 140312
rect 582010 129648 582066 129704
rect 600042 151408 600098 151464
rect 599858 150320 599914 150376
rect 599950 149368 600006 149424
rect 599858 148280 599914 148336
rect 599950 147328 600006 147384
rect 599858 146240 599914 146296
rect 600042 145288 600098 145344
rect 599950 144200 600006 144256
rect 600042 143248 600098 143304
rect 599950 142160 600006 142216
rect 599858 141208 599914 141264
rect 600042 140120 600098 140176
rect 599858 139168 599914 139224
rect 599950 138116 599952 138136
rect 599952 138116 600004 138136
rect 600004 138116 600006 138136
rect 599950 138080 600006 138116
rect 599858 137128 599914 137184
rect 599950 136040 600006 136096
rect 600042 135088 600098 135144
rect 582286 134136 582342 134192
rect 599858 134000 599914 134056
rect 599950 133048 600006 133104
rect 600042 131960 600098 132016
rect 599858 131008 599914 131064
rect 599950 129920 600006 129976
rect 599858 128968 599914 129024
rect 582194 128152 582250 128208
rect 599950 127880 600006 127936
rect 599858 126928 599914 126984
rect 599766 124888 599822 124944
rect 581918 122032 581974 122088
rect 581826 90208 581882 90264
rect 581734 77968 581790 78024
rect 581642 74976 581698 75032
rect 581550 71984 581606 72040
rect 581182 67360 581238 67416
rect 581090 64368 581146 64424
rect 582102 88576 582158 88632
rect 582010 87080 582066 87136
rect 599950 125840 600006 125896
rect 600042 123800 600098 123856
rect 599858 122848 599914 122904
rect 599950 121760 600006 121816
rect 600042 120808 600098 120864
rect 599950 119720 600006 119776
rect 582286 93200 582342 93256
rect 582194 85584 582250 85640
rect 581918 84088 581974 84144
rect 581826 56752 581882 56808
rect 582194 61240 582250 61296
rect 582102 59744 582158 59800
rect 599858 118768 599914 118824
rect 600042 117680 600098 117736
rect 599950 116728 600006 116784
rect 599858 115640 599914 115696
rect 599950 114688 600006 114744
rect 599858 112648 599914 112704
rect 599950 111560 600006 111616
rect 600226 110608 600282 110664
rect 599306 109520 599362 109576
rect 599950 107480 600006 107536
rect 599950 100408 600006 100464
rect 582286 58248 582342 58304
rect 582010 55256 582066 55312
rect 580906 53760 580962 53816
rect 600318 108568 600374 108624
rect 600594 106528 600650 106584
rect 600410 105440 600466 105496
rect 600502 102448 600558 102504
rect 600870 104488 600926 104544
rect 600686 103400 600742 103456
rect 600778 101360 600834 101416
rect 575846 43560 575902 43616
rect 577962 43424 578018 43480
rect 586426 43288 586482 43344
rect 575662 43152 575718 43208
rect 622490 87896 622546 87952
rect 623226 88848 623282 88904
rect 623410 86944 623466 87000
rect 628286 95920 628342 95976
rect 640522 95684 640524 95704
rect 640524 95684 640576 95704
rect 640576 95684 640578 95704
rect 640522 95648 640578 95684
rect 627918 94424 627974 94480
rect 627274 93472 627330 93528
rect 626446 92520 626502 92576
rect 625894 91568 625950 91624
rect 623962 90616 624018 90672
rect 623778 89664 623834 89720
rect 623502 85992 623558 86048
rect 623318 85040 623374 85096
rect 623134 84088 623190 84144
rect 622122 83136 622178 83192
rect 622306 82184 622362 82240
rect 622490 81368 622546 81424
rect 642730 92656 642786 92712
rect 645858 89664 645914 89720
rect 646042 87080 646098 87136
rect 653954 92520 654010 92576
rect 655334 93336 655390 93392
rect 654046 91432 654102 91488
rect 653126 90616 653182 90672
rect 656990 90344 657046 90400
rect 662234 95512 662290 95568
rect 657358 94696 657414 94752
rect 663246 93744 663302 93800
rect 663430 93064 663486 93120
rect 663522 92248 663578 92304
rect 662142 88712 662198 88768
rect 663522 91024 663578 91080
rect 663614 90344 663670 90400
rect 663430 89528 663486 89584
rect 646134 84632 646190 84688
rect 645950 82184 646006 82240
rect 661130 47504 661186 47560
rect 666742 168544 666798 168600
rect 666742 165144 666798 165200
rect 666742 163512 666798 163568
rect 666742 160112 666798 160168
rect 666742 158344 666798 158400
rect 666742 154944 666798 155000
rect 666742 153312 666798 153368
rect 666742 149912 666798 149968
rect 666742 148144 666798 148200
rect 666742 144880 666798 144936
rect 666742 143112 666798 143168
rect 666742 139712 666798 139768
rect 666742 132912 666798 132968
rect 666742 129512 666798 129568
rect 666650 127880 666706 127936
rect 666650 124480 666706 124536
rect 666650 122848 666706 122904
rect 666650 119448 666706 119504
rect 667110 205944 667166 206000
rect 671894 217096 671950 217152
rect 670698 193976 670754 194032
rect 670698 190576 670754 190632
rect 670698 178744 670754 178800
rect 670698 175344 670754 175400
rect 670698 138080 670754 138136
rect 670698 134680 670754 134736
rect 676034 896280 676090 896336
rect 676126 895192 676182 895248
rect 676034 893852 676090 893888
rect 676034 893832 676036 893852
rect 676036 893832 676088 893852
rect 676088 893832 676090 893852
rect 676034 893036 676090 893072
rect 676034 893016 676036 893036
rect 676036 893016 676088 893036
rect 676088 893016 676090 893036
rect 679622 892608 679678 892664
rect 676034 892200 676090 892256
rect 679346 891792 679402 891848
rect 679162 891384 679218 891440
rect 676034 890976 676090 891032
rect 676034 890568 676090 890624
rect 675942 888936 675998 888992
rect 678978 890160 679034 890216
rect 676034 888528 676090 888584
rect 676034 887712 676090 887768
rect 675942 887304 675998 887360
rect 679070 888120 679126 888176
rect 679254 889752 679310 889808
rect 679438 889344 679494 889400
rect 679530 884992 679586 885048
rect 675114 788296 675170 788352
rect 675114 787208 675170 787264
rect 675114 786664 675170 786720
rect 671986 178744 672042 178800
rect 673826 745320 673882 745376
rect 672078 173576 672134 173632
rect 672170 168544 672226 168600
rect 674562 745184 674618 745240
rect 674746 734848 674802 734904
rect 674286 687112 674342 687168
rect 672262 163512 672318 163568
rect 673550 554648 673606 554704
rect 672354 158344 672410 158400
rect 675390 742872 675446 742928
rect 675390 742464 675446 742520
rect 675482 741648 675538 741704
rect 675390 739744 675446 739800
rect 675390 739064 675446 739120
rect 675390 738656 675446 738712
rect 675390 737976 675446 738032
rect 675206 733352 675262 733408
rect 675482 699352 675538 699408
rect 675758 716488 675814 716544
rect 675850 716080 675906 716136
rect 675942 715672 675998 715728
rect 676034 715264 676090 715320
rect 676034 714876 676090 714912
rect 676034 714856 676036 714876
rect 676036 714856 676088 714876
rect 676088 714856 676090 714876
rect 676034 714484 676036 714504
rect 676036 714484 676088 714504
rect 676088 714484 676090 714504
rect 676034 714448 676090 714484
rect 676034 714060 676090 714096
rect 676034 714040 676036 714060
rect 676036 714040 676088 714060
rect 676088 714040 676090 714060
rect 676034 713632 676090 713688
rect 675850 713224 675906 713280
rect 675942 712816 675998 712872
rect 676034 712408 676090 712464
rect 676034 711592 676090 711648
rect 676034 710776 676090 710832
rect 675942 710368 675998 710424
rect 678978 709960 679034 710016
rect 675758 709144 675814 709200
rect 675666 708736 675722 708792
rect 676034 708328 676090 708384
rect 676034 707920 676090 707976
rect 676034 707512 676090 707568
rect 676034 706288 676090 706344
rect 676034 705100 676036 705120
rect 676036 705100 676088 705120
rect 676088 705100 676090 705120
rect 676034 705064 676090 705100
rect 675574 699216 675630 699272
rect 675114 698264 675170 698320
rect 675758 697176 675814 697232
rect 675114 695544 675170 695600
rect 675114 694728 675170 694784
rect 675114 694592 675170 694648
rect 675758 692960 675814 693016
rect 675758 690104 675814 690160
rect 675206 685752 675262 685808
rect 674286 571512 674342 571568
rect 674654 610136 674710 610192
rect 676126 677912 676182 677968
rect 676126 676416 676182 676472
rect 676218 671064 676274 671120
rect 676034 670928 676090 670984
rect 678978 670248 679034 670304
rect 676126 669840 676182 669896
rect 676034 669332 676036 669352
rect 676036 669332 676088 669352
rect 676088 669332 676090 669352
rect 676034 669296 676090 669332
rect 676310 669432 676366 669488
rect 676218 668208 676274 668264
rect 675298 668072 675354 668128
rect 678978 667392 679034 667448
rect 676218 666984 676274 667040
rect 676034 666032 676090 666088
rect 676034 665216 676090 665272
rect 679162 678816 679218 678872
rect 679162 666984 679218 667040
rect 679070 666576 679126 666632
rect 676126 664944 676182 665000
rect 676034 664400 676090 664456
rect 676034 663176 676090 663232
rect 676034 662768 676090 662824
rect 678978 660864 679034 660920
rect 678978 660048 679034 660104
rect 675390 652840 675446 652896
rect 675482 652160 675538 652216
rect 675390 651616 675446 651672
rect 675390 649168 675446 649224
rect 675390 638424 675446 638480
rect 675298 610000 675354 610056
rect 675666 638152 675722 638208
rect 678978 626048 679034 626104
rect 676310 625640 676366 625696
rect 676034 625504 676090 625560
rect 675942 623872 675998 623928
rect 676218 624824 676274 624880
rect 676126 624416 676182 624472
rect 675942 623464 675998 623520
rect 676126 622784 676182 622840
rect 676034 621424 676090 621480
rect 676310 622376 676366 622432
rect 676218 621968 676274 622024
rect 676034 620200 676090 620256
rect 679070 619928 679126 619984
rect 676034 618568 676090 618624
rect 676034 618196 676036 618216
rect 676036 618196 676088 618216
rect 676088 618196 676090 618216
rect 676034 618160 676090 618196
rect 676034 617752 676090 617808
rect 676218 616700 676220 616720
rect 676220 616700 676272 616720
rect 676272 616700 676274 616720
rect 676218 616664 676274 616700
rect 679070 615848 679126 615904
rect 679070 615032 679126 615088
rect 675298 608096 675354 608152
rect 675298 607280 675354 607336
rect 675298 605104 675354 605160
rect 675206 604968 675262 605024
rect 675206 604424 675262 604480
rect 675206 601840 675262 601896
rect 676126 580896 676182 580952
rect 676310 580488 676366 580544
rect 676218 580100 676274 580136
rect 676218 580080 676220 580100
rect 676220 580080 676272 580100
rect 676272 580080 676274 580100
rect 676218 579692 676274 579728
rect 676218 579672 676220 579692
rect 676220 579672 676272 579692
rect 676272 579672 676274 579692
rect 676034 579028 676036 579048
rect 676036 579028 676088 579048
rect 676088 579028 676090 579048
rect 676034 578992 676090 579028
rect 676218 578468 676274 578504
rect 676218 578448 676220 578468
rect 676220 578448 676272 578468
rect 676272 578448 676274 578468
rect 676126 578040 676182 578096
rect 676218 577224 676274 577280
rect 676034 576136 676090 576192
rect 675942 575320 675998 575376
rect 678978 575184 679034 575240
rect 676034 574504 676090 574560
rect 675574 573280 675630 573336
rect 676034 572872 676090 572928
rect 676034 572464 676090 572520
rect 676034 572056 676090 572112
rect 678978 570696 679034 570752
rect 678978 569880 679034 569936
rect 675482 562672 675538 562728
rect 675298 562264 675354 562320
rect 675482 561176 675538 561232
rect 675298 554920 675354 554976
rect 677506 546488 677562 546544
rect 675390 489232 675446 489288
rect 675482 487192 675538 487248
rect 675114 485968 675170 486024
rect 675942 543292 675998 543348
rect 675942 539560 675998 539616
rect 676218 535880 676274 535936
rect 676034 535712 676036 535732
rect 676036 535712 676088 535732
rect 676088 535712 676090 535732
rect 676034 535676 676090 535712
rect 675850 534452 675906 534508
rect 675758 528332 675814 528388
rect 676034 534080 676036 534100
rect 676036 534080 676088 534100
rect 676088 534080 676090 534100
rect 676034 534044 676090 534080
rect 677414 533432 677470 533488
rect 676034 532752 676090 532808
rect 675942 532004 675998 532060
rect 675758 491544 675814 491600
rect 675758 491408 675814 491464
rect 675666 491272 675722 491328
rect 675666 487600 675722 487656
rect 675758 486784 675814 486840
rect 676126 532616 676182 532672
rect 676034 531596 676090 531652
rect 676034 527924 676090 527980
rect 676034 526292 676090 526348
rect 676218 531392 676274 531448
rect 675942 492088 675998 492144
rect 676034 491700 676090 491736
rect 676034 491680 676036 491700
rect 676036 491680 676088 491700
rect 676088 491680 676090 491700
rect 676034 491272 676090 491328
rect 679162 543632 679218 543688
rect 678978 535064 679034 535120
rect 679070 533024 679126 533080
rect 679070 530576 679126 530632
rect 678978 530168 679034 530224
rect 679346 543496 679402 543552
rect 679254 533840 679310 533896
rect 679254 530984 679310 531040
rect 679438 529760 679494 529816
rect 679346 529352 679402 529408
rect 679162 528944 679218 529000
rect 677598 527720 677654 527776
rect 677506 527312 677562 527368
rect 678978 525680 679034 525736
rect 678978 524864 679034 524920
rect 676034 490048 676090 490104
rect 679438 490456 679494 490512
rect 676034 489640 676090 489696
rect 675942 488416 675998 488472
rect 675850 486376 675906 486432
rect 675574 484744 675630 484800
rect 675850 484336 675906 484392
rect 676034 485560 676090 485616
rect 675942 483928 675998 483984
rect 676034 483520 676090 483576
rect 676034 483112 676090 483168
rect 675942 482704 675998 482760
rect 676034 482296 676090 482352
rect 676034 481888 676090 481944
rect 676034 480700 676036 480720
rect 676036 480700 676088 480720
rect 676088 480700 676090 480720
rect 672446 153312 672502 153368
rect 676034 480664 676090 480700
rect 675850 403028 675906 403064
rect 675850 403008 675852 403028
rect 675852 403008 675904 403028
rect 675904 403008 675906 403028
rect 675942 402600 675998 402656
rect 675298 401376 675354 401432
rect 672538 148144 672594 148200
rect 671986 114280 672042 114336
rect 666926 107480 666982 107536
rect 672262 105848 672318 105904
rect 672170 104080 672226 104136
rect 672630 127880 672686 127936
rect 676034 400968 676090 401024
rect 676310 403688 676366 403744
rect 676218 403280 676274 403336
rect 679162 488008 679218 488064
rect 679622 488824 679678 488880
rect 677486 402056 677542 402112
rect 676034 400152 676090 400208
rect 676034 399336 676090 399392
rect 675758 398520 675814 398576
rect 676126 398792 676182 398848
rect 676034 398112 676090 398168
rect 675942 397704 675998 397760
rect 676034 397296 676090 397352
rect 676034 396888 676090 396944
rect 675942 396072 675998 396128
rect 675850 395664 675906 395720
rect 675850 395256 675906 395312
rect 675942 394848 675998 394904
rect 676126 396344 676182 396400
rect 676034 394440 676090 394496
rect 676034 394032 676090 394088
rect 678978 393488 679034 393544
rect 678978 392672 679034 392728
rect 675666 357060 675722 357096
rect 675666 357040 675668 357060
rect 675668 357040 675720 357060
rect 675720 357040 675722 357060
rect 672814 143112 672870 143168
rect 675850 358672 675906 358728
rect 675758 356632 675814 356688
rect 675942 358264 675998 358320
rect 676034 357856 676090 357912
rect 676034 356224 676090 356280
rect 676034 355428 676090 355464
rect 676034 355408 676036 355428
rect 676036 355408 676088 355428
rect 676088 355408 676090 355428
rect 676034 354612 676090 354648
rect 676034 354592 676036 354612
rect 676036 354592 676088 354612
rect 676088 354592 676090 354612
rect 676034 354184 676090 354240
rect 675390 353776 675446 353832
rect 675298 351736 675354 351792
rect 676034 353368 676090 353424
rect 676034 352960 676090 353016
rect 675942 352552 675998 352608
rect 675850 352144 675906 352200
rect 676034 351328 676090 351384
rect 675942 350920 675998 350976
rect 675850 350512 675906 350568
rect 676034 350104 676090 350160
rect 676034 349696 676090 349752
rect 675942 349288 675998 349344
rect 675850 348880 675906 348936
rect 676034 347268 676090 347304
rect 676034 347248 676036 347268
rect 676036 347248 676088 347268
rect 676088 347248 676090 347268
rect 676310 313520 676366 313576
rect 676126 313112 676182 313168
rect 676034 312452 676090 312488
rect 676034 312432 676036 312452
rect 676036 312432 676088 312452
rect 676088 312432 676090 312452
rect 676218 312704 676274 312760
rect 676218 311908 676274 311944
rect 676218 311888 676220 311908
rect 676220 311888 676272 311908
rect 676272 311888 676274 311908
rect 676034 311652 676036 311672
rect 676036 311652 676088 311672
rect 676088 311652 676090 311672
rect 676034 311616 676090 311652
rect 676218 311092 676274 311128
rect 676218 311072 676220 311092
rect 676220 311072 676272 311092
rect 676272 311072 676274 311092
rect 672906 138400 672962 138456
rect 676218 310684 676274 310720
rect 676218 310664 676220 310684
rect 676220 310664 676272 310684
rect 676272 310664 676274 310684
rect 676218 310276 676274 310312
rect 676218 310256 676220 310276
rect 676220 310256 676272 310276
rect 676272 310256 676274 310276
rect 676218 309868 676274 309904
rect 676218 309848 676220 309868
rect 676220 309848 676272 309868
rect 676272 309848 676274 309868
rect 676218 309460 676274 309496
rect 676218 309440 676220 309460
rect 676220 309440 676272 309460
rect 676272 309440 676274 309460
rect 676034 309188 676090 309224
rect 676034 309168 676036 309188
rect 676036 309168 676088 309188
rect 676088 309168 676090 309188
rect 676034 308760 676090 308816
rect 675298 308352 675354 308408
rect 676034 307944 676090 308000
rect 675390 307128 675446 307184
rect 676126 307400 676182 307456
rect 676034 306720 676090 306776
rect 676034 306312 676090 306368
rect 676034 305904 676090 305960
rect 676126 305360 676182 305416
rect 676126 304952 676182 305008
rect 676034 304680 676090 304736
rect 676126 304136 676182 304192
rect 676034 303864 676090 303920
rect 678978 303320 679034 303376
rect 678978 302504 679034 302560
rect 676126 268504 676182 268560
rect 676034 267824 676090 267880
rect 676218 268116 676274 268152
rect 676218 268096 676220 268116
rect 676220 268096 676272 268116
rect 676272 268096 676274 268116
rect 678978 267688 679034 267744
rect 675666 267008 675722 267064
rect 676034 266636 676036 266656
rect 676036 266636 676088 266656
rect 676088 266636 676090 266656
rect 676034 266600 676090 266636
rect 676034 266192 676090 266248
rect 679070 266056 679126 266112
rect 675758 265376 675814 265432
rect 675666 260480 675722 260536
rect 675666 260072 675722 260128
rect 679162 265240 679218 265296
rect 676034 264152 676090 264208
rect 675850 263336 675906 263392
rect 676126 263608 676182 263664
rect 676034 262928 676090 262984
rect 676126 262384 676182 262440
rect 676034 262112 676090 262168
rect 676034 261704 676090 261760
rect 675942 260888 675998 260944
rect 676126 261160 676182 261216
rect 676126 259548 676182 259584
rect 676126 259528 676128 259548
rect 676128 259528 676180 259548
rect 676180 259528 676182 259548
rect 676034 259256 676090 259312
rect 676034 258848 676090 258904
rect 678978 258304 679034 258360
rect 678978 257488 679034 257544
rect 675666 222264 675722 222320
rect 675022 221448 675078 221504
rect 673090 216824 673146 216880
rect 672998 132912 673054 132968
rect 673274 216552 673330 216608
rect 674838 204856 674894 204912
rect 674930 176840 674986 176896
rect 675574 221856 675630 221912
rect 675390 221040 675446 221096
rect 675850 223488 675906 223544
rect 675942 223080 675998 223136
rect 676034 222672 676090 222728
rect 675758 220632 675814 220688
rect 675942 220224 675998 220280
rect 675482 218592 675538 218648
rect 675574 206216 675630 206272
rect 676034 219408 676090 219464
rect 676034 219000 676090 219056
rect 676034 218184 676090 218240
rect 676034 217776 676090 217832
rect 675942 217368 675998 217424
rect 675850 216960 675906 217016
rect 676034 216552 676090 216608
rect 675942 216144 675998 216200
rect 675850 215736 675906 215792
rect 675758 215328 675814 215384
rect 676034 214920 676090 214976
rect 676034 214512 676090 214568
rect 675942 214104 675998 214160
rect 675758 213696 675814 213752
rect 676034 212084 676090 212120
rect 676034 212064 676036 212084
rect 676036 212064 676088 212084
rect 676088 212064 676090 212084
rect 675390 205944 675446 206000
rect 675850 178472 675906 178528
rect 675298 177248 675354 177304
rect 675942 178064 675998 178120
rect 676034 177656 676090 177712
rect 676034 176432 676090 176488
rect 675942 176044 675998 176080
rect 675942 176024 675944 176044
rect 675944 176024 675996 176044
rect 675996 176024 675998 176044
rect 676034 175616 676090 175672
rect 675390 175208 675446 175264
rect 676034 174800 676090 174856
rect 675758 174392 675814 174448
rect 675574 173168 675630 173224
rect 675666 171536 675722 171592
rect 676034 173984 676090 174040
rect 676034 173576 676090 173632
rect 676034 172760 676090 172816
rect 675942 172352 675998 172408
rect 675942 171944 675998 172000
rect 676034 171148 676090 171184
rect 676034 171128 676036 171148
rect 676036 171128 676088 171148
rect 676088 171128 676090 171148
rect 676034 170720 676090 170776
rect 675942 170312 675998 170368
rect 675942 169904 675998 169960
rect 676034 169496 676090 169552
rect 675942 169088 675998 169144
rect 676034 168680 676090 168736
rect 676034 167068 676090 167104
rect 676034 167048 676036 167068
rect 676036 167048 676088 167068
rect 676088 167048 676090 167068
rect 676126 133048 676182 133104
rect 676034 132912 676090 132968
rect 676218 132640 676274 132696
rect 676034 132096 676090 132152
rect 676034 131708 676090 131744
rect 676034 131688 676036 131708
rect 676036 131688 676088 131708
rect 676088 131688 676090 131708
rect 676218 131452 676220 131472
rect 676220 131452 676272 131472
rect 676272 131452 676274 131472
rect 676218 131416 676274 131452
rect 676034 130892 676090 130928
rect 676034 130872 676036 130892
rect 676036 130872 676088 130892
rect 676088 130872 676090 130892
rect 675298 130464 675354 130520
rect 676034 130076 676090 130112
rect 676034 130056 676036 130076
rect 676036 130056 676088 130076
rect 676088 130056 676090 130076
rect 675758 129648 675814 129704
rect 676218 129412 676220 129432
rect 676220 129412 676272 129432
rect 676272 129412 676274 129432
rect 676218 129376 676274 129412
rect 676034 128832 676090 128888
rect 675942 128424 675998 128480
rect 675574 128016 675630 128072
rect 672722 122848 672778 122904
rect 672446 109248 672502 109304
rect 675298 125976 675354 126032
rect 675206 125568 675262 125624
rect 672354 102448 672410 102504
rect 676034 127608 676090 127664
rect 675942 127200 675998 127256
rect 676034 126792 676090 126848
rect 676034 126384 676090 126440
rect 675942 125160 675998 125216
rect 675942 124752 675998 124808
rect 675942 124344 675998 124400
rect 676034 123936 676090 123992
rect 675942 123528 675998 123584
rect 676218 121644 676274 121680
rect 676218 121624 676220 121644
rect 676220 121624 676272 121644
rect 676272 121624 676274 121644
rect 672078 100816 672134 100872
rect 666558 48456 666614 48512
rect 665178 47368 665234 47424
rect 549258 40976 549314 41032
rect 229374 6160 229430 6216
<< metal3 >>
rect 483565 1004730 483631 1004733
rect 483565 1004728 483644 1004730
rect 483565 1004672 483570 1004728
rect 483626 1004672 483644 1004728
rect 483565 1004670 483644 1004672
rect 483565 1004667 483631 1004670
tri 81502 983518 82144 984160 se
rect 82144 984060 87144 997762
rect 82144 983518 86502 984060
rect 81502 982718 86502 983518
tri 86502 983418 87144 984060 nw
rect 133544 983518 138544 997772
rect 133502 983382 138544 983518
rect 184944 983518 189944 997736
rect 221000 995620 235279 997736
rect 221000 993820 221400 995620
rect 234879 993820 235279 995620
rect 221000 993420 235279 993820
tri 221000 983518 230902 993420 ne
rect 230902 983518 235279 993420
rect 235579 984141 237779 997736
tri 235579 983518 236202 984141 ne
rect 236202 983518 237779 984141
rect 237978 984242 240178 997736
tri 237978 983868 238352 984242 ne
rect 238352 983868 240178 984242
rect 240478 995620 254800 997736
rect 240478 993820 240878 995620
rect 254357 993820 254800 995620
rect 240478 992116 254800 993820
rect 240478 984242 246202 992116
tri 240478 983868 240852 984242 ne
rect 240852 983868 246202 984242
tri 237779 983518 238129 983868 sw
tri 238352 983518 238702 983868 ne
rect 238702 983518 240178 983868
tri 240178 983518 240528 983868 sw
tri 240852 983518 241202 983868 ne
rect 184944 983452 190502 983518
rect 133502 982718 138502 983382
rect 185502 982718 190502 983452
rect 230902 982718 235902 983518
rect 236202 982718 238402 983518
rect 238702 982718 240902 983518
rect 241202 982718 246202 983868
tri 246202 983518 254800 992116 nw
rect 273600 995620 287879 997754
rect 273600 993820 274000 995620
rect 287479 993820 287879 995620
rect 273600 992520 287879 993820
tri 273600 983518 282602 992520 ne
rect 282602 983795 287879 992520
rect 282602 982718 287602 983795
tri 287602 983518 287879 983795 nw
rect 288179 983795 290379 997754
tri 287979 983518 288179 983718 se
rect 288179 983518 290102 983795
tri 290102 983518 290379 983795 nw
rect 290578 983694 292778 997754
tri 290402 983518 290578 983694 se
rect 290578 983518 292602 983694
tri 292602 983518 292778 983694 nw
rect 293078 995620 307400 997754
rect 293078 993820 293478 995620
rect 306957 993820 307400 995620
rect 293078 993016 307400 993820
rect 293078 983518 297902 993016
tri 297902 983518 307400 993016 nw
rect 375400 995620 389679 997722
rect 375400 993820 375800 995620
rect 389279 993820 389679 995620
rect 375400 992420 389679 993820
tri 375400 983518 384302 992420 ne
rect 384302 983895 389679 992420
rect 287902 982718 290102 983518
rect 290402 982718 292602 983518
rect 292902 982718 297902 983518
rect 384302 982718 389302 983895
tri 389302 983518 389679 983895 nw
rect 389979 983895 392179 997722
tri 389699 983518 389979 983798 se
rect 389979 983794 392078 983895
tri 392078 983794 392179 983895 nw
rect 392378 983794 394578 997722
rect 389979 983518 391802 983794
tri 391802 983518 392078 983794 nw
tri 392102 983518 392378 983794 se
rect 392378 983518 394302 983794
tri 394302 983518 394578 983794 nw
rect 394878 995620 409200 997722
rect 394878 993820 395278 995620
rect 408757 993820 409200 995620
rect 394878 993116 409200 993820
rect 394878 983518 399602 993116
tri 399602 983518 409200 993116 nw
rect 478744 983518 483744 997704
rect 389602 982718 391802 983518
rect 392102 982718 394302 983518
rect 394602 982718 399602 983518
rect 478702 983384 483744 983518
rect 530144 984064 535144 997792
tri 530144 983506 530702 984064 ne
rect 530702 983518 535144 984064
tri 535144 983518 535702 984076 sw
rect 478702 982718 483702 983384
rect 530702 982718 535702 983518
rect 575700 983678 580479 995092
tri 575700 983476 575902 983678 ne
rect 575902 983518 580479 983678
tri 580479 983518 580702 983741 sw
rect 575902 982718 580702 983518
rect 585678 983700 590458 995092
tri 585678 983476 585902 983700 ne
rect 585902 983518 590458 983700
tri 590458 983518 590702 983762 sw
rect 631944 983518 636944 997846
rect 585902 982718 590702 983518
rect 631902 983374 636944 983518
rect 631902 982718 636902 983374
rect 39764 963960 63464 965144
tri 63464 963960 64648 965144 sw
rect 39764 960144 65308 963960
tri 63325 958961 64508 960144 ne
rect 64508 958960 65308 960144
rect 649308 961656 650108 961702
rect 649308 956702 677806 961656
rect 650016 956656 677806 956702
rect 64508 926940 65308 927360
rect 46756 922560 65308 926940
rect 46756 922151 64552 922560
rect 649308 922502 650108 923302
tri 650108 922502 650908 923302 sw
rect 649308 918502 670780 922502
tri 649926 917700 650728 918502 ne
rect 650728 917700 670780 918502
rect 64508 916900 65308 917361
rect 46756 912560 65308 916900
rect 46756 912100 64560 912560
rect 649308 912449 650108 913302
tri 650108 912449 650961 913302 sw
rect 649308 908502 670788 912449
tri 649934 907660 650776 908502 ne
rect 650776 907660 670788 908502
rect 676029 897154 676095 897157
rect 676029 897152 676292 897154
rect 676029 897096 676034 897152
rect 676090 897096 676292 897152
rect 676029 897094 676292 897096
rect 676029 897091 676095 897094
rect 675937 896746 676003 896749
rect 675937 896744 676292 896746
rect 675937 896688 675942 896744
rect 675998 896688 676292 896744
rect 675937 896686 676292 896688
rect 675937 896683 676003 896686
rect 676029 896338 676095 896341
rect 676029 896336 676292 896338
rect 676029 896280 676034 896336
rect 676090 896280 676292 896336
rect 676029 896278 676292 896280
rect 676029 896275 676095 896278
rect 676121 895250 676187 895253
rect 676262 895250 676322 895492
rect 676121 895248 676322 895250
rect 676121 895192 676126 895248
rect 676182 895192 676322 895248
rect 676121 895190 676322 895192
rect 676121 895187 676187 895190
rect 675845 894706 675911 894709
rect 675845 894704 676292 894706
rect 675845 894648 675850 894704
rect 675906 894648 676292 894704
rect 675845 894646 676292 894648
rect 675845 894643 675911 894646
rect 676029 893890 676095 893893
rect 676029 893888 676292 893890
rect 676029 893832 676034 893888
rect 676090 893832 676292 893888
rect 676029 893830 676292 893832
rect 676029 893827 676095 893830
rect 676029 893074 676095 893077
rect 676029 893072 676292 893074
rect 676029 893016 676034 893072
rect 676090 893016 676292 893072
rect 676029 893014 676292 893016
rect 676029 893011 676095 893014
rect 679617 892666 679683 892669
rect 679604 892664 679683 892666
rect 679604 892608 679622 892664
rect 679678 892608 679683 892664
rect 679604 892606 679683 892608
rect 679617 892603 679683 892606
rect 676029 892258 676095 892261
rect 676029 892256 676292 892258
rect 676029 892200 676034 892256
rect 676090 892200 676292 892256
rect 676029 892198 676292 892200
rect 676029 892195 676095 892198
rect 679341 891850 679407 891853
rect 679341 891848 679420 891850
rect 679341 891792 679346 891848
rect 679402 891792 679420 891848
rect 679341 891790 679420 891792
rect 679341 891787 679407 891790
rect 679157 891442 679223 891445
rect 679157 891440 679236 891442
rect 679157 891384 679162 891440
rect 679218 891384 679236 891440
rect 679157 891382 679236 891384
rect 679157 891379 679223 891382
rect 676029 891034 676095 891037
rect 676029 891032 676292 891034
rect 676029 890976 676034 891032
rect 676090 890976 676292 891032
rect 676029 890974 676292 890976
rect 676029 890971 676095 890974
rect 676029 890626 676095 890629
rect 676029 890624 676292 890626
rect 676029 890568 676034 890624
rect 676090 890568 676292 890624
rect 676029 890566 676292 890568
rect 676029 890563 676095 890566
rect 678973 890218 679039 890221
rect 678973 890216 679052 890218
rect 678973 890160 678978 890216
rect 679034 890160 679052 890216
rect 678973 890158 679052 890160
rect 678973 890155 679039 890158
rect 679249 889810 679315 889813
rect 679236 889808 679315 889810
rect 679236 889752 679254 889808
rect 679310 889752 679315 889808
rect 679236 889750 679315 889752
rect 679249 889747 679315 889750
rect 679433 889402 679499 889405
rect 679420 889400 679499 889402
rect 679420 889344 679438 889400
rect 679494 889344 679499 889400
rect 679420 889342 679499 889344
rect 679433 889339 679499 889342
rect 675937 888994 676003 888997
rect 675937 888992 676292 888994
rect 675937 888936 675942 888992
rect 675998 888936 676292 888992
rect 675937 888934 676292 888936
rect 675937 888931 676003 888934
rect 676029 888586 676095 888589
rect 676029 888584 676292 888586
rect 676029 888528 676034 888584
rect 676090 888528 676292 888584
rect 676029 888526 676292 888528
rect 676029 888523 676095 888526
rect 679065 888178 679131 888181
rect 679052 888176 679131 888178
rect 679052 888120 679070 888176
rect 679126 888120 679131 888176
rect 679052 888118 679131 888120
rect 679065 888115 679131 888118
rect 676029 887770 676095 887773
rect 676029 887768 676292 887770
rect 676029 887712 676034 887768
rect 676090 887712 676292 887768
rect 676029 887710 676292 887712
rect 676029 887707 676095 887710
rect 675937 887362 676003 887365
rect 675937 887360 676292 887362
rect 675937 887304 675942 887360
rect 675998 887304 676292 887360
rect 675937 887302 676292 887304
rect 675937 887299 676003 887302
rect 679206 886684 679266 886924
rect 679198 886620 679204 886684
rect 679268 886620 679274 886684
rect 684542 886108 684602 886516
rect 679198 885804 679204 885868
rect 679268 885804 679274 885868
rect 679206 885700 679266 885804
rect 679198 884988 679204 885052
rect 679268 885050 679274 885052
rect 679525 885050 679591 885053
rect 679268 885048 679591 885050
rect 679268 884992 679530 885048
rect 679586 884992 679591 885048
rect 679268 884990 679591 884992
rect 679268 884988 679274 884990
rect 679525 884987 679591 884990
rect 655697 868866 655763 868869
rect 649950 868864 655763 868866
rect 649950 868808 655702 868864
rect 655758 868808 655763 868864
rect 649950 868806 655763 868808
rect 649950 868246 650010 868806
rect 655697 868803 655763 868806
rect 655513 867642 655579 867645
rect 649950 867640 655579 867642
rect 649950 867584 655518 867640
rect 655574 867584 655579 867640
rect 649950 867582 655579 867584
rect 649950 867064 650010 867582
rect 655513 867579 655579 867582
rect 655421 866554 655487 866557
rect 649950 866552 655487 866554
rect 649950 866496 655426 866552
rect 655482 866496 655487 866552
rect 649950 866494 655487 866496
rect 649950 865882 650010 866494
rect 655421 866491 655487 866494
rect 655605 865330 655671 865333
rect 649950 865328 655671 865330
rect 649950 865272 655610 865328
rect 655666 865272 655671 865328
rect 649950 865270 655671 865272
rect 649950 864700 650010 865270
rect 655605 865267 655671 865270
rect 655789 863834 655855 863837
rect 649950 863832 655855 863834
rect 649950 863776 655794 863832
rect 655850 863776 655855 863832
rect 649950 863774 655855 863776
rect 649950 863518 650010 863774
rect 655789 863771 655855 863774
rect 656801 862610 656867 862613
rect 649950 862608 656867 862610
rect 649950 862552 656806 862608
rect 656862 862552 656867 862608
rect 649950 862550 656867 862552
rect 649950 862336 650010 862550
rect 656801 862547 656867 862550
tri 64006 842458 64508 842960 se
rect 64508 842458 65308 842960
rect 49892 838160 65308 842458
rect 49892 837678 64152 838160
tri 64152 837678 64634 838160 nw
rect 649308 833301 650108 834080
tri 64027 832479 64508 832960 se
rect 64508 832479 65308 832960
rect 49892 828160 65308 832479
rect 649308 829280 667192 833301
rect 649858 828521 667192 829280
rect 49892 828159 64634 828160
rect 49892 827699 64174 828159
tri 64174 827699 64634 828159 nw
rect 649308 823322 650108 824080
rect 649308 819280 667192 823322
rect 649858 818542 667192 819280
rect 41781 817730 41847 817733
rect 41492 817728 41847 817730
rect 41492 817672 41786 817728
rect 41842 817672 41847 817728
rect 41492 817670 41847 817672
rect 41781 817667 41847 817670
rect 41781 817322 41847 817325
rect 41492 817320 41847 817322
rect 41492 817264 41786 817320
rect 41842 817264 41847 817320
rect 41492 817262 41847 817264
rect 41781 817259 41847 817262
rect 41781 816914 41847 816917
rect 41492 816912 41847 816914
rect 41492 816856 41786 816912
rect 41842 816856 41847 816912
rect 41492 816854 41847 816856
rect 41781 816851 41847 816854
rect 44589 816132 44659 816135
rect 41594 816130 44668 816132
rect 41594 816072 44594 816130
rect 44589 816070 44594 816072
rect 44654 816072 44668 816130
rect 44654 816070 44659 816072
rect 44589 816065 44659 816070
rect 43621 815282 43687 815285
rect 41492 815280 43687 815282
rect 41492 815224 43626 815280
rect 43682 815224 43687 815280
rect 41492 815222 43687 815224
rect 43621 815219 43687 815222
rect 41781 814602 41847 814605
rect 59261 814602 59327 814605
rect 41781 814600 59327 814602
rect 41781 814544 41786 814600
rect 41842 814544 59266 814600
rect 59322 814544 59327 814600
rect 41781 814542 59327 814544
rect 41781 814539 41847 814542
rect 59261 814539 59327 814542
rect 44681 814468 44751 814473
rect 44681 814466 44686 814468
rect 41600 814408 44686 814466
rect 44746 814466 44751 814468
rect 44746 814408 44758 814466
rect 41600 814406 44758 814408
rect 44681 814403 44751 814406
rect 44773 813676 44843 813681
rect 44773 813670 44778 813676
rect 41600 813616 44778 813670
rect 44838 813670 44843 813676
rect 44838 813616 44864 813670
rect 41600 813610 44864 813616
rect 43437 813242 43503 813245
rect 41492 813240 43503 813242
rect 41492 813184 43442 813240
rect 43498 813184 43503 813240
rect 41492 813182 43503 813184
rect 43437 813179 43503 813182
rect 42701 812834 42767 812837
rect 41492 812832 42767 812834
rect 41492 812776 42706 812832
rect 42762 812776 42767 812832
rect 41492 812774 42767 812776
rect 42701 812771 42767 812774
rect 43069 812426 43135 812429
rect 41492 812424 43135 812426
rect 41492 812368 43074 812424
rect 43130 812368 43135 812424
rect 41492 812366 43135 812368
rect 43069 812363 43135 812366
rect 42793 812018 42859 812021
rect 41492 812016 42859 812018
rect 41492 811960 42798 812016
rect 42854 811960 42859 812016
rect 41492 811958 42859 811960
rect 42793 811955 42859 811958
rect 42885 811610 42951 811613
rect 41492 811608 42951 811610
rect 41492 811552 42890 811608
rect 42946 811552 42951 811608
rect 41492 811550 42951 811552
rect 42885 811547 42951 811550
rect 42241 811202 42307 811205
rect 41492 811200 42307 811202
rect 41492 811144 42246 811200
rect 42302 811144 42307 811200
rect 41492 811142 42307 811144
rect 42241 811139 42307 811142
rect 43713 810794 43779 810797
rect 41492 810792 43779 810794
rect 41492 810736 43718 810792
rect 43774 810736 43779 810792
rect 41492 810734 43779 810736
rect 43713 810731 43779 810734
rect 43805 810386 43871 810389
rect 41492 810384 43871 810386
rect 41492 810328 43810 810384
rect 43866 810328 43871 810384
rect 41492 810326 43871 810328
rect 43805 810323 43871 810326
rect 43897 809978 43963 809981
rect 41492 809976 43963 809978
rect 41492 809920 43902 809976
rect 43958 809920 43963 809976
rect 41492 809918 43963 809920
rect 43897 809915 43963 809918
rect 42609 809570 42675 809573
rect 41492 809568 42675 809570
rect 41492 809512 42614 809568
rect 42670 809512 42675 809568
rect 41492 809510 42675 809512
rect 42609 809507 42675 809510
rect 41965 809162 42031 809165
rect 41492 809160 42031 809162
rect 41492 809104 41970 809160
rect 42026 809104 42031 809160
rect 41492 809102 42031 809104
rect 41965 809099 42031 809102
rect 41873 808754 41939 808757
rect 41492 808752 41939 808754
rect 41492 808696 41878 808752
rect 41934 808696 41939 808752
rect 41492 808694 41939 808696
rect 41873 808691 41939 808694
rect 41781 808346 41847 808349
rect 41492 808344 41847 808346
rect 41492 808288 41786 808344
rect 41842 808288 41847 808344
rect 41492 808286 41847 808288
rect 41781 808283 41847 808286
rect 41822 807938 41828 807940
rect 41492 807878 41828 807938
rect 41822 807876 41828 807878
rect 41892 807876 41898 807940
rect 41781 807530 41847 807533
rect 41492 807528 41847 807530
rect 41492 807472 41786 807528
rect 41842 807472 41847 807528
rect 41492 807470 41847 807472
rect 41781 807467 41847 807470
rect 30422 806684 30482 807092
rect 41781 806306 41847 806309
rect 42333 806306 42399 806309
rect 41492 806304 42399 806306
rect 41492 806248 41786 806304
rect 41842 806248 42338 806304
rect 42394 806248 42399 806304
rect 41492 806246 42399 806248
rect 41781 806243 41847 806246
rect 42333 806243 42399 806246
rect 41873 795020 41939 795021
rect 41822 795018 41828 795020
rect 41782 794958 41828 795018
rect 41892 795016 41939 795020
rect 41934 794960 41939 795016
rect 41822 794956 41828 794958
rect 41892 794956 41939 794960
rect 41873 794955 41939 794956
rect 58249 790938 58315 790941
rect 58249 790936 64706 790938
rect 58249 790880 58254 790936
rect 58310 790880 64706 790936
rect 58249 790878 64706 790880
rect 58249 790875 58315 790878
rect 64646 790304 64706 790878
rect 58525 789306 58591 789309
rect 58525 789304 64706 789306
rect 58525 789248 58530 789304
rect 58586 789248 64706 789304
rect 58525 789246 64706 789248
rect 58525 789243 58591 789246
rect 64646 789122 64706 789246
rect 58065 788490 58131 788493
rect 58065 788488 64706 788490
rect 58065 788432 58070 788488
rect 58126 788432 64706 788488
rect 58065 788430 64706 788432
rect 58065 788427 58131 788430
rect 64646 787940 64706 788430
rect 674966 788292 674972 788356
rect 675036 788354 675042 788356
rect 675109 788354 675175 788357
rect 675036 788352 675175 788354
rect 675036 788296 675114 788352
rect 675170 788296 675175 788352
rect 675036 788294 675175 788296
rect 675036 788292 675042 788294
rect 675109 788291 675175 788294
rect 59261 787402 59327 787405
rect 59261 787400 64706 787402
rect 59261 787344 59266 787400
rect 59322 787344 64706 787400
rect 59261 787342 64706 787344
rect 59261 787339 59327 787342
rect 64646 786758 64706 787342
rect 674598 787204 674604 787268
rect 674668 787266 674674 787268
rect 675109 787266 675175 787269
rect 674668 787264 675175 787266
rect 674668 787208 675114 787264
rect 675170 787208 675175 787264
rect 674668 787206 675175 787208
rect 674668 787204 674674 787206
rect 675109 787203 675175 787206
rect 674782 786660 674788 786724
rect 674852 786722 674858 786724
rect 675109 786722 675175 786725
rect 674852 786720 675175 786722
rect 674852 786664 675114 786720
rect 675170 786664 675175 786720
rect 674852 786662 675175 786664
rect 674852 786660 674858 786662
rect 675109 786659 675175 786662
rect 58525 786178 58591 786181
rect 58525 786176 64706 786178
rect 58525 786120 58530 786176
rect 58586 786120 64706 786176
rect 58525 786118 64706 786120
rect 58525 786115 58591 786118
rect 64646 785576 64706 786118
rect 58433 784954 58499 784957
rect 58433 784952 64706 784954
rect 58433 784896 58438 784952
rect 58494 784896 64706 784952
rect 58433 784894 64706 784896
rect 58433 784891 58499 784894
rect 64646 784394 64706 784894
rect 649950 778426 650010 778824
rect 655421 778426 655487 778429
rect 649950 778424 655487 778426
rect 649950 778368 655426 778424
rect 655482 778368 655487 778424
rect 649950 778366 655487 778368
rect 655421 778363 655487 778366
rect 649950 777066 650010 777642
rect 655605 777066 655671 777069
rect 649950 777064 655671 777066
rect 649950 777008 655610 777064
rect 655666 777008 655671 777064
rect 649950 777006 655671 777008
rect 655605 777003 655671 777006
rect 649950 775978 650010 776460
rect 655789 775978 655855 775981
rect 649950 775976 655855 775978
rect 649950 775920 655794 775976
rect 655850 775920 655855 775976
rect 649950 775918 655855 775920
rect 655789 775915 655855 775918
rect 655513 775570 655579 775573
rect 649950 775568 655579 775570
rect 649950 775512 655518 775568
rect 655574 775512 655579 775568
rect 649950 775510 655579 775512
rect 649950 775278 650010 775510
rect 655513 775507 655579 775510
rect 41505 774754 41571 774757
rect 656525 774754 656591 774757
rect 41462 774752 41571 774754
rect 41462 774696 41510 774752
rect 41566 774696 41571 774752
rect 41462 774691 41571 774696
rect 649950 774752 656591 774754
rect 649950 774696 656530 774752
rect 656586 774696 656591 774752
rect 649950 774694 656591 774696
rect 41462 774452 41522 774691
rect 649950 774096 650010 774694
rect 656525 774691 656591 774694
rect 41462 773941 41522 774044
rect 41462 773936 41571 773941
rect 41462 773880 41510 773936
rect 41566 773880 41571 773936
rect 41462 773878 41571 773880
rect 41505 773875 41571 773878
rect 41462 773533 41522 773636
rect 41462 773528 41571 773533
rect 654961 773530 655027 773533
rect 41462 773472 41510 773528
rect 41566 773472 41571 773528
rect 41462 773470 41571 773472
rect 41505 773467 41571 773470
rect 649950 773528 655027 773530
rect 649950 773472 654966 773528
rect 655022 773472 655027 773528
rect 649950 773470 655027 773472
rect 44589 773314 44659 773319
rect 41620 773254 44594 773314
rect 44654 773254 44668 773314
rect 44589 773249 44659 773254
rect 44589 772932 44659 772935
rect 41620 772930 44668 772932
rect 41620 772872 44594 772930
rect 44589 772870 44594 772872
rect 44654 772872 44668 772930
rect 649950 772914 650010 773470
rect 654961 773467 655027 773470
rect 44654 772870 44659 772872
rect 44589 772865 44659 772870
rect 43621 772442 43687 772445
rect 41492 772440 43687 772442
rect 41492 772384 43626 772440
rect 43682 772384 43687 772440
rect 41492 772382 43687 772384
rect 43621 772379 43687 772382
rect 43713 772034 43779 772037
rect 41492 772032 43779 772034
rect 41492 771976 43718 772032
rect 43774 771976 43779 772032
rect 41492 771974 43779 771976
rect 43713 771971 43779 771974
rect 44681 771680 44751 771683
rect 41596 771678 44758 771680
rect 41596 771620 44686 771678
rect 44681 771618 44686 771620
rect 44746 771620 44758 771678
rect 44746 771618 44751 771620
rect 44681 771613 44751 771618
rect 44681 771268 44751 771273
rect 44681 771266 44686 771268
rect 41596 771208 44686 771266
rect 44746 771266 44751 771268
rect 44746 771208 44758 771266
rect 41596 771206 44758 771208
rect 44681 771203 44751 771206
rect 44773 770888 44843 770893
rect 41596 770828 44778 770888
rect 44838 770828 44864 770888
rect 44773 770823 44843 770828
rect 44773 770476 44843 770481
rect 44773 770470 44778 770476
rect 41596 770416 44778 770470
rect 44838 770470 44843 770476
rect 44838 770416 44864 770470
rect 41596 770410 44864 770416
rect 44081 769994 44147 769997
rect 41492 769992 44147 769994
rect 41492 769936 44086 769992
rect 44142 769936 44147 769992
rect 41492 769934 44147 769936
rect 44081 769931 44147 769934
rect 42333 769586 42399 769589
rect 41492 769584 42399 769586
rect 41492 769528 42338 769584
rect 42394 769528 42399 769584
rect 41492 769526 42399 769528
rect 42333 769523 42399 769526
rect 43621 769178 43687 769181
rect 41492 769176 43687 769178
rect 41492 769120 43626 769176
rect 43682 769120 43687 769176
rect 41492 769118 43687 769120
rect 43621 769115 43687 769118
rect 43069 768770 43135 768773
rect 41492 768768 43135 768770
rect 41492 768712 43074 768768
rect 43130 768712 43135 768768
rect 41492 768710 43135 768712
rect 43069 768707 43135 768710
rect 42701 768362 42767 768365
rect 41492 768360 42767 768362
rect 41492 768304 42706 768360
rect 42762 768304 42767 768360
rect 41492 768302 42767 768304
rect 42701 768299 42767 768302
rect 38334 767821 38394 767924
rect 38285 767816 38394 767821
rect 38285 767760 38290 767816
rect 38346 767760 38394 767816
rect 38285 767758 38394 767760
rect 38285 767755 38351 767758
rect 38150 767413 38210 767516
rect 38150 767408 38259 767413
rect 38150 767352 38198 767408
rect 38254 767352 38259 767408
rect 38150 767350 38259 767352
rect 38193 767347 38259 767350
rect 43897 767138 43963 767141
rect 41492 767136 43963 767138
rect 41492 767080 43902 767136
rect 43958 767080 43963 767136
rect 41492 767078 43963 767080
rect 43897 767075 43963 767078
rect 43805 766730 43871 766733
rect 41492 766728 43871 766730
rect 41492 766672 43810 766728
rect 43866 766672 43871 766728
rect 41492 766670 43871 766672
rect 43805 766667 43871 766670
rect 43161 766322 43227 766325
rect 41492 766320 43227 766322
rect 41492 766264 43166 766320
rect 43222 766264 43227 766320
rect 41492 766262 43227 766264
rect 43161 766259 43227 766262
rect 43253 765914 43319 765917
rect 41492 765912 43319 765914
rect 41492 765856 43258 765912
rect 43314 765856 43319 765912
rect 41492 765854 43319 765856
rect 43253 765851 43319 765854
rect 42425 765506 42491 765509
rect 41492 765504 42491 765506
rect 41492 765448 42430 765504
rect 42486 765448 42491 765504
rect 41492 765446 42491 765448
rect 42425 765443 42491 765446
rect 41462 764965 41522 765068
rect 41462 764960 41571 764965
rect 41462 764904 41510 764960
rect 41566 764904 41571 764960
rect 41462 764902 41571 764904
rect 41505 764899 41571 764902
rect 38518 764557 38578 764660
rect 38518 764552 38627 764557
rect 38518 764496 38566 764552
rect 38622 764496 38627 764552
rect 38518 764494 38627 764496
rect 38561 764491 38627 764494
rect 41462 764146 41522 764252
rect 41597 764146 41663 764149
rect 41462 764144 41663 764146
rect 41462 764088 41602 764144
rect 41658 764088 41663 764144
rect 41462 764086 41663 764088
rect 41597 764083 41663 764086
rect 30422 763436 30482 763844
rect 41462 762922 41522 763028
rect 41597 762922 41663 762925
rect 41462 762920 41663 762922
rect 41462 762864 41602 762920
rect 41658 762864 41663 762920
rect 41462 762862 41663 762864
rect 41597 762859 41663 762862
rect 58433 747690 58499 747693
rect 58433 747688 64706 747690
rect 58433 747632 58438 747688
rect 58494 747632 64706 747688
rect 58433 747630 64706 747632
rect 58433 747627 58499 747630
rect 64646 747082 64706 747630
rect 59261 746466 59327 746469
rect 59261 746464 64706 746466
rect 59261 746408 59266 746464
rect 59322 746408 64706 746464
rect 59261 746406 64706 746408
rect 59261 746403 59327 746406
rect 64646 745900 64706 746406
rect 673821 745378 673887 745381
rect 676806 745378 676812 745380
rect 673821 745376 676812 745378
rect 673821 745320 673826 745376
rect 673882 745320 676812 745376
rect 673821 745318 676812 745320
rect 673821 745315 673887 745318
rect 676806 745316 676812 745318
rect 676876 745316 676882 745380
rect 674557 745242 674623 745245
rect 676622 745242 676628 745244
rect 674557 745240 676628 745242
rect 674557 745184 674562 745240
rect 674618 745184 676628 745240
rect 674557 745182 676628 745184
rect 674557 745179 674623 745182
rect 676622 745180 676628 745182
rect 676692 745180 676698 745244
rect 58433 744970 58499 744973
rect 58433 744968 64706 744970
rect 58433 744912 58438 744968
rect 58494 744912 64706 744968
rect 58433 744910 64706 744912
rect 58433 744907 58499 744910
rect 64646 744718 64706 744910
rect 58525 744154 58591 744157
rect 58525 744152 64706 744154
rect 58525 744096 58530 744152
rect 58586 744096 64706 744152
rect 58525 744094 64706 744096
rect 58525 744091 58591 744094
rect 64646 743536 64706 744094
rect 674046 742868 674052 742932
rect 674116 742930 674122 742932
rect 675385 742930 675451 742933
rect 674116 742928 675451 742930
rect 674116 742872 675390 742928
rect 675446 742872 675451 742928
rect 674116 742870 675451 742872
rect 674116 742868 674122 742870
rect 675385 742867 675451 742870
rect 673862 742460 673868 742524
rect 673932 742522 673938 742524
rect 675385 742522 675451 742525
rect 673932 742520 675451 742522
rect 673932 742464 675390 742520
rect 675446 742464 675451 742520
rect 673932 742462 675451 742464
rect 673932 742460 673938 742462
rect 675385 742459 675451 742462
rect 57973 742386 58039 742389
rect 57973 742384 64706 742386
rect 57973 742328 57978 742384
rect 58034 742328 64706 742384
rect 57973 742326 64706 742328
rect 57973 742323 58039 742326
rect 58433 741842 58499 741845
rect 58433 741840 64706 741842
rect 58433 741784 58438 741840
rect 58494 741784 64706 741840
rect 58433 741782 64706 741784
rect 58433 741779 58499 741782
rect 64646 741172 64706 741782
rect 674230 741644 674236 741708
rect 674300 741706 674306 741708
rect 675477 741706 675543 741709
rect 674300 741704 675543 741706
rect 674300 741648 675482 741704
rect 675538 741648 675543 741704
rect 674300 741646 675543 741648
rect 674300 741644 674306 741646
rect 675477 741643 675543 741646
rect 675150 739740 675156 739804
rect 675220 739802 675226 739804
rect 675385 739802 675451 739805
rect 675220 739800 675451 739802
rect 675220 739744 675390 739800
rect 675446 739744 675451 739800
rect 675220 739742 675451 739744
rect 675220 739740 675226 739742
rect 675385 739739 675451 739742
rect 673678 739060 673684 739124
rect 673748 739122 673754 739124
rect 675385 739122 675451 739125
rect 673748 739120 675451 739122
rect 673748 739064 675390 739120
rect 675446 739064 675451 739120
rect 673748 739062 675451 739064
rect 673748 739060 673754 739062
rect 675385 739059 675451 739062
rect 674414 738652 674420 738716
rect 674484 738714 674490 738716
rect 675385 738714 675451 738717
rect 674484 738712 675451 738714
rect 674484 738656 675390 738712
rect 675446 738656 675451 738712
rect 674484 738654 675451 738656
rect 674484 738652 674490 738654
rect 675385 738651 675451 738654
rect 675385 738036 675451 738037
rect 675334 738034 675340 738036
rect 675294 737974 675340 738034
rect 675404 738032 675451 738036
rect 675446 737976 675451 738032
rect 675334 737972 675340 737974
rect 675404 737972 675451 737976
rect 675385 737971 675451 737972
rect 674741 734906 674807 734909
rect 674741 734904 675218 734906
rect 674741 734848 674746 734904
rect 674802 734848 675218 734904
rect 674741 734846 675218 734848
rect 674741 734843 674807 734846
rect 649950 734362 650010 734402
rect 655697 734362 655763 734365
rect 649950 734360 655763 734362
rect 649950 734304 655702 734360
rect 655758 734304 655763 734360
rect 649950 734302 655763 734304
rect 655697 734299 655763 734302
rect 675158 733413 675218 734846
rect 675158 733408 675267 733413
rect 675158 733352 675206 733408
rect 675262 733352 675267 733408
rect 675158 733350 675267 733352
rect 675201 733347 675267 733350
rect 649950 732730 650010 733220
rect 655881 732730 655947 732733
rect 649950 732728 655947 732730
rect 649950 732672 655886 732728
rect 655942 732672 655947 732728
rect 649950 732670 655947 732672
rect 655881 732667 655947 732670
rect 649950 731506 650010 732038
rect 655513 731506 655579 731509
rect 649950 731504 655579 731506
rect 649950 731448 655518 731504
rect 655574 731448 655579 731504
rect 649950 731446 655579 731448
rect 655513 731443 655579 731446
rect 655973 731370 656039 731373
rect 649950 731368 656039 731370
rect 41462 731098 41522 731340
rect 649950 731312 655978 731368
rect 656034 731312 656039 731368
rect 649950 731310 656039 731312
rect 44301 731098 44367 731101
rect 41462 731096 44367 731098
rect 41462 731040 44306 731096
rect 44362 731040 44367 731096
rect 41462 731038 44367 731040
rect 44301 731035 44367 731038
rect 41462 730690 41522 730932
rect 649950 730856 650010 731310
rect 655973 731307 656039 731310
rect 673494 730764 673500 730828
rect 673564 730826 673570 730828
rect 674598 730826 674604 730828
rect 673564 730766 674604 730826
rect 673564 730764 673570 730766
rect 674598 730764 674604 730766
rect 674668 730764 674674 730828
rect 44123 730690 44189 730693
rect 41462 730688 44189 730690
rect 41462 730632 44128 730688
rect 44184 730632 44189 730688
rect 41462 730630 44189 730632
rect 44123 730627 44189 730630
rect 41462 730282 41522 730524
rect 43897 730282 43963 730285
rect 655145 730282 655211 730285
rect 41462 730280 43963 730282
rect 41462 730224 43902 730280
rect 43958 730224 43963 730280
rect 41462 730222 43963 730224
rect 43897 730219 43963 730222
rect 649950 730280 655211 730282
rect 649950 730224 655150 730280
rect 655206 730224 655211 730280
rect 649950 730222 655211 730224
rect 44589 730114 44659 730119
rect 41590 730054 44594 730114
rect 44654 730054 44668 730114
rect 44589 730049 44659 730054
rect 44589 729732 44659 729735
rect 41590 729730 44668 729732
rect 41590 729672 44594 729730
rect 44589 729670 44594 729672
rect 44654 729672 44668 729730
rect 649950 729674 650010 730222
rect 655145 730219 655211 730222
rect 44654 729670 44659 729672
rect 44589 729665 44659 729670
rect 41505 729466 41571 729469
rect 41462 729464 41571 729466
rect 41462 729408 41510 729464
rect 41566 729408 41571 729464
rect 41462 729403 41571 729408
rect 41462 729300 41522 729403
rect 44301 729194 44367 729197
rect 59629 729194 59695 729197
rect 44301 729192 59695 729194
rect 44301 729136 44306 729192
rect 44362 729136 59634 729192
rect 59690 729136 59695 729192
rect 44301 729134 59695 729136
rect 44301 729131 44367 729134
rect 59629 729131 59695 729134
rect 44133 729058 44199 729061
rect 59261 729058 59327 729061
rect 44133 729056 59327 729058
rect 44133 729000 44138 729056
rect 44194 729000 59266 729056
rect 59322 729000 59327 729056
rect 44133 728998 59327 729000
rect 44133 728995 44199 728998
rect 59261 728995 59327 728998
rect 43713 728922 43779 728925
rect 41492 728920 43779 728922
rect 41492 728864 43718 728920
rect 43774 728864 43779 728920
rect 41492 728862 43779 728864
rect 43713 728859 43779 728862
rect 43897 728922 43963 728925
rect 59445 728922 59511 728925
rect 43897 728920 59511 728922
rect 43897 728864 43902 728920
rect 43958 728864 59450 728920
rect 59506 728864 59511 728920
rect 43897 728862 59511 728864
rect 43897 728859 43963 728862
rect 59445 728859 59511 728862
rect 656065 728650 656131 728653
rect 651330 728648 656131 728650
rect 651330 728592 656070 728648
rect 656126 728592 656131 728648
rect 651330 728590 656131 728592
rect 651330 728514 651390 728590
rect 656065 728587 656131 728590
rect 44681 728480 44751 728483
rect 41570 728478 44758 728480
rect 41570 728420 44686 728478
rect 44681 728418 44686 728420
rect 44746 728420 44758 728478
rect 649950 728454 651390 728514
rect 44746 728418 44751 728420
rect 44681 728413 44751 728418
rect 44681 728068 44751 728073
rect 44681 728066 44686 728068
rect 41570 728008 44686 728066
rect 44746 728066 44751 728068
rect 44746 728008 44758 728066
rect 41570 728006 44758 728008
rect 44681 728003 44751 728006
rect 44773 727688 44843 727693
rect 41570 727628 44778 727688
rect 44838 727628 44864 727688
rect 44773 727623 44843 727628
rect 44773 727276 44843 727281
rect 44773 727270 44778 727276
rect 41570 727216 44778 727270
rect 44838 727270 44843 727276
rect 44838 727216 44864 727270
rect 41570 727210 44864 727216
rect 43161 726882 43227 726885
rect 41492 726880 43227 726882
rect 41492 726824 43166 726880
rect 43222 726824 43227 726880
rect 41492 726822 43227 726824
rect 43161 726819 43227 726822
rect 43345 726474 43411 726477
rect 41492 726472 43411 726474
rect 41492 726416 43350 726472
rect 43406 726416 43411 726472
rect 41492 726414 43411 726416
rect 43345 726411 43411 726414
rect 43805 726066 43871 726069
rect 41492 726064 43871 726066
rect 41492 726008 43810 726064
rect 43866 726008 43871 726064
rect 41492 726006 43871 726008
rect 43805 726003 43871 726006
rect 43989 725658 44055 725661
rect 41492 725656 44055 725658
rect 41492 725600 43994 725656
rect 44050 725600 44055 725656
rect 41492 725598 44055 725600
rect 43989 725595 44055 725598
rect 43897 725250 43963 725253
rect 41492 725248 43963 725250
rect 41492 725192 43902 725248
rect 43958 725192 43963 725248
rect 41492 725190 43963 725192
rect 43897 725187 43963 725190
rect 41781 724842 41847 724845
rect 41492 724840 41847 724842
rect 41492 724784 41786 724840
rect 41842 724784 41847 724840
rect 41492 724782 41847 724784
rect 41781 724779 41847 724782
rect 44081 724434 44147 724437
rect 41492 724432 44147 724434
rect 41492 724376 44086 724432
rect 44142 724376 44147 724432
rect 41492 724374 44147 724376
rect 44081 724371 44147 724374
rect 43437 724026 43503 724029
rect 41492 724024 43503 724026
rect 41492 723968 43442 724024
rect 43498 723968 43503 724024
rect 41492 723966 43503 723968
rect 43437 723963 43503 723966
rect 41462 723349 41522 723588
rect 41413 723344 41522 723349
rect 41413 723288 41418 723344
rect 41474 723288 41522 723344
rect 41413 723286 41522 723288
rect 41413 723283 41479 723286
rect 42241 723210 42307 723213
rect 41492 723208 42307 723210
rect 41492 723152 42246 723208
rect 42302 723152 42307 723208
rect 41492 723150 42307 723152
rect 42241 723147 42307 723150
rect 42701 722802 42767 722805
rect 41492 722800 42767 722802
rect 41492 722744 42706 722800
rect 42762 722744 42767 722800
rect 41492 722742 42767 722744
rect 42701 722739 42767 722742
rect 43253 722394 43319 722397
rect 41492 722392 43319 722394
rect 41492 722336 43258 722392
rect 43314 722336 43319 722392
rect 41492 722334 43319 722336
rect 43253 722331 43319 722334
rect 42333 721986 42399 721989
rect 41492 721984 42399 721986
rect 41492 721928 42338 721984
rect 42394 721928 42399 721984
rect 41492 721926 42399 721928
rect 42333 721923 42399 721926
rect 43621 721578 43687 721581
rect 41492 721576 43687 721578
rect 41492 721520 43626 721576
rect 43682 721520 43687 721576
rect 41492 721518 43687 721520
rect 43621 721515 43687 721518
rect 41462 720901 41522 721140
rect 41462 720896 41571 720901
rect 41462 720840 41510 720896
rect 41566 720840 41571 720896
rect 41462 720838 41571 720840
rect 41505 720835 41571 720838
rect 29870 720324 29930 720732
rect 41462 719677 41522 719916
rect 41462 719672 41571 719677
rect 41462 719616 41510 719672
rect 41566 719616 41571 719672
rect 41462 719614 41571 719616
rect 41505 719611 41571 719614
rect 675753 716546 675819 716549
rect 675753 716544 676292 716546
rect 675753 716488 675758 716544
rect 675814 716488 676292 716544
rect 675753 716486 676292 716488
rect 675753 716483 675819 716486
rect 675845 716138 675911 716141
rect 675845 716136 676292 716138
rect 675845 716080 675850 716136
rect 675906 716080 676292 716136
rect 675845 716078 676292 716080
rect 675845 716075 675911 716078
rect 675937 715730 676003 715733
rect 675937 715728 676292 715730
rect 675937 715672 675942 715728
rect 675998 715672 676292 715728
rect 675937 715670 676292 715672
rect 675937 715667 676003 715670
rect 676029 715322 676095 715325
rect 676029 715320 676292 715322
rect 676029 715264 676034 715320
rect 676090 715264 676292 715320
rect 676029 715262 676292 715264
rect 676029 715259 676095 715262
rect 676029 714914 676095 714917
rect 676029 714912 676292 714914
rect 676029 714856 676034 714912
rect 676090 714856 676292 714912
rect 676029 714854 676292 714856
rect 676029 714851 676095 714854
rect 676029 714506 676095 714509
rect 676029 714504 676292 714506
rect 676029 714448 676034 714504
rect 676090 714448 676292 714504
rect 676029 714446 676292 714448
rect 676029 714443 676095 714446
rect 676029 714098 676095 714101
rect 676029 714096 676292 714098
rect 676029 714040 676034 714096
rect 676090 714040 676292 714096
rect 676029 714038 676292 714040
rect 676029 714035 676095 714038
rect 676029 713690 676095 713693
rect 676029 713688 676292 713690
rect 676029 713632 676034 713688
rect 676090 713632 676292 713688
rect 676029 713630 676292 713632
rect 676029 713627 676095 713630
rect 675845 713282 675911 713285
rect 675845 713280 676292 713282
rect 675845 713224 675850 713280
rect 675906 713224 676292 713280
rect 675845 713222 676292 713224
rect 675845 713219 675911 713222
rect 675937 712874 676003 712877
rect 675937 712872 676292 712874
rect 675937 712816 675942 712872
rect 675998 712816 676292 712872
rect 675937 712814 676292 712816
rect 675937 712811 676003 712814
rect 676029 712466 676095 712469
rect 676029 712464 676292 712466
rect 676029 712408 676034 712464
rect 676090 712408 676292 712464
rect 676029 712406 676292 712408
rect 676029 712403 676095 712406
rect 674598 711996 674604 712060
rect 674668 712058 674674 712060
rect 674668 711998 676292 712058
rect 674668 711996 674674 711998
rect 676029 711650 676095 711653
rect 676029 711648 676292 711650
rect 676029 711592 676034 711648
rect 676090 711592 676292 711648
rect 676029 711590 676292 711592
rect 676029 711587 676095 711590
rect 674782 711180 674788 711244
rect 674852 711242 674858 711244
rect 674852 711182 676292 711242
rect 674852 711180 674858 711182
rect 676029 710834 676095 710837
rect 676029 710832 676292 710834
rect 676029 710776 676034 710832
rect 676090 710776 676292 710832
rect 676029 710774 676292 710776
rect 676029 710771 676095 710774
rect 675937 710426 676003 710429
rect 675937 710424 676292 710426
rect 675937 710368 675942 710424
rect 675998 710368 676292 710424
rect 675937 710366 676292 710368
rect 675937 710363 676003 710366
rect 678973 710018 679039 710021
rect 678973 710016 679052 710018
rect 678973 709960 678978 710016
rect 679034 709960 679052 710016
rect 678973 709958 679052 709960
rect 678973 709955 679039 709958
rect 673494 709548 673500 709612
rect 673564 709610 673570 709612
rect 673564 709550 676292 709610
rect 673564 709548 673570 709550
rect 675753 709202 675819 709205
rect 675753 709200 676292 709202
rect 675753 709144 675758 709200
rect 675814 709144 676292 709200
rect 675753 709142 676292 709144
rect 675753 709139 675819 709142
rect 675661 708794 675727 708797
rect 675661 708792 676292 708794
rect 675661 708736 675666 708792
rect 675722 708736 676292 708792
rect 675661 708734 676292 708736
rect 675661 708731 675727 708734
rect 676029 708386 676095 708389
rect 676029 708384 676292 708386
rect 676029 708328 676034 708384
rect 676090 708328 676292 708384
rect 676029 708326 676292 708328
rect 676029 708323 676095 708326
rect 676029 707978 676095 707981
rect 676029 707976 676292 707978
rect 676029 707920 676034 707976
rect 676090 707920 676292 707976
rect 676029 707918 676292 707920
rect 676029 707915 676095 707918
rect 676029 707570 676095 707573
rect 676029 707568 676292 707570
rect 676029 707512 676034 707568
rect 676090 707512 676292 707568
rect 676029 707510 676292 707512
rect 676029 707507 676095 707510
rect 676070 707236 676076 707300
rect 676140 707236 676146 707300
rect 676078 707162 676138 707236
rect 676078 707102 676292 707162
rect 676070 706828 676076 706892
rect 676140 706828 676146 706892
rect 676078 706754 676138 706828
rect 676078 706694 676292 706754
rect 676029 706346 676095 706349
rect 676029 706344 676292 706346
rect 676029 706288 676034 706344
rect 676090 706288 676292 706344
rect 676029 706286 676292 706288
rect 676029 706283 676095 706286
rect 684542 705500 684602 705908
rect 676029 705122 676095 705125
rect 676029 705120 676292 705122
rect 676029 705064 676034 705120
rect 676090 705064 676292 705120
rect 676029 705062 676292 705064
rect 676029 705059 676095 705062
rect 59353 704442 59419 704445
rect 59353 704440 64706 704442
rect 59353 704384 59358 704440
rect 59414 704384 64706 704440
rect 59353 704382 64706 704384
rect 59353 704379 59419 704382
rect 64646 703860 64706 704382
rect 59261 703354 59327 703357
rect 59261 703352 64706 703354
rect 59261 703296 59266 703352
rect 59322 703296 64706 703352
rect 59261 703294 64706 703296
rect 59261 703291 59327 703294
rect 64646 702678 64706 703294
rect 58525 702130 58591 702133
rect 58525 702128 64706 702130
rect 58525 702072 58530 702128
rect 58586 702072 64706 702128
rect 58525 702070 64706 702072
rect 58525 702067 58591 702070
rect 64646 701496 64706 702070
rect 59445 700906 59511 700909
rect 59445 700904 64706 700906
rect 59445 700848 59450 700904
rect 59506 700848 64706 700904
rect 59445 700846 64706 700848
rect 59445 700843 59511 700846
rect 64646 700314 64706 700846
rect 59629 699682 59695 699685
rect 59629 699680 64706 699682
rect 59629 699624 59634 699680
rect 59690 699624 64706 699680
rect 59629 699622 64706 699624
rect 59629 699619 59695 699622
rect 64646 699132 64706 699622
rect 675477 699410 675543 699413
rect 676990 699410 676996 699412
rect 675477 699408 676996 699410
rect 675477 699352 675482 699408
rect 675538 699352 676996 699408
rect 675477 699350 676996 699352
rect 675477 699347 675543 699350
rect 676990 699348 676996 699350
rect 677060 699348 677066 699412
rect 675569 699274 675635 699277
rect 676806 699274 676812 699276
rect 675569 699272 676812 699274
rect 675569 699216 675574 699272
rect 675630 699216 676812 699272
rect 675569 699214 676812 699216
rect 675569 699211 675635 699214
rect 676806 699212 676812 699214
rect 676876 699212 676882 699276
rect 673494 698260 673500 698324
rect 673564 698322 673570 698324
rect 675109 698322 675175 698325
rect 673564 698320 675175 698322
rect 673564 698264 675114 698320
rect 675170 698264 675175 698320
rect 673564 698262 675175 698264
rect 673564 698260 673570 698262
rect 675109 698259 675175 698262
rect 59169 698186 59235 698189
rect 59169 698184 64706 698186
rect 59169 698128 59174 698184
rect 59230 698128 64706 698184
rect 59169 698126 64706 698128
rect 59169 698123 59235 698126
rect 64646 697950 64706 698126
rect 675753 697234 675819 697237
rect 676070 697234 676076 697236
rect 675753 697232 676076 697234
rect 675753 697176 675758 697232
rect 675814 697176 676076 697232
rect 675753 697174 676076 697176
rect 675753 697171 675819 697174
rect 676070 697172 676076 697174
rect 676140 697172 676146 697236
rect 674966 695540 674972 695604
rect 675036 695602 675042 695604
rect 675109 695602 675175 695605
rect 675036 695600 675175 695602
rect 675036 695544 675114 695600
rect 675170 695544 675175 695600
rect 675036 695542 675175 695544
rect 675036 695540 675042 695542
rect 675109 695539 675175 695542
rect 674598 694724 674604 694788
rect 674668 694786 674674 694788
rect 675109 694786 675175 694789
rect 674668 694784 675175 694786
rect 674668 694728 675114 694784
rect 675170 694728 675175 694784
rect 674668 694726 675175 694728
rect 674668 694724 674674 694726
rect 675109 694723 675175 694726
rect 674782 694588 674788 694652
rect 674852 694650 674858 694652
rect 675109 694650 675175 694653
rect 674852 694648 675175 694650
rect 674852 694592 675114 694648
rect 675170 694592 675175 694648
rect 674852 694590 675175 694592
rect 674852 694588 674858 694590
rect 675109 694587 675175 694590
rect 675753 693018 675819 693021
rect 677174 693018 677180 693020
rect 675753 693016 677180 693018
rect 675753 692960 675758 693016
rect 675814 692960 677180 693016
rect 675753 692958 677180 692960
rect 675753 692955 675819 692958
rect 677174 692956 677180 692958
rect 677244 692956 677250 693020
rect 675753 690162 675819 690165
rect 676622 690162 676628 690164
rect 675753 690160 676628 690162
rect 675753 690104 675758 690160
rect 675814 690104 676628 690160
rect 675753 690102 676628 690104
rect 675753 690099 675819 690102
rect 676622 690100 676628 690102
rect 676692 690100 676698 690164
rect 649950 689482 650010 689980
rect 655605 689482 655671 689485
rect 649950 689480 655671 689482
rect 649950 689424 655610 689480
rect 655666 689424 655671 689480
rect 649950 689422 655671 689424
rect 655605 689419 655671 689422
rect 41505 688394 41571 688397
rect 41462 688392 41571 688394
rect 41462 688336 41510 688392
rect 41566 688336 41571 688392
rect 41462 688331 41571 688336
rect 41462 688092 41522 688331
rect 649950 688258 650010 688798
rect 655789 688258 655855 688261
rect 649950 688256 655855 688258
rect 649950 688200 655794 688256
rect 655850 688200 655855 688256
rect 649950 688198 655855 688200
rect 655789 688195 655855 688198
rect 41781 687714 41847 687717
rect 41492 687712 41847 687714
rect 41492 687656 41786 687712
rect 41842 687656 41847 687712
rect 41492 687654 41847 687656
rect 41781 687651 41847 687654
rect 41781 687306 41847 687309
rect 41492 687304 41847 687306
rect 41492 687248 41786 687304
rect 41842 687248 41847 687304
rect 41492 687246 41847 687248
rect 649950 687306 650010 687616
rect 655421 687306 655487 687309
rect 649950 687304 655487 687306
rect 649950 687248 655426 687304
rect 655482 687248 655487 687304
rect 649950 687246 655487 687248
rect 41781 687243 41847 687246
rect 655421 687243 655487 687246
rect 673862 687108 673868 687172
rect 673932 687170 673938 687172
rect 674281 687170 674347 687173
rect 673932 687168 674347 687170
rect 673932 687112 674286 687168
rect 674342 687112 674347 687168
rect 673932 687110 674347 687112
rect 673932 687108 673938 687110
rect 674281 687107 674347 687110
rect 655973 687034 656039 687037
rect 649950 687032 656039 687034
rect 649950 686976 655978 687032
rect 656034 686976 656039 687032
rect 649950 686974 656039 686976
rect 44589 686914 44659 686919
rect 41590 686854 44594 686914
rect 44654 686854 44668 686914
rect 44589 686849 44659 686854
rect 44589 686532 44659 686535
rect 41590 686530 44668 686532
rect 41590 686472 44594 686530
rect 44589 686470 44594 686472
rect 44654 686472 44668 686530
rect 44654 686470 44659 686472
rect 44589 686465 44659 686470
rect 649950 686434 650010 686974
rect 655973 686971 656039 686974
rect 43713 686082 43779 686085
rect 41492 686080 43779 686082
rect 41492 686024 43718 686080
rect 43774 686024 43779 686080
rect 41492 686022 43779 686024
rect 43713 686019 43779 686022
rect 654225 685810 654291 685813
rect 649950 685808 654291 685810
rect 649950 685752 654230 685808
rect 654286 685752 654291 685808
rect 649950 685750 654291 685752
rect 43069 685674 43135 685677
rect 41492 685672 43135 685674
rect 41492 685616 43074 685672
rect 43130 685616 43135 685672
rect 41492 685614 43135 685616
rect 43069 685611 43135 685614
rect 44681 685280 44751 685283
rect 41590 685278 44758 685280
rect 41590 685220 44686 685278
rect 44681 685218 44686 685220
rect 44746 685220 44758 685278
rect 649950 685252 650010 685750
rect 654225 685747 654291 685750
rect 674046 685748 674052 685812
rect 674116 685810 674122 685812
rect 675201 685810 675267 685813
rect 674116 685808 675267 685810
rect 674116 685752 675206 685808
rect 675262 685752 675267 685808
rect 674116 685750 675267 685752
rect 674116 685748 674122 685750
rect 675201 685747 675267 685750
rect 44746 685218 44751 685220
rect 44681 685213 44751 685218
rect 44681 684868 44751 684873
rect 44681 684866 44686 684868
rect 41590 684808 44686 684866
rect 44746 684866 44751 684868
rect 44746 684808 44758 684866
rect 41590 684806 44758 684808
rect 44681 684803 44751 684806
rect 44773 684488 44843 684493
rect 41590 684428 44778 684488
rect 44838 684428 44864 684488
rect 654133 684450 654199 684453
rect 649950 684448 654199 684450
rect 44773 684423 44843 684428
rect 649950 684392 654138 684448
rect 654194 684392 654199 684448
rect 649950 684390 654199 684392
rect 44773 684076 44843 684081
rect 44773 684070 44778 684076
rect 41590 684016 44778 684070
rect 44838 684070 44843 684076
rect 649950 684070 650010 684390
rect 654133 684387 654199 684390
rect 44838 684016 44864 684070
rect 41590 684010 44864 684016
rect 43253 683634 43319 683637
rect 41492 683632 43319 683634
rect 41492 683576 43258 683632
rect 43314 683576 43319 683632
rect 41492 683574 43319 683576
rect 43253 683571 43319 683574
rect 42241 683226 42307 683229
rect 41492 683224 42307 683226
rect 41492 683168 42246 683224
rect 42302 683168 42307 683224
rect 41492 683166 42307 683168
rect 42241 683163 42307 683166
rect 43529 682818 43595 682821
rect 41492 682816 43595 682818
rect 41492 682760 43534 682816
rect 43590 682760 43595 682816
rect 41492 682758 43595 682760
rect 43529 682755 43595 682758
rect 43437 682410 43503 682413
rect 41492 682408 43503 682410
rect 41492 682352 43442 682408
rect 43498 682352 43503 682408
rect 41492 682350 43503 682352
rect 43437 682347 43503 682350
rect 41873 682002 41939 682005
rect 41492 682000 41939 682002
rect 41492 681944 41878 682000
rect 41934 681944 41939 682000
rect 41492 681942 41939 681944
rect 41873 681939 41939 681942
rect 41462 681458 41522 681564
rect 41689 681458 41755 681461
rect 41462 681456 41755 681458
rect 41462 681400 41694 681456
rect 41750 681400 41755 681456
rect 41462 681398 41755 681400
rect 41689 681395 41755 681398
rect 42333 681186 42399 681189
rect 41492 681184 42399 681186
rect 41492 681128 42338 681184
rect 42394 681128 42399 681184
rect 41492 681126 42399 681128
rect 42333 681123 42399 681126
rect 43713 680778 43779 680781
rect 41492 680776 43779 680778
rect 41492 680720 43718 680776
rect 43774 680720 43779 680776
rect 41492 680718 43779 680720
rect 43713 680715 43779 680718
rect 42057 680370 42123 680373
rect 41492 680368 42123 680370
rect 41492 680312 42062 680368
rect 42118 680312 42123 680368
rect 41492 680310 42123 680312
rect 42057 680307 42123 680310
rect 674230 680308 674236 680372
rect 674300 680370 674306 680372
rect 674966 680370 674972 680372
rect 674300 680310 674972 680370
rect 674300 680308 674306 680310
rect 674966 680308 674972 680310
rect 675036 680308 675042 680372
rect 676622 680308 676628 680372
rect 676692 680370 676698 680372
rect 677358 680370 677364 680372
rect 676692 680310 677364 680370
rect 676692 680308 676698 680310
rect 677358 680308 677364 680310
rect 677428 680308 677434 680372
rect 43621 679962 43687 679965
rect 41492 679960 43687 679962
rect 41492 679904 43626 679960
rect 43682 679904 43687 679960
rect 41492 679902 43687 679904
rect 43621 679899 43687 679902
rect 42425 679554 42491 679557
rect 41492 679552 42491 679554
rect 41492 679496 42430 679552
rect 42486 679496 42491 679552
rect 41492 679494 42491 679496
rect 42425 679491 42491 679494
rect 30606 679012 30666 679116
rect 30598 678948 30604 679012
rect 30668 678948 30674 679012
rect 674046 678812 674052 678876
rect 674116 678874 674122 678876
rect 679157 678874 679223 678877
rect 674116 678872 679223 678874
rect 674116 678816 679162 678872
rect 679218 678816 679223 678872
rect 674116 678814 679223 678816
rect 674116 678812 674122 678814
rect 679157 678811 679223 678814
rect 41781 678738 41847 678741
rect 41492 678736 41847 678738
rect 41492 678680 41786 678736
rect 41842 678680 41847 678736
rect 41492 678678 41847 678680
rect 41781 678675 41847 678678
rect 41781 678330 41847 678333
rect 41492 678328 41847 678330
rect 41492 678272 41786 678328
rect 41842 678272 41847 678328
rect 41492 678270 41847 678272
rect 41781 678267 41847 678270
rect 676121 677972 676187 677973
rect 676070 677908 676076 677972
rect 676140 677970 676187 677972
rect 676140 677968 676232 677970
rect 676182 677912 676232 677968
rect 676140 677910 676232 677912
rect 676140 677908 676187 677910
rect 676121 677907 676187 677908
rect 41462 677786 41522 677892
rect 41462 677726 41890 677786
rect 30422 677076 30482 677484
rect 41830 676970 41890 677726
rect 41462 676910 41890 676970
rect 41462 676562 41522 676910
rect 60774 676562 60780 676564
rect 41462 676502 60780 676562
rect 60774 676500 60780 676502
rect 60844 676500 60850 676564
rect 676121 676476 676187 676477
rect 676070 676474 676076 676476
rect 676030 676414 676076 676474
rect 676140 676472 676187 676476
rect 676182 676416 676187 676472
rect 676070 676412 676076 676414
rect 676140 676412 676187 676416
rect 676121 676411 676187 676412
rect 5441 676290 5507 676293
rect 5441 676288 5550 676290
rect 5441 676232 5446 676288
rect 5502 676232 5550 676288
rect 5441 676227 5550 676232
rect 5490 676157 5550 676227
rect 5490 676152 5599 676157
rect 5490 676096 5538 676152
rect 5594 676096 5599 676152
rect 5490 676094 5599 676096
rect 5533 676091 5599 676094
rect 30557 676020 30623 676021
rect 30557 676018 30604 676020
rect 30512 676016 30604 676018
rect 30512 675960 30562 676016
rect 30512 675958 30604 675960
rect 30557 675956 30604 675958
rect 30668 675956 30674 676020
rect 30557 675955 30623 675956
rect 674230 674052 674236 674116
rect 674300 674114 674306 674116
rect 674966 674114 674972 674116
rect 674300 674054 674972 674114
rect 674300 674052 674306 674054
rect 674966 674052 674972 674054
rect 675036 674052 675042 674116
rect 676262 671125 676322 671364
rect 676213 671120 676322 671125
rect 676213 671064 676218 671120
rect 676274 671064 676322 671120
rect 676213 671062 676322 671064
rect 676213 671059 676279 671062
rect 676029 670986 676095 670989
rect 676029 670984 676292 670986
rect 676029 670928 676034 670984
rect 676090 670928 676292 670984
rect 676029 670926 676292 670928
rect 676029 670923 676095 670926
rect 42057 670714 42123 670717
rect 42558 670714 42564 670716
rect 42057 670712 42564 670714
rect 42057 670656 42062 670712
rect 42118 670656 42564 670712
rect 42057 670654 42564 670656
rect 42057 670651 42123 670654
rect 42558 670652 42564 670654
rect 42628 670652 42634 670716
rect 679022 670309 679082 670548
rect 678973 670304 679082 670309
rect 678973 670248 678978 670304
rect 679034 670248 679082 670304
rect 678973 670246 679082 670248
rect 678973 670243 679039 670246
rect 676121 669898 676187 669901
rect 676262 669898 676322 670140
rect 676121 669896 676322 669898
rect 676121 669840 676126 669896
rect 676182 669840 676322 669896
rect 676121 669838 676322 669840
rect 676121 669835 676187 669838
rect 676262 669493 676322 669732
rect 676262 669488 676371 669493
rect 676262 669432 676310 669488
rect 676366 669432 676371 669488
rect 676262 669430 676371 669432
rect 676305 669427 676371 669430
rect 676029 669354 676095 669357
rect 676029 669352 676292 669354
rect 676029 669296 676034 669352
rect 676090 669296 676292 669352
rect 676029 669294 676292 669296
rect 676029 669291 676095 669294
rect 676630 668676 676690 668916
rect 676622 668612 676628 668676
rect 676692 668612 676698 668676
rect 676262 668269 676322 668508
rect 676213 668264 676322 668269
rect 676213 668208 676218 668264
rect 676274 668208 676322 668264
rect 676213 668206 676322 668208
rect 676213 668203 676279 668206
rect 675293 668130 675359 668133
rect 675293 668128 676292 668130
rect 675293 668072 675298 668128
rect 675354 668072 676292 668128
rect 675293 668070 676292 668072
rect 675293 668067 675359 668070
rect 679022 667453 679082 667692
rect 678973 667448 679082 667453
rect 678973 667392 678978 667448
rect 679034 667392 679082 667448
rect 678973 667390 679082 667392
rect 678973 667387 679039 667390
rect 676262 667045 676322 667284
rect 676213 667040 676322 667045
rect 676213 666984 676218 667040
rect 676274 666984 676322 667040
rect 676213 666982 676322 666984
rect 679157 667042 679223 667045
rect 679157 667040 679266 667042
rect 679157 666984 679162 667040
rect 679218 666984 679266 667040
rect 676213 666979 676279 666982
rect 679157 666979 679266 666984
rect 679206 666876 679266 666979
rect 679065 666634 679131 666637
rect 679022 666632 679131 666634
rect 679022 666576 679070 666632
rect 679126 666576 679131 666632
rect 679022 666571 679131 666576
rect 679022 666468 679082 666571
rect 676029 666090 676095 666093
rect 676029 666088 676292 666090
rect 676029 666032 676034 666088
rect 676090 666032 676292 666088
rect 676029 666030 676292 666032
rect 676029 666027 676095 666030
rect 675150 665620 675156 665684
rect 675220 665682 675226 665684
rect 675220 665622 676292 665682
rect 675220 665620 675226 665622
rect 676029 665274 676095 665277
rect 676029 665272 676292 665274
rect 676029 665216 676034 665272
rect 676090 665216 676292 665272
rect 676029 665214 676292 665216
rect 676029 665211 676095 665214
rect 42558 665076 42564 665140
rect 42628 665138 42634 665140
rect 43253 665138 43319 665141
rect 42628 665136 43319 665138
rect 42628 665080 43258 665136
rect 43314 665080 43319 665136
rect 42628 665078 43319 665080
rect 42628 665076 42634 665078
rect 43253 665075 43319 665078
rect 676121 665002 676187 665005
rect 676121 665000 676322 665002
rect 676121 664944 676126 665000
rect 676182 664944 676322 665000
rect 676121 664942 676322 664944
rect 676121 664939 676187 664942
rect 676262 664836 676322 664942
rect 676029 664458 676095 664461
rect 676029 664456 676292 664458
rect 676029 664400 676034 664456
rect 676090 664400 676292 664456
rect 676029 664398 676292 664400
rect 676029 664395 676095 664398
rect 673678 663988 673684 664052
rect 673748 664050 673754 664052
rect 673748 663990 676292 664050
rect 673748 663988 673754 663990
rect 674414 663580 674420 663644
rect 674484 663642 674490 663644
rect 674484 663582 676292 663642
rect 674484 663580 674490 663582
rect 676029 663234 676095 663237
rect 676029 663232 676292 663234
rect 676029 663176 676034 663232
rect 676090 663176 676292 663232
rect 676029 663174 676292 663176
rect 676029 663171 676095 663174
rect 676029 662826 676095 662829
rect 676029 662824 676292 662826
rect 676029 662768 676034 662824
rect 676090 662768 676292 662824
rect 676029 662766 676292 662768
rect 676029 662763 676095 662766
rect 675702 662356 675708 662420
rect 675772 662418 675778 662420
rect 675772 662358 676292 662418
rect 675772 662356 675778 662358
rect 676990 662084 676996 662148
rect 677060 662084 677066 662148
rect 676998 661980 677058 662084
rect 676806 661676 676812 661740
rect 676876 661676 676882 661740
rect 676814 661572 676874 661676
rect 60641 661194 60707 661197
rect 60641 661192 64706 661194
rect 60641 661136 60646 661192
rect 60702 661136 64706 661192
rect 60641 661134 64706 661136
rect 60641 661131 60707 661134
rect 64646 660638 64706 661134
rect 679022 660925 679082 661164
rect 678973 660920 679082 660925
rect 678973 660864 678978 660920
rect 679034 660864 679082 660920
rect 678973 660862 679082 660864
rect 678973 660859 679039 660862
rect 684542 660348 684602 660756
rect 678973 660106 679039 660109
rect 678973 660104 679082 660106
rect 678973 660048 678978 660104
rect 679034 660048 679082 660104
rect 678973 660043 679082 660048
rect 679022 659940 679082 660043
rect 58525 659562 58591 659565
rect 58525 659560 64706 659562
rect 58525 659504 58530 659560
rect 58586 659504 64706 659560
rect 58525 659502 64706 659504
rect 58525 659499 58591 659502
rect 64646 659456 64706 659502
rect 58433 658882 58499 658885
rect 58433 658880 64706 658882
rect 58433 658824 58438 658880
rect 58494 658824 64706 658880
rect 58433 658822 64706 658824
rect 58433 658819 58499 658822
rect 64646 658274 64706 658822
rect 58617 657658 58683 657661
rect 58617 657656 64706 657658
rect 58617 657600 58622 657656
rect 58678 657600 64706 657656
rect 58617 657598 64706 657600
rect 58617 657595 58683 657598
rect 64646 657092 64706 657598
rect 58985 656570 59051 656573
rect 58985 656568 64706 656570
rect 58985 656512 58990 656568
rect 59046 656512 64706 656568
rect 58985 656510 64706 656512
rect 58985 656507 59051 656510
rect 64646 655910 64706 656510
rect 58433 655346 58499 655349
rect 58433 655344 64706 655346
rect 58433 655288 58438 655344
rect 58494 655288 64706 655344
rect 58433 655286 64706 655288
rect 58433 655283 58499 655286
rect 64646 654728 64706 655286
rect 673862 652836 673868 652900
rect 673932 652898 673938 652900
rect 675385 652898 675451 652901
rect 673932 652896 675451 652898
rect 673932 652840 675390 652896
rect 675446 652840 675451 652896
rect 673932 652838 675451 652840
rect 673932 652836 673938 652838
rect 675385 652835 675451 652838
rect 674046 652156 674052 652220
rect 674116 652218 674122 652220
rect 675477 652218 675543 652221
rect 674116 652216 675543 652218
rect 674116 652160 675482 652216
rect 675538 652160 675543 652216
rect 674116 652158 675543 652160
rect 674116 652156 674122 652158
rect 675477 652155 675543 652158
rect 674230 651612 674236 651676
rect 674300 651674 674306 651676
rect 675385 651674 675451 651677
rect 674300 651672 675451 651674
rect 674300 651616 675390 651672
rect 675446 651616 675451 651672
rect 674300 651614 675451 651616
rect 674300 651612 674306 651614
rect 675385 651611 675451 651614
rect 675150 649164 675156 649228
rect 675220 649226 675226 649228
rect 675385 649226 675451 649229
rect 675220 649224 675451 649226
rect 675220 649168 675390 649224
rect 675446 649168 675451 649224
rect 675220 649166 675451 649168
rect 675220 649164 675226 649166
rect 675385 649163 675451 649166
rect 41781 644942 41847 644945
rect 41492 644940 41847 644942
rect 41492 644884 41786 644940
rect 41842 644884 41847 644940
rect 41492 644882 41847 644884
rect 41781 644879 41847 644882
rect 41505 644738 41571 644741
rect 41462 644736 41571 644738
rect 41462 644680 41510 644736
rect 41566 644680 41571 644736
rect 41462 644675 41571 644680
rect 41462 644504 41522 644675
rect 41781 644126 41847 644129
rect 41492 644124 41847 644126
rect 41492 644068 41786 644124
rect 41842 644068 41847 644124
rect 41492 644066 41847 644068
rect 41781 644063 41847 644066
rect 44589 643714 44659 643719
rect 41582 643654 44594 643714
rect 44654 643654 44668 643714
rect 44589 643649 44659 643654
rect 44589 643332 44659 643335
rect 41582 643330 44668 643332
rect 41582 643272 44594 643330
rect 44589 643270 44594 643272
rect 44654 643272 44668 643330
rect 44654 643270 44659 643272
rect 44589 643265 44659 643270
rect 649950 643242 650010 643558
rect 655513 643242 655579 643245
rect 649950 643240 655579 643242
rect 649950 643184 655518 643240
rect 655574 643184 655579 643240
rect 649950 643182 655579 643184
rect 655513 643179 655579 643182
rect 43989 643106 44055 643109
rect 41462 643104 44055 643106
rect 41462 643048 43994 643104
rect 44050 643048 44055 643104
rect 41462 643046 44055 643048
rect 41462 642872 41522 643046
rect 43989 643043 44055 643046
rect 41462 642290 41522 642464
rect 43897 642290 43963 642293
rect 41462 642288 43963 642290
rect 41462 642232 43902 642288
rect 43958 642232 43963 642288
rect 41462 642230 43963 642232
rect 43897 642227 43963 642230
rect 44681 642080 44751 642083
rect 41564 642078 44758 642080
rect 41564 642020 44686 642078
rect 44681 642018 44686 642020
rect 44746 642020 44758 642078
rect 44746 642018 44751 642020
rect 44681 642013 44751 642018
rect 649950 641882 650010 642376
rect 655973 641882 656039 641885
rect 649950 641880 656039 641882
rect 649950 641824 655978 641880
rect 656034 641824 656039 641880
rect 649950 641822 656039 641824
rect 655973 641819 656039 641822
rect 44681 641668 44751 641673
rect 44681 641666 44686 641668
rect 41564 641608 44686 641666
rect 44746 641666 44751 641668
rect 44746 641608 44758 641666
rect 41564 641606 44758 641608
rect 44681 641603 44751 641606
rect 44773 641288 44843 641293
rect 41564 641228 44778 641288
rect 44838 641228 44864 641288
rect 44773 641223 44843 641228
rect 44773 640876 44843 640881
rect 44773 640870 44778 640876
rect 41564 640816 44778 640870
rect 44838 640870 44843 640876
rect 44838 640816 44864 640870
rect 41564 640810 44864 640816
rect 649950 640658 650010 641194
rect 656157 640658 656223 640661
rect 649950 640656 656223 640658
rect 649950 640600 656162 640656
rect 656218 640600 656223 640656
rect 649950 640598 656223 640600
rect 656157 640595 656223 640598
rect 41462 640386 41522 640424
rect 43069 640386 43135 640389
rect 41462 640384 43135 640386
rect 41462 640328 43074 640384
rect 43130 640328 43135 640384
rect 41462 640326 43135 640328
rect 43069 640323 43135 640326
rect 655697 640250 655763 640253
rect 649950 640248 655763 640250
rect 649950 640192 655702 640248
rect 655758 640192 655763 640248
rect 649950 640190 655763 640192
rect 41462 639842 41522 640016
rect 649950 640012 650010 640190
rect 655697 640187 655763 640190
rect 42333 639842 42399 639845
rect 41462 639840 42399 639842
rect 41462 639784 42338 639840
rect 42394 639784 42399 639840
rect 41462 639782 42399 639784
rect 42333 639779 42399 639782
rect 41462 639434 41522 639608
rect 44081 639434 44147 639437
rect 654409 639434 654475 639437
rect 41462 639432 44147 639434
rect 41462 639376 44086 639432
rect 44142 639376 44147 639432
rect 41462 639374 44147 639376
rect 44081 639371 44147 639374
rect 649950 639432 654475 639434
rect 649950 639376 654414 639432
rect 654470 639376 654475 639432
rect 649950 639374 654475 639376
rect 41462 639026 41522 639200
rect 43161 639026 43227 639029
rect 41462 639024 43227 639026
rect 41462 638968 43166 639024
rect 43222 638968 43227 639024
rect 41462 638966 43227 638968
rect 43161 638963 43227 638966
rect 649950 638830 650010 639374
rect 654409 639371 654475 639374
rect 41462 638618 41522 638792
rect 43621 638618 43687 638621
rect 41462 638616 43687 638618
rect 41462 638560 43626 638616
rect 43682 638560 43687 638616
rect 41462 638558 43687 638560
rect 43621 638555 43687 638558
rect 675385 638482 675451 638485
rect 675385 638480 675586 638482
rect 675385 638424 675390 638480
rect 675446 638424 675586 638480
rect 675385 638422 675586 638424
rect 675385 638419 675451 638422
rect 41462 638210 41522 638384
rect 42241 638210 42307 638213
rect 656433 638210 656499 638213
rect 41462 638208 42307 638210
rect 41462 638152 42246 638208
rect 42302 638152 42307 638208
rect 41462 638150 42307 638152
rect 42241 638147 42307 638150
rect 649950 638208 656499 638210
rect 649950 638152 656438 638208
rect 656494 638152 656499 638208
rect 649950 638150 656499 638152
rect 675526 638210 675586 638422
rect 675661 638210 675727 638213
rect 675526 638208 675727 638210
rect 675526 638152 675666 638208
rect 675722 638152 675727 638208
rect 675526 638150 675727 638152
rect 30238 637805 30298 637976
rect 30189 637800 30298 637805
rect 30189 637744 30194 637800
rect 30250 637744 30298 637800
rect 30189 637742 30298 637744
rect 30189 637739 30255 637742
rect 649950 637648 650010 638150
rect 656433 638147 656499 638150
rect 675661 638147 675727 638150
rect 30054 637397 30114 637568
rect 30054 637392 30163 637397
rect 30054 637336 30102 637392
rect 30158 637336 30163 637392
rect 30054 637334 30163 637336
rect 30097 637331 30163 637334
rect 41462 636986 41522 637160
rect 42701 636986 42767 636989
rect 41462 636984 42767 636986
rect 41462 636928 42706 636984
rect 42762 636928 42767 636984
rect 41462 636926 42767 636928
rect 42701 636923 42767 636926
rect 41462 636578 41522 636752
rect 43253 636578 43319 636581
rect 41462 636576 43319 636578
rect 41462 636520 43258 636576
rect 43314 636520 43319 636576
rect 41462 636518 43319 636520
rect 43253 636515 43319 636518
rect 41462 636170 41522 636344
rect 43437 636170 43503 636173
rect 41462 636168 43503 636170
rect 41462 636112 43442 636168
rect 43498 636112 43503 636168
rect 41462 636110 43503 636112
rect 43437 636107 43503 636110
rect 41462 635762 41522 635936
rect 43713 635762 43779 635765
rect 41462 635760 43779 635762
rect 41462 635704 43718 635760
rect 43774 635704 43779 635760
rect 41462 635702 43779 635704
rect 43713 635699 43779 635702
rect 41462 635354 41522 635528
rect 43345 635354 43411 635357
rect 41462 635352 43411 635354
rect 41462 635296 43350 635352
rect 43406 635296 43411 635352
rect 41462 635294 43411 635296
rect 43345 635291 43411 635294
rect 38518 634949 38578 635120
rect 38469 634944 38578 634949
rect 38469 634888 38474 634944
rect 38530 634888 38578 634944
rect 38469 634886 38578 634888
rect 38469 634883 38535 634886
rect 41462 634541 41522 634712
rect 41462 634536 41571 634541
rect 41462 634480 41510 634536
rect 41566 634480 41571 634536
rect 41462 634478 41571 634480
rect 41505 634475 41571 634478
rect 30422 633896 30482 634304
rect 41462 633317 41522 633488
rect 41462 633312 41571 633317
rect 41462 633256 41510 633312
rect 41566 633256 41571 633312
rect 41462 633254 41571 633256
rect 41505 633251 41571 633254
rect 674966 633056 674972 633120
rect 675036 633118 675042 633120
rect 676070 633118 676076 633120
rect 675036 633058 676076 633118
rect 675036 633056 675042 633058
rect 676070 633056 676076 633058
rect 676140 633056 676146 633120
rect 24761 632634 24827 632637
rect 30097 632634 30163 632637
rect 24761 632632 30163 632634
rect 24761 632576 24766 632632
rect 24822 632576 30102 632632
rect 30158 632576 30163 632632
rect 24761 632574 30163 632576
rect 24761 632571 24827 632574
rect 30097 632571 30163 632574
rect 42425 627468 42491 627469
rect 42374 627466 42380 627468
rect 42334 627406 42380 627466
rect 42444 627464 42491 627468
rect 42486 627408 42491 627464
rect 42374 627404 42380 627406
rect 42444 627404 42491 627408
rect 42425 627403 42491 627404
rect 43478 626996 43484 627060
rect 43548 627058 43554 627060
rect 43621 627058 43687 627061
rect 43548 627056 43687 627058
rect 43548 627000 43626 627056
rect 43682 627000 43687 627056
rect 43548 626998 43687 627000
rect 43548 626996 43554 626998
rect 43621 626995 43687 626998
rect 679022 626109 679082 626348
rect 678973 626104 679082 626109
rect 678973 626048 678978 626104
rect 679034 626048 679082 626104
rect 678973 626046 679082 626048
rect 678973 626043 679039 626046
rect 676262 625701 676322 625940
rect 676262 625696 676371 625701
rect 676262 625640 676310 625696
rect 676366 625640 676371 625696
rect 676262 625638 676371 625640
rect 676305 625635 676371 625638
rect 676029 625562 676095 625565
rect 676029 625560 676292 625562
rect 676029 625504 676034 625560
rect 676090 625504 676292 625560
rect 676029 625502 676292 625504
rect 676029 625499 676095 625502
rect 676262 624885 676322 625124
rect 676213 624880 676322 624885
rect 676213 624824 676218 624880
rect 676274 624824 676322 624880
rect 676213 624822 676322 624824
rect 676213 624819 676279 624822
rect 676121 624474 676187 624477
rect 676262 624474 676322 624716
rect 676121 624472 676322 624474
rect 676121 624416 676126 624472
rect 676182 624416 676322 624472
rect 676121 624414 676322 624416
rect 676121 624411 676187 624414
rect 676622 624412 676628 624476
rect 676692 624412 676698 624476
rect 676630 624308 676690 624412
rect 675937 623930 676003 623933
rect 675937 623928 676292 623930
rect 675937 623872 675942 623928
rect 675998 623872 676292 623928
rect 675937 623870 676292 623872
rect 675937 623867 676003 623870
rect 675937 623522 676003 623525
rect 675937 623520 676292 623522
rect 675937 623464 675942 623520
rect 675998 623464 676292 623520
rect 675937 623462 676292 623464
rect 675937 623459 676003 623462
rect 676121 622842 676187 622845
rect 676262 622842 676322 623084
rect 676121 622840 676322 622842
rect 676121 622784 676126 622840
rect 676182 622784 676322 622840
rect 676121 622782 676322 622784
rect 676121 622779 676187 622782
rect 676262 622437 676322 622676
rect 676262 622432 676371 622437
rect 676262 622376 676310 622432
rect 676366 622376 676371 622432
rect 676262 622374 676371 622376
rect 676305 622371 676371 622374
rect 43069 622162 43135 622165
rect 43478 622162 43484 622164
rect 43069 622160 43484 622162
rect 43069 622104 43074 622160
rect 43130 622104 43484 622160
rect 43069 622102 43484 622104
rect 43069 622099 43135 622102
rect 43478 622100 43484 622102
rect 43548 622100 43554 622164
rect 676262 622029 676322 622268
rect 676213 622024 676322 622029
rect 676213 621968 676218 622024
rect 676274 621968 676322 622024
rect 676213 621966 676322 621968
rect 676213 621963 676279 621966
rect 674782 621828 674788 621892
rect 674852 621890 674858 621892
rect 674852 621830 676292 621890
rect 674852 621828 674858 621830
rect 676029 621482 676095 621485
rect 676029 621480 676292 621482
rect 676029 621424 676034 621480
rect 676090 621424 676292 621480
rect 676029 621422 676292 621424
rect 676029 621419 676095 621422
rect 673494 621012 673500 621076
rect 673564 621074 673570 621076
rect 673564 621014 676292 621074
rect 673564 621012 673570 621014
rect 42333 620940 42399 620941
rect 42333 620938 42380 620940
rect 42288 620936 42380 620938
rect 42288 620880 42338 620936
rect 42288 620878 42380 620880
rect 42333 620876 42380 620878
rect 42444 620876 42450 620940
rect 42333 620875 42399 620876
rect 674414 620604 674420 620668
rect 674484 620666 674490 620668
rect 674484 620606 676292 620666
rect 674484 620604 674490 620606
rect 676029 620258 676095 620261
rect 676029 620256 676292 620258
rect 676029 620200 676034 620256
rect 676090 620200 676292 620256
rect 676029 620198 676292 620200
rect 676029 620195 676095 620198
rect 679065 619986 679131 619989
rect 679022 619984 679131 619986
rect 679022 619928 679070 619984
rect 679126 619928 679131 619984
rect 679022 619923 679131 619928
rect 679022 619820 679082 619923
rect 674966 619380 674972 619444
rect 675036 619442 675042 619444
rect 675036 619382 676292 619442
rect 675036 619380 675042 619382
rect 674598 618972 674604 619036
rect 674668 619034 674674 619036
rect 674668 618974 676292 619034
rect 674668 618972 674674 618974
rect 676029 618626 676095 618629
rect 676029 618624 676292 618626
rect 676029 618568 676034 618624
rect 676090 618568 676292 618624
rect 676029 618566 676292 618568
rect 676029 618563 676095 618566
rect 676029 618218 676095 618221
rect 676029 618216 676292 618218
rect 676029 618160 676034 618216
rect 676090 618160 676292 618216
rect 676029 618158 676292 618160
rect 676029 618155 676095 618158
rect 58157 617810 58223 617813
rect 676029 617810 676095 617813
rect 58157 617808 64706 617810
rect 58157 617752 58162 617808
rect 58218 617752 64706 617808
rect 58157 617750 64706 617752
rect 58157 617747 58223 617750
rect 64646 617416 64706 617750
rect 676029 617808 676292 617810
rect 676029 617752 676034 617808
rect 676090 617752 676292 617808
rect 676029 617750 676292 617752
rect 676029 617747 676095 617750
rect 677174 617476 677180 617540
rect 677244 617476 677250 617540
rect 677182 617372 677242 617476
rect 677358 617068 677364 617132
rect 677428 617068 677434 617132
rect 677366 616964 677426 617068
rect 58525 616858 58591 616861
rect 58525 616856 64706 616858
rect 58525 616800 58530 616856
rect 58586 616800 64706 616856
rect 58525 616798 64706 616800
rect 58525 616795 58591 616798
rect 64646 616234 64706 616798
rect 676213 616722 676279 616725
rect 676213 616720 676322 616722
rect 676213 616664 676218 616720
rect 676274 616664 676322 616720
rect 676213 616659 676322 616664
rect 676262 616556 676322 616659
rect 679022 615909 679082 616148
rect 679022 615904 679131 615909
rect 679022 615848 679070 615904
rect 679126 615848 679131 615904
rect 679022 615846 679131 615848
rect 679065 615843 679131 615846
rect 58525 615498 58591 615501
rect 58525 615496 64706 615498
rect 58525 615440 58530 615496
rect 58586 615440 64706 615496
rect 58525 615438 64706 615440
rect 58525 615435 58591 615438
rect 64646 615052 64706 615438
rect 679022 615332 679082 615740
rect 679065 615090 679131 615093
rect 679022 615088 679131 615090
rect 679022 615032 679070 615088
rect 679126 615032 679131 615088
rect 679022 615027 679131 615032
rect 679022 614924 679082 615027
rect 58157 614546 58223 614549
rect 58157 614544 64706 614546
rect 58157 614488 58162 614544
rect 58218 614488 64706 614544
rect 58157 614486 64706 614488
rect 58157 614483 58223 614486
rect 64646 613870 64706 614486
rect 57973 612642 58039 612645
rect 64646 612642 64706 612688
rect 57973 612640 64706 612642
rect 57973 612584 57978 612640
rect 58034 612584 64706 612640
rect 57973 612582 64706 612584
rect 57973 612579 58039 612582
rect 57973 612098 58039 612101
rect 57973 612096 64706 612098
rect 57973 612040 57978 612096
rect 58034 612040 64706 612096
rect 57973 612038 64706 612040
rect 57973 612035 58039 612038
rect 64646 611506 64706 612038
rect 674649 610194 674715 610197
rect 677174 610194 677180 610196
rect 674649 610192 677180 610194
rect 674649 610136 674654 610192
rect 674710 610136 677180 610192
rect 674649 610134 677180 610136
rect 674649 610131 674715 610134
rect 677174 610132 677180 610134
rect 677244 610132 677250 610196
rect 675293 610058 675359 610061
rect 677358 610058 677364 610060
rect 675293 610056 677364 610058
rect 675293 610000 675298 610056
rect 675354 610000 677364 610056
rect 675293 609998 677364 610000
rect 675293 609995 675359 609998
rect 677358 609996 677364 609998
rect 677428 609996 677434 610060
rect 673678 608092 673684 608156
rect 673748 608154 673754 608156
rect 675293 608154 675359 608157
rect 673748 608152 675359 608154
rect 673748 608096 675298 608152
rect 675354 608096 675359 608152
rect 673748 608094 675359 608096
rect 673748 608092 673754 608094
rect 675293 608091 675359 608094
rect 673494 607276 673500 607340
rect 673564 607338 673570 607340
rect 675293 607338 675359 607341
rect 673564 607336 675359 607338
rect 673564 607280 675298 607336
rect 675354 607280 675359 607336
rect 673564 607278 675359 607280
rect 673564 607276 673570 607278
rect 675293 607275 675359 607278
rect 674782 605100 674788 605164
rect 674852 605162 674858 605164
rect 675293 605162 675359 605165
rect 674852 605160 675359 605162
rect 674852 605104 675298 605160
rect 675354 605104 675359 605160
rect 674852 605102 675359 605104
rect 674852 605100 674858 605102
rect 675293 605099 675359 605102
rect 674966 604964 674972 605028
rect 675036 605026 675042 605028
rect 675201 605026 675267 605029
rect 675036 605024 675267 605026
rect 675036 604968 675206 605024
rect 675262 604968 675267 605024
rect 675036 604966 675267 604968
rect 675036 604964 675042 604966
rect 675201 604963 675267 604966
rect 674598 604420 674604 604484
rect 674668 604482 674674 604484
rect 675201 604482 675267 604485
rect 674668 604480 675267 604482
rect 674668 604424 675206 604480
rect 675262 604424 675267 604480
rect 674668 604422 675267 604424
rect 674668 604420 674674 604422
rect 675201 604419 675267 604422
rect 674414 601836 674420 601900
rect 674484 601898 674490 601900
rect 675201 601898 675267 601901
rect 674484 601896 675267 601898
rect 674484 601840 675206 601896
rect 675262 601840 675267 601896
rect 674484 601838 675267 601840
rect 674484 601836 674490 601838
rect 675201 601835 675267 601838
rect 41781 601762 41847 601765
rect 41492 601760 41847 601762
rect 41492 601704 41786 601760
rect 41842 601704 41847 601760
rect 41492 601702 41847 601704
rect 41781 601699 41847 601702
rect 41505 601490 41571 601493
rect 43897 601490 43963 601493
rect 41505 601488 43963 601490
rect 41505 601432 41510 601488
rect 41566 601432 43902 601488
rect 43958 601432 43963 601488
rect 41505 601430 43963 601432
rect 41505 601427 41571 601430
rect 43897 601427 43963 601430
rect 41462 601082 41522 601324
rect 42701 601082 42767 601085
rect 41462 601080 42767 601082
rect 41462 601024 42706 601080
rect 42762 601024 42767 601080
rect 41462 601022 42767 601024
rect 42701 601019 42767 601022
rect 41462 600674 41522 600916
rect 43069 600674 43135 600677
rect 41462 600672 43135 600674
rect 41462 600616 43074 600672
rect 43130 600616 43135 600672
rect 41462 600614 43135 600616
rect 43069 600611 43135 600614
rect 44589 600514 44659 600519
rect 41582 600454 44594 600514
rect 44654 600454 44668 600514
rect 44589 600449 44659 600454
rect 44589 600132 44659 600135
rect 41582 600130 44668 600132
rect 41582 600072 44594 600130
rect 44589 600070 44594 600072
rect 44654 600072 44668 600130
rect 44654 600070 44659 600072
rect 44589 600065 44659 600070
rect 41505 599858 41571 599861
rect 41462 599856 41571 599858
rect 41462 599800 41510 599856
rect 41566 599800 41571 599856
rect 41462 599795 41571 599800
rect 41462 599692 41522 599795
rect 43897 599314 43963 599317
rect 41492 599312 43963 599314
rect 41492 599256 43902 599312
rect 43958 599256 43963 599312
rect 41492 599254 43963 599256
rect 43897 599251 43963 599254
rect 42701 599178 42767 599181
rect 59261 599178 59327 599181
rect 42701 599176 59327 599178
rect 42701 599120 42706 599176
rect 42762 599120 59266 599176
rect 59322 599120 59327 599176
rect 42701 599118 59327 599120
rect 42701 599115 42767 599118
rect 59261 599115 59327 599118
rect 43069 599042 43135 599045
rect 59445 599042 59511 599045
rect 43069 599040 59511 599042
rect 43069 598984 43074 599040
rect 43130 598984 59450 599040
rect 59506 598984 59511 599040
rect 43069 598982 59511 598984
rect 43069 598979 43135 598982
rect 59445 598979 59511 598982
rect 44681 598880 44751 598883
rect 41530 598878 44758 598880
rect 41530 598820 44686 598878
rect 44681 598818 44686 598820
rect 44746 598820 44758 598878
rect 44746 598818 44751 598820
rect 44681 598813 44751 598818
rect 44681 598468 44751 598473
rect 44681 598466 44686 598468
rect 41530 598408 44686 598466
rect 44746 598466 44751 598468
rect 44746 598408 44758 598466
rect 41530 598406 44758 598408
rect 44681 598403 44751 598406
rect 44773 598088 44843 598093
rect 41530 598028 44778 598088
rect 44838 598028 44864 598088
rect 44773 598023 44843 598028
rect 649950 597818 650010 598336
rect 655881 597818 655947 597821
rect 649950 597816 655947 597818
rect 649950 597760 655886 597816
rect 655942 597760 655947 597816
rect 649950 597758 655947 597760
rect 655881 597755 655947 597758
rect 44773 597676 44843 597681
rect 44773 597670 44778 597676
rect 41530 597616 44778 597670
rect 44838 597670 44843 597676
rect 44838 597616 44864 597670
rect 41530 597610 44864 597616
rect 44081 597274 44147 597277
rect 41492 597272 44147 597274
rect 41492 597216 44086 597272
rect 44142 597216 44147 597272
rect 41492 597214 44147 597216
rect 44081 597211 44147 597214
rect 43161 596866 43227 596869
rect 41492 596864 43227 596866
rect 41492 596808 43166 596864
rect 43222 596808 43227 596864
rect 41492 596806 43227 596808
rect 43161 596803 43227 596806
rect 649950 596594 650010 597154
rect 655697 596594 655763 596597
rect 649950 596592 655763 596594
rect 649950 596536 655702 596592
rect 655758 596536 655763 596592
rect 649950 596534 655763 596536
rect 655697 596531 655763 596534
rect 43713 596458 43779 596461
rect 41492 596456 43779 596458
rect 41492 596400 43718 596456
rect 43774 596400 43779 596456
rect 41492 596398 43779 596400
rect 43713 596395 43779 596398
rect 43989 596050 44055 596053
rect 41492 596048 44055 596050
rect 41492 595992 43994 596048
rect 44050 595992 44055 596048
rect 41492 595990 44055 595992
rect 43989 595987 44055 595990
rect 43345 595642 43411 595645
rect 41492 595640 43411 595642
rect 41492 595584 43350 595640
rect 43406 595584 43411 595640
rect 41492 595582 43411 595584
rect 43345 595579 43411 595582
rect 649950 595506 650010 595972
rect 655789 595506 655855 595509
rect 649950 595504 655855 595506
rect 649950 595448 655794 595504
rect 655850 595448 655855 595504
rect 649950 595446 655855 595448
rect 655789 595443 655855 595446
rect 655421 595370 655487 595373
rect 649950 595368 655487 595370
rect 649950 595312 655426 595368
rect 655482 595312 655487 595368
rect 649950 595310 655487 595312
rect 41781 595234 41847 595237
rect 41492 595232 41847 595234
rect 41492 595176 41786 595232
rect 41842 595176 41847 595232
rect 41492 595174 41847 595176
rect 41781 595171 41847 595174
rect 42425 594826 42491 594829
rect 41492 594824 42491 594826
rect 41492 594768 42430 594824
rect 42486 594768 42491 594824
rect 649950 594790 650010 595310
rect 655421 595307 655487 595310
rect 41492 594766 42491 594768
rect 42425 594763 42491 594766
rect 43437 594418 43503 594421
rect 41492 594416 43503 594418
rect 41492 594360 43442 594416
rect 43498 594360 43503 594416
rect 41492 594358 43503 594360
rect 43437 594355 43503 594358
rect 656801 594282 656867 594285
rect 649950 594280 656867 594282
rect 649950 594224 656806 594280
rect 656862 594224 656867 594280
rect 649950 594222 656867 594224
rect 43529 594010 43595 594013
rect 41492 594008 43595 594010
rect 41492 593952 43534 594008
rect 43590 593952 43595 594008
rect 41492 593950 43595 593952
rect 43529 593947 43595 593950
rect 649950 593608 650010 594222
rect 656801 594219 656867 594222
rect 38518 593333 38578 593572
rect 38518 593328 38627 593333
rect 38518 593272 38566 593328
rect 38622 593272 38627 593328
rect 38518 593270 38627 593272
rect 38561 593267 38627 593270
rect 43805 593194 43871 593197
rect 41492 593192 43871 593194
rect 41492 593136 43810 593192
rect 43866 593136 43871 593192
rect 41492 593134 43871 593136
rect 43805 593131 43871 593134
rect 655605 593058 655671 593061
rect 649950 593056 655671 593058
rect 649950 593000 655610 593056
rect 655666 593000 655671 593056
rect 649950 592998 655671 593000
rect 44081 592786 44147 592789
rect 41492 592784 44147 592786
rect 41492 592728 44086 592784
rect 44142 592728 44147 592784
rect 41492 592726 44147 592728
rect 44081 592723 44147 592726
rect 649950 592426 650010 592998
rect 655605 592995 655671 592998
rect 43621 592378 43687 592381
rect 41492 592376 43687 592378
rect 41492 592320 43626 592376
rect 43682 592320 43687 592376
rect 41492 592318 43687 592320
rect 43621 592315 43687 592318
rect 43161 591970 43227 591973
rect 41492 591968 43227 591970
rect 41492 591912 43166 591968
rect 43222 591912 43227 591968
rect 41492 591910 43227 591912
rect 43161 591907 43227 591910
rect 41462 591293 41522 591532
rect 41462 591288 41571 591293
rect 41462 591232 41510 591288
rect 41566 591232 41571 591288
rect 41462 591230 41571 591232
rect 41505 591227 41571 591230
rect 30422 590716 30482 591124
rect 41462 590069 41522 590308
rect 41462 590064 41571 590069
rect 41462 590008 41510 590064
rect 41566 590008 41571 590064
rect 41462 590006 41571 590008
rect 41505 590003 41571 590006
rect 43069 585308 43135 585309
rect 43069 585304 43116 585308
rect 43180 585306 43186 585308
rect 43069 585248 43074 585304
rect 43069 585244 43116 585248
rect 43180 585246 43226 585306
rect 43180 585244 43186 585246
rect 43069 585243 43135 585244
rect 43345 583810 43411 583813
rect 43529 583810 43595 583813
rect 43345 583808 43595 583810
rect 43345 583752 43350 583808
rect 43406 583752 43534 583808
rect 43590 583752 43595 583808
rect 43345 583750 43595 583752
rect 43345 583747 43411 583750
rect 43529 583747 43595 583750
rect 43069 581364 43135 581365
rect 43069 581362 43116 581364
rect 43024 581360 43116 581362
rect 43024 581304 43074 581360
rect 43024 581302 43116 581304
rect 43069 581300 43116 581302
rect 43180 581300 43186 581364
rect 43069 581299 43135 581300
rect 676121 580954 676187 580957
rect 676262 580954 676322 581060
rect 676121 580952 676322 580954
rect 676121 580896 676126 580952
rect 676182 580896 676322 580952
rect 676121 580894 676322 580896
rect 676121 580891 676187 580894
rect 676262 580549 676322 580652
rect 676262 580544 676371 580549
rect 676262 580488 676310 580544
rect 676366 580488 676371 580544
rect 676262 580486 676371 580488
rect 676305 580483 676371 580486
rect 676262 580141 676322 580244
rect 676213 580136 676322 580141
rect 676213 580080 676218 580136
rect 676274 580080 676322 580136
rect 676213 580078 676322 580080
rect 676213 580075 676279 580078
rect 676262 579733 676322 579836
rect 676213 579728 676322 579733
rect 676213 579672 676218 579728
rect 676274 579672 676322 579728
rect 676213 579670 676322 579672
rect 676213 579667 676279 579670
rect 676070 579260 676076 579324
rect 676140 579322 676146 579324
rect 676262 579322 676322 579428
rect 676140 579262 676322 579322
rect 676140 579260 676146 579262
rect 676029 579050 676095 579053
rect 676029 579048 676292 579050
rect 676029 578992 676034 579048
rect 676090 578992 676292 579048
rect 676029 578990 676292 578992
rect 676029 578987 676095 578990
rect 676262 578509 676322 578612
rect 676213 578504 676322 578509
rect 676213 578448 676218 578504
rect 676274 578448 676322 578504
rect 676213 578446 676322 578448
rect 676213 578443 676279 578446
rect 676121 578098 676187 578101
rect 676262 578098 676322 578204
rect 676121 578096 676322 578098
rect 676121 578040 676126 578096
rect 676182 578040 676322 578096
rect 676121 578038 676322 578040
rect 676121 578035 676187 578038
rect 676630 577692 676690 577796
rect 676622 577628 676628 577692
rect 676692 577628 676698 577692
rect 676262 577285 676322 577388
rect 676213 577280 676322 577285
rect 676213 577224 676218 577280
rect 676274 577224 676322 577280
rect 676213 577222 676322 577224
rect 676213 577219 676279 577222
rect 676814 576876 676874 576980
rect 676806 576812 676812 576876
rect 676876 576812 676882 576876
rect 674230 576540 674236 576604
rect 674300 576602 674306 576604
rect 674300 576542 676292 576602
rect 674300 576540 674306 576542
rect 676029 576194 676095 576197
rect 676029 576192 676292 576194
rect 676029 576136 676034 576192
rect 676090 576136 676292 576192
rect 676029 576134 676292 576136
rect 676029 576131 676095 576134
rect 673862 575724 673868 575788
rect 673932 575786 673938 575788
rect 673932 575726 676292 575786
rect 673932 575724 673938 575726
rect 675937 575378 676003 575381
rect 675937 575376 676292 575378
rect 675937 575320 675942 575376
rect 675998 575320 676292 575376
rect 675937 575318 676292 575320
rect 675937 575315 676003 575318
rect 678973 575242 679039 575245
rect 678973 575240 679082 575242
rect 678973 575184 678978 575240
rect 679034 575184 679082 575240
rect 678973 575179 679082 575184
rect 679022 574940 679082 575179
rect 58525 574834 58591 574837
rect 58525 574832 64706 574834
rect 58525 574776 58530 574832
rect 58586 574776 64706 574832
rect 58525 574774 64706 574776
rect 58525 574771 58591 574774
rect 64646 574194 64706 574774
rect 676029 574562 676095 574565
rect 676029 574560 676292 574562
rect 676029 574504 676034 574560
rect 676090 574504 676292 574560
rect 676029 574502 676292 574504
rect 676029 574499 676095 574502
rect 674046 574092 674052 574156
rect 674116 574154 674122 574156
rect 674116 574094 676292 574154
rect 674116 574092 674122 574094
rect 675150 573684 675156 573748
rect 675220 573746 675226 573748
rect 675220 573686 676292 573746
rect 675220 573684 675226 573686
rect 59353 573610 59419 573613
rect 59353 573608 64706 573610
rect 59353 573552 59358 573608
rect 59414 573552 64706 573608
rect 59353 573550 64706 573552
rect 59353 573547 59419 573550
rect 64646 573012 64706 573550
rect 675569 573338 675635 573341
rect 675569 573336 676292 573338
rect 675569 573280 675574 573336
rect 675630 573280 676292 573336
rect 675569 573278 676292 573280
rect 675569 573275 675635 573278
rect 676029 572930 676095 572933
rect 676029 572928 676292 572930
rect 676029 572872 676034 572928
rect 676090 572872 676292 572928
rect 676029 572870 676292 572872
rect 676029 572867 676095 572870
rect 676029 572522 676095 572525
rect 676029 572520 676292 572522
rect 676029 572464 676034 572520
rect 676090 572464 676292 572520
rect 676029 572462 676292 572464
rect 676029 572459 676095 572462
rect 60641 572386 60707 572389
rect 60641 572384 64706 572386
rect 60641 572328 60646 572384
rect 60702 572328 64706 572384
rect 60641 572326 64706 572328
rect 60641 572323 60707 572326
rect 64646 571830 64706 572326
rect 676029 572114 676095 572117
rect 676029 572112 676292 572114
rect 676029 572056 676034 572112
rect 676090 572056 676292 572112
rect 676029 572054 676292 572056
rect 676029 572051 676095 572054
rect 677174 571916 677180 571980
rect 677244 571916 677250 571980
rect 677182 571676 677242 571916
rect 674281 571570 674347 571573
rect 676990 571570 676996 571572
rect 674281 571568 676996 571570
rect 674281 571512 674286 571568
rect 674342 571512 676996 571568
rect 674281 571510 676996 571512
rect 674281 571507 674347 571510
rect 676990 571508 676996 571510
rect 677060 571508 677066 571572
rect 677358 571508 677364 571572
rect 677428 571508 677434 571572
rect 59445 571298 59511 571301
rect 59445 571296 64706 571298
rect 59445 571240 59450 571296
rect 59506 571240 64706 571296
rect 677366 571268 677426 571508
rect 59445 571238 64706 571240
rect 59445 571235 59511 571238
rect 64646 570648 64706 571238
rect 679022 570757 679082 570860
rect 678973 570752 679082 570757
rect 678973 570696 678978 570752
rect 679034 570696 679082 570752
rect 678973 570694 679082 570696
rect 678973 570691 679039 570694
rect 58709 570074 58775 570077
rect 58709 570072 64706 570074
rect 58709 570016 58714 570072
rect 58770 570016 64706 570072
rect 684542 570044 684602 570452
rect 58709 570014 64706 570016
rect 58709 570011 58775 570014
rect 64646 569466 64706 570014
rect 678973 569938 679039 569941
rect 678973 569936 679082 569938
rect 678973 569880 678978 569936
rect 679034 569880 679082 569936
rect 678973 569875 679082 569880
rect 679022 569636 679082 569875
rect 59261 568578 59327 568581
rect 59261 568576 64706 568578
rect 59261 568520 59266 568576
rect 59322 568520 64706 568576
rect 59261 568518 64706 568520
rect 59261 568515 59327 568518
rect 64646 568284 64706 568518
rect 674046 562668 674052 562732
rect 674116 562730 674122 562732
rect 675477 562730 675543 562733
rect 674116 562728 675543 562730
rect 674116 562672 675482 562728
rect 675538 562672 675543 562728
rect 674116 562670 675543 562672
rect 674116 562668 674122 562670
rect 675477 562667 675543 562670
rect 675150 562260 675156 562324
rect 675220 562322 675226 562324
rect 675293 562322 675359 562325
rect 675220 562320 675359 562322
rect 675220 562264 675298 562320
rect 675354 562264 675359 562320
rect 675220 562262 675359 562264
rect 675220 562260 675226 562262
rect 675293 562259 675359 562262
rect 674230 561172 674236 561236
rect 674300 561234 674306 561236
rect 675477 561234 675543 561237
rect 674300 561232 675543 561234
rect 674300 561176 675482 561232
rect 675538 561176 675543 561232
rect 674300 561174 675543 561176
rect 674300 561172 674306 561174
rect 675477 561171 675543 561174
rect 41505 558786 41571 558789
rect 41462 558784 41571 558786
rect 41462 558728 41510 558784
rect 41566 558728 41571 558784
rect 41462 558723 41571 558728
rect 41462 558484 41522 558723
rect 41505 558378 41571 558381
rect 41462 558376 41571 558378
rect 41462 558320 41510 558376
rect 41566 558320 41571 558376
rect 41462 558315 41571 558320
rect 41462 558076 41522 558315
rect 41462 557565 41522 557668
rect 41462 557560 41571 557565
rect 41462 557504 41510 557560
rect 41566 557504 41571 557560
rect 41462 557502 41571 557504
rect 41505 557499 41571 557502
rect 44589 557314 44659 557319
rect 41574 557254 44594 557314
rect 44654 557254 44668 557314
rect 44589 557249 44659 557254
rect 44589 556932 44659 556935
rect 41574 556930 44668 556932
rect 41574 556872 44594 556930
rect 44589 556870 44594 556872
rect 44654 556872 44668 556930
rect 44654 556870 44659 556872
rect 44589 556865 44659 556870
rect 43897 556474 43963 556477
rect 41492 556472 43963 556474
rect 41492 556416 43902 556472
rect 43958 556416 43963 556472
rect 41492 556414 43963 556416
rect 43897 556411 43963 556414
rect 42558 556066 42564 556068
rect 41492 556006 42564 556066
rect 42558 556004 42564 556006
rect 42628 556004 42634 556068
rect 44681 555680 44751 555683
rect 41552 555678 44758 555680
rect 38150 555525 38210 555628
rect 41552 555620 44686 555678
rect 44681 555618 44686 555620
rect 44746 555620 44758 555678
rect 44746 555618 44751 555620
rect 44681 555613 44751 555618
rect 38101 555520 38210 555525
rect 38101 555464 38106 555520
rect 38162 555464 38210 555520
rect 38101 555462 38210 555464
rect 38101 555459 38167 555462
rect 44681 555268 44751 555273
rect 44681 555266 44686 555268
rect 41552 555208 44686 555266
rect 44746 555266 44751 555268
rect 44746 555208 44758 555266
rect 41552 555206 44758 555208
rect 44681 555203 44751 555206
rect 675293 554980 675359 554981
rect 675293 554976 675340 554980
rect 675404 554978 675410 554980
rect 675293 554920 675298 554976
rect 675293 554916 675340 554920
rect 675404 554918 675450 554978
rect 675404 554916 675410 554918
rect 675293 554915 675359 554916
rect 44773 554888 44843 554893
rect 41552 554828 44778 554888
rect 44838 554828 44864 554888
rect 44773 554823 44843 554828
rect 673545 554706 673611 554709
rect 675334 554706 675340 554708
rect 673545 554704 675340 554706
rect 673545 554648 673550 554704
rect 673606 554648 675340 554704
rect 673545 554646 675340 554648
rect 673545 554643 673611 554646
rect 675334 554644 675340 554646
rect 675404 554644 675410 554708
rect 44773 554476 44843 554481
rect 44773 554470 44778 554476
rect 41552 554416 44778 554470
rect 44838 554470 44843 554476
rect 44838 554416 44864 554470
rect 41552 554410 44864 554416
rect 41462 553890 41522 553996
rect 41638 553890 41644 553892
rect 41462 553830 41644 553890
rect 41638 553828 41644 553830
rect 41708 553828 41714 553892
rect 43345 553618 43411 553621
rect 41492 553616 43411 553618
rect 41492 553560 43350 553616
rect 43406 553560 43411 553616
rect 41492 553558 43411 553560
rect 43345 553555 43411 553558
rect 649950 553346 650010 553914
rect 655605 553346 655671 553349
rect 649950 553344 655671 553346
rect 649950 553288 655610 553344
rect 655666 553288 655671 553344
rect 649950 553286 655671 553288
rect 655605 553283 655671 553286
rect 42926 553210 42932 553212
rect 41492 553150 42932 553210
rect 42926 553148 42932 553150
rect 42996 553148 43002 553212
rect 42190 552802 42196 552804
rect 41492 552742 42196 552802
rect 42190 552740 42196 552742
rect 42260 552740 42266 552804
rect 42374 552394 42380 552396
rect 41492 552334 42380 552394
rect 42374 552332 42380 552334
rect 42444 552332 42450 552396
rect 649950 552122 650010 552732
rect 655421 552122 655487 552125
rect 649950 552120 655487 552122
rect 649950 552064 655426 552120
rect 655482 552064 655487 552120
rect 649950 552062 655487 552064
rect 655421 552059 655487 552062
rect 41781 551986 41847 551989
rect 41492 551984 41847 551986
rect 41492 551928 41786 551984
rect 41842 551928 41847 551984
rect 41492 551926 41847 551928
rect 41781 551923 41847 551926
rect 42006 551578 42012 551580
rect 41492 551518 42012 551578
rect 42006 551516 42012 551518
rect 42076 551516 42082 551580
rect 41462 551036 41522 551140
rect 41454 550972 41460 551036
rect 41524 550972 41530 551036
rect 649950 551034 650010 551550
rect 655513 551034 655579 551037
rect 649950 551032 655579 551034
rect 649950 550976 655518 551032
rect 655574 550976 655579 551032
rect 649950 550974 655579 550976
rect 655513 550971 655579 550974
rect 655973 550898 656039 550901
rect 649950 550896 656039 550898
rect 649950 550840 655978 550896
rect 656034 550840 656039 550896
rect 649950 550838 656039 550840
rect 41822 550762 41828 550764
rect 41492 550702 41828 550762
rect 41822 550700 41828 550702
rect 41892 550700 41898 550764
rect 649950 550368 650010 550838
rect 655973 550835 656039 550838
rect 43161 550354 43227 550357
rect 41492 550352 43227 550354
rect 41492 550296 43166 550352
rect 43222 550296 43227 550352
rect 41492 550294 43227 550296
rect 43161 550291 43227 550294
rect 41462 549810 41522 549916
rect 41597 549810 41663 549813
rect 41462 549808 41663 549810
rect 41462 549752 41602 549808
rect 41658 549752 41663 549808
rect 41462 549750 41663 549752
rect 41597 549747 41663 549750
rect 41462 549405 41522 549508
rect 41413 549400 41522 549405
rect 41413 549344 41418 549400
rect 41474 549344 41522 549400
rect 41413 549342 41522 549344
rect 41413 549339 41479 549342
rect 654225 549266 654291 549269
rect 649950 549264 654291 549266
rect 649950 549208 654230 549264
rect 654286 549208 654291 549264
rect 649950 549206 654291 549208
rect 649950 549186 650010 549206
rect 654225 549203 654291 549206
rect 41462 548997 41522 549100
rect 41462 548992 41571 548997
rect 41462 548936 41510 548992
rect 41566 548936 41571 548992
rect 41462 548934 41571 548936
rect 41505 548931 41571 548934
rect 41462 548589 41522 548692
rect 41462 548584 41571 548589
rect 654133 548586 654199 548589
rect 41462 548528 41510 548584
rect 41566 548528 41571 548584
rect 41462 548526 41571 548528
rect 41505 548523 41571 548526
rect 649950 548584 654199 548586
rect 649950 548528 654138 548584
rect 654194 548528 654199 548584
rect 649950 548526 654199 548528
rect 41462 548181 41522 548284
rect 41462 548176 41571 548181
rect 41462 548120 41510 548176
rect 41566 548120 41571 548176
rect 41462 548118 41571 548120
rect 41505 548115 41571 548118
rect 649950 548004 650010 548526
rect 654133 548523 654199 548526
rect 30422 547468 30482 547876
rect 41462 546957 41522 547060
rect 41462 546952 41571 546957
rect 41462 546896 41510 546952
rect 41566 546896 41571 546952
rect 41462 546894 41571 546896
rect 41505 546891 41571 546894
rect 674414 546484 674420 546548
rect 674484 546546 674490 546548
rect 677501 546546 677567 546549
rect 674484 546544 677567 546546
rect 674484 546488 677506 546544
rect 677562 546488 677567 546544
rect 674484 546486 677567 546488
rect 674484 546484 674490 546486
rect 677501 546483 677567 546486
rect 38101 546410 38167 546413
rect 39982 546410 39988 546412
rect 38101 546408 39988 546410
rect 38101 546352 38106 546408
rect 38162 546352 39988 546408
rect 38101 546350 39988 546352
rect 38101 546347 38167 546350
rect 39982 546348 39988 546350
rect 40052 546348 40058 546412
rect 674598 543628 674604 543692
rect 674668 543690 674674 543692
rect 679157 543690 679223 543693
rect 674668 543688 679223 543690
rect 674668 543632 679162 543688
rect 679218 543632 679223 543688
rect 674668 543630 679223 543632
rect 674668 543628 674674 543630
rect 679157 543627 679223 543630
rect 673494 543492 673500 543556
rect 673564 543554 673570 543556
rect 679341 543554 679407 543557
rect 673564 543552 679407 543554
rect 673564 543496 679346 543552
rect 679402 543496 679407 543552
rect 673564 543494 679407 543496
rect 673564 543492 673570 543494
rect 679341 543491 679407 543494
rect 675937 543350 676003 543353
rect 676070 543350 676076 543352
rect 675937 543348 676076 543350
rect 675937 543292 675942 543348
rect 675998 543292 676076 543348
rect 675937 543290 676076 543292
rect 675937 543287 676003 543290
rect 676070 543288 676076 543290
rect 676140 543288 676146 543352
rect 675937 539620 676003 539621
rect 675886 539618 675892 539620
rect 675846 539558 675892 539618
rect 675956 539616 676003 539620
rect 675998 539560 676003 539616
rect 675886 539556 675892 539558
rect 675956 539556 676003 539560
rect 675937 539555 676003 539556
rect 42374 538732 42380 538796
rect 42444 538794 42450 538796
rect 43345 538794 43411 538797
rect 42444 538792 43411 538794
rect 42444 538736 43350 538792
rect 43406 538736 43411 538792
rect 42444 538734 43411 538736
rect 42444 538732 42450 538734
rect 43345 538731 43411 538734
rect 676262 535941 676322 536112
rect 676213 535936 676322 535941
rect 676213 535880 676218 535936
rect 676274 535880 676322 535936
rect 676213 535878 676322 535880
rect 676213 535875 676279 535878
rect 41822 535740 41828 535804
rect 41892 535802 41898 535804
rect 42241 535802 42307 535805
rect 41892 535800 42307 535802
rect 41892 535744 42246 535800
rect 42302 535744 42307 535800
rect 41892 535742 42307 535744
rect 41892 535740 41898 535742
rect 42241 535739 42307 535742
rect 676029 535734 676095 535737
rect 676029 535732 676292 535734
rect 676029 535676 676034 535732
rect 676090 535676 676292 535732
rect 676029 535674 676292 535676
rect 676029 535671 676095 535674
rect 679022 535125 679082 535296
rect 678973 535120 679082 535125
rect 678973 535064 678978 535120
rect 679034 535064 679082 535120
rect 678973 535062 679082 535064
rect 678973 535059 679039 535062
rect 675886 534986 675892 534988
rect 675872 534926 675892 534986
rect 675886 534924 675892 534926
rect 675956 534986 675962 534988
rect 675956 534926 676322 534986
rect 675956 534924 675962 534926
rect 676262 534888 676322 534926
rect 675845 534510 675911 534513
rect 675845 534508 676292 534510
rect 675845 534452 675850 534508
rect 675906 534452 676292 534508
rect 675845 534450 676292 534452
rect 675845 534447 675911 534450
rect 676029 534102 676095 534105
rect 676029 534100 676292 534102
rect 676029 534044 676034 534100
rect 676090 534044 676292 534100
rect 676029 534042 676292 534044
rect 676029 534039 676095 534042
rect 673678 533836 673684 533900
rect 673748 533898 673754 533900
rect 679249 533898 679315 533901
rect 673748 533896 679315 533898
rect 673748 533840 679254 533896
rect 679310 533840 679315 533896
rect 673748 533838 679315 533840
rect 673748 533836 673754 533838
rect 679249 533835 679315 533838
rect 677366 533493 677426 533664
rect 676622 533428 676628 533492
rect 676692 533428 676698 533492
rect 677366 533488 677475 533493
rect 677366 533432 677414 533488
rect 677470 533432 677475 533488
rect 677366 533430 677475 533432
rect 676630 533276 676690 533428
rect 677409 533427 677475 533430
rect 42190 533020 42196 533084
rect 42260 533082 42266 533084
rect 43069 533082 43135 533085
rect 42260 533080 43135 533082
rect 42260 533024 43074 533080
rect 43130 533024 43135 533080
rect 42260 533022 43135 533024
rect 42260 533020 42266 533022
rect 43069 533019 43135 533022
rect 674966 533020 674972 533084
rect 675036 533082 675042 533084
rect 679065 533082 679131 533085
rect 675036 533080 679131 533082
rect 675036 533024 679070 533080
rect 679126 533024 679131 533080
rect 675036 533022 679131 533024
rect 675036 533020 675042 533022
rect 679065 533019 679131 533022
rect 41638 532884 41644 532948
rect 41708 532946 41714 532948
rect 41708 532886 42442 532946
rect 41708 532884 41714 532886
rect 42382 532813 42442 532886
rect 41454 532748 41460 532812
rect 41524 532810 41530 532812
rect 42149 532810 42215 532813
rect 41524 532808 42215 532810
rect 41524 532752 42154 532808
rect 42210 532752 42215 532808
rect 41524 532750 42215 532752
rect 42382 532808 42491 532813
rect 42382 532752 42430 532808
rect 42486 532752 42491 532808
rect 42382 532750 42491 532752
rect 41524 532748 41530 532750
rect 42149 532747 42215 532750
rect 42425 532747 42491 532750
rect 674782 532748 674788 532812
rect 674852 532810 674858 532812
rect 676029 532810 676095 532813
rect 674852 532808 676095 532810
rect 674852 532752 676034 532808
rect 676090 532752 676095 532808
rect 674852 532750 676095 532752
rect 674852 532748 674858 532750
rect 676029 532747 676095 532750
rect 676121 532674 676187 532677
rect 676262 532674 676322 532848
rect 676121 532672 676322 532674
rect 676121 532616 676126 532672
rect 676182 532616 676322 532672
rect 676121 532614 676322 532616
rect 676121 532611 676187 532614
rect 676806 532612 676812 532676
rect 676876 532612 676882 532676
rect 676814 532470 676874 532612
rect 676322 532440 676874 532470
rect 676322 532410 676844 532440
rect 675937 532062 676003 532065
rect 675937 532060 676292 532062
rect 675937 532004 675942 532060
rect 675998 532004 676292 532060
rect 675937 532002 676292 532004
rect 675937 531999 676003 532002
rect 59445 531722 59511 531725
rect 59445 531720 64706 531722
rect 59445 531664 59450 531720
rect 59506 531664 64706 531720
rect 59445 531662 64706 531664
rect 59445 531659 59511 531662
rect 64646 531172 64706 531662
rect 676029 531654 676095 531657
rect 676029 531652 676292 531654
rect 676029 531596 676034 531652
rect 676090 531596 676292 531652
rect 676029 531594 676292 531596
rect 676029 531591 676095 531594
rect 676213 531450 676279 531453
rect 676213 531448 676322 531450
rect 676213 531392 676218 531448
rect 676274 531392 676322 531448
rect 676213 531387 676322 531392
rect 676262 531216 676322 531387
rect 679249 531042 679315 531045
rect 679206 531040 679315 531042
rect 679206 530984 679254 531040
rect 679310 530984 679315 531040
rect 679206 530979 679315 530984
rect 679206 530808 679266 530979
rect 42926 530708 42932 530772
rect 42996 530770 43002 530772
rect 43161 530770 43227 530773
rect 42996 530768 43227 530770
rect 42996 530712 43166 530768
rect 43222 530712 43227 530768
rect 42996 530710 43227 530712
rect 42996 530708 43002 530710
rect 43161 530707 43227 530710
rect 59261 530634 59327 530637
rect 679065 530634 679131 530637
rect 59261 530632 64706 530634
rect 59261 530576 59266 530632
rect 59322 530576 64706 530632
rect 59261 530574 64706 530576
rect 59261 530571 59327 530574
rect 42006 530164 42012 530228
rect 42076 530226 42082 530228
rect 42333 530226 42399 530229
rect 42076 530224 42399 530226
rect 42076 530168 42338 530224
rect 42394 530168 42399 530224
rect 42076 530166 42399 530168
rect 42076 530164 42082 530166
rect 42333 530163 42399 530166
rect 64646 529990 64706 530574
rect 679022 530632 679131 530634
rect 679022 530576 679070 530632
rect 679126 530576 679131 530632
rect 679022 530571 679131 530576
rect 679022 530400 679082 530571
rect 678973 530226 679039 530229
rect 678973 530224 679082 530226
rect 678973 530168 678978 530224
rect 679034 530168 679082 530224
rect 678973 530163 679082 530168
rect 679022 529992 679082 530163
rect 679433 529818 679499 529821
rect 679390 529816 679499 529818
rect 679390 529760 679438 529816
rect 679494 529760 679499 529816
rect 679390 529755 679499 529760
rect 679390 529584 679450 529755
rect 58525 529410 58591 529413
rect 679341 529410 679407 529413
rect 58525 529408 64706 529410
rect 58525 529352 58530 529408
rect 58586 529352 64706 529408
rect 58525 529350 64706 529352
rect 58525 529347 58591 529350
rect 64646 528808 64706 529350
rect 679341 529408 679450 529410
rect 679341 529352 679346 529408
rect 679402 529352 679450 529408
rect 679341 529347 679450 529352
rect 679390 529176 679450 529347
rect 679157 529002 679223 529005
rect 679157 529000 679266 529002
rect 679157 528944 679162 529000
rect 679218 528944 679266 529000
rect 679157 528939 679266 528944
rect 679206 528768 679266 528939
rect 675753 528390 675819 528393
rect 675753 528388 676292 528390
rect 675753 528332 675758 528388
rect 675814 528332 676292 528388
rect 675753 528330 676292 528332
rect 675753 528327 675819 528330
rect 58341 528186 58407 528189
rect 58341 528184 64706 528186
rect 58341 528128 58346 528184
rect 58402 528128 64706 528184
rect 58341 528126 64706 528128
rect 58341 528123 58407 528126
rect 64646 527626 64706 528126
rect 676029 527982 676095 527985
rect 676029 527980 676292 527982
rect 676029 527924 676034 527980
rect 676090 527924 676292 527980
rect 676029 527922 676292 527924
rect 676029 527919 676095 527922
rect 677593 527778 677659 527781
rect 677550 527776 677659 527778
rect 677550 527720 677598 527776
rect 677654 527720 677659 527776
rect 677550 527715 677659 527720
rect 677550 527544 677610 527715
rect 677501 527370 677567 527373
rect 677501 527368 677610 527370
rect 677501 527312 677506 527368
rect 677562 527312 677610 527368
rect 677501 527307 677610 527312
rect 677550 527136 677610 527307
rect 60641 527098 60707 527101
rect 60641 527096 64706 527098
rect 60641 527040 60646 527096
rect 60702 527040 64706 527096
rect 60641 527038 64706 527040
rect 60641 527035 60707 527038
rect 64646 526444 64706 527038
rect 676990 526900 676996 526964
rect 677060 526900 677066 526964
rect 676998 526728 677058 526900
rect 676029 526350 676095 526353
rect 676029 526348 676292 526350
rect 676029 526292 676034 526348
rect 676090 526292 676292 526348
rect 676029 526290 676292 526292
rect 676029 526287 676095 526290
rect 59353 525874 59419 525877
rect 59353 525872 64706 525874
rect 59353 525816 59358 525872
rect 59414 525816 64706 525872
rect 59353 525814 64706 525816
rect 59353 525811 59419 525814
rect 64646 525262 64706 525814
rect 679022 525741 679082 525912
rect 678973 525736 679082 525741
rect 678973 525680 678978 525736
rect 679034 525680 679082 525736
rect 678973 525678 679082 525680
rect 678973 525675 679039 525678
rect 684542 525096 684602 525504
rect 678973 524922 679039 524925
rect 678973 524920 679082 524922
rect 678973 524864 678978 524920
rect 679034 524864 679082 524920
rect 678973 524859 679082 524864
rect 679022 524688 679082 524859
rect 649308 518701 650108 518748
rect 649308 513948 667116 518701
rect 650058 513921 667116 513948
rect 649308 508722 650108 508748
rect 649308 503948 667124 508722
rect 650066 503942 667124 503948
tri 63960 497858 64508 498406 se
rect 64508 497858 65308 498406
rect 52228 493606 65308 497858
rect 52228 493078 64012 493606
tri 64012 493078 64540 493606 nw
rect 675937 492146 676003 492149
rect 675937 492144 676292 492146
rect 675937 492088 675942 492144
rect 675998 492088 676292 492144
rect 675937 492086 676292 492088
rect 675937 492083 676003 492086
rect 676029 491738 676095 491741
rect 676029 491736 676292 491738
rect 676029 491680 676034 491736
rect 676090 491680 676292 491736
rect 676029 491678 676292 491680
rect 676029 491675 676095 491678
rect 675753 491602 675819 491605
rect 675753 491600 675954 491602
rect 675753 491544 675758 491600
rect 675814 491544 675954 491600
rect 675753 491542 675954 491544
rect 675753 491539 675819 491542
rect 674046 491404 674052 491468
rect 674116 491466 674122 491468
rect 675753 491466 675819 491469
rect 674116 491464 675819 491466
rect 674116 491408 675758 491464
rect 675814 491408 675819 491464
rect 674116 491406 675819 491408
rect 674116 491404 674122 491406
rect 675753 491403 675819 491406
rect 674230 491268 674236 491332
rect 674300 491330 674306 491332
rect 675661 491330 675727 491333
rect 674300 491328 675727 491330
rect 674300 491272 675666 491328
rect 675722 491272 675727 491328
rect 674300 491270 675727 491272
rect 674300 491268 674306 491270
rect 675661 491267 675727 491270
rect 675894 490922 675954 491542
rect 676029 491330 676095 491333
rect 676029 491328 676292 491330
rect 676029 491272 676034 491328
rect 676090 491272 676292 491328
rect 676029 491270 676292 491272
rect 676029 491267 676095 491270
rect 675894 490862 676292 490922
rect 679433 490514 679499 490517
rect 679420 490512 679499 490514
rect 679420 490456 679438 490512
rect 679494 490456 679499 490512
rect 679420 490454 679499 490456
rect 679433 490451 679499 490454
rect 676029 490106 676095 490109
rect 676029 490104 676292 490106
rect 676029 490048 676034 490104
rect 676090 490048 676292 490104
rect 676029 490046 676292 490048
rect 676029 490043 676095 490046
rect 676029 489698 676095 489701
rect 676029 489696 676292 489698
rect 676029 489640 676034 489696
rect 676090 489640 676292 489696
rect 676029 489638 676292 489640
rect 676029 489635 676095 489638
rect 675385 489290 675451 489293
rect 675385 489288 676292 489290
rect 675385 489232 675390 489288
rect 675446 489232 676292 489288
rect 675385 489230 676292 489232
rect 675385 489227 675451 489230
rect 679617 488882 679683 488885
rect 679604 488880 679683 488882
rect 679604 488824 679622 488880
rect 679678 488824 679683 488880
rect 679604 488822 679683 488824
rect 679617 488819 679683 488822
rect 675937 488474 676003 488477
rect 675937 488472 676292 488474
rect 675937 488416 675942 488472
rect 675998 488416 676292 488472
rect 675937 488414 676292 488416
rect 675937 488411 676003 488414
tri 63982 487879 64508 488405 se
rect 64508 487879 65308 488406
rect 679157 488066 679223 488069
rect 679157 488064 679236 488066
rect 679157 488008 679162 488064
rect 679218 488008 679236 488064
rect 679157 488006 679236 488008
rect 679157 488003 679223 488006
rect 52236 483606 65308 487879
rect 675661 487658 675727 487661
rect 675661 487656 676292 487658
rect 675661 487600 675666 487656
rect 675722 487600 676292 487656
rect 675661 487598 676292 487600
rect 675661 487595 675727 487598
rect 675477 487250 675543 487253
rect 675477 487248 676292 487250
rect 675477 487192 675482 487248
rect 675538 487192 676292 487248
rect 675477 487190 676292 487192
rect 675477 487187 675543 487190
rect 675753 486842 675819 486845
rect 675753 486840 676292 486842
rect 675753 486784 675758 486840
rect 675814 486784 676292 486840
rect 675753 486782 676292 486784
rect 675753 486779 675819 486782
rect 675845 486434 675911 486437
rect 675845 486432 676292 486434
rect 675845 486376 675850 486432
rect 675906 486376 676292 486432
rect 675845 486374 676292 486376
rect 675845 486371 675911 486374
rect 675109 486026 675175 486029
rect 675109 486024 676292 486026
rect 675109 485968 675114 486024
rect 675170 485968 676292 486024
rect 675109 485966 676292 485968
rect 675109 485963 675175 485966
rect 676029 485618 676095 485621
rect 676029 485616 676292 485618
rect 676029 485560 676034 485616
rect 676090 485560 676292 485616
rect 676029 485558 676292 485560
rect 676029 485555 676095 485558
rect 675150 485148 675156 485212
rect 675220 485210 675226 485212
rect 675220 485150 676292 485210
rect 675220 485148 675226 485150
rect 675569 484802 675635 484805
rect 675569 484800 676292 484802
rect 675569 484744 675574 484800
rect 675630 484744 676292 484800
rect 675569 484742 676292 484744
rect 675569 484739 675635 484742
rect 675845 484394 675911 484397
rect 675845 484392 676292 484394
rect 675845 484336 675850 484392
rect 675906 484336 676292 484392
rect 675845 484334 676292 484336
rect 675845 484331 675911 484334
rect 675937 483986 676003 483989
rect 675937 483984 676292 483986
rect 675937 483928 675942 483984
rect 675998 483928 676292 483984
rect 675937 483926 676292 483928
rect 675937 483923 676003 483926
rect 52236 483099 64041 483606
tri 64041 483099 64548 483606 nw
rect 676029 483578 676095 483581
rect 676029 483576 676292 483578
rect 676029 483520 676034 483576
rect 676090 483520 676292 483576
rect 676029 483518 676292 483520
rect 676029 483515 676095 483518
rect 676029 483170 676095 483173
rect 676029 483168 676292 483170
rect 676029 483112 676034 483168
rect 676090 483112 676292 483168
rect 676029 483110 676292 483112
rect 676029 483107 676095 483110
rect 675937 482762 676003 482765
rect 675937 482760 676292 482762
rect 675937 482704 675942 482760
rect 675998 482704 676292 482760
rect 675937 482702 676292 482704
rect 675937 482699 676003 482702
rect 676029 482354 676095 482357
rect 676029 482352 676292 482354
rect 676029 482296 676034 482352
rect 676090 482296 676292 482352
rect 676029 482294 676292 482296
rect 676029 482291 676095 482294
rect 676029 481946 676095 481949
rect 676029 481944 676292 481946
rect 676029 481888 676034 481944
rect 676090 481888 676292 481944
rect 676029 481886 676292 481888
rect 676029 481883 676095 481886
rect 684542 481100 684602 481508
rect 676029 480722 676095 480725
rect 676029 480720 676292 480722
rect 676029 480664 676034 480720
rect 676090 480664 676292 480720
rect 676029 480662 676292 480664
rect 676029 480659 676095 480662
rect 649308 474700 650108 474948
rect 649308 470148 670778 474700
rect 650042 469900 670778 470148
rect 649308 464649 650108 464948
rect 649308 460148 670778 464649
rect 650042 459860 670778 460148
rect 42425 455970 42491 455973
rect 42558 455970 42564 455972
rect 42425 455968 42564 455970
rect 42425 455912 42430 455968
rect 42486 455912 42564 455968
rect 42425 455910 42564 455912
rect 42425 455907 42491 455910
rect 42558 455908 42564 455910
rect 42628 455908 42634 455972
tri 63842 455740 64508 456406 se
rect 64508 455740 65308 456406
rect 46742 451606 65308 455740
rect 46742 450951 63927 451606
tri 63927 450951 64582 451606 nw
rect 42425 450804 42491 450805
rect 42374 450802 42380 450804
rect 42334 450742 42380 450802
rect 42444 450800 42491 450804
rect 42486 450744 42491 450800
rect 42374 450740 42380 450742
rect 42444 450740 42491 450744
rect 42425 450739 42491 450740
rect 42425 445908 42491 445909
rect 42374 445844 42380 445908
rect 42444 445906 42491 445908
rect 42444 445904 42536 445906
rect 42486 445848 42536 445904
rect 42444 445846 42536 445848
rect 42444 445844 42491 445846
rect 42425 445843 42491 445844
tri 63802 445700 64508 446406 se
rect 64508 445700 65308 446406
rect 46768 441606 65308 445700
rect 46768 440900 63858 441606
tri 63858 440900 64564 441606 nw
rect 42425 440740 42491 440741
rect 42374 440738 42380 440740
rect 42334 440678 42380 440738
rect 42444 440736 42491 440740
rect 42486 440680 42491 440736
rect 42374 440676 42380 440678
rect 42444 440676 42491 440680
rect 42425 440675 42491 440676
rect 41781 430946 41847 430949
rect 41492 430944 41847 430946
rect 41492 430888 41786 430944
rect 41842 430888 41847 430944
rect 41492 430886 41847 430888
rect 41781 430883 41847 430886
rect 41781 430538 41847 430541
rect 41492 430536 41847 430538
rect 41492 430480 41786 430536
rect 41842 430480 41847 430536
rect 41492 430478 41847 430480
rect 41781 430475 41847 430478
rect 650068 430348 663976 430501
rect 42057 430130 42123 430133
rect 41492 430128 42123 430130
rect 41492 430072 42062 430128
rect 42118 430072 42123 430128
rect 41492 430070 42123 430072
rect 42057 430067 42123 430070
rect 44589 429714 44659 429719
rect 41590 429654 44594 429714
rect 44654 429654 44668 429714
rect 44589 429649 44659 429654
rect 44589 429332 44659 429335
rect 41590 429330 44668 429332
rect 41590 429272 44594 429330
rect 44589 429270 44594 429272
rect 44654 429272 44668 429330
rect 44654 429270 44659 429272
rect 44589 429265 44659 429270
rect 42374 428906 42380 428908
rect 41492 428846 42380 428906
rect 42374 428844 42380 428846
rect 42444 428844 42450 428908
rect 43713 428498 43779 428501
rect 41492 428496 43779 428498
rect 41492 428440 43718 428496
rect 43774 428440 43779 428496
rect 41492 428438 43779 428440
rect 43713 428435 43779 428438
rect 42049 428314 42115 428317
rect 42049 428312 45102 428314
rect 42049 428256 42054 428312
rect 42110 428256 45102 428312
rect 42049 428254 45102 428256
rect 42049 428251 42115 428254
rect 30097 428090 30163 428093
rect 30084 428088 30163 428090
rect 30084 428032 30102 428088
rect 30158 428032 30163 428088
rect 44680 428090 44752 428096
rect 45042 428090 45102 428254
rect 59261 428090 59327 428093
rect 44680 428084 44758 428090
rect 44680 428080 44686 428084
rect 30084 428030 30163 428032
rect 30097 428027 30163 428030
rect 41560 428024 44686 428080
rect 44746 428024 44758 428084
rect 45042 428088 59327 428090
rect 45042 428032 59266 428088
rect 59322 428032 59327 428088
rect 45042 428030 59327 428032
rect 59261 428027 59327 428030
rect 41560 428020 44758 428024
rect 44681 428019 44751 428020
rect 59445 427954 59511 427957
rect 45046 427952 59511 427954
rect 45046 427896 59450 427952
rect 59506 427896 59511 427952
rect 45046 427894 59511 427896
rect 41781 427874 41847 427877
rect 45046 427874 45106 427894
rect 59445 427891 59511 427894
rect 41781 427872 45106 427874
rect 41781 427816 41786 427872
rect 41842 427816 45106 427872
rect 41781 427814 45106 427816
rect 41781 427811 41847 427814
rect 30005 427682 30071 427685
rect 30005 427680 30084 427682
rect 30005 427624 30010 427680
rect 30066 427624 30084 427680
rect 44681 427668 44751 427673
rect 44681 427666 44686 427668
rect 30005 427622 30084 427624
rect 30005 427619 30071 427622
rect 41560 427608 44686 427666
rect 44746 427666 44751 427668
rect 44746 427608 44758 427666
rect 41560 427606 44758 427608
rect 44681 427603 44751 427606
rect 44773 427288 44843 427293
rect 41560 427228 44778 427288
rect 44838 427228 44864 427288
rect 44773 427223 44843 427228
rect 44773 426876 44843 426881
rect 44773 426870 44778 426876
rect 41560 426816 44778 426870
rect 44838 426870 44843 426876
rect 44838 426816 44864 426870
rect 41560 426810 44864 426816
rect 43437 426458 43503 426461
rect 41492 426456 43503 426458
rect 41492 426400 43442 426456
rect 43498 426400 43503 426456
rect 41492 426398 43503 426400
rect 43437 426395 43503 426398
rect 42333 426050 42399 426053
rect 41492 426048 42399 426050
rect 41492 425992 42338 426048
rect 42394 425992 42399 426048
rect 41492 425990 42399 425992
rect 42333 425987 42399 425990
rect 42701 425642 42767 425645
rect 41492 425640 42767 425642
rect 41492 425584 42706 425640
rect 42762 425584 42767 425640
rect 41492 425582 42767 425584
rect 42701 425579 42767 425582
rect 649308 425562 663976 430348
rect 649308 425548 650108 425562
rect 43529 425234 43595 425237
rect 41492 425232 43595 425234
rect 41492 425176 43534 425232
rect 43590 425176 43595 425232
rect 41492 425174 43595 425176
rect 43529 425171 43595 425174
rect 43621 424826 43687 424829
rect 41492 424824 43687 424826
rect 41492 424768 43626 424824
rect 43682 424768 43687 424824
rect 41492 424766 43687 424768
rect 43621 424763 43687 424766
rect 42241 424418 42307 424421
rect 41492 424416 42307 424418
rect 41492 424360 42246 424416
rect 42302 424360 42307 424416
rect 41492 424358 42307 424360
rect 42241 424355 42307 424358
rect 43897 424010 43963 424013
rect 41492 424008 43963 424010
rect 41492 423952 43902 424008
rect 43958 423952 43963 424008
rect 41492 423950 43963 423952
rect 43897 423947 43963 423950
rect 43805 423602 43871 423605
rect 41492 423600 43871 423602
rect 41492 423544 43810 423600
rect 43866 423544 43871 423600
rect 41492 423542 43871 423544
rect 43805 423539 43871 423542
rect 43989 423194 44055 423197
rect 41492 423192 44055 423194
rect 41492 423136 43994 423192
rect 44050 423136 44055 423192
rect 41492 423134 44055 423136
rect 43989 423131 44055 423134
rect 41873 422786 41939 422789
rect 41492 422784 41939 422786
rect 41492 422728 41878 422784
rect 41934 422728 41939 422784
rect 41492 422726 41939 422728
rect 41873 422723 41939 422726
rect 41965 422378 42031 422381
rect 41492 422376 42031 422378
rect 41492 422320 41970 422376
rect 42026 422320 42031 422376
rect 41492 422318 42031 422320
rect 41965 422315 42031 422318
rect 44081 421970 44147 421973
rect 41492 421968 44147 421970
rect 41492 421912 44086 421968
rect 44142 421912 44147 421968
rect 41492 421910 44147 421912
rect 44081 421907 44147 421910
rect 43345 421562 43411 421565
rect 41492 421560 43411 421562
rect 41492 421504 43350 421560
rect 43406 421504 43411 421560
rect 41492 421502 43411 421504
rect 43345 421499 43411 421502
rect 43253 421154 43319 421157
rect 41492 421152 43319 421154
rect 41492 421096 43258 421152
rect 43314 421096 43319 421152
rect 41492 421094 43319 421096
rect 43253 421091 43319 421094
rect 41781 420746 41847 420749
rect 41492 420744 41847 420746
rect 41492 420688 41786 420744
rect 41842 420688 41847 420744
rect 41492 420686 41847 420688
rect 41781 420683 41847 420686
rect 650058 420348 663966 420522
rect 30422 419900 30482 420308
rect 41781 419522 41847 419525
rect 41492 419520 41847 419522
rect 41492 419464 41786 419520
rect 41842 419464 41847 419520
rect 41492 419462 41847 419464
rect 41781 419459 41847 419462
rect 649308 415742 663966 420348
rect 649308 415548 650108 415742
rect 58157 404154 58223 404157
rect 58157 404152 64706 404154
rect 58157 404096 58162 404152
rect 58218 404096 64706 404152
rect 58157 404094 64706 404096
rect 58157 404091 58223 404094
rect 64646 403550 64706 404094
rect 676262 403749 676322 403852
rect 676262 403744 676371 403749
rect 676262 403688 676310 403744
rect 676366 403688 676371 403744
rect 676262 403686 676371 403688
rect 676305 403683 676371 403686
rect 676262 403341 676322 403444
rect 676213 403336 676322 403341
rect 676213 403280 676218 403336
rect 676274 403280 676322 403336
rect 676213 403278 676322 403280
rect 676213 403275 676279 403278
rect 675845 403066 675911 403069
rect 675845 403064 676292 403066
rect 675845 403008 675850 403064
rect 675906 403008 676292 403064
rect 675845 403006 676292 403008
rect 675845 403003 675911 403006
rect 58157 402930 58223 402933
rect 58157 402928 64706 402930
rect 58157 402872 58162 402928
rect 58218 402872 64706 402928
rect 58157 402870 64706 402872
rect 58157 402867 58223 402870
rect 64646 402368 64706 402870
rect 675937 402658 676003 402661
rect 675926 402656 676292 402658
rect 675926 402600 675942 402656
rect 675998 402600 676292 402656
rect 675926 402598 676292 402600
rect 675937 402595 676003 402598
rect 675150 402188 675156 402252
rect 675220 402250 675226 402252
rect 675220 402190 676292 402250
rect 675220 402188 675226 402190
rect 677481 402114 677547 402117
rect 677481 402112 677590 402114
rect 677481 402056 677486 402112
rect 677542 402056 677590 402112
rect 677481 402051 677590 402056
rect 677530 401812 677590 402051
rect 675293 401434 675359 401437
rect 675293 401432 676292 401434
rect 675293 401376 675298 401432
rect 675354 401376 676292 401432
rect 675293 401374 676292 401376
rect 675293 401371 675359 401374
rect 58893 400754 58959 400757
rect 64646 400754 64706 401186
rect 676029 401026 676095 401029
rect 676029 401024 676292 401026
rect 676029 400968 676034 401024
rect 676090 400968 676292 401024
rect 676029 400966 676292 400968
rect 676029 400963 676095 400966
rect 58893 400752 64706 400754
rect 58893 400696 58898 400752
rect 58954 400696 64706 400752
rect 58893 400694 64706 400696
rect 58893 400691 58959 400694
rect 674966 400556 674972 400620
rect 675036 400618 675042 400620
rect 675036 400558 676292 400618
rect 675036 400556 675042 400558
rect 676029 400210 676095 400213
rect 676006 400208 676292 400210
rect 676006 400152 676034 400208
rect 676090 400152 676292 400208
rect 676006 400150 676292 400152
rect 676029 400147 676095 400150
rect 59261 400074 59327 400077
rect 59261 400072 64706 400074
rect 59261 400016 59266 400072
rect 59322 400016 64706 400072
rect 59261 400014 64706 400016
rect 59261 400011 59327 400014
rect 64646 400004 64706 400014
rect 674782 399740 674788 399804
rect 674852 399802 674858 399804
rect 674852 399742 676292 399802
rect 674852 399740 674858 399742
rect 58157 399394 58223 399397
rect 676029 399394 676095 399397
rect 58157 399392 64706 399394
rect 58157 399336 58162 399392
rect 58218 399336 64706 399392
rect 58157 399334 64706 399336
rect 58157 399331 58223 399334
rect 64646 398822 64706 399334
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 676121 398850 676187 398853
rect 676262 398850 676322 398956
rect 676121 398848 676322 398850
rect 676121 398792 676126 398848
rect 676182 398792 676322 398848
rect 676121 398790 676322 398792
rect 676121 398787 676187 398790
rect 675753 398578 675819 398581
rect 675753 398576 676292 398578
rect 675753 398520 675758 398576
rect 675814 398520 676292 398576
rect 675753 398518 676292 398520
rect 675753 398515 675819 398518
rect 59445 398306 59511 398309
rect 59445 398304 64706 398306
rect 59445 398248 59450 398304
rect 59506 398248 64706 398304
rect 59445 398246 64706 398248
rect 59445 398243 59511 398246
rect 64646 397640 64706 398246
rect 676029 398170 676095 398173
rect 676029 398168 676292 398170
rect 676029 398112 676034 398168
rect 676090 398112 676292 398168
rect 676029 398110 676292 398112
rect 676029 398107 676095 398110
rect 675937 397762 676003 397765
rect 675937 397760 676292 397762
rect 675937 397704 675942 397760
rect 675998 397704 676292 397760
rect 675937 397702 676292 397704
rect 675937 397699 676003 397702
rect 676029 397354 676095 397357
rect 676029 397352 676292 397354
rect 676029 397296 676034 397352
rect 676090 397296 676292 397352
rect 676029 397294 676292 397296
rect 676029 397291 676095 397294
rect 676029 396946 676095 396949
rect 676029 396944 676292 396946
rect 676029 396888 676034 396944
rect 676090 396888 676292 396944
rect 676029 396886 676292 396888
rect 676029 396883 676095 396886
rect 676121 396402 676187 396405
rect 676262 396402 676322 396508
rect 676121 396400 676322 396402
rect 676121 396344 676126 396400
rect 676182 396344 676322 396400
rect 676121 396342 676322 396344
rect 676121 396339 676187 396342
rect 675937 396130 676003 396133
rect 675937 396128 676292 396130
rect 675937 396072 675942 396128
rect 675998 396072 676292 396128
rect 675937 396070 676292 396072
rect 675937 396067 676003 396070
rect 675845 395722 675911 395725
rect 675845 395720 676292 395722
rect 675845 395664 675850 395720
rect 675906 395664 676292 395720
rect 675845 395662 676292 395664
rect 675845 395659 675911 395662
rect 675845 395314 675911 395317
rect 675845 395312 676292 395314
rect 675845 395256 675850 395312
rect 675906 395256 676292 395312
rect 675845 395254 676292 395256
rect 675845 395251 675911 395254
rect 675937 394906 676003 394909
rect 675937 394904 676292 394906
rect 675937 394848 675942 394904
rect 675998 394848 676292 394904
rect 675937 394846 676292 394848
rect 675937 394843 676003 394846
rect 676029 394498 676095 394501
rect 676029 394496 676292 394498
rect 676029 394440 676034 394496
rect 676090 394440 676292 394496
rect 676029 394438 676292 394440
rect 676029 394435 676095 394438
rect 676029 394090 676095 394093
rect 676029 394088 676292 394090
rect 676029 394032 676034 394088
rect 676090 394032 676292 394088
rect 676029 394030 676292 394032
rect 676029 394027 676095 394030
rect 679022 393549 679082 393652
rect 678973 393544 679082 393549
rect 678973 393488 678978 393544
rect 679034 393488 679082 393544
rect 678973 393486 679082 393488
rect 678973 393483 679039 393486
rect 684542 392836 684602 393244
rect 678973 392730 679039 392733
rect 678973 392728 679082 392730
rect 678973 392672 678978 392728
rect 679034 392672 679082 392728
rect 678973 392667 679082 392672
rect 679022 392428 679082 392667
rect 41781 387698 41847 387701
rect 41492 387696 41847 387698
rect 41492 387640 41786 387696
rect 41842 387640 41847 387696
rect 41492 387638 41847 387640
rect 41781 387635 41847 387638
rect 41505 387562 41571 387565
rect 41462 387560 41571 387562
rect 41462 387504 41510 387560
rect 41566 387504 41571 387560
rect 41462 387499 41571 387504
rect 41462 387260 41522 387499
rect 41462 386749 41522 386852
rect 41462 386744 41571 386749
rect 41462 386688 41510 386744
rect 41566 386688 41571 386744
rect 41462 386686 41571 386688
rect 41505 386683 41571 386686
rect 44589 386514 44659 386519
rect 41560 386454 44594 386514
rect 44654 386454 44668 386514
rect 44589 386449 44659 386454
rect 44589 386132 44659 386135
rect 41560 386130 44668 386132
rect 41560 386072 44594 386130
rect 44589 386070 44594 386072
rect 44654 386072 44668 386130
rect 44654 386070 44659 386072
rect 44589 386065 44659 386070
rect 43713 385658 43779 385661
rect 41492 385656 43779 385658
rect 41492 385600 43718 385656
rect 43774 385600 43779 385656
rect 41492 385598 43779 385600
rect 43713 385595 43779 385598
rect 43529 385250 43595 385253
rect 41492 385248 43595 385250
rect 41492 385192 43534 385248
rect 43590 385192 43595 385248
rect 41492 385190 43595 385192
rect 43529 385187 43595 385190
rect 44681 384880 44751 384883
rect 41548 384878 44758 384880
rect 41548 384820 44686 384878
rect 44681 384818 44686 384820
rect 44746 384820 44758 384878
rect 44746 384818 44751 384820
rect 44681 384813 44751 384818
rect 44681 384468 44751 384473
rect 44681 384466 44686 384468
rect 41548 384408 44686 384466
rect 44746 384466 44751 384468
rect 44746 384408 44758 384466
rect 41548 384406 44758 384408
rect 44681 384403 44751 384406
rect 44773 384088 44843 384093
rect 41548 384028 44778 384088
rect 44838 384028 44864 384088
rect 44773 384023 44843 384028
rect 44773 383676 44843 383681
rect 44773 383670 44778 383676
rect 41548 383616 44778 383670
rect 44838 383670 44843 383676
rect 44838 383616 44864 383670
rect 41548 383610 44864 383616
rect 43437 383210 43503 383213
rect 41492 383208 43503 383210
rect 41492 383152 43442 383208
rect 43498 383152 43503 383208
rect 41492 383150 43503 383152
rect 43437 383147 43503 383150
rect 42701 382802 42767 382805
rect 41492 382800 42767 382802
rect 41492 382744 42706 382800
rect 42762 382744 42767 382800
rect 41492 382742 42767 382744
rect 42701 382739 42767 382742
rect 43713 382394 43779 382397
rect 41492 382392 43779 382394
rect 41492 382336 43718 382392
rect 43774 382336 43779 382392
rect 41492 382334 43779 382336
rect 43713 382331 43779 382334
rect 43069 381986 43135 381989
rect 41492 381984 43135 381986
rect 41492 381928 43074 381984
rect 43130 381928 43135 381984
rect 41492 381926 43135 381928
rect 43069 381923 43135 381926
rect 43253 381578 43319 381581
rect 41492 381576 43319 381578
rect 41492 381520 43258 381576
rect 43314 381520 43319 381576
rect 41492 381518 43319 381520
rect 43253 381515 43319 381518
rect 38150 381037 38210 381140
rect 38150 381032 38259 381037
rect 38150 380976 38198 381032
rect 38254 380976 38259 381032
rect 38150 380974 38259 380976
rect 38193 380971 38259 380974
rect 43713 380762 43779 380765
rect 41492 380760 43779 380762
rect 41492 380704 43718 380760
rect 43774 380704 43779 380760
rect 41492 380702 43779 380704
rect 43713 380699 43779 380702
rect 43897 380354 43963 380357
rect 41492 380352 43963 380354
rect 41492 380296 43902 380352
rect 43958 380296 43963 380352
rect 41492 380294 43963 380296
rect 43897 380291 43963 380294
rect 41965 379946 42031 379949
rect 41492 379944 42031 379946
rect 41492 379888 41970 379944
rect 42026 379888 42031 379944
rect 41492 379886 42031 379888
rect 41965 379883 42031 379886
rect 43161 379538 43227 379541
rect 41492 379536 43227 379538
rect 41492 379480 43166 379536
rect 43222 379480 43227 379536
rect 41492 379478 43227 379480
rect 43161 379475 43227 379478
rect 43437 379130 43503 379133
rect 41492 379128 43503 379130
rect 41492 379072 43442 379128
rect 43498 379072 43503 379128
rect 41492 379070 43503 379072
rect 43437 379067 43503 379070
rect 41462 378586 41522 378692
rect 41597 378586 41663 378589
rect 41462 378584 41663 378586
rect 41462 378528 41602 378584
rect 41658 378528 41663 378584
rect 41462 378526 41663 378528
rect 41597 378523 41663 378526
rect 41462 378181 41522 378284
rect 41413 378176 41522 378181
rect 41413 378120 41418 378176
rect 41474 378120 41522 378176
rect 41413 378118 41522 378120
rect 41413 378115 41479 378118
rect 41462 377773 41522 377876
rect 41462 377768 41571 377773
rect 41462 377712 41510 377768
rect 41566 377712 41571 377768
rect 41462 377710 41571 377712
rect 41505 377707 41571 377710
rect 41781 377498 41847 377501
rect 41492 377496 41847 377498
rect 41492 377440 41786 377496
rect 41842 377440 41847 377496
rect 41492 377438 41847 377440
rect 41781 377435 41847 377438
rect 30422 376652 30482 377060
rect 41781 376274 41847 376277
rect 41492 376272 41847 376274
rect 41492 376216 41786 376272
rect 41842 376216 41847 376272
rect 41492 376214 41847 376216
rect 41781 376211 41847 376214
rect 655697 374506 655763 374509
rect 649950 374504 655763 374506
rect 649950 374448 655702 374504
rect 655758 374448 655763 374504
rect 649950 374446 655763 374448
rect 649950 373892 650010 374446
rect 655697 374443 655763 374446
rect 655513 373282 655579 373285
rect 649950 373280 655579 373282
rect 649950 373224 655518 373280
rect 655574 373224 655579 373280
rect 649950 373222 655579 373224
rect 649950 372710 650010 373222
rect 655513 373219 655579 373222
rect 655421 372194 655487 372197
rect 649950 372192 655487 372194
rect 649950 372136 655426 372192
rect 655482 372136 655487 372192
rect 649950 372134 655487 372136
rect 649950 371528 650010 372134
rect 655421 372131 655487 372134
rect 654501 370970 654567 370973
rect 649950 370968 654567 370970
rect 649950 370912 654506 370968
rect 654562 370912 654567 370968
rect 649950 370910 654567 370912
rect 649950 370346 650010 370910
rect 654501 370907 654567 370910
rect 58157 360906 58223 360909
rect 58157 360904 64706 360906
rect 58157 360848 58162 360904
rect 58218 360848 64706 360904
rect 58157 360846 64706 360848
rect 58157 360843 58223 360846
rect 64646 360328 64706 360846
rect 58341 359818 58407 359821
rect 58341 359816 64706 359818
rect 58341 359760 58346 359816
rect 58402 359760 64706 359816
rect 58341 359758 64706 359760
rect 58341 359755 58407 359758
rect 64646 359146 64706 359758
rect 675845 358730 675911 358733
rect 675845 358728 676292 358730
rect 675845 358672 675850 358728
rect 675906 358672 676292 358728
rect 675845 358670 676292 358672
rect 675845 358667 675911 358670
rect 675937 358322 676003 358325
rect 675937 358320 676292 358322
rect 675937 358264 675942 358320
rect 675998 358264 676292 358320
rect 675937 358262 676292 358264
rect 675937 358259 676003 358262
rect 58617 357506 58683 357509
rect 64646 357506 64706 357964
rect 676029 357914 676095 357917
rect 676029 357912 676292 357914
rect 676029 357856 676034 357912
rect 676090 357856 676292 357912
rect 676029 357854 676292 357856
rect 676029 357851 676095 357854
rect 675150 357506 675156 357508
rect 58617 357504 64706 357506
rect 58617 357448 58622 357504
rect 58678 357448 64706 357504
rect 58617 357446 64706 357448
rect 675140 357446 675156 357506
rect 58617 357443 58683 357446
rect 675150 357444 675156 357446
rect 675220 357506 675226 357508
rect 675220 357446 676292 357506
rect 675220 357444 675226 357446
rect 58525 357370 58591 357373
rect 58525 357368 64706 357370
rect 58525 357312 58530 357368
rect 58586 357312 64706 357368
rect 58525 357310 64706 357312
rect 58525 357307 58591 357310
rect 64646 356782 64706 357310
rect 675661 357098 675727 357101
rect 675661 357096 676292 357098
rect 675661 357040 675666 357096
rect 675722 357040 676292 357096
rect 675661 357038 676292 357040
rect 675661 357035 675727 357038
rect 675753 356690 675819 356693
rect 675753 356688 676292 356690
rect 675753 356632 675758 356688
rect 675814 356632 676292 356688
rect 675753 356630 676292 356632
rect 675753 356627 675819 356630
rect 676029 356282 676095 356285
rect 676029 356280 676292 356282
rect 676029 356224 676034 356280
rect 676090 356224 676292 356280
rect 676029 356222 676292 356224
rect 676029 356219 676095 356222
rect 58065 356010 58131 356013
rect 58065 356008 64706 356010
rect 58065 355952 58070 356008
rect 58126 355952 64706 356008
rect 58065 355950 64706 355952
rect 58065 355947 58131 355950
rect 64646 355600 64706 355950
rect 674966 355812 674972 355876
rect 675036 355874 675042 355876
rect 675036 355814 676292 355874
rect 675036 355812 675042 355814
rect 676029 355466 676095 355469
rect 676029 355464 676292 355466
rect 676029 355408 676034 355464
rect 676090 355408 676292 355464
rect 676029 355406 676292 355408
rect 676029 355403 676095 355406
rect 59353 355058 59419 355061
rect 59353 355056 64706 355058
rect 59353 355000 59358 355056
rect 59414 355000 64706 355056
rect 59353 354998 64706 355000
rect 59353 354995 59419 354998
rect 64646 354418 64706 354998
rect 674782 354996 674788 355060
rect 674852 355058 674858 355060
rect 674852 354998 676292 355058
rect 674852 354996 674858 354998
rect 676029 354650 676095 354653
rect 676029 354648 676292 354650
rect 676029 354592 676034 354648
rect 676090 354592 676292 354648
rect 676029 354590 676292 354592
rect 676029 354587 676095 354590
rect 676029 354242 676095 354245
rect 676029 354240 676292 354242
rect 676029 354184 676034 354240
rect 676090 354184 676292 354240
rect 676029 354182 676292 354184
rect 676029 354179 676095 354182
rect 675385 353834 675451 353837
rect 675385 353832 676292 353834
rect 675385 353776 675390 353832
rect 675446 353776 676292 353832
rect 675385 353774 676292 353776
rect 675385 353771 675451 353774
rect 676029 353426 676095 353429
rect 676029 353424 676292 353426
rect 676029 353368 676034 353424
rect 676090 353368 676292 353424
rect 676029 353366 676292 353368
rect 676029 353363 676095 353366
rect 676029 353018 676095 353021
rect 676029 353016 676292 353018
rect 676029 352960 676034 353016
rect 676090 352960 676292 353016
rect 676029 352958 676292 352960
rect 676029 352955 676095 352958
rect 675937 352610 676003 352613
rect 675937 352608 676292 352610
rect 675937 352552 675942 352608
rect 675998 352552 676292 352608
rect 675937 352550 676292 352552
rect 675937 352547 676003 352550
rect 675845 352202 675911 352205
rect 675845 352200 676292 352202
rect 675845 352144 675850 352200
rect 675906 352144 676292 352200
rect 675845 352142 676292 352144
rect 675845 352139 675911 352142
rect 675293 351794 675359 351797
rect 675293 351792 676292 351794
rect 675293 351736 675298 351792
rect 675354 351736 676292 351792
rect 675293 351734 676292 351736
rect 675293 351731 675359 351734
rect 676029 351386 676095 351389
rect 676029 351384 676292 351386
rect 676029 351328 676034 351384
rect 676090 351328 676292 351384
rect 676029 351326 676292 351328
rect 676029 351323 676095 351326
rect 675937 350978 676003 350981
rect 675937 350976 676292 350978
rect 675937 350920 675942 350976
rect 675998 350920 676292 350976
rect 675937 350918 676292 350920
rect 675937 350915 676003 350918
rect 675845 350570 675911 350573
rect 675845 350568 676292 350570
rect 675845 350512 675850 350568
rect 675906 350512 676292 350568
rect 675845 350510 676292 350512
rect 675845 350507 675911 350510
rect 676029 350162 676095 350165
rect 676029 350160 676292 350162
rect 676029 350104 676034 350160
rect 676090 350104 676292 350160
rect 676029 350102 676292 350104
rect 676029 350099 676095 350102
rect 676029 349754 676095 349757
rect 676029 349752 676292 349754
rect 676029 349696 676034 349752
rect 676090 349696 676292 349752
rect 676029 349694 676292 349696
rect 676029 349691 676095 349694
rect 675937 349346 676003 349349
rect 675937 349344 676292 349346
rect 675937 349288 675942 349344
rect 675998 349288 676292 349344
rect 675937 349286 676292 349288
rect 675937 349283 676003 349286
rect 675845 348938 675911 348941
rect 675845 348936 676292 348938
rect 675845 348880 675850 348936
rect 675906 348880 676292 348936
rect 675845 348878 676292 348880
rect 675845 348875 675911 348878
rect 676078 348470 676292 348530
rect 676078 347309 676138 348470
rect 679022 347684 679082 348092
rect 676029 347306 676138 347309
rect 675948 347304 676292 347306
rect 675948 347248 676034 347304
rect 676090 347248 676292 347304
rect 675948 347246 676292 347248
rect 676029 347243 676095 347246
rect 41462 344317 41522 344556
rect 41462 344312 41571 344317
rect 41462 344256 41510 344312
rect 41566 344256 41571 344312
rect 41462 344254 41571 344256
rect 41505 344251 41571 344254
rect 41462 343909 41522 344148
rect 41462 343904 41571 343909
rect 41462 343848 41510 343904
rect 41566 343848 41571 343904
rect 41462 343846 41571 343848
rect 41505 343843 41571 343846
rect 41462 343501 41522 343740
rect 41462 343496 41571 343501
rect 41462 343440 41510 343496
rect 41566 343440 41571 343496
rect 41462 343438 41571 343440
rect 41505 343435 41571 343438
rect 44588 343314 44660 343320
rect 41590 343254 44594 343314
rect 44654 343254 44668 343314
rect 44588 343248 44660 343254
rect 44589 342932 44659 342935
rect 41590 342930 44668 342932
rect 41590 342872 44594 342930
rect 44589 342870 44594 342872
rect 44654 342872 44668 342930
rect 44654 342870 44659 342872
rect 44589 342865 44659 342870
rect 41505 342682 41571 342685
rect 41462 342680 41571 342682
rect 41462 342624 41510 342680
rect 41566 342624 41571 342680
rect 41462 342619 41571 342624
rect 41462 342516 41522 342619
rect 43345 342138 43411 342141
rect 41492 342136 43411 342138
rect 41492 342080 43350 342136
rect 43406 342080 43411 342136
rect 41492 342078 43411 342080
rect 43345 342075 43411 342078
rect 44681 341680 44751 341683
rect 41522 341678 44758 341680
rect 41522 341620 44686 341678
rect 44681 341618 44686 341620
rect 44746 341620 44758 341678
rect 44746 341618 44751 341620
rect 44681 341613 44751 341618
rect 44681 341268 44751 341273
rect 44681 341266 44686 341268
rect 41522 341208 44686 341266
rect 44746 341266 44751 341268
rect 44746 341208 44758 341266
rect 41522 341206 44758 341208
rect 44681 341203 44751 341206
rect 44773 340888 44843 340893
rect 41522 340828 44778 340888
rect 44838 340828 44864 340888
rect 44773 340823 44843 340828
rect 44773 340476 44843 340481
rect 44773 340470 44778 340476
rect 41522 340416 44778 340470
rect 44838 340470 44843 340476
rect 44838 340416 44864 340470
rect 41522 340410 44864 340416
rect 32814 339829 32874 340068
rect 32814 339824 32923 339829
rect 33041 339826 33107 339829
rect 32814 339768 32862 339824
rect 32918 339768 32923 339824
rect 32814 339766 32923 339768
rect 32857 339763 32923 339766
rect 32998 339824 33107 339826
rect 32998 339768 33046 339824
rect 33102 339768 33107 339824
rect 32998 339763 33107 339768
rect 32998 339660 33058 339763
rect 41462 339010 41522 339252
rect 41638 339010 41644 339012
rect 41462 338950 41644 339010
rect 41638 338948 41644 338950
rect 41708 338948 41714 339012
rect 42006 338874 42012 338876
rect 41492 338814 42012 338874
rect 42006 338812 42012 338814
rect 42076 338812 42082 338876
rect 43161 338466 43227 338469
rect 41492 338464 43227 338466
rect 41492 338408 43166 338464
rect 43222 338408 43227 338464
rect 41492 338406 43227 338408
rect 43161 338403 43227 338406
rect 41781 338058 41847 338061
rect 41492 338056 41847 338058
rect 41492 338000 41786 338056
rect 41842 338000 41847 338056
rect 41492 337998 41847 338000
rect 41781 337995 41847 337998
rect 41822 337650 41828 337652
rect 41492 337590 41828 337650
rect 41822 337588 41828 337590
rect 41892 337588 41898 337652
rect 41462 336973 41522 337212
rect 41462 336968 41571 336973
rect 41462 336912 41510 336968
rect 41566 336912 41571 336968
rect 41462 336910 41571 336912
rect 41505 336907 41571 336910
rect 41462 336565 41522 336804
rect 41413 336560 41522 336565
rect 41413 336504 41418 336560
rect 41474 336504 41522 336560
rect 41413 336502 41522 336504
rect 41413 336499 41479 336502
rect 42333 336426 42399 336429
rect 41492 336424 42399 336426
rect 41492 336368 42338 336424
rect 42394 336368 42399 336424
rect 41492 336366 42399 336368
rect 42333 336363 42399 336366
rect 43253 336018 43319 336021
rect 41492 336016 43319 336018
rect 41492 335960 43258 336016
rect 43314 335960 43319 336016
rect 41492 335958 43319 335960
rect 43253 335955 43319 335958
rect 42701 335610 42767 335613
rect 41492 335608 42767 335610
rect 41492 335552 42706 335608
rect 42762 335552 42767 335608
rect 41492 335550 42767 335552
rect 42701 335547 42767 335550
rect 43621 335202 43687 335205
rect 41492 335200 43687 335202
rect 41492 335144 43626 335200
rect 43682 335144 43687 335200
rect 41492 335142 43687 335144
rect 43621 335139 43687 335142
rect 43437 334794 43503 334797
rect 41492 334792 43503 334794
rect 41492 334736 43442 334792
rect 43498 334736 43503 334792
rect 41492 334734 43503 334736
rect 43437 334731 43503 334734
rect 41462 334114 41522 334356
rect 41597 334114 41663 334117
rect 41462 334112 41663 334114
rect 41462 334056 41602 334112
rect 41658 334056 41663 334112
rect 41462 334054 41663 334056
rect 41597 334051 41663 334054
rect 30422 333540 30482 333948
rect 41462 332890 41522 333132
rect 41597 332890 41663 332893
rect 41462 332888 41663 332890
rect 41462 332832 41602 332888
rect 41658 332832 41663 332888
rect 41462 332830 41663 332832
rect 41597 332827 41663 332830
rect 655513 329898 655579 329901
rect 649950 329896 655579 329898
rect 649950 329840 655518 329896
rect 655574 329840 655579 329896
rect 649950 329838 655579 329840
rect 32857 329762 32923 329765
rect 42190 329762 42196 329764
rect 32857 329760 42196 329762
rect 32857 329704 32862 329760
rect 32918 329704 42196 329760
rect 32857 329702 42196 329704
rect 32857 329699 32923 329702
rect 42190 329700 42196 329702
rect 42260 329700 42266 329764
rect 649950 329234 650010 329838
rect 655513 329835 655579 329838
rect 655605 328266 655671 328269
rect 649950 328264 655671 328266
rect 649950 328208 655610 328264
rect 655666 328208 655671 328264
rect 649950 328206 655671 328208
rect 649950 328052 650010 328206
rect 655605 328203 655671 328206
rect 655421 327450 655487 327453
rect 649950 327448 655487 327450
rect 649950 327392 655426 327448
rect 655482 327392 655487 327448
rect 649950 327390 655487 327392
rect 649950 326870 650010 327390
rect 655421 327387 655487 327390
rect 649950 325682 650010 325688
rect 655973 325682 656039 325685
rect 649950 325680 656039 325682
rect 649950 325624 655978 325680
rect 656034 325624 656039 325680
rect 649950 325622 656039 325624
rect 655973 325619 656039 325622
rect 58433 317386 58499 317389
rect 58433 317384 64706 317386
rect 58433 317328 58438 317384
rect 58494 317328 64706 317384
rect 58433 317326 64706 317328
rect 58433 317323 58499 317326
rect 64646 317106 64706 317326
rect 58157 316570 58223 316573
rect 58157 316568 64706 316570
rect 58157 316512 58162 316568
rect 58218 316512 64706 316568
rect 58157 316510 64706 316512
rect 58157 316507 58223 316510
rect 64646 315924 64706 316510
rect 41965 315620 42031 315621
rect 41965 315616 42012 315620
rect 42076 315618 42082 315620
rect 41965 315560 41970 315616
rect 41965 315556 42012 315560
rect 42076 315558 42122 315618
rect 42076 315556 42082 315558
rect 41965 315555 42031 315556
rect 58341 314802 58407 314805
rect 58341 314800 64706 314802
rect 58341 314744 58346 314800
rect 58402 314744 64706 314800
rect 58341 314742 64706 314744
rect 58341 314739 58407 314742
rect 58525 314122 58591 314125
rect 58525 314120 64706 314122
rect 58525 314064 58530 314120
rect 58586 314064 64706 314120
rect 58525 314062 64706 314064
rect 58525 314059 58591 314062
rect 42149 313852 42215 313853
rect 42149 313850 42196 313852
rect 42104 313848 42196 313850
rect 42104 313792 42154 313848
rect 42104 313790 42196 313792
rect 42149 313788 42196 313790
rect 42260 313788 42266 313852
rect 42149 313787 42215 313788
rect 64646 313560 64706 314062
rect 676262 313581 676322 313684
rect 676262 313576 676371 313581
rect 676262 313520 676310 313576
rect 676366 313520 676371 313576
rect 676262 313518 676371 313520
rect 676305 313515 676371 313518
rect 41781 313172 41847 313173
rect 41781 313168 41828 313172
rect 41892 313170 41898 313172
rect 676121 313170 676187 313173
rect 676262 313170 676322 313276
rect 41781 313112 41786 313168
rect 41781 313108 41828 313112
rect 41892 313110 41938 313170
rect 676121 313168 676322 313170
rect 676121 313112 676126 313168
rect 676182 313112 676322 313168
rect 676121 313110 676322 313112
rect 41892 313108 41898 313110
rect 41781 313107 41847 313108
rect 676121 313107 676187 313110
rect 58157 313034 58223 313037
rect 58157 313032 64706 313034
rect 58157 312976 58162 313032
rect 58218 312976 64706 313032
rect 58157 312974 64706 312976
rect 58157 312971 58223 312974
rect 64646 312378 64706 312974
rect 676262 312765 676322 312868
rect 676213 312760 676322 312765
rect 676213 312704 676218 312760
rect 676274 312704 676322 312760
rect 676213 312702 676322 312704
rect 676213 312699 676279 312702
rect 676029 312490 676095 312493
rect 676029 312488 676292 312490
rect 676029 312432 676034 312488
rect 676090 312432 676292 312488
rect 676029 312430 676292 312432
rect 676029 312427 676095 312430
rect 41638 312292 41644 312356
rect 41708 312354 41714 312356
rect 41781 312354 41847 312357
rect 41708 312352 41847 312354
rect 41708 312296 41786 312352
rect 41842 312296 41847 312352
rect 41708 312294 41847 312296
rect 41708 312292 41714 312294
rect 41781 312291 41847 312294
rect 676262 311949 676322 312052
rect 676213 311944 676322 311949
rect 676213 311888 676218 311944
rect 676274 311888 676322 311944
rect 676213 311886 676322 311888
rect 676213 311883 676279 311886
rect 58525 311810 58591 311813
rect 58525 311808 64706 311810
rect 58525 311752 58530 311808
rect 58586 311752 64706 311808
rect 58525 311750 64706 311752
rect 58525 311747 58591 311750
rect 64646 311196 64706 311750
rect 676029 311674 676095 311677
rect 676029 311672 676292 311674
rect 676029 311616 676034 311672
rect 676090 311616 676292 311672
rect 676029 311614 676292 311616
rect 676029 311611 676095 311614
rect 676262 311133 676322 311236
rect 676213 311128 676322 311133
rect 676213 311072 676218 311128
rect 676274 311072 676322 311128
rect 676213 311070 676322 311072
rect 676213 311067 676279 311070
rect 676262 310725 676322 310828
rect 676213 310720 676322 310725
rect 676213 310664 676218 310720
rect 676274 310664 676322 310720
rect 676213 310662 676322 310664
rect 676213 310659 676279 310662
rect 676262 310317 676322 310420
rect 676213 310312 676322 310317
rect 676213 310256 676218 310312
rect 676274 310256 676322 310312
rect 676213 310254 676322 310256
rect 676213 310251 676279 310254
rect 676262 309909 676322 310012
rect 676213 309904 676322 309909
rect 676213 309848 676218 309904
rect 676274 309848 676322 309904
rect 676213 309846 676322 309848
rect 676213 309843 676279 309846
rect 676262 309501 676322 309604
rect 676213 309496 676322 309501
rect 676213 309440 676218 309496
rect 676274 309440 676322 309496
rect 676213 309438 676322 309440
rect 676213 309435 676279 309438
rect 676029 309226 676095 309229
rect 676029 309224 676292 309226
rect 676029 309168 676034 309224
rect 676090 309168 676292 309224
rect 676029 309166 676292 309168
rect 676029 309163 676095 309166
rect 676029 308818 676095 308821
rect 676029 308816 676292 308818
rect 676029 308760 676034 308816
rect 676090 308760 676292 308816
rect 676029 308758 676292 308760
rect 676029 308755 676095 308758
rect 675293 308410 675359 308413
rect 675293 308408 676292 308410
rect 675293 308352 675298 308408
rect 675354 308352 676292 308408
rect 675293 308350 676292 308352
rect 675293 308347 675359 308350
rect 676029 308002 676095 308005
rect 676029 308000 676292 308002
rect 676029 307944 676034 308000
rect 676090 307944 676292 308000
rect 676029 307942 676292 307944
rect 676029 307939 676095 307942
rect 676121 307458 676187 307461
rect 676262 307458 676322 307564
rect 676121 307456 676322 307458
rect 676121 307400 676126 307456
rect 676182 307400 676322 307456
rect 676121 307398 676322 307400
rect 676121 307395 676187 307398
rect 675385 307186 675451 307189
rect 675385 307184 676292 307186
rect 675385 307128 675390 307184
rect 675446 307128 676292 307184
rect 675385 307126 676292 307128
rect 675385 307123 675451 307126
rect 676029 306778 676095 306781
rect 676029 306776 676292 306778
rect 676029 306720 676034 306776
rect 676090 306720 676292 306776
rect 676029 306718 676292 306720
rect 676029 306715 676095 306718
rect 676029 306370 676095 306373
rect 676029 306368 676292 306370
rect 676029 306312 676034 306368
rect 676090 306312 676292 306368
rect 676029 306310 676292 306312
rect 676029 306307 676095 306310
rect 676029 305962 676095 305965
rect 676029 305960 676292 305962
rect 676029 305904 676034 305960
rect 676090 305904 676292 305960
rect 676029 305902 676292 305904
rect 676029 305899 676095 305902
rect 676121 305418 676187 305421
rect 676262 305418 676322 305524
rect 676121 305416 676322 305418
rect 676121 305360 676126 305416
rect 676182 305360 676322 305416
rect 676121 305358 676322 305360
rect 676121 305355 676187 305358
rect 676121 305010 676187 305013
rect 676262 305010 676322 305116
rect 676121 305008 676322 305010
rect 676121 304952 676126 305008
rect 676182 304952 676322 305008
rect 676121 304950 676322 304952
rect 676121 304947 676187 304950
rect 676029 304738 676095 304741
rect 676029 304736 676292 304738
rect 676029 304680 676034 304736
rect 676090 304680 676292 304736
rect 676029 304678 676292 304680
rect 676029 304675 676095 304678
rect 676121 304194 676187 304197
rect 676262 304194 676322 304300
rect 676121 304192 676322 304194
rect 676121 304136 676126 304192
rect 676182 304136 676322 304192
rect 676121 304134 676322 304136
rect 676121 304131 676187 304134
rect 676029 303922 676095 303925
rect 676029 303920 676292 303922
rect 676029 303864 676034 303920
rect 676090 303864 676292 303920
rect 676029 303862 676292 303864
rect 676029 303859 676095 303862
rect 679022 303381 679082 303484
rect 655513 303378 655579 303381
rect 649950 303376 655579 303378
rect 649950 303320 655518 303376
rect 655574 303320 655579 303376
rect 649950 303318 655579 303320
rect 649950 302776 650010 303318
rect 655513 303315 655579 303318
rect 678973 303376 679082 303381
rect 678973 303320 678978 303376
rect 679034 303320 679082 303376
rect 678973 303318 679082 303320
rect 678973 303315 679039 303318
rect 684542 302668 684602 303076
rect 678973 302562 679039 302565
rect 678973 302560 679082 302562
rect 678973 302504 678978 302560
rect 679034 302504 679082 302560
rect 678973 302499 679082 302504
rect 679022 302260 679082 302499
rect 655697 302154 655763 302157
rect 649950 302152 655763 302154
rect 649950 302096 655702 302152
rect 655758 302096 655763 302152
rect 649950 302094 655763 302096
rect 649950 301594 650010 302094
rect 655697 302091 655763 302094
rect 41781 301338 41847 301341
rect 41492 301336 41847 301338
rect 41492 301280 41786 301336
rect 41842 301280 41847 301336
rect 41492 301278 41847 301280
rect 41781 301275 41847 301278
rect 41873 300930 41939 300933
rect 41492 300928 41939 300930
rect 41492 300872 41878 300928
rect 41934 300872 41939 300928
rect 41492 300870 41939 300872
rect 41873 300867 41939 300870
rect 655421 300794 655487 300797
rect 649950 300792 655487 300794
rect 649950 300736 655426 300792
rect 655482 300736 655487 300792
rect 649950 300734 655487 300736
rect 42701 300522 42767 300525
rect 41492 300520 42767 300522
rect 41492 300464 42706 300520
rect 42762 300464 42767 300520
rect 41492 300462 42767 300464
rect 42701 300459 42767 300462
rect 649950 300412 650010 300734
rect 655421 300731 655487 300734
rect 44589 300114 44659 300119
rect 41586 300054 44594 300114
rect 44654 300054 44668 300114
rect 44589 300049 44659 300054
rect 44589 299732 44659 299735
rect 41586 299730 44668 299732
rect 41586 299672 44594 299730
rect 44589 299670 44594 299672
rect 44654 299672 44668 299730
rect 44654 299670 44659 299672
rect 44589 299665 44659 299670
rect 41781 299298 41847 299301
rect 41492 299296 41847 299298
rect 41492 299240 41786 299296
rect 41842 299240 41847 299296
rect 41492 299238 41847 299240
rect 41781 299235 41847 299238
rect 43069 298890 43135 298893
rect 41492 298888 43135 298890
rect 41492 298832 43074 298888
rect 43130 298832 43135 298888
rect 41492 298830 43135 298832
rect 43069 298827 43135 298830
rect 649950 298754 650010 299230
rect 655053 298754 655119 298757
rect 649950 298752 655119 298754
rect 649950 298696 655058 298752
rect 655114 298696 655119 298752
rect 649950 298694 655119 298696
rect 655053 298691 655119 298694
rect 44681 298480 44751 298483
rect 41586 298478 44758 298480
rect 41586 298420 44686 298478
rect 44681 298418 44686 298420
rect 44746 298420 44758 298478
rect 44746 298418 44751 298420
rect 44681 298413 44751 298418
rect 42701 298210 42767 298213
rect 58433 298210 58499 298213
rect 42701 298208 58499 298210
rect 42701 298152 42706 298208
rect 42762 298152 58438 298208
rect 58494 298152 58499 298208
rect 42701 298150 58499 298152
rect 42701 298147 42767 298150
rect 58433 298147 58499 298150
rect 44681 298068 44751 298073
rect 44681 298066 44686 298068
rect 41586 298008 44686 298066
rect 44746 298066 44751 298068
rect 44746 298008 44758 298066
rect 41586 298006 44758 298008
rect 44681 298003 44751 298006
rect 44773 297688 44843 297693
rect 41586 297628 44778 297688
rect 44838 297628 44864 297688
rect 44773 297623 44843 297628
rect 649950 297530 650010 298048
rect 656157 297530 656223 297533
rect 649950 297528 656223 297530
rect 649950 297472 656162 297528
rect 656218 297472 656223 297528
rect 649950 297470 656223 297472
rect 656157 297467 656223 297470
rect 44773 297276 44843 297281
rect 44773 297270 44778 297276
rect 41586 297216 44778 297270
rect 44838 297270 44843 297276
rect 44838 297216 44864 297270
rect 41586 297210 44864 297216
rect 41822 296850 41828 296852
rect 41492 296790 41828 296850
rect 41822 296788 41828 296790
rect 41892 296788 41898 296852
rect 43621 296442 43687 296445
rect 41492 296440 43687 296442
rect 41492 296384 43626 296440
rect 43682 296384 43687 296440
rect 41492 296382 43687 296384
rect 43621 296379 43687 296382
rect 649950 296306 650010 296866
rect 655789 296306 655855 296309
rect 649950 296304 655855 296306
rect 649950 296248 655794 296304
rect 655850 296248 655855 296304
rect 649950 296246 655855 296248
rect 655789 296243 655855 296246
rect 43253 296034 43319 296037
rect 41492 296032 43319 296034
rect 41492 295976 43258 296032
rect 43314 295976 43319 296032
rect 41492 295974 43319 295976
rect 43253 295971 43319 295974
rect 43713 295626 43779 295629
rect 41492 295624 43779 295626
rect 41492 295568 43718 295624
rect 43774 295568 43779 295624
rect 41492 295566 43779 295568
rect 43713 295563 43779 295566
rect 58525 295490 58591 295493
rect 64646 295490 64706 295684
rect 58525 295488 64706 295490
rect 58525 295432 58530 295488
rect 58586 295432 64706 295488
rect 58525 295430 64706 295432
rect 58525 295427 58591 295430
rect 649950 295354 650010 295684
rect 655973 295354 656039 295357
rect 649950 295352 656039 295354
rect 649950 295296 655978 295352
rect 656034 295296 656039 295352
rect 649950 295294 656039 295296
rect 655973 295291 656039 295294
rect 43529 295218 43595 295221
rect 41492 295216 43595 295218
rect 41492 295160 43534 295216
rect 43590 295160 43595 295216
rect 41492 295158 43595 295160
rect 43529 295155 43595 295158
rect 41873 294810 41939 294813
rect 41492 294808 41939 294810
rect 41492 294752 41878 294808
rect 41934 294752 41939 294808
rect 41492 294750 41939 294752
rect 41873 294747 41939 294750
rect 43897 294402 43963 294405
rect 41492 294400 43963 294402
rect 41492 294344 43902 294400
rect 43958 294344 43963 294400
rect 41492 294342 43963 294344
rect 43897 294339 43963 294342
rect 42425 293994 42491 293997
rect 41492 293992 42491 293994
rect 41492 293936 42430 293992
rect 42486 293936 42491 293992
rect 41492 293934 42491 293936
rect 42425 293931 42491 293934
rect 58341 293994 58407 293997
rect 64646 293994 64706 294502
rect 58341 293992 64706 293994
rect 58341 293936 58346 293992
rect 58402 293936 64706 293992
rect 58341 293934 64706 293936
rect 649950 293994 650010 294502
rect 655605 293994 655671 293997
rect 649950 293992 655671 293994
rect 649950 293936 655610 293992
rect 655666 293936 655671 293992
rect 649950 293934 655671 293936
rect 58341 293931 58407 293934
rect 655605 293931 655671 293934
rect 43989 293586 44055 293589
rect 41492 293584 44055 293586
rect 41492 293528 43994 293584
rect 44050 293528 44055 293584
rect 41492 293526 44055 293528
rect 43989 293523 44055 293526
rect 43161 293178 43227 293181
rect 41492 293176 43227 293178
rect 41492 293120 43166 293176
rect 43222 293120 43227 293176
rect 41492 293118 43227 293120
rect 43161 293115 43227 293118
rect 30005 292770 30071 292773
rect 59445 292770 59511 292773
rect 64646 292770 64706 293320
rect 30005 292768 30084 292770
rect 30005 292712 30010 292768
rect 30066 292712 30084 292768
rect 30005 292710 30084 292712
rect 59445 292768 64706 292770
rect 59445 292712 59450 292768
rect 59506 292712 64706 292768
rect 59445 292710 64706 292712
rect 649950 292770 650010 293320
rect 655421 292770 655487 292773
rect 649950 292768 655487 292770
rect 649950 292712 655426 292768
rect 655482 292712 655487 292768
rect 649950 292710 655487 292712
rect 30005 292707 30071 292710
rect 59445 292707 59511 292710
rect 655421 292707 655487 292710
rect 58433 292498 58499 292501
rect 58433 292496 64706 292498
rect 58433 292440 58438 292496
rect 58494 292440 64706 292496
rect 58433 292438 64706 292440
rect 58433 292435 58499 292438
rect 44081 292362 44147 292365
rect 41492 292360 44147 292362
rect 41492 292304 44086 292360
rect 44142 292304 44147 292360
rect 41492 292302 44147 292304
rect 44081 292299 44147 292302
rect 64646 292138 64706 292438
rect 41781 291954 41847 291957
rect 41492 291952 41847 291954
rect 41492 291896 41786 291952
rect 41842 291896 41847 291952
rect 41492 291894 41847 291896
rect 41781 291891 41847 291894
rect 41781 291546 41847 291549
rect 41492 291544 41847 291546
rect 41492 291488 41786 291544
rect 41842 291488 41847 291544
rect 41492 291486 41847 291488
rect 41781 291483 41847 291486
rect 57881 291546 57947 291549
rect 649950 291546 650010 292138
rect 655513 291546 655579 291549
rect 57881 291544 64706 291546
rect 57881 291488 57886 291544
rect 57942 291488 64706 291544
rect 57881 291486 64706 291488
rect 649950 291544 655579 291546
rect 649950 291488 655518 291544
rect 655574 291488 655579 291544
rect 649950 291486 655579 291488
rect 57881 291483 57947 291486
rect 61837 291138 61903 291141
rect 41492 291136 61903 291138
rect 41492 291080 61842 291136
rect 61898 291080 61903 291136
rect 41492 291078 61903 291080
rect 61837 291075 61903 291078
rect 64646 290956 64706 291486
rect 655513 291483 655579 291486
rect 50981 290730 51047 290733
rect 41492 290728 51047 290730
rect 41492 290672 50986 290728
rect 51042 290672 51047 290728
rect 41492 290670 51047 290672
rect 50981 290667 51047 290670
rect 649950 290458 650010 290956
rect 655697 290458 655763 290461
rect 649950 290456 655763 290458
rect 649950 290400 655702 290456
rect 655758 290400 655763 290456
rect 649950 290398 655763 290400
rect 655697 290395 655763 290398
rect 48589 289914 48655 289917
rect 41492 289912 48655 289914
rect 41492 289856 48594 289912
rect 48650 289856 48655 289912
rect 41492 289854 48655 289856
rect 48589 289851 48655 289854
rect 58525 289778 58591 289781
rect 58525 289776 64706 289778
rect 58525 289720 58530 289776
rect 58586 289720 64706 289776
rect 58525 289718 64706 289720
rect 58525 289715 58591 289718
rect 649950 289234 650010 289774
rect 654133 289234 654199 289237
rect 649950 289232 654199 289234
rect 649950 289176 654138 289232
rect 654194 289176 654199 289232
rect 649950 289174 654199 289176
rect 654133 289171 654199 289174
rect 57973 288010 58039 288013
rect 64646 288010 64706 288592
rect 57973 288008 64706 288010
rect 57973 287952 57978 288008
rect 58034 287952 64706 288008
rect 57973 287950 64706 287952
rect 649950 288010 650010 288592
rect 654133 288010 654199 288013
rect 649950 288008 654199 288010
rect 649950 287952 654138 288008
rect 654194 287952 654199 288008
rect 649950 287950 654199 287952
rect 57973 287947 58039 287950
rect 654133 287947 654199 287950
rect 58525 287194 58591 287197
rect 64646 287194 64706 287410
rect 649766 287406 651390 287466
rect 651330 287330 651390 287406
rect 656801 287330 656867 287333
rect 651330 287328 656867 287330
rect 651330 287272 656806 287328
rect 656862 287272 656867 287328
rect 651330 287270 656867 287272
rect 656801 287267 656867 287270
rect 58525 287192 64706 287194
rect 58525 287136 58530 287192
rect 58586 287136 64706 287192
rect 58525 287134 64706 287136
rect 58525 287131 58591 287134
rect 57973 285698 58039 285701
rect 64646 285698 64706 286228
rect 57973 285696 64706 285698
rect 57973 285640 57978 285696
rect 58034 285640 64706 285696
rect 57973 285638 64706 285640
rect 649950 285698 650010 286228
rect 655237 285698 655303 285701
rect 649950 285696 655303 285698
rect 649950 285640 655242 285696
rect 655298 285640 655303 285696
rect 649950 285638 655303 285640
rect 57973 285635 58039 285638
rect 655237 285635 655303 285638
rect 58525 284474 58591 284477
rect 64646 284474 64706 285046
rect 649950 284746 650010 285046
rect 654501 284746 654567 284749
rect 649950 284744 654567 284746
rect 649950 284688 654506 284744
rect 654562 284688 654567 284744
rect 649950 284686 654567 284688
rect 654501 284683 654567 284686
rect 58525 284472 64706 284474
rect 58525 284416 58530 284472
rect 58586 284416 64706 284472
rect 58525 284414 64706 284416
rect 58525 284411 58591 284414
rect 57973 283250 58039 283253
rect 64646 283250 64706 283864
rect 649950 283658 650010 283864
rect 654225 283658 654291 283661
rect 649950 283656 654291 283658
rect 649950 283600 654230 283656
rect 654286 283600 654291 283656
rect 649950 283598 654291 283600
rect 654225 283595 654291 283598
rect 57973 283248 64706 283250
rect 57973 283192 57978 283248
rect 58034 283192 64706 283248
rect 57973 283190 64706 283192
rect 57973 283187 58039 283190
rect 59261 282162 59327 282165
rect 64646 282162 64706 282682
rect 59261 282160 64706 282162
rect 59261 282104 59266 282160
rect 59322 282104 64706 282160
rect 59261 282102 64706 282104
rect 649950 282162 650010 282682
rect 655237 282162 655303 282165
rect 649950 282160 655303 282162
rect 649950 282104 655242 282160
rect 655298 282104 655303 282160
rect 649950 282102 655303 282104
rect 59261 282099 59327 282102
rect 655237 282099 655303 282102
rect 59537 280938 59603 280941
rect 64646 280938 64706 281500
rect 59537 280936 64706 280938
rect 59537 280880 59542 280936
rect 59598 280880 64706 280936
rect 59537 280878 64706 280880
rect 649950 280938 650010 281500
rect 654133 280938 654199 280941
rect 649950 280936 654199 280938
rect 649950 280880 654138 280936
rect 654194 280880 654199 280936
rect 649950 280878 654199 280880
rect 59537 280875 59603 280878
rect 654133 280875 654199 280878
rect 59353 279714 59419 279717
rect 64646 279714 64706 280318
rect 59353 279712 64706 279714
rect 59353 279656 59358 279712
rect 59414 279656 64706 279712
rect 59353 279654 64706 279656
rect 649950 279714 650010 280318
rect 654869 279714 654935 279717
rect 649950 279712 654935 279714
rect 649950 279656 654874 279712
rect 654930 279656 654935 279712
rect 649950 279654 654935 279656
rect 59353 279651 59419 279654
rect 654869 279651 654935 279654
rect 60774 275980 60780 276044
rect 60844 276042 60850 276044
rect 63401 276042 63467 276045
rect 60844 276040 63467 276042
rect 60844 275984 63406 276040
rect 63462 275984 63467 276040
rect 60844 275982 63467 275984
rect 60844 275980 60850 275982
rect 63401 275979 63467 275982
rect 397361 275906 397427 275909
rect 609605 275906 609671 275909
rect 397361 275904 609671 275906
rect 397361 275848 397366 275904
rect 397422 275848 609610 275904
rect 609666 275848 609671 275904
rect 397361 275846 609671 275848
rect 397361 275843 397427 275846
rect 609605 275843 609671 275846
rect 396257 275770 396323 275773
rect 607213 275770 607279 275773
rect 396257 275768 607279 275770
rect 396257 275712 396262 275768
rect 396318 275712 607218 275768
rect 607274 275712 607279 275768
rect 396257 275710 607279 275712
rect 396257 275707 396323 275710
rect 607213 275707 607279 275710
rect 398925 275634 398991 275637
rect 614297 275634 614363 275637
rect 398925 275632 614363 275634
rect 398925 275576 398930 275632
rect 398986 275576 614302 275632
rect 614358 275576 614363 275632
rect 398925 275574 614363 275576
rect 398925 275571 398991 275574
rect 614297 275571 614363 275574
rect 398465 275498 398531 275501
rect 613101 275498 613167 275501
rect 398465 275496 613167 275498
rect 398465 275440 398470 275496
rect 398526 275440 613106 275496
rect 613162 275440 613167 275496
rect 398465 275438 613167 275440
rect 398465 275435 398531 275438
rect 613101 275435 613167 275438
rect 401133 275362 401199 275365
rect 620185 275362 620251 275365
rect 401133 275360 620251 275362
rect 401133 275304 401138 275360
rect 401194 275304 620190 275360
rect 620246 275304 620251 275360
rect 401133 275302 620251 275304
rect 401133 275299 401199 275302
rect 620185 275299 620251 275302
rect 399845 275226 399911 275229
rect 616689 275226 616755 275229
rect 399845 275224 616755 275226
rect 399845 275168 399850 275224
rect 399906 275168 616694 275224
rect 616750 275168 616755 275224
rect 399845 275166 616755 275168
rect 399845 275163 399911 275166
rect 616689 275163 616755 275166
rect 401961 275090 402027 275093
rect 621381 275090 621447 275093
rect 401961 275088 621447 275090
rect 401961 275032 401966 275088
rect 402022 275032 621386 275088
rect 621442 275032 621447 275088
rect 401961 275030 621447 275032
rect 401961 275027 402027 275030
rect 621381 275027 621447 275030
rect 402513 274954 402579 274957
rect 623773 274954 623839 274957
rect 402513 274952 623839 274954
rect 402513 274896 402518 274952
rect 402574 274896 623778 274952
rect 623834 274896 623839 274952
rect 402513 274894 623839 274896
rect 402513 274891 402579 274894
rect 623773 274891 623839 274894
rect 405181 274818 405247 274821
rect 630857 274818 630923 274821
rect 405181 274816 630923 274818
rect 405181 274760 405186 274816
rect 405242 274760 630862 274816
rect 630918 274760 630923 274816
rect 405181 274758 630923 274760
rect 405181 274755 405247 274758
rect 630857 274755 630923 274758
rect 408309 274682 408375 274685
rect 639137 274682 639203 274685
rect 408309 274680 639203 274682
rect 408309 274624 408314 274680
rect 408370 274624 639142 274680
rect 639198 274624 639203 274680
rect 408309 274622 639203 274624
rect 408309 274619 408375 274622
rect 639137 274619 639203 274622
rect 407849 274546 407915 274549
rect 637941 274546 638007 274549
rect 407849 274544 638007 274546
rect 407849 274488 407854 274544
rect 407910 274488 637946 274544
rect 638002 274488 638007 274544
rect 407849 274486 638007 274488
rect 407849 274483 407915 274486
rect 637941 274483 638007 274486
rect 395797 274410 395863 274413
rect 606017 274410 606083 274413
rect 395797 274408 606083 274410
rect 395797 274352 395802 274408
rect 395858 274352 606022 274408
rect 606078 274352 606083 274408
rect 395797 274350 606083 274352
rect 395797 274347 395863 274350
rect 606017 274347 606083 274350
rect 393589 274274 393655 274277
rect 600129 274274 600195 274277
rect 393589 274272 600195 274274
rect 393589 274216 393594 274272
rect 393650 274216 600134 274272
rect 600190 274216 600195 274272
rect 393589 274214 600195 274216
rect 393589 274211 393655 274214
rect 600129 274211 600195 274214
rect 106089 273186 106155 273189
rect 207473 273186 207539 273189
rect 106089 273184 207539 273186
rect 106089 273128 106094 273184
rect 106150 273128 207478 273184
rect 207534 273128 207539 273184
rect 106089 273126 207539 273128
rect 106089 273123 106155 273126
rect 207473 273123 207539 273126
rect 364057 273186 364123 273189
rect 522113 273186 522179 273189
rect 364057 273184 522179 273186
rect 364057 273128 364062 273184
rect 364118 273128 522118 273184
rect 522174 273128 522179 273184
rect 364057 273126 522179 273128
rect 364057 273123 364123 273126
rect 522113 273123 522179 273126
rect 103697 273050 103763 273053
rect 207013 273050 207079 273053
rect 103697 273048 207079 273050
rect 103697 272992 103702 273048
rect 103758 272992 207018 273048
rect 207074 272992 207079 273048
rect 103697 272990 207079 272992
rect 103697 272987 103763 272990
rect 207013 272987 207079 272990
rect 366909 273050 366975 273053
rect 529197 273050 529263 273053
rect 366909 273048 529263 273050
rect 366909 272992 366914 273048
rect 366970 272992 529202 273048
rect 529258 272992 529263 273048
rect 366909 272990 529263 272992
rect 366909 272987 366975 272990
rect 529197 272987 529263 272990
rect 96613 272914 96679 272917
rect 204345 272914 204411 272917
rect 96613 272912 204411 272914
rect 96613 272856 96618 272912
rect 96674 272856 204350 272912
rect 204406 272856 204411 272912
rect 96613 272854 204411 272856
rect 96613 272851 96679 272854
rect 204345 272851 204411 272854
rect 368657 272914 368723 272917
rect 533889 272914 533955 272917
rect 368657 272912 533955 272914
rect 368657 272856 368662 272912
rect 368718 272856 533894 272912
rect 533950 272856 533955 272912
rect 368657 272854 533955 272856
rect 368657 272851 368723 272854
rect 533889 272851 533955 272854
rect 99005 272778 99071 272781
rect 204805 272778 204871 272781
rect 99005 272776 204871 272778
rect 99005 272720 99010 272776
rect 99066 272720 204810 272776
rect 204866 272720 204871 272776
rect 99005 272718 204871 272720
rect 99005 272715 99071 272718
rect 204805 272715 204871 272718
rect 369669 272778 369735 272781
rect 536281 272778 536347 272781
rect 369669 272776 536347 272778
rect 369669 272720 369674 272776
rect 369730 272720 536286 272776
rect 536342 272720 536347 272776
rect 369669 272718 536347 272720
rect 369669 272715 369735 272718
rect 536281 272715 536347 272718
rect 88333 272642 88399 272645
rect 201217 272642 201283 272645
rect 88333 272640 201283 272642
rect 88333 272584 88338 272640
rect 88394 272584 201222 272640
rect 201278 272584 201283 272640
rect 88333 272582 201283 272584
rect 88333 272579 88399 272582
rect 201217 272579 201283 272582
rect 372613 272642 372679 272645
rect 540973 272642 541039 272645
rect 372613 272640 541039 272642
rect 372613 272584 372618 272640
rect 372674 272584 540978 272640
rect 541034 272584 541039 272640
rect 372613 272582 541039 272584
rect 372613 272579 372679 272582
rect 540973 272579 541039 272582
rect 90725 272506 90791 272509
rect 201677 272506 201743 272509
rect 90725 272504 201743 272506
rect 90725 272448 90730 272504
rect 90786 272448 201682 272504
rect 201738 272448 201743 272504
rect 90725 272446 201743 272448
rect 90725 272443 90791 272446
rect 201677 272443 201743 272446
rect 372429 272506 372495 272509
rect 543365 272506 543431 272509
rect 372429 272504 543431 272506
rect 372429 272448 372434 272504
rect 372490 272448 543370 272504
rect 543426 272448 543431 272504
rect 372429 272446 543431 272448
rect 372429 272443 372495 272446
rect 543365 272443 543431 272446
rect 80053 272370 80119 272373
rect 196893 272370 196959 272373
rect 80053 272368 196959 272370
rect 80053 272312 80058 272368
rect 80114 272312 196898 272368
rect 196954 272312 196959 272368
rect 80053 272310 196959 272312
rect 80053 272307 80119 272310
rect 196893 272307 196959 272310
rect 380709 272370 380775 272373
rect 565813 272370 565879 272373
rect 380709 272368 565879 272370
rect 380709 272312 380714 272368
rect 380770 272312 565818 272368
rect 565874 272312 565879 272368
rect 380709 272310 565879 272312
rect 380709 272307 380775 272310
rect 565813 272307 565879 272310
rect 83641 272234 83707 272237
rect 199101 272234 199167 272237
rect 83641 272232 199167 272234
rect 83641 272176 83646 272232
rect 83702 272176 199106 272232
rect 199162 272176 199167 272232
rect 83641 272174 199167 272176
rect 83641 272171 83707 272174
rect 199101 272171 199167 272174
rect 395429 272234 395495 272237
rect 604821 272234 604887 272237
rect 395429 272232 604887 272234
rect 395429 272176 395434 272232
rect 395490 272176 604826 272232
rect 604882 272176 604887 272232
rect 395429 272174 604887 272176
rect 395429 272171 395495 272174
rect 604821 272171 604887 272174
rect 81249 272098 81315 272101
rect 198089 272098 198155 272101
rect 81249 272096 198155 272098
rect 81249 272040 81254 272096
rect 81310 272040 198094 272096
rect 198150 272040 198155 272096
rect 81249 272038 198155 272040
rect 81249 272035 81315 272038
rect 198089 272035 198155 272038
rect 404721 272098 404787 272101
rect 629661 272098 629727 272101
rect 404721 272096 629727 272098
rect 404721 272040 404726 272096
rect 404782 272040 629666 272096
rect 629722 272040 629727 272096
rect 404721 272038 629727 272040
rect 404721 272035 404787 272038
rect 629661 272035 629727 272038
rect 70577 271962 70643 271965
rect 194133 271962 194199 271965
rect 70577 271960 194199 271962
rect 70577 271904 70582 271960
rect 70638 271904 194138 271960
rect 194194 271904 194199 271960
rect 70577 271902 194199 271904
rect 70577 271899 70643 271902
rect 194133 271899 194199 271902
rect 410517 271962 410583 271965
rect 645025 271962 645091 271965
rect 410517 271960 645091 271962
rect 410517 271904 410522 271960
rect 410578 271904 645030 271960
rect 645086 271904 645091 271960
rect 410517 271902 645091 271904
rect 410517 271899 410583 271902
rect 645025 271899 645091 271902
rect 69381 271826 69447 271829
rect 193673 271826 193739 271829
rect 69381 271824 193739 271826
rect 69381 271768 69386 271824
rect 69442 271768 193678 271824
rect 193734 271768 193739 271824
rect 69381 271766 193739 271768
rect 69381 271763 69447 271766
rect 193673 271763 193739 271766
rect 410057 271826 410123 271829
rect 643829 271826 643895 271829
rect 410057 271824 643895 271826
rect 410057 271768 410062 271824
rect 410118 271768 643834 271824
rect 643890 271768 643895 271824
rect 410057 271766 643895 271768
rect 410057 271763 410123 271766
rect 643829 271763 643895 271766
rect 111977 271690 112043 271693
rect 209221 271690 209287 271693
rect 111977 271688 209287 271690
rect 111977 271632 111982 271688
rect 112038 271632 209226 271688
rect 209282 271632 209287 271688
rect 111977 271630 209287 271632
rect 111977 271627 112043 271630
rect 209221 271627 209287 271630
rect 361021 271690 361087 271693
rect 512637 271690 512703 271693
rect 361021 271688 512703 271690
rect 361021 271632 361026 271688
rect 361082 271632 512642 271688
rect 512698 271632 512703 271688
rect 361021 271630 512703 271632
rect 361021 271627 361087 271630
rect 512637 271627 512703 271630
rect 115473 271554 115539 271557
rect 210601 271554 210667 271557
rect 115473 271552 210667 271554
rect 115473 271496 115478 271552
rect 115534 271496 210606 271552
rect 210662 271496 210667 271552
rect 115473 271494 210667 271496
rect 115473 271491 115539 271494
rect 210601 271491 210667 271494
rect 358905 271554 358971 271557
rect 507945 271554 508011 271557
rect 358905 271552 508011 271554
rect 358905 271496 358910 271552
rect 358966 271496 507950 271552
rect 508006 271496 508011 271552
rect 358905 271494 508011 271496
rect 358905 271491 358971 271494
rect 507945 271491 508011 271494
rect 110781 271418 110847 271421
rect 209681 271418 209747 271421
rect 110781 271416 209747 271418
rect 110781 271360 110786 271416
rect 110842 271360 209686 271416
rect 209742 271360 209747 271416
rect 110781 271358 209747 271360
rect 110781 271355 110847 271358
rect 209681 271355 209747 271358
rect 357985 271418 358051 271421
rect 505553 271418 505619 271421
rect 357985 271416 505619 271418
rect 357985 271360 357990 271416
rect 358046 271360 505558 271416
rect 505614 271360 505619 271416
rect 357985 271358 505619 271360
rect 357985 271355 358051 271358
rect 505553 271355 505619 271358
rect 117865 271282 117931 271285
rect 212349 271282 212415 271285
rect 117865 271280 212415 271282
rect 117865 271224 117870 271280
rect 117926 271224 212354 271280
rect 212410 271224 212415 271280
rect 117865 271222 212415 271224
rect 117865 271219 117931 271222
rect 212349 271219 212415 271222
rect 355317 271282 355383 271285
rect 498469 271282 498535 271285
rect 355317 271280 498535 271282
rect 355317 271224 355322 271280
rect 355378 271224 498474 271280
rect 498530 271224 498535 271280
rect 355317 271222 498535 271224
rect 355317 271219 355383 271222
rect 498469 271219 498535 271222
rect 122557 271146 122623 271149
rect 213269 271146 213335 271149
rect 122557 271144 213335 271146
rect 122557 271088 122562 271144
rect 122618 271088 213274 271144
rect 213330 271088 213335 271144
rect 122557 271086 213335 271088
rect 122557 271083 122623 271086
rect 213269 271083 213335 271086
rect 353017 271146 353083 271149
rect 491385 271146 491451 271149
rect 353017 271144 491451 271146
rect 353017 271088 353022 271144
rect 353078 271088 491390 271144
rect 491446 271088 491451 271144
rect 353017 271086 491451 271088
rect 353017 271083 353083 271086
rect 491385 271083 491451 271086
rect 41638 270404 41644 270468
rect 41708 270466 41714 270468
rect 41781 270466 41847 270469
rect 41708 270464 41847 270466
rect 41708 270408 41786 270464
rect 41842 270408 41847 270464
rect 41708 270406 41847 270408
rect 41708 270404 41714 270406
rect 41781 270403 41847 270406
rect 120257 270466 120323 270469
rect 212809 270466 212875 270469
rect 120257 270464 212875 270466
rect 120257 270408 120262 270464
rect 120318 270408 212814 270464
rect 212870 270408 212875 270464
rect 120257 270406 212875 270408
rect 120257 270403 120323 270406
rect 212809 270403 212875 270406
rect 362861 270466 362927 270469
rect 518525 270466 518591 270469
rect 362861 270464 518591 270466
rect 362861 270408 362866 270464
rect 362922 270408 518530 270464
rect 518586 270408 518591 270464
rect 362861 270406 518591 270408
rect 362861 270403 362927 270406
rect 518525 270403 518591 270406
rect 107193 270330 107259 270333
rect 208393 270330 208459 270333
rect 107193 270328 208459 270330
rect 107193 270272 107198 270328
rect 107254 270272 208398 270328
rect 208454 270272 208459 270328
rect 107193 270270 208459 270272
rect 107193 270267 107259 270270
rect 208393 270267 208459 270270
rect 362033 270330 362099 270333
rect 516225 270330 516291 270333
rect 362033 270328 516291 270330
rect 362033 270272 362038 270328
rect 362094 270272 516230 270328
rect 516286 270272 516291 270328
rect 362033 270270 516291 270272
rect 362033 270267 362099 270270
rect 516225 270267 516291 270270
rect 101305 270194 101371 270197
rect 205265 270194 205331 270197
rect 101305 270192 205331 270194
rect 101305 270136 101310 270192
rect 101366 270136 205270 270192
rect 205326 270136 205331 270192
rect 101305 270134 205331 270136
rect 101305 270131 101371 270134
rect 205265 270131 205331 270134
rect 365529 270194 365595 270197
rect 525609 270194 525675 270197
rect 365529 270192 525675 270194
rect 365529 270136 365534 270192
rect 365590 270136 525614 270192
rect 525670 270136 525675 270192
rect 365529 270134 525675 270136
rect 365529 270131 365595 270134
rect 525609 270131 525675 270134
rect 100109 270058 100175 270061
rect 205725 270058 205791 270061
rect 100109 270056 205791 270058
rect 100109 270000 100114 270056
rect 100170 270000 205730 270056
rect 205786 270000 205791 270056
rect 100109 269998 205791 270000
rect 100109 269995 100175 269998
rect 205725 269995 205791 269998
rect 370037 270058 370103 270061
rect 537477 270058 537543 270061
rect 370037 270056 537543 270058
rect 370037 270000 370042 270056
rect 370098 270000 537482 270056
rect 537538 270000 537543 270056
rect 370037 269998 537543 270000
rect 370037 269995 370103 269998
rect 537477 269995 537543 269998
rect 93025 269922 93091 269925
rect 203057 269922 203123 269925
rect 93025 269920 203123 269922
rect 93025 269864 93030 269920
rect 93086 269864 203062 269920
rect 203118 269864 203123 269920
rect 93025 269862 203123 269864
rect 93025 269859 93091 269862
rect 203057 269859 203123 269862
rect 370865 269922 370931 269925
rect 539869 269922 539935 269925
rect 370865 269920 539935 269922
rect 370865 269864 370870 269920
rect 370926 269864 539874 269920
rect 539930 269864 539935 269920
rect 370865 269862 539935 269864
rect 370865 269859 370931 269862
rect 539869 269859 539935 269862
rect 85941 269786 86007 269789
rect 199929 269786 199995 269789
rect 85941 269784 199995 269786
rect 85941 269728 85946 269784
rect 86002 269728 199934 269784
rect 199990 269728 199995 269784
rect 85941 269726 199995 269728
rect 85941 269723 86007 269726
rect 199929 269723 199995 269726
rect 376661 269786 376727 269789
rect 555233 269786 555299 269789
rect 376661 269784 555299 269786
rect 376661 269728 376666 269784
rect 376722 269728 555238 269784
rect 555294 269728 555299 269784
rect 376661 269726 555299 269728
rect 376661 269723 376727 269726
rect 555233 269723 555299 269726
rect 84745 269650 84811 269653
rect 199009 269650 199075 269653
rect 84745 269648 199075 269650
rect 84745 269592 84750 269648
rect 84806 269592 199014 269648
rect 199070 269592 199075 269648
rect 84745 269590 199075 269592
rect 84745 269587 84811 269590
rect 199009 269587 199075 269590
rect 381997 269650 382063 269653
rect 569401 269650 569467 269653
rect 381997 269648 569467 269650
rect 381997 269592 382002 269648
rect 382058 269592 569406 269648
rect 569462 269592 569467 269648
rect 381997 269590 569467 269592
rect 381997 269587 382063 269590
rect 569401 269587 569467 269590
rect 78857 269514 78923 269517
rect 197721 269514 197787 269517
rect 78857 269512 197787 269514
rect 78857 269456 78862 269512
rect 78918 269456 197726 269512
rect 197782 269456 197787 269512
rect 78857 269454 197787 269456
rect 78857 269451 78923 269454
rect 197721 269451 197787 269454
rect 391381 269514 391447 269517
rect 594241 269514 594307 269517
rect 391381 269512 594307 269514
rect 391381 269456 391386 269512
rect 391442 269456 594246 269512
rect 594302 269456 594307 269512
rect 391381 269454 594307 269456
rect 391381 269451 391447 269454
rect 594241 269451 594307 269454
rect 77661 269378 77727 269381
rect 196801 269378 196867 269381
rect 77661 269376 196867 269378
rect 77661 269320 77666 269376
rect 77722 269320 196806 269376
rect 196862 269320 196867 269376
rect 77661 269318 196867 269320
rect 77661 269315 77727 269318
rect 196801 269315 196867 269318
rect 403433 269378 403499 269381
rect 626073 269378 626139 269381
rect 403433 269376 626139 269378
rect 403433 269320 403438 269376
rect 403494 269320 626078 269376
rect 626134 269320 626139 269376
rect 403433 269318 626139 269320
rect 403433 269315 403499 269318
rect 626073 269315 626139 269318
rect 76465 269242 76531 269245
rect 196341 269242 196407 269245
rect 76465 269240 196407 269242
rect 76465 269184 76470 269240
rect 76526 269184 196346 269240
rect 196402 269184 196407 269240
rect 76465 269182 196407 269184
rect 76465 269179 76531 269182
rect 196341 269179 196407 269182
rect 406101 269242 406167 269245
rect 633249 269242 633315 269245
rect 406101 269240 633315 269242
rect 406101 269184 406106 269240
rect 406162 269184 633254 269240
rect 633310 269184 633315 269240
rect 406101 269182 633315 269184
rect 406101 269179 406167 269182
rect 633249 269179 633315 269182
rect 71773 269106 71839 269109
rect 194593 269106 194659 269109
rect 71773 269104 194659 269106
rect 71773 269048 71778 269104
rect 71834 269048 194598 269104
rect 194654 269048 194659 269104
rect 71773 269046 194659 269048
rect 71773 269043 71839 269046
rect 194593 269043 194659 269046
rect 410977 269106 411043 269109
rect 646221 269106 646287 269109
rect 410977 269104 646287 269106
rect 410977 269048 410982 269104
rect 411038 269048 646226 269104
rect 646282 269048 646287 269104
rect 410977 269046 646287 269048
rect 410977 269043 411043 269046
rect 646221 269043 646287 269046
rect 128537 268970 128603 268973
rect 216397 268970 216463 268973
rect 128537 268968 216463 268970
rect 128537 268912 128542 268968
rect 128598 268912 216402 268968
rect 216458 268912 216463 268968
rect 128537 268910 216463 268912
rect 128537 268907 128603 268910
rect 216397 268907 216463 268910
rect 357525 268970 357591 268973
rect 504357 268970 504423 268973
rect 357525 268968 504423 268970
rect 357525 268912 357530 268968
rect 357586 268912 504362 268968
rect 504418 268912 504423 268968
rect 357525 268910 504423 268912
rect 357525 268907 357591 268910
rect 504357 268907 504423 268910
rect 146201 268834 146267 268837
rect 221733 268834 221799 268837
rect 146201 268832 221799 268834
rect 146201 268776 146206 268832
rect 146262 268776 221738 268832
rect 221794 268776 221799 268832
rect 146201 268774 221799 268776
rect 146201 268771 146267 268774
rect 221733 268771 221799 268774
rect 356605 268834 356671 268837
rect 501965 268834 502031 268837
rect 356605 268832 502031 268834
rect 356605 268776 356610 268832
rect 356666 268776 501970 268832
rect 502026 268776 502031 268832
rect 356605 268774 502031 268776
rect 356605 268771 356671 268774
rect 501965 268771 502031 268774
rect 150985 268698 151051 268701
rect 223941 268698 224007 268701
rect 150985 268696 224007 268698
rect 150985 268640 150990 268696
rect 151046 268640 223946 268696
rect 224002 268640 224007 268696
rect 150985 268638 224007 268640
rect 150985 268635 151051 268638
rect 223941 268635 224007 268638
rect 354857 268698 354923 268701
rect 497273 268698 497339 268701
rect 354857 268696 497339 268698
rect 354857 268640 354862 268696
rect 354918 268640 497278 268696
rect 497334 268640 497339 268696
rect 354857 268638 497339 268640
rect 354857 268635 354923 268638
rect 497273 268635 497339 268638
rect 158069 268562 158135 268565
rect 226609 268562 226675 268565
rect 158069 268560 226675 268562
rect 158069 268504 158074 268560
rect 158130 268504 226614 268560
rect 226670 268504 226675 268560
rect 158069 268502 226675 268504
rect 158069 268499 158135 268502
rect 226609 268499 226675 268502
rect 353937 268562 354003 268565
rect 494881 268562 494947 268565
rect 353937 268560 494947 268562
rect 353937 268504 353942 268560
rect 353998 268504 494886 268560
rect 494942 268504 494947 268560
rect 353937 268502 494947 268504
rect 353937 268499 354003 268502
rect 494881 268499 494947 268502
rect 676121 268562 676187 268565
rect 676262 268562 676322 268668
rect 676121 268560 676322 268562
rect 676121 268504 676126 268560
rect 676182 268504 676322 268560
rect 676121 268502 676322 268504
rect 676121 268499 676187 268502
rect 159265 268426 159331 268429
rect 227529 268426 227595 268429
rect 159265 268424 227595 268426
rect 159265 268368 159270 268424
rect 159326 268368 227534 268424
rect 227590 268368 227595 268424
rect 159265 268366 227595 268368
rect 159265 268363 159331 268366
rect 227529 268363 227595 268366
rect 352189 268426 352255 268429
rect 490189 268426 490255 268429
rect 352189 268424 490255 268426
rect 352189 268368 352194 268424
rect 352250 268368 490194 268424
rect 490250 268368 490255 268424
rect 352189 268366 490255 268368
rect 352189 268363 352255 268366
rect 490189 268363 490255 268366
rect 195973 268290 196039 268293
rect 202137 268290 202203 268293
rect 195973 268288 202203 268290
rect 195973 268232 195978 268288
rect 196034 268232 202142 268288
rect 202198 268232 202203 268288
rect 195973 268230 202203 268232
rect 195973 268227 196039 268230
rect 202137 268227 202203 268230
rect 365989 268290 366055 268293
rect 372061 268290 372127 268293
rect 365989 268288 372127 268290
rect 365989 268232 365994 268288
rect 366050 268232 372066 268288
rect 372122 268232 372127 268288
rect 365989 268230 372127 268232
rect 365989 268227 366055 268230
rect 372061 268227 372127 268230
rect 676262 268157 676322 268260
rect 676213 268152 676322 268157
rect 676213 268096 676218 268152
rect 676274 268096 676322 268152
rect 676213 268094 676322 268096
rect 676213 268091 676279 268094
rect 676029 267882 676095 267885
rect 676029 267880 676292 267882
rect 676029 267824 676034 267880
rect 676090 267824 676292 267880
rect 676029 267822 676292 267824
rect 676029 267819 676095 267822
rect 405641 267746 405707 267749
rect 441797 267746 441863 267749
rect 405641 267744 441863 267746
rect 405641 267688 405646 267744
rect 405702 267688 441802 267744
rect 441858 267688 441863 267744
rect 405641 267686 441863 267688
rect 405641 267683 405707 267686
rect 441797 267683 441863 267686
rect 678973 267746 679039 267749
rect 678973 267744 679082 267746
rect 678973 267688 678978 267744
rect 679034 267688 679082 267744
rect 678973 267683 679082 267688
rect 402973 267610 403039 267613
rect 455965 267610 456031 267613
rect 402973 267608 456031 267610
rect 402973 267552 402978 267608
rect 403034 267552 455970 267608
rect 456026 267552 456031 267608
rect 402973 267550 456031 267552
rect 402973 267547 403039 267550
rect 455965 267547 456031 267550
rect 397637 267474 397703 267477
rect 472525 267474 472591 267477
rect 397637 267472 472591 267474
rect 397637 267416 397642 267472
rect 397698 267416 472530 267472
rect 472586 267416 472591 267472
rect 679022 267444 679082 267683
rect 397637 267414 472591 267416
rect 397637 267411 397703 267414
rect 472525 267411 472591 267414
rect 406929 267338 406995 267341
rect 485037 267338 485103 267341
rect 406929 267336 485103 267338
rect 406929 267280 406934 267336
rect 406990 267280 485042 267336
rect 485098 267280 485103 267336
rect 406929 267278 485103 267280
rect 406929 267275 406995 267278
rect 485037 267275 485103 267278
rect 386965 267202 387031 267205
rect 582373 267202 582439 267205
rect 386965 267200 582439 267202
rect 386965 267144 386970 267200
rect 387026 267144 582378 267200
rect 582434 267144 582439 267200
rect 386965 267142 582439 267144
rect 386965 267139 387031 267142
rect 582373 267139 582439 267142
rect 389633 267066 389699 267069
rect 589457 267066 589523 267069
rect 389633 267064 589523 267066
rect 389633 267008 389638 267064
rect 389694 267008 589462 267064
rect 589518 267008 589523 267064
rect 389633 267006 589523 267008
rect 389633 267003 389699 267006
rect 589457 267003 589523 267006
rect 675661 267066 675727 267069
rect 675661 267064 676292 267066
rect 675661 267008 675666 267064
rect 675722 267008 676292 267064
rect 675661 267006 676292 267008
rect 675661 267003 675727 267006
rect 390461 266930 390527 266933
rect 591849 266930 591915 266933
rect 390461 266928 591915 266930
rect 390461 266872 390466 266928
rect 390522 266872 591854 266928
rect 591910 266872 591915 266928
rect 390461 266870 591915 266872
rect 390461 266867 390527 266870
rect 591849 266867 591915 266870
rect 391841 266794 391907 266797
rect 595345 266794 595411 266797
rect 391841 266792 595411 266794
rect 391841 266736 391846 266792
rect 391902 266736 595350 266792
rect 595406 266736 595411 266792
rect 391841 266734 595411 266736
rect 391841 266731 391907 266734
rect 595345 266731 595411 266734
rect 393129 266658 393195 266661
rect 598933 266658 598999 266661
rect 393129 266656 598999 266658
rect 393129 266600 393134 266656
rect 393190 266600 598938 266656
rect 598994 266600 598999 266656
rect 393129 266598 598999 266600
rect 393129 266595 393195 266598
rect 598933 266595 598999 266598
rect 676029 266658 676095 266661
rect 676029 266656 676292 266658
rect 676029 266600 676034 266656
rect 676090 266600 676292 266656
rect 676029 266598 676292 266600
rect 676029 266595 676095 266598
rect 394509 266522 394575 266525
rect 602429 266522 602495 266525
rect 394509 266520 602495 266522
rect 394509 266464 394514 266520
rect 394570 266464 602434 266520
rect 602490 266464 602495 266520
rect 394509 266462 602495 266464
rect 394509 266459 394575 266462
rect 602429 266459 602495 266462
rect 676029 266250 676095 266253
rect 676029 266248 676292 266250
rect 676029 266192 676034 266248
rect 676090 266192 676292 266248
rect 676029 266190 676292 266192
rect 676029 266187 676095 266190
rect 679065 266114 679131 266117
rect 679022 266112 679131 266114
rect 679022 266056 679070 266112
rect 679126 266056 679131 266112
rect 679022 266051 679131 266056
rect 679022 265812 679082 266051
rect 675753 265434 675819 265437
rect 675753 265432 676292 265434
rect 675753 265376 675758 265432
rect 675814 265376 676292 265432
rect 675753 265374 676292 265376
rect 675753 265371 675819 265374
rect 679157 265298 679223 265301
rect 679157 265296 679266 265298
rect 679157 265240 679162 265296
rect 679218 265240 679266 265296
rect 679157 265235 679266 265240
rect 679206 264996 679266 265235
rect 675150 264618 675156 264620
rect 675146 264558 675156 264618
rect 675150 264556 675156 264558
rect 675220 264618 675226 264620
rect 675220 264558 676292 264618
rect 675220 264556 675226 264558
rect 676029 264210 676095 264213
rect 676029 264208 676292 264210
rect 676029 264152 676034 264208
rect 676090 264152 676292 264208
rect 676029 264150 676292 264152
rect 676029 264147 676095 264150
rect 676121 263666 676187 263669
rect 676262 263666 676322 263772
rect 676121 263664 676322 263666
rect 676121 263608 676126 263664
rect 676182 263608 676322 263664
rect 676121 263606 676322 263608
rect 676121 263603 676187 263606
rect 675845 263394 675911 263397
rect 675845 263392 676292 263394
rect 675845 263336 675850 263392
rect 675906 263336 676292 263392
rect 675845 263334 676292 263336
rect 675845 263331 675911 263334
rect 676029 262986 676095 262989
rect 676029 262984 676292 262986
rect 676029 262928 676034 262984
rect 676090 262928 676292 262984
rect 676029 262926 676292 262928
rect 676029 262923 676095 262926
rect 676121 262442 676187 262445
rect 676262 262442 676322 262548
rect 676121 262440 676322 262442
rect 676121 262384 676126 262440
rect 676182 262384 676322 262440
rect 676121 262382 676322 262384
rect 676121 262379 676187 262382
rect 676029 262170 676095 262173
rect 676029 262168 676292 262170
rect 676029 262112 676034 262168
rect 676090 262112 676292 262168
rect 676029 262110 676292 262112
rect 676029 262107 676095 262110
rect 676029 261762 676095 261765
rect 676029 261760 676292 261762
rect 676029 261704 676034 261760
rect 676090 261704 676292 261760
rect 676029 261702 676292 261704
rect 676029 261699 676095 261702
rect 676121 261218 676187 261221
rect 676262 261218 676322 261324
rect 676121 261216 676322 261218
rect 676121 261160 676126 261216
rect 676182 261160 676322 261216
rect 676121 261158 676322 261160
rect 676121 261155 676187 261158
rect 675937 260946 676003 260949
rect 675937 260944 676292 260946
rect 675937 260888 675942 260944
rect 675998 260888 676292 260944
rect 675937 260886 676292 260888
rect 675937 260883 676003 260886
rect 675661 260538 675727 260541
rect 675661 260536 676292 260538
rect 675661 260480 675666 260536
rect 675722 260480 676292 260536
rect 675661 260478 676292 260480
rect 675661 260475 675727 260478
rect 675661 260130 675727 260133
rect 675661 260128 676292 260130
rect 675661 260072 675666 260128
rect 675722 260072 676292 260128
rect 675661 260070 676292 260072
rect 675661 260067 675727 260070
rect 676121 259586 676187 259589
rect 676262 259586 676322 259692
rect 676121 259584 676322 259586
rect 676121 259528 676126 259584
rect 676182 259528 676322 259584
rect 676121 259526 676322 259528
rect 676121 259523 676187 259526
rect 676029 259314 676095 259317
rect 676029 259312 676292 259314
rect 676029 259256 676034 259312
rect 676090 259256 676292 259312
rect 676029 259254 676292 259256
rect 676029 259251 676095 259254
rect 676029 258906 676095 258909
rect 676029 258904 676292 258906
rect 676029 258848 676034 258904
rect 676090 258848 676292 258904
rect 676029 258846 676292 258848
rect 676029 258843 676095 258846
rect 184933 258634 184999 258637
rect 184933 258632 191820 258634
rect 184933 258576 184938 258632
rect 184994 258576 191820 258632
rect 184933 258574 191820 258576
rect 184933 258571 184999 258574
rect 679022 258365 679082 258468
rect 678973 258360 679082 258365
rect 678973 258304 678978 258360
rect 679034 258304 679082 258360
rect 678973 258302 679082 258304
rect 678973 258299 679039 258302
rect 41781 258090 41847 258093
rect 41492 258088 41847 258090
rect 41492 258032 41786 258088
rect 41842 258032 41847 258088
rect 41492 258030 41847 258032
rect 41781 258027 41847 258030
rect 41505 257954 41571 257957
rect 41462 257952 41571 257954
rect 41462 257896 41510 257952
rect 41566 257896 41571 257952
rect 41462 257891 41571 257896
rect 41462 257652 41522 257891
rect 684542 257652 684602 258060
rect 41505 257546 41571 257549
rect 41462 257544 41571 257546
rect 41462 257488 41510 257544
rect 41566 257488 41571 257544
rect 41462 257483 41571 257488
rect 678973 257546 679039 257549
rect 678973 257544 679082 257546
rect 678973 257488 678978 257544
rect 679034 257488 679082 257544
rect 678973 257483 679082 257488
rect 41462 257244 41522 257483
rect 679022 257244 679082 257483
rect 44589 256914 44659 256919
rect 41534 256854 44594 256914
rect 44654 256854 44668 256914
rect 44589 256849 44659 256854
rect 44589 256532 44659 256535
rect 41550 256530 44668 256532
rect 41550 256472 44594 256530
rect 44589 256470 44594 256472
rect 44654 256472 44668 256530
rect 44654 256470 44659 256472
rect 44589 256465 44659 256470
rect 43713 256050 43779 256053
rect 41492 256048 43779 256050
rect 41492 255992 43718 256048
rect 43774 255992 43779 256048
rect 41492 255990 43779 255992
rect 43713 255987 43779 255990
rect 42241 255642 42307 255645
rect 41492 255640 42307 255642
rect 41492 255584 42246 255640
rect 42302 255584 42307 255640
rect 41492 255582 42307 255584
rect 42241 255579 42307 255582
rect 44681 255280 44751 255283
rect 41564 255278 44758 255280
rect 41564 255220 44686 255278
rect 44681 255218 44686 255220
rect 44746 255220 44758 255278
rect 44746 255218 44751 255220
rect 44681 255213 44751 255218
rect 44681 254868 44751 254873
rect 44681 254866 44686 254868
rect 41572 254808 44686 254866
rect 44746 254866 44751 254868
rect 44746 254808 44758 254866
rect 41572 254806 44758 254808
rect 44681 254803 44751 254806
rect 44773 254488 44843 254493
rect 41576 254428 44778 254488
rect 44838 254428 44864 254488
rect 44773 254423 44843 254428
rect 44773 254076 44843 254081
rect 44773 254070 44778 254076
rect 41568 254016 44778 254070
rect 44838 254070 44843 254076
rect 44838 254016 44864 254070
rect 41568 254010 44864 254016
rect 42333 253602 42399 253605
rect 41492 253600 42399 253602
rect 41492 253544 42338 253600
rect 42394 253544 42399 253600
rect 41492 253542 42399 253544
rect 42333 253539 42399 253542
rect 43805 253194 43871 253197
rect 41492 253192 43871 253194
rect 41492 253136 43810 253192
rect 43866 253136 43871 253192
rect 41492 253134 43871 253136
rect 43805 253131 43871 253134
rect 416773 252786 416839 252789
rect 412436 252784 416839 252786
rect 41462 252650 41522 252756
rect 412436 252728 416778 252784
rect 416834 252728 416839 252784
rect 412436 252726 416839 252728
rect 416773 252723 416839 252726
rect 41638 252650 41644 252652
rect 41462 252590 41644 252650
rect 41638 252588 41644 252590
rect 41708 252588 41714 252652
rect 43253 252378 43319 252381
rect 41492 252376 43319 252378
rect 41492 252320 43258 252376
rect 43314 252320 43319 252376
rect 41492 252318 43319 252320
rect 43253 252315 43319 252318
rect 43529 251970 43595 251973
rect 41492 251968 43595 251970
rect 41492 251912 43534 251968
rect 43590 251912 43595 251968
rect 41492 251910 43595 251912
rect 43529 251907 43595 251910
rect 30054 251429 30114 251532
rect 30054 251424 30163 251429
rect 30054 251368 30102 251424
rect 30158 251368 30163 251424
rect 30054 251366 30163 251368
rect 30097 251363 30163 251366
rect 43621 251154 43687 251157
rect 41492 251152 43687 251154
rect 41492 251096 43626 251152
rect 43682 251096 43687 251152
rect 41492 251094 43687 251096
rect 43621 251091 43687 251094
rect 43713 250746 43779 250749
rect 41492 250744 43779 250746
rect 41492 250688 43718 250744
rect 43774 250688 43779 250744
rect 41492 250686 43779 250688
rect 43713 250683 43779 250686
rect 43989 250338 44055 250341
rect 41492 250336 44055 250338
rect 41492 250280 43994 250336
rect 44050 250280 44055 250336
rect 41492 250278 44055 250280
rect 43989 250275 44055 250278
rect 42701 249930 42767 249933
rect 41492 249928 42767 249930
rect 41492 249872 42706 249928
rect 42762 249872 42767 249928
rect 41492 249870 42767 249872
rect 42701 249867 42767 249870
rect 43069 249522 43135 249525
rect 416773 249522 416839 249525
rect 41492 249520 43135 249522
rect 41492 249464 43074 249520
rect 43130 249464 43135 249520
rect 41492 249462 43135 249464
rect 412436 249520 416839 249522
rect 412436 249464 416778 249520
rect 416834 249464 416839 249520
rect 412436 249462 416839 249464
rect 43069 249459 43135 249462
rect 416773 249459 416839 249462
rect 38150 248981 38210 249084
rect 38101 248976 38210 248981
rect 38101 248920 38106 248976
rect 38162 248920 38210 248976
rect 38101 248918 38210 248920
rect 38101 248915 38167 248918
rect 38150 248573 38210 248676
rect 38150 248568 38259 248573
rect 38150 248512 38198 248568
rect 38254 248512 38259 248568
rect 38150 248510 38259 248512
rect 38193 248507 38259 248510
rect 41462 248165 41522 248268
rect 41462 248160 41571 248165
rect 41462 248104 41510 248160
rect 41566 248104 41571 248160
rect 41462 248102 41571 248104
rect 41505 248099 41571 248102
rect 184933 248026 184999 248029
rect 184933 248024 191820 248026
rect 184933 247968 184938 248024
rect 184994 247968 191820 248024
rect 184933 247966 191820 247968
rect 184933 247963 184999 247966
rect 41462 247757 41522 247860
rect 41413 247752 41522 247757
rect 41413 247696 41418 247752
rect 41474 247696 41522 247752
rect 41413 247694 41522 247696
rect 41413 247691 41479 247694
rect 41462 247349 41522 247452
rect 41413 247344 41522 247349
rect 41413 247288 41418 247344
rect 41474 247288 41522 247344
rect 41413 247286 41522 247288
rect 41413 247283 41479 247286
rect 41462 246533 41522 246636
rect 41462 246528 41571 246533
rect 41462 246472 41510 246528
rect 41566 246472 41571 246528
rect 41462 246470 41571 246472
rect 41505 246467 41571 246470
rect 416773 246394 416839 246397
rect 412436 246392 416839 246394
rect 412436 246336 416778 246392
rect 416834 246336 416839 246392
rect 412436 246334 416839 246336
rect 416773 246331 416839 246334
rect 418061 243130 418127 243133
rect 412436 243128 418127 243130
rect 412436 243072 418066 243128
rect 418122 243072 418127 243128
rect 412436 243070 418127 243072
rect 418061 243067 418127 243070
rect 418153 240002 418219 240005
rect 412436 240000 418219 240002
rect 412436 239944 418158 240000
rect 418214 239944 418219 240000
rect 412436 239942 418219 239944
rect 418153 239939 418219 239942
rect 184933 237418 184999 237421
rect 184933 237416 191820 237418
rect 184933 237360 184938 237416
rect 184994 237360 191820 237416
rect 184933 237358 191820 237360
rect 184933 237355 184999 237358
rect 418429 236738 418495 236741
rect 412436 236736 418495 236738
rect 412436 236680 418434 236736
rect 418490 236680 418495 236736
rect 412436 236678 418495 236680
rect 418429 236675 418495 236678
rect 418521 233610 418587 233613
rect 412436 233608 418587 233610
rect 412436 233552 418526 233608
rect 418582 233552 418587 233608
rect 412436 233550 418587 233552
rect 418521 233547 418587 233550
rect 84653 228986 84719 228989
rect 206185 228986 206251 228989
rect 84653 228984 206251 228986
rect 84653 228928 84658 228984
rect 84714 228928 206190 228984
rect 206246 228928 206251 228984
rect 84653 228926 206251 228928
rect 84653 228923 84719 228926
rect 206185 228923 206251 228926
rect 207013 228986 207079 228989
rect 210785 228986 210851 228989
rect 207013 228984 210851 228986
rect 207013 228928 207018 228984
rect 207074 228928 210790 228984
rect 210846 228928 210851 228984
rect 207013 228926 210851 228928
rect 207013 228923 207079 228926
rect 210785 228923 210851 228926
rect 384757 228986 384823 228989
rect 507393 228986 507459 228989
rect 384757 228984 507459 228986
rect 384757 228928 384762 228984
rect 384818 228928 507398 228984
rect 507454 228928 507459 228984
rect 384757 228926 507459 228928
rect 384757 228923 384823 228926
rect 507393 228923 507459 228926
rect 88057 228850 88123 228853
rect 207565 228850 207631 228853
rect 88057 228848 207631 228850
rect 88057 228792 88062 228848
rect 88118 228792 207570 228848
rect 207626 228792 207631 228848
rect 88057 228790 207631 228792
rect 88057 228787 88123 228790
rect 207565 228787 207631 228790
rect 245653 228850 245719 228853
rect 261385 228850 261451 228853
rect 245653 228848 261451 228850
rect 245653 228792 245658 228848
rect 245714 228792 261390 228848
rect 261446 228792 261451 228848
rect 245653 228790 261451 228792
rect 245653 228787 245719 228790
rect 261385 228787 261451 228790
rect 382641 228850 382707 228853
rect 503805 228850 503871 228853
rect 382641 228848 503871 228850
rect 382641 228792 382646 228848
rect 382702 228792 503810 228848
rect 503866 228792 503871 228848
rect 382641 228790 503871 228792
rect 382641 228787 382707 228790
rect 503805 228787 503871 228790
rect 86309 228714 86375 228717
rect 207197 228714 207263 228717
rect 86309 228712 207263 228714
rect 86309 228656 86314 228712
rect 86370 228656 207202 228712
rect 207258 228656 207263 228712
rect 86309 228654 207263 228656
rect 86309 228651 86375 228654
rect 207197 228651 207263 228654
rect 386873 228714 386939 228717
rect 512177 228714 512243 228717
rect 386873 228712 512243 228714
rect 386873 228656 386878 228712
rect 386934 228656 512182 228712
rect 512238 228656 512243 228712
rect 386873 228654 512243 228656
rect 386873 228651 386939 228654
rect 512177 228651 512243 228654
rect 82721 228578 82787 228581
rect 205817 228578 205883 228581
rect 82721 228576 205883 228578
rect 82721 228520 82726 228576
rect 82782 228520 205822 228576
rect 205878 228520 205883 228576
rect 82721 228518 205883 228520
rect 82721 228515 82787 228518
rect 205817 228515 205883 228518
rect 237005 228578 237071 228581
rect 259637 228578 259703 228581
rect 237005 228576 259703 228578
rect 237005 228520 237010 228576
rect 237066 228520 259642 228576
rect 259698 228520 259703 228576
rect 237005 228518 259703 228520
rect 237005 228515 237071 228518
rect 259637 228515 259703 228518
rect 390093 228578 390159 228581
rect 518985 228578 519051 228581
rect 390093 228576 519051 228578
rect 390093 228520 390098 228576
rect 390154 228520 518990 228576
rect 519046 228520 519051 228576
rect 390093 228518 519051 228520
rect 390093 228515 390159 228518
rect 518985 228515 519051 228518
rect 77937 228442 78003 228445
rect 203333 228442 203399 228445
rect 77937 228440 203399 228442
rect 77937 228384 77942 228440
rect 77998 228384 203338 228440
rect 203394 228384 203399 228440
rect 77937 228382 203399 228384
rect 77937 228379 78003 228382
rect 203333 228379 203399 228382
rect 236729 228442 236795 228445
rect 262489 228442 262555 228445
rect 236729 228440 262555 228442
rect 236729 228384 236734 228440
rect 236790 228384 262494 228440
rect 262550 228384 262555 228440
rect 236729 228382 262555 228384
rect 236729 228379 236795 228382
rect 262489 228379 262555 228382
rect 392209 228442 392275 228445
rect 525057 228442 525123 228445
rect 392209 228440 525123 228442
rect 392209 228384 392214 228440
rect 392270 228384 525062 228440
rect 525118 228384 525123 228440
rect 392209 228382 525123 228384
rect 392209 228379 392275 228382
rect 525057 228379 525123 228382
rect 76281 228306 76347 228309
rect 202965 228306 203031 228309
rect 76281 228304 203031 228306
rect 76281 228248 76286 228304
rect 76342 228248 202970 228304
rect 203026 228248 203031 228304
rect 76281 228246 203031 228248
rect 76281 228243 76347 228246
rect 202965 228243 203031 228246
rect 225965 228306 226031 228309
rect 266077 228306 266143 228309
rect 225965 228304 266143 228306
rect 225965 228248 225970 228304
rect 226026 228248 266082 228304
rect 266138 228248 266143 228304
rect 225965 228246 266143 228248
rect 225965 228243 226031 228246
rect 266077 228243 266143 228246
rect 394417 228306 394483 228309
rect 530117 228306 530183 228309
rect 394417 228304 530183 228306
rect 394417 228248 394422 228304
rect 394478 228248 530122 228304
rect 530178 228248 530183 228304
rect 394417 228246 530183 228248
rect 394417 228243 394483 228246
rect 530117 228243 530183 228246
rect 71221 228170 71287 228173
rect 200481 228170 200547 228173
rect 71221 228168 200547 228170
rect 71221 228112 71226 228168
rect 71282 228112 200486 228168
rect 200542 228112 200547 228168
rect 71221 228110 200547 228112
rect 71221 228107 71287 228110
rect 200481 228107 200547 228110
rect 219249 228170 219315 228173
rect 263225 228170 263291 228173
rect 219249 228168 263291 228170
rect 219249 228112 219254 228168
rect 219310 228112 263230 228168
rect 263286 228112 263291 228168
rect 219249 228110 263291 228112
rect 219249 228107 219315 228110
rect 263225 228107 263291 228110
rect 396533 228170 396599 228173
rect 534901 228170 534967 228173
rect 396533 228168 534967 228170
rect 396533 228112 396538 228168
rect 396594 228112 534906 228168
rect 534962 228112 534967 228168
rect 396533 228110 534967 228112
rect 396533 228107 396599 228110
rect 534901 228107 534967 228110
rect 64505 228034 64571 228037
rect 197629 228034 197695 228037
rect 64505 228032 197695 228034
rect 64505 227976 64510 228032
rect 64566 227976 197634 228032
rect 197690 227976 197695 228032
rect 64505 227974 197695 227976
rect 64505 227971 64571 227974
rect 197629 227971 197695 227974
rect 220721 228034 220787 228037
rect 264237 228034 264303 228037
rect 220721 228032 264303 228034
rect 220721 227976 220726 228032
rect 220782 227976 264242 228032
rect 264298 227976 264303 228032
rect 220721 227974 264303 227976
rect 220721 227971 220787 227974
rect 264237 227971 264303 227974
rect 398649 228034 398715 228037
rect 538305 228034 538371 228037
rect 398649 228032 538371 228034
rect 398649 227976 398654 228032
rect 398710 227976 538310 228032
rect 538366 227976 538371 228032
rect 398649 227974 538371 227976
rect 398649 227971 398715 227974
rect 538305 227971 538371 227974
rect 62665 227898 62731 227901
rect 197261 227898 197327 227901
rect 62665 227896 197327 227898
rect 62665 227840 62670 227896
rect 62726 227840 197266 227896
rect 197322 227840 197327 227896
rect 62665 227838 197327 227840
rect 62665 227835 62731 227838
rect 197261 227835 197327 227838
rect 217593 227898 217659 227901
rect 262857 227898 262923 227901
rect 217593 227896 262923 227898
rect 217593 227840 217598 227896
rect 217654 227840 262862 227896
rect 262918 227840 262923 227896
rect 217593 227838 262923 227840
rect 217593 227835 217659 227838
rect 262857 227835 262923 227838
rect 399753 227898 399819 227901
rect 542721 227898 542787 227901
rect 399753 227896 542787 227898
rect 399753 227840 399758 227896
rect 399814 227840 542726 227896
rect 542782 227840 542787 227896
rect 399753 227838 542787 227840
rect 399753 227835 399819 227838
rect 542721 227835 542787 227838
rect 57605 227762 57671 227765
rect 194777 227762 194843 227765
rect 57605 227760 194843 227762
rect 57605 227704 57610 227760
rect 57666 227704 194782 227760
rect 194838 227704 194843 227760
rect 57605 227702 194843 227704
rect 57605 227699 57671 227702
rect 194777 227699 194843 227702
rect 212349 227762 212415 227765
rect 260373 227762 260439 227765
rect 212349 227760 260439 227762
rect 212349 227704 212354 227760
rect 212410 227704 260378 227760
rect 260434 227704 260439 227760
rect 212349 227702 260439 227704
rect 212349 227699 212415 227702
rect 260373 227699 260439 227702
rect 403985 227762 404051 227765
rect 552565 227762 552631 227765
rect 403985 227760 552631 227762
rect 403985 227704 403990 227760
rect 404046 227704 552570 227760
rect 552626 227704 552631 227760
rect 403985 227702 552631 227704
rect 403985 227699 404051 227702
rect 552565 227699 552631 227702
rect 56041 227626 56107 227629
rect 194409 227626 194475 227629
rect 56041 227624 194475 227626
rect 56041 227568 56046 227624
rect 56102 227568 194414 227624
rect 194470 227568 194475 227624
rect 56041 227566 194475 227568
rect 56041 227563 56107 227566
rect 194409 227563 194475 227566
rect 210785 227626 210851 227629
rect 260005 227626 260071 227629
rect 210785 227624 260071 227626
rect 210785 227568 210790 227624
rect 210846 227568 260010 227624
rect 260066 227568 260071 227624
rect 210785 227566 260071 227568
rect 210785 227563 210851 227566
rect 260005 227563 260071 227566
rect 411161 227626 411227 227629
rect 569309 227626 569375 227629
rect 411161 227624 569375 227626
rect 411161 227568 411166 227624
rect 411222 227568 569314 227624
rect 569370 227568 569375 227624
rect 411161 227566 569375 227568
rect 411161 227563 411227 227566
rect 569309 227563 569375 227566
rect 93025 227490 93091 227493
rect 210049 227490 210115 227493
rect 93025 227488 210115 227490
rect 93025 227432 93030 227488
rect 93086 227432 210054 227488
rect 210110 227432 210115 227488
rect 93025 227430 210115 227432
rect 93025 227427 93091 227430
rect 210049 227427 210115 227430
rect 379789 227490 379855 227493
rect 495341 227490 495407 227493
rect 379789 227488 495407 227490
rect 379789 227432 379794 227488
rect 379850 227432 495346 227488
rect 495402 227432 495407 227488
rect 379789 227430 495407 227432
rect 379789 227427 379855 227430
rect 495341 227427 495407 227430
rect 94773 227354 94839 227357
rect 210417 227354 210483 227357
rect 94773 227352 210483 227354
rect 94773 227296 94778 227352
rect 94834 227296 210422 227352
rect 210478 227296 210483 227352
rect 94773 227294 210483 227296
rect 94773 227291 94839 227294
rect 210417 227291 210483 227294
rect 380157 227354 380223 227357
rect 496169 227354 496235 227357
rect 380157 227352 496235 227354
rect 380157 227296 380162 227352
rect 380218 227296 496174 227352
rect 496230 227296 496235 227352
rect 380157 227294 496235 227296
rect 380157 227291 380223 227294
rect 496169 227291 496235 227294
rect 101489 227218 101555 227221
rect 213269 227218 213335 227221
rect 101489 227216 213335 227218
rect 101489 227160 101494 227216
rect 101550 227160 213274 227216
rect 213330 227160 213335 227216
rect 101489 227158 213335 227160
rect 101489 227155 101555 227158
rect 213269 227155 213335 227158
rect 377305 227218 377371 227221
rect 489729 227218 489795 227221
rect 377305 227216 489795 227218
rect 377305 227160 377310 227216
rect 377366 227160 489734 227216
rect 489790 227160 489795 227216
rect 377305 227158 489795 227160
rect 377305 227155 377371 227158
rect 489729 227155 489795 227158
rect 99833 227082 99899 227085
rect 212901 227082 212967 227085
rect 99833 227080 212967 227082
rect 99833 227024 99838 227080
rect 99894 227024 212906 227080
rect 212962 227024 212967 227080
rect 99833 227022 212967 227024
rect 99833 227019 99899 227022
rect 212901 227019 212967 227022
rect 259177 227082 259243 227085
rect 261753 227082 261819 227085
rect 259177 227080 261819 227082
rect 259177 227024 259182 227080
rect 259238 227024 261758 227080
rect 261814 227024 261819 227080
rect 259177 227022 261819 227024
rect 259177 227019 259243 227022
rect 261753 227019 261819 227022
rect 376937 227082 377003 227085
rect 488901 227082 488967 227085
rect 376937 227080 488967 227082
rect 376937 227024 376942 227080
rect 376998 227024 488906 227080
rect 488962 227024 488967 227080
rect 376937 227022 488967 227024
rect 376937 227019 377003 227022
rect 488901 227019 488967 227022
rect 106549 226946 106615 226949
rect 215753 226946 215819 226949
rect 106549 226944 215819 226946
rect 106549 226888 106554 226944
rect 106610 226888 215758 226944
rect 215814 226888 215819 226944
rect 106549 226886 215819 226888
rect 106549 226883 106615 226886
rect 215753 226883 215819 226886
rect 113081 226810 113147 226813
rect 218605 226810 218671 226813
rect 113081 226808 218671 226810
rect 113081 226752 113086 226808
rect 113142 226752 218610 226808
rect 218666 226752 218671 226808
rect 113081 226750 218671 226752
rect 113081 226747 113147 226750
rect 218605 226747 218671 226750
rect 201677 226538 201743 226541
rect 208669 226538 208735 226541
rect 201677 226536 208735 226538
rect 201677 226480 201682 226536
rect 201738 226480 208674 226536
rect 208730 226480 208735 226536
rect 201677 226478 208735 226480
rect 201677 226475 201743 226478
rect 208669 226475 208735 226478
rect 109033 226266 109099 226269
rect 215385 226266 215451 226269
rect 109033 226264 215451 226266
rect 109033 226208 109038 226264
rect 109094 226208 215390 226264
rect 215446 226208 215451 226264
rect 109033 226206 215451 226208
rect 109033 226203 109099 226206
rect 215385 226203 215451 226206
rect 397361 226266 397427 226269
rect 513465 226266 513531 226269
rect 397361 226264 513531 226266
rect 397361 226208 397366 226264
rect 397422 226208 513470 226264
rect 513526 226208 513531 226264
rect 397361 226206 513531 226208
rect 397361 226203 397427 226206
rect 513465 226203 513531 226206
rect 103973 226130 104039 226133
rect 213637 226130 213703 226133
rect 103973 226128 213703 226130
rect 103973 226072 103978 226128
rect 104034 226072 213642 226128
rect 213698 226072 213703 226128
rect 103973 226070 213703 226072
rect 103973 226067 104039 226070
rect 213637 226067 213703 226070
rect 389357 226130 389423 226133
rect 518709 226130 518775 226133
rect 389357 226128 518775 226130
rect 389357 226072 389362 226128
rect 389418 226072 518714 226128
rect 518770 226072 518775 226128
rect 389357 226070 518775 226072
rect 389357 226067 389423 226070
rect 518709 226067 518775 226070
rect 41638 225932 41644 225996
rect 41708 225994 41714 225996
rect 41781 225994 41847 225997
rect 41708 225992 41847 225994
rect 41708 225936 41786 225992
rect 41842 225936 41847 225992
rect 41708 225934 41847 225936
rect 41708 225932 41714 225934
rect 41781 225931 41847 225934
rect 98913 225994 98979 225997
rect 211153 225994 211219 225997
rect 98913 225992 211219 225994
rect 98913 225936 98918 225992
rect 98974 225936 211158 225992
rect 211214 225936 211219 225992
rect 98913 225934 211219 225936
rect 98913 225931 98979 225934
rect 211153 225931 211219 225934
rect 390461 225994 390527 225997
rect 520825 225994 520891 225997
rect 390461 225992 520891 225994
rect 390461 225936 390466 225992
rect 390522 225936 520830 225992
rect 520886 225936 520891 225992
rect 390461 225934 520891 225936
rect 390461 225931 390527 225934
rect 520825 225931 520891 225934
rect 102041 225858 102107 225861
rect 212533 225858 212599 225861
rect 102041 225856 212599 225858
rect 102041 225800 102046 225856
rect 102102 225800 212538 225856
rect 212594 225800 212599 225856
rect 102041 225798 212599 225800
rect 102041 225795 102107 225798
rect 212533 225795 212599 225798
rect 391565 225858 391631 225861
rect 523401 225858 523467 225861
rect 391565 225856 523467 225858
rect 391565 225800 391570 225856
rect 391626 225800 523406 225856
rect 523462 225800 523467 225856
rect 391565 225798 523467 225800
rect 391565 225795 391631 225798
rect 523401 225795 523467 225798
rect 83825 225722 83891 225725
rect 205081 225722 205147 225725
rect 83825 225720 205147 225722
rect 83825 225664 83830 225720
rect 83886 225664 205086 225720
rect 205142 225664 205147 225720
rect 83825 225662 205147 225664
rect 83825 225659 83891 225662
rect 205081 225659 205147 225662
rect 392577 225722 392643 225725
rect 525793 225722 525859 225725
rect 392577 225720 525859 225722
rect 392577 225664 392582 225720
rect 392638 225664 525798 225720
rect 525854 225664 525859 225720
rect 392577 225662 525859 225664
rect 392577 225659 392643 225662
rect 525793 225659 525859 225662
rect 80421 225586 80487 225589
rect 203701 225586 203767 225589
rect 80421 225584 203767 225586
rect 80421 225528 80426 225584
rect 80482 225528 203706 225584
rect 203762 225528 203767 225584
rect 80421 225526 203767 225528
rect 80421 225523 80487 225526
rect 203701 225523 203767 225526
rect 394785 225586 394851 225589
rect 530669 225586 530735 225589
rect 394785 225584 530735 225586
rect 394785 225528 394790 225584
rect 394846 225528 530674 225584
rect 530730 225528 530735 225584
rect 394785 225526 530735 225528
rect 394785 225523 394851 225526
rect 530669 225523 530735 225526
rect 77109 225450 77175 225453
rect 202229 225450 202295 225453
rect 77109 225448 202295 225450
rect 77109 225392 77114 225448
rect 77170 225392 202234 225448
rect 202290 225392 202295 225448
rect 77109 225390 202295 225392
rect 77109 225387 77175 225390
rect 202229 225387 202295 225390
rect 397913 225450 397979 225453
rect 538857 225450 538923 225453
rect 397913 225448 538923 225450
rect 397913 225392 397918 225448
rect 397974 225392 538862 225448
rect 538918 225392 538923 225448
rect 397913 225390 538923 225392
rect 397913 225387 397979 225390
rect 538857 225387 538923 225390
rect 70393 225314 70459 225317
rect 199377 225314 199443 225317
rect 70393 225312 199443 225314
rect 70393 225256 70398 225312
rect 70454 225256 199382 225312
rect 199438 225256 199443 225312
rect 70393 225254 199443 225256
rect 70393 225251 70459 225254
rect 199377 225251 199443 225254
rect 401133 225314 401199 225317
rect 545757 225314 545823 225317
rect 401133 225312 545823 225314
rect 401133 225256 401138 225312
rect 401194 225256 545762 225312
rect 545818 225256 545823 225312
rect 401133 225254 545823 225256
rect 401133 225251 401199 225254
rect 545757 225251 545823 225254
rect 63309 225178 63375 225181
rect 196525 225178 196591 225181
rect 63309 225176 196591 225178
rect 63309 225120 63314 225176
rect 63370 225120 196530 225176
rect 196586 225120 196591 225176
rect 63309 225118 196591 225120
rect 63309 225115 63375 225118
rect 196525 225115 196591 225118
rect 405457 225178 405523 225181
rect 556061 225178 556127 225181
rect 405457 225176 556127 225178
rect 405457 225120 405462 225176
rect 405518 225120 556066 225176
rect 556122 225120 556127 225176
rect 405457 225118 556127 225120
rect 405457 225115 405523 225118
rect 556061 225115 556127 225118
rect 58617 225042 58683 225045
rect 194041 225042 194107 225045
rect 58617 225040 194107 225042
rect 58617 224984 58622 225040
rect 58678 224984 194046 225040
rect 194102 224984 194107 225040
rect 58617 224982 194107 224984
rect 58617 224979 58683 224982
rect 194041 224979 194107 224982
rect 406469 225042 406535 225045
rect 559097 225042 559163 225045
rect 406469 225040 559163 225042
rect 406469 224984 406474 225040
rect 406530 224984 559102 225040
rect 559158 224984 559163 225040
rect 406469 224982 559163 224984
rect 406469 224979 406535 224982
rect 559097 224979 559163 224982
rect 56869 224906 56935 224909
rect 193673 224906 193739 224909
rect 56869 224904 193739 224906
rect 56869 224848 56874 224904
rect 56930 224848 193678 224904
rect 193734 224848 193739 224904
rect 56869 224846 193739 224848
rect 56869 224843 56935 224846
rect 193673 224843 193739 224846
rect 410793 224906 410859 224909
rect 568573 224906 568639 224909
rect 410793 224904 568639 224906
rect 410793 224848 410798 224904
rect 410854 224848 568578 224904
rect 568634 224848 568639 224904
rect 410793 224846 568639 224848
rect 410793 224843 410859 224846
rect 568573 224843 568639 224846
rect 112437 224770 112503 224773
rect 216857 224770 216923 224773
rect 112437 224768 216923 224770
rect 112437 224712 112442 224768
rect 112498 224712 216862 224768
rect 216918 224712 216923 224768
rect 112437 224710 216923 224712
rect 112437 224707 112503 224710
rect 216857 224707 216923 224710
rect 372245 224770 372311 224773
rect 478505 224770 478571 224773
rect 372245 224768 478571 224770
rect 372245 224712 372250 224768
rect 372306 224712 478510 224768
rect 478566 224712 478571 224768
rect 372245 224710 478571 224712
rect 372245 224707 372311 224710
rect 478505 224707 478571 224710
rect 115749 224634 115815 224637
rect 218237 224634 218303 224637
rect 115749 224632 218303 224634
rect 115749 224576 115754 224632
rect 115810 224576 218242 224632
rect 218298 224576 218303 224632
rect 115749 224574 218303 224576
rect 115749 224571 115815 224574
rect 218237 224571 218303 224574
rect 373717 224634 373783 224637
rect 481909 224634 481975 224637
rect 373717 224632 481975 224634
rect 373717 224576 373722 224632
rect 373778 224576 481914 224632
rect 481970 224576 481975 224632
rect 373717 224574 481975 224576
rect 373717 224571 373783 224574
rect 481909 224571 481975 224574
rect 117497 224498 117563 224501
rect 219341 224498 219407 224501
rect 117497 224496 219407 224498
rect 117497 224440 117502 224496
rect 117558 224440 219346 224496
rect 219402 224440 219407 224496
rect 117497 224438 219407 224440
rect 117497 224435 117563 224438
rect 219341 224435 219407 224438
rect 370865 224498 370931 224501
rect 475101 224498 475167 224501
rect 370865 224496 475167 224498
rect 370865 224440 370870 224496
rect 370926 224440 475106 224496
rect 475162 224440 475167 224496
rect 370865 224438 475167 224440
rect 370865 224435 370931 224438
rect 475101 224435 475167 224438
rect 120809 224362 120875 224365
rect 220813 224362 220879 224365
rect 120809 224360 220879 224362
rect 120809 224304 120814 224360
rect 120870 224304 220818 224360
rect 220874 224304 220879 224360
rect 120809 224302 220879 224304
rect 120809 224299 120875 224302
rect 220813 224299 220879 224302
rect 369393 224362 369459 224365
rect 471973 224362 472039 224365
rect 369393 224360 472039 224362
rect 369393 224304 369398 224360
rect 369454 224304 471978 224360
rect 472034 224304 472039 224360
rect 369393 224302 472039 224304
rect 369393 224299 369459 224302
rect 471973 224299 472039 224302
rect 160093 224226 160159 224229
rect 207933 224226 207999 224229
rect 160093 224224 207999 224226
rect 160093 224168 160098 224224
rect 160154 224168 207938 224224
rect 207994 224168 207999 224224
rect 160093 224166 207999 224168
rect 160093 224163 160159 224166
rect 207933 224163 207999 224166
rect 172421 224090 172487 224093
rect 206553 224090 206619 224093
rect 172421 224088 206619 224090
rect 172421 224032 172426 224088
rect 172482 224032 206558 224088
rect 206614 224032 206619 224088
rect 172421 224030 206619 224032
rect 172421 224027 172487 224030
rect 206553 224027 206619 224030
rect 103145 223546 103211 223549
rect 214373 223546 214439 223549
rect 103145 223544 214439 223546
rect 103145 223488 103150 223544
rect 103206 223488 214378 223544
rect 214434 223488 214439 223544
rect 103145 223486 214439 223488
rect 103145 223483 103211 223486
rect 214373 223483 214439 223486
rect 375097 223546 375163 223549
rect 483841 223546 483907 223549
rect 375097 223544 483907 223546
rect 375097 223488 375102 223544
rect 375158 223488 483846 223544
rect 483902 223488 483907 223544
rect 375097 223486 483907 223488
rect 375097 223483 375163 223486
rect 483841 223483 483907 223486
rect 675845 223546 675911 223549
rect 675845 223544 676292 223546
rect 675845 223488 675850 223544
rect 675906 223488 676292 223544
rect 675845 223486 676292 223488
rect 675845 223483 675911 223486
rect 98085 223410 98151 223413
rect 211889 223410 211955 223413
rect 98085 223408 211955 223410
rect 98085 223352 98090 223408
rect 98146 223352 211894 223408
rect 211950 223352 211955 223408
rect 98085 223350 211955 223352
rect 98085 223347 98151 223350
rect 211889 223347 211955 223350
rect 378317 223410 378383 223413
rect 491937 223410 492003 223413
rect 378317 223408 492003 223410
rect 378317 223352 378322 223408
rect 378378 223352 491942 223408
rect 491998 223352 492003 223408
rect 378317 223350 492003 223352
rect 378317 223347 378383 223350
rect 491937 223347 492003 223350
rect 96429 223274 96495 223277
rect 211521 223274 211587 223277
rect 96429 223272 211587 223274
rect 96429 223216 96434 223272
rect 96490 223216 211526 223272
rect 211582 223216 211587 223272
rect 96429 223214 211587 223216
rect 96429 223211 96495 223214
rect 211521 223211 211587 223214
rect 378685 223274 378751 223277
rect 491385 223274 491451 223277
rect 378685 223272 491451 223274
rect 378685 223216 378690 223272
rect 378746 223216 491390 223272
rect 491446 223216 491451 223272
rect 378685 223214 491451 223216
rect 378685 223211 378751 223214
rect 491385 223211 491451 223214
rect 79593 223138 79659 223141
rect 204345 223138 204411 223141
rect 79593 223136 204411 223138
rect 79593 223080 79598 223136
rect 79654 223080 204350 223136
rect 204406 223080 204411 223136
rect 79593 223078 204411 223080
rect 79593 223075 79659 223078
rect 204345 223075 204411 223078
rect 381169 223138 381235 223141
rect 498653 223138 498719 223141
rect 381169 223136 498719 223138
rect 381169 223080 381174 223136
rect 381230 223080 498658 223136
rect 498714 223080 498719 223136
rect 381169 223078 498719 223080
rect 381169 223075 381235 223078
rect 498653 223075 498719 223078
rect 675937 223138 676003 223141
rect 675937 223136 676292 223138
rect 675937 223080 675942 223136
rect 675998 223080 676292 223136
rect 675937 223078 676292 223080
rect 675937 223075 676003 223078
rect 72877 223002 72943 223005
rect 201493 223002 201559 223005
rect 72877 223000 201559 223002
rect 72877 222944 72882 223000
rect 72938 222944 201498 223000
rect 201554 222944 201559 223000
rect 72877 222942 201559 222944
rect 72877 222939 72943 222942
rect 201493 222939 201559 222942
rect 383653 223002 383719 223005
rect 504817 223002 504883 223005
rect 383653 223000 504883 223002
rect 383653 222944 383658 223000
rect 383714 222944 504822 223000
rect 504878 222944 504883 223000
rect 383653 222942 504883 222944
rect 383653 222939 383719 222942
rect 504817 222939 504883 222942
rect 74441 222866 74507 222869
rect 201861 222866 201927 222869
rect 74441 222864 201927 222866
rect 74441 222808 74446 222864
rect 74502 222808 201866 222864
rect 201922 222808 201927 222864
rect 74441 222806 201927 222808
rect 74441 222803 74507 222806
rect 201861 222803 201927 222806
rect 381537 222866 381603 222869
rect 500217 222866 500283 222869
rect 381537 222864 500283 222866
rect 381537 222808 381542 222864
rect 381598 222808 500222 222864
rect 500278 222808 500283 222864
rect 381537 222806 500283 222808
rect 381537 222803 381603 222806
rect 500217 222803 500283 222806
rect 66161 222730 66227 222733
rect 198641 222730 198707 222733
rect 66161 222728 198707 222730
rect 66161 222672 66166 222728
rect 66222 222672 198646 222728
rect 198702 222672 198707 222728
rect 66161 222670 198707 222672
rect 66161 222667 66227 222670
rect 198641 222667 198707 222670
rect 330937 222730 331003 222733
rect 381077 222730 381143 222733
rect 330937 222728 381143 222730
rect 330937 222672 330942 222728
rect 330998 222672 381082 222728
rect 381138 222672 381143 222728
rect 330937 222670 381143 222672
rect 330937 222667 331003 222670
rect 381077 222667 381143 222670
rect 385861 222730 385927 222733
rect 509601 222730 509667 222733
rect 385861 222728 509667 222730
rect 385861 222672 385866 222728
rect 385922 222672 509606 222728
rect 509662 222672 509667 222728
rect 385861 222670 509667 222672
rect 385861 222667 385927 222670
rect 509601 222667 509667 222670
rect 676029 222730 676095 222733
rect 676029 222728 676292 222730
rect 676029 222672 676034 222728
rect 676090 222672 676292 222728
rect 676029 222670 676292 222672
rect 676029 222667 676095 222670
rect 67817 222594 67883 222597
rect 199009 222594 199075 222597
rect 67817 222592 199075 222594
rect 67817 222536 67822 222592
rect 67878 222536 199014 222592
rect 199070 222536 199075 222592
rect 67817 222534 199075 222536
rect 67817 222531 67883 222534
rect 199009 222531 199075 222534
rect 332317 222594 332383 222597
rect 384297 222594 384363 222597
rect 332317 222592 384363 222594
rect 332317 222536 332322 222592
rect 332378 222536 384302 222592
rect 384358 222536 384363 222592
rect 332317 222534 384363 222536
rect 332317 222531 332383 222534
rect 384297 222531 384363 222534
rect 387977 222594 388043 222597
rect 514661 222594 514727 222597
rect 387977 222592 514727 222594
rect 387977 222536 387982 222592
rect 388038 222536 514666 222592
rect 514722 222536 514727 222592
rect 387977 222534 514727 222536
rect 387977 222531 388043 222534
rect 514661 222531 514727 222534
rect 61101 222458 61167 222461
rect 196157 222458 196223 222461
rect 61101 222456 196223 222458
rect 61101 222400 61106 222456
rect 61162 222400 196162 222456
rect 196218 222400 196223 222456
rect 61101 222398 196223 222400
rect 61101 222395 61167 222398
rect 196157 222395 196223 222398
rect 333053 222458 333119 222461
rect 383653 222458 383719 222461
rect 333053 222456 383719 222458
rect 333053 222400 333058 222456
rect 333114 222400 383658 222456
rect 383714 222400 383719 222456
rect 333053 222398 383719 222400
rect 333053 222395 333119 222398
rect 383653 222395 383719 222398
rect 388989 222458 389055 222461
rect 517053 222458 517119 222461
rect 388989 222456 517119 222458
rect 388989 222400 388994 222456
rect 389050 222400 517058 222456
rect 517114 222400 517119 222456
rect 388989 222398 517119 222400
rect 388989 222395 389055 222398
rect 517053 222395 517119 222398
rect 59169 222322 59235 222325
rect 195789 222322 195855 222325
rect 59169 222320 195855 222322
rect 59169 222264 59174 222320
rect 59230 222264 195794 222320
rect 195850 222264 195855 222320
rect 59169 222262 195855 222264
rect 59169 222259 59235 222262
rect 195789 222259 195855 222262
rect 333789 222322 333855 222325
rect 387701 222322 387767 222325
rect 333789 222320 387767 222322
rect 333789 222264 333794 222320
rect 333850 222264 387706 222320
rect 387762 222264 387767 222320
rect 333789 222262 387767 222264
rect 333789 222259 333855 222262
rect 387701 222259 387767 222262
rect 391197 222322 391263 222325
rect 522205 222322 522271 222325
rect 391197 222320 522271 222322
rect 391197 222264 391202 222320
rect 391258 222264 522210 222320
rect 522266 222264 522271 222320
rect 391197 222262 522271 222264
rect 391197 222259 391263 222262
rect 522205 222259 522271 222262
rect 675661 222322 675727 222325
rect 675661 222320 676292 222322
rect 675661 222264 675666 222320
rect 675722 222264 676292 222320
rect 675661 222262 676292 222264
rect 675661 222259 675727 222262
rect 54385 222186 54451 222189
rect 193305 222186 193371 222189
rect 54385 222184 193371 222186
rect 54385 222128 54390 222184
rect 54446 222128 193310 222184
rect 193366 222128 193371 222184
rect 54385 222126 193371 222128
rect 54385 222123 54451 222126
rect 193305 222123 193371 222126
rect 335905 222186 335971 222189
rect 390185 222186 390251 222189
rect 335905 222184 390251 222186
rect 335905 222128 335910 222184
rect 335966 222128 390190 222184
rect 390246 222128 390251 222184
rect 335905 222126 390251 222128
rect 335905 222123 335971 222126
rect 390185 222123 390251 222126
rect 393313 222186 393379 222189
rect 527265 222186 527331 222189
rect 393313 222184 527331 222186
rect 393313 222128 393318 222184
rect 393374 222128 527270 222184
rect 527326 222128 527331 222184
rect 393313 222126 527331 222128
rect 393313 222123 393379 222126
rect 527265 222123 527331 222126
rect 104801 222050 104867 222053
rect 214741 222050 214807 222053
rect 104801 222048 214807 222050
rect 104801 221992 104806 222048
rect 104862 221992 214746 222048
rect 214802 221992 214807 222048
rect 104801 221990 214807 221992
rect 104801 221987 104867 221990
rect 214741 221987 214807 221990
rect 375833 222050 375899 222053
rect 486325 222050 486391 222053
rect 375833 222048 486391 222050
rect 375833 221992 375838 222048
rect 375894 221992 486330 222048
rect 486386 221992 486391 222048
rect 375833 221990 486391 221992
rect 375833 221987 375899 221990
rect 486325 221987 486391 221990
rect 109861 221914 109927 221917
rect 217225 221914 217291 221917
rect 109861 221912 217291 221914
rect 109861 221856 109866 221912
rect 109922 221856 217230 221912
rect 217286 221856 217291 221912
rect 109861 221854 217291 221856
rect 109861 221851 109927 221854
rect 217225 221851 217291 221854
rect 338757 221914 338823 221917
rect 396901 221914 396967 221917
rect 338757 221912 396967 221914
rect 338757 221856 338762 221912
rect 338818 221856 396906 221912
rect 396962 221856 396967 221912
rect 338757 221854 396967 221856
rect 338757 221851 338823 221854
rect 396901 221851 396967 221854
rect 675569 221914 675635 221917
rect 675569 221912 676292 221914
rect 675569 221856 675574 221912
rect 675630 221856 676292 221912
rect 675569 221854 676292 221856
rect 675569 221851 675635 221854
rect 111609 221778 111675 221781
rect 217317 221778 217383 221781
rect 111609 221776 217383 221778
rect 111609 221720 111614 221776
rect 111670 221720 217322 221776
rect 217378 221720 217383 221776
rect 111609 221718 217383 221720
rect 111609 221715 111675 221718
rect 217317 221715 217383 221718
rect 335813 221778 335879 221781
rect 388529 221778 388595 221781
rect 335813 221776 388595 221778
rect 335813 221720 335818 221776
rect 335874 221720 388534 221776
rect 388590 221720 388595 221776
rect 335813 221718 388595 221720
rect 335813 221715 335879 221718
rect 388529 221715 388595 221718
rect 564341 221778 564407 221781
rect 564341 221776 574110 221778
rect 564341 221720 564346 221776
rect 564402 221720 574110 221776
rect 564341 221718 574110 221720
rect 564341 221715 564407 221718
rect 119981 221642 120047 221645
rect 221457 221642 221523 221645
rect 119981 221640 221523 221642
rect 119981 221584 119986 221640
rect 120042 221584 221462 221640
rect 221518 221584 221523 221640
rect 119981 221582 221523 221584
rect 119981 221579 120047 221582
rect 221457 221579 221523 221582
rect 334525 221642 334591 221645
rect 386781 221642 386847 221645
rect 334525 221640 386847 221642
rect 334525 221584 334530 221640
rect 334586 221584 386786 221640
rect 386842 221584 386847 221640
rect 334525 221582 386847 221584
rect 334525 221579 334591 221582
rect 386781 221579 386847 221582
rect 567101 221642 567167 221645
rect 574050 221642 574110 221718
rect 574369 221642 574435 221645
rect 567101 221640 573834 221642
rect 567101 221584 567106 221640
rect 567162 221584 573834 221640
rect 567101 221582 573834 221584
rect 574050 221640 574435 221642
rect 574050 221584 574374 221640
rect 574430 221584 574435 221640
rect 574050 221582 574435 221584
rect 567101 221579 567167 221582
rect 121361 221506 121427 221509
rect 221825 221506 221891 221509
rect 121361 221504 221891 221506
rect 121361 221448 121366 221504
rect 121422 221448 221830 221504
rect 221886 221448 221891 221504
rect 121361 221446 221891 221448
rect 121361 221443 121427 221446
rect 221825 221443 221891 221446
rect 564525 221506 564591 221509
rect 573541 221506 573607 221509
rect 564525 221504 573607 221506
rect 564525 221448 564530 221504
rect 564586 221448 573546 221504
rect 573602 221448 573607 221504
rect 564525 221446 573607 221448
rect 573774 221506 573834 221582
rect 574369 221579 574435 221582
rect 575197 221506 575263 221509
rect 573774 221504 575263 221506
rect 573774 221448 575202 221504
rect 575258 221448 575263 221504
rect 573774 221446 575263 221448
rect 564525 221443 564591 221446
rect 573541 221443 573607 221446
rect 575197 221443 575263 221446
rect 675017 221506 675083 221509
rect 675017 221504 676292 221506
rect 675017 221448 675022 221504
rect 675078 221448 676292 221504
rect 675017 221446 676292 221448
rect 675017 221443 675083 221446
rect 118325 221370 118391 221373
rect 220445 221370 220511 221373
rect 118325 221368 220511 221370
rect 118325 221312 118330 221368
rect 118386 221312 220450 221368
rect 220506 221312 220511 221368
rect 118325 221310 220511 221312
rect 118325 221307 118391 221310
rect 220445 221307 220511 221310
rect 507393 221370 507459 221373
rect 624325 221370 624391 221373
rect 507393 221368 624391 221370
rect 507393 221312 507398 221368
rect 507454 221312 624330 221368
rect 624386 221312 624391 221368
rect 507393 221310 624391 221312
rect 507393 221307 507459 221310
rect 624325 221307 624391 221310
rect 495341 221234 495407 221237
rect 622485 221234 622551 221237
rect 495341 221232 622551 221234
rect 495341 221176 495346 221232
rect 495402 221176 622490 221232
rect 622546 221176 622551 221232
rect 495341 221174 622551 221176
rect 495341 221171 495407 221174
rect 622485 221171 622551 221174
rect 500217 221098 500283 221101
rect 637849 221098 637915 221101
rect 500217 221096 637915 221098
rect 500217 221040 500222 221096
rect 500278 221040 637854 221096
rect 637910 221040 637915 221096
rect 500217 221038 637915 221040
rect 500217 221035 500283 221038
rect 637849 221035 637915 221038
rect 675385 221098 675451 221101
rect 675385 221096 676292 221098
rect 675385 221040 675390 221096
rect 675446 221040 676292 221096
rect 675385 221038 676292 221040
rect 675385 221035 675451 221038
rect 491385 220962 491451 220965
rect 493041 220962 493107 220965
rect 636929 220962 636995 220965
rect 491385 220960 636995 220962
rect 491385 220904 491390 220960
rect 491446 220904 493046 220960
rect 493102 220904 636934 220960
rect 636990 220904 636995 220960
rect 491385 220902 636995 220904
rect 491385 220899 491451 220902
rect 493041 220899 493107 220902
rect 636929 220899 636995 220902
rect 675753 220690 675819 220693
rect 675753 220688 676292 220690
rect 675753 220632 675758 220688
rect 675814 220632 676292 220688
rect 675753 220630 676292 220632
rect 675753 220627 675819 220630
rect 675937 220282 676003 220285
rect 675937 220280 676292 220282
rect 675937 220224 675942 220280
rect 675998 220224 676292 220280
rect 675937 220222 676292 220224
rect 675937 220219 676003 220222
rect 675150 219812 675156 219876
rect 675220 219874 675226 219876
rect 675220 219814 676292 219874
rect 675220 219812 675226 219814
rect 676029 219466 676095 219469
rect 676029 219464 676292 219466
rect 676029 219408 676034 219464
rect 676090 219408 676292 219464
rect 676029 219406 676292 219408
rect 676029 219403 676095 219406
rect 676029 219058 676095 219061
rect 676029 219056 676292 219058
rect 676029 219000 676034 219056
rect 676090 219000 676292 219056
rect 676029 218998 676292 219000
rect 676029 218995 676095 218998
rect 675477 218650 675543 218653
rect 675477 218648 676292 218650
rect 675477 218592 675482 218648
rect 675538 218592 676292 218648
rect 675477 218590 676292 218592
rect 675477 218587 675543 218590
rect 676029 218242 676095 218245
rect 676029 218240 676292 218242
rect 676029 218184 676034 218240
rect 676090 218184 676292 218240
rect 676029 218182 676292 218184
rect 676029 218179 676095 218182
rect 676029 217834 676095 217837
rect 676029 217832 676292 217834
rect 676029 217776 676034 217832
rect 676090 217776 676292 217832
rect 676029 217774 676292 217776
rect 676029 217771 676095 217774
rect 675937 217426 676003 217429
rect 675937 217424 676292 217426
rect 675937 217368 675942 217424
rect 675998 217368 676292 217424
rect 675937 217366 676292 217368
rect 675937 217363 676003 217366
rect 63401 217290 63467 217293
rect 652753 217290 652819 217293
rect 63401 217288 652819 217290
rect 63401 217232 63406 217288
rect 63462 217232 652758 217288
rect 652814 217232 652819 217288
rect 63401 217230 652819 217232
rect 63401 217227 63467 217230
rect 652753 217227 652819 217230
rect 671889 217154 671955 217157
rect 47280 217152 671955 217154
rect 47280 217146 671894 217152
rect 47280 217094 47298 217146
rect 47293 217086 47298 217094
rect 47358 217096 671894 217146
rect 671950 217096 671955 217152
rect 47358 217094 671955 217096
rect 47358 217086 47363 217094
rect 671889 217091 671955 217094
rect 47293 217081 47363 217086
rect 675845 217018 675911 217021
rect 675845 217016 676292 217018
rect 675845 216960 675850 217016
rect 675906 216960 676292 217016
rect 675845 216958 676292 216960
rect 675845 216955 675911 216958
rect 47385 216882 47455 216885
rect 673085 216882 673151 216885
rect 47370 216880 673151 216882
rect 47370 216822 47390 216880
rect 47385 216820 47390 216822
rect 47450 216824 673090 216880
rect 673146 216824 673151 216880
rect 47450 216822 673151 216824
rect 47450 216820 47455 216822
rect 47385 216815 47455 216820
rect 673085 216819 673151 216822
rect 673269 216610 673335 216613
rect 47458 216608 673335 216610
rect 47458 216604 673274 216608
rect 47458 216550 47482 216604
rect 47477 216544 47482 216550
rect 47542 216552 673274 216604
rect 673330 216552 673335 216608
rect 47542 216550 673335 216552
rect 47542 216544 47547 216550
rect 673269 216547 673335 216550
rect 676029 216610 676095 216613
rect 676029 216608 676292 216610
rect 676029 216552 676034 216608
rect 676090 216552 676292 216608
rect 676029 216550 676292 216552
rect 676029 216547 676095 216550
rect 47477 216539 47547 216544
rect 582281 216202 582347 216205
rect 576380 216200 582347 216202
rect 576380 216144 582286 216200
rect 582342 216144 582347 216200
rect 576380 216142 582347 216144
rect 582281 216139 582347 216142
rect 675937 216202 676003 216205
rect 675937 216200 676292 216202
rect 675937 216144 675942 216200
rect 675998 216144 676292 216200
rect 675937 216142 676292 216144
rect 675937 216139 676003 216142
rect 675845 215794 675911 215797
rect 675845 215792 676292 215794
rect 675845 215736 675850 215792
rect 675906 215736 676292 215792
rect 675845 215734 676292 215736
rect 675845 215731 675911 215734
rect 675753 215386 675819 215389
rect 675753 215384 676292 215386
rect 675753 215328 675758 215384
rect 675814 215328 676292 215384
rect 675753 215326 676292 215328
rect 675753 215323 675819 215326
rect 41689 215114 41755 215117
rect 41462 215112 41755 215114
rect 41462 215056 41694 215112
rect 41750 215056 41755 215112
rect 41462 215054 41755 215056
rect 41462 214948 41522 215054
rect 41689 215051 41755 215054
rect 676029 214978 676095 214981
rect 676029 214976 676292 214978
rect 676029 214920 676034 214976
rect 676090 214920 676292 214976
rect 676029 214918 676292 214920
rect 676029 214915 676095 214918
rect 41505 214706 41571 214709
rect 582281 214706 582347 214709
rect 41462 214704 41571 214706
rect 41462 214648 41510 214704
rect 41566 214648 41571 214704
rect 41462 214643 41571 214648
rect 576380 214704 582347 214706
rect 576380 214648 582286 214704
rect 582342 214648 582347 214704
rect 576380 214646 582347 214648
rect 582281 214643 582347 214646
rect 41462 214540 41522 214643
rect 676029 214570 676095 214573
rect 676029 214568 676292 214570
rect 676029 214512 676034 214568
rect 676090 214512 676292 214568
rect 676029 214510 676292 214512
rect 676029 214507 676095 214510
rect 41413 214298 41479 214301
rect 41413 214296 41522 214298
rect 41413 214240 41418 214296
rect 41474 214240 41522 214296
rect 41413 214235 41522 214240
rect 41462 214132 41522 214235
rect 675937 214162 676003 214165
rect 675937 214160 676292 214162
rect 675937 214104 675942 214160
rect 675998 214104 676292 214160
rect 675937 214102 676292 214104
rect 675937 214099 676003 214102
rect 675753 213754 675819 213757
rect 675753 213752 676292 213754
rect 44587 213712 44653 213715
rect 41540 213710 44670 213712
rect 41540 213654 44592 213710
rect 44648 213654 44670 213710
rect 675753 213696 675758 213752
rect 675814 213696 676292 213752
rect 675753 213694 676292 213696
rect 675753 213691 675819 213694
rect 41540 213652 44670 213654
rect 44587 213649 44653 213652
rect 47477 213312 47547 213313
rect 41476 213308 47554 213312
rect 41476 213252 47482 213308
rect 47477 213248 47482 213252
rect 47542 213252 47554 213308
rect 676078 213286 676292 213346
rect 47542 213248 47547 213252
rect 47477 213243 47547 213248
rect 580257 213210 580323 213213
rect 576380 213208 580323 213210
rect 576380 213152 580262 213208
rect 580318 213152 580323 213208
rect 576380 213150 580323 213152
rect 580257 213147 580323 213150
rect 42333 212938 42399 212941
rect 41492 212936 42399 212938
rect 41492 212880 42338 212936
rect 42394 212880 42399 212936
rect 41492 212878 42399 212880
rect 42333 212875 42399 212878
rect 41505 212666 41571 212669
rect 41462 212664 41571 212666
rect 41462 212608 41510 212664
rect 41566 212608 41571 212664
rect 41462 212603 41571 212608
rect 41462 212500 41522 212603
rect 676078 212125 676138 213286
rect 679022 212500 679082 212908
rect 676029 212122 676138 212125
rect 675948 212120 676292 212122
rect 44683 212078 44749 212081
rect 41556 212076 44760 212078
rect 41556 212020 44688 212076
rect 44744 212020 44760 212076
rect 675948 212064 676034 212120
rect 676090 212064 676292 212120
rect 675948 212062 676292 212064
rect 676029 212059 676095 212062
rect 41556 212018 44760 212020
rect 44683 212015 44749 212018
rect 580073 211714 580139 211717
rect 576380 211712 580139 211714
rect 47293 211680 47363 211685
rect 41510 211620 47298 211680
rect 47358 211620 47374 211680
rect 576380 211656 580078 211712
rect 580134 211656 580139 211712
rect 576380 211654 580139 211656
rect 580073 211651 580139 211654
rect 47293 211615 47363 211620
rect 44773 211268 44839 211271
rect 41552 211266 44850 211268
rect 41552 211210 44778 211266
rect 44834 211210 44850 211266
rect 41552 211208 44850 211210
rect 44773 211205 44839 211208
rect 47385 210870 47455 210871
rect 41502 210866 47462 210870
rect 41502 210810 47390 210866
rect 47385 210806 47390 210810
rect 47450 210810 47462 210866
rect 47450 210806 47455 210810
rect 47385 210801 47455 210806
rect 37782 210221 37842 210460
rect 37782 210216 37891 210221
rect 582281 210218 582347 210221
rect 37782 210160 37830 210216
rect 37886 210160 37891 210216
rect 37782 210158 37891 210160
rect 576380 210216 582347 210218
rect 576380 210160 582286 210216
rect 582342 210160 582347 210216
rect 576380 210158 582347 210160
rect 37825 210155 37891 210158
rect 582281 210155 582347 210158
rect 37966 209813 38026 210052
rect 37966 209808 38075 209813
rect 37966 209752 38014 209808
rect 38070 209752 38075 209808
rect 37966 209750 38075 209752
rect 38009 209747 38075 209750
rect 38334 209405 38394 209644
rect 600037 209538 600103 209541
rect 600037 209536 606556 209538
rect 600037 209480 600042 209536
rect 600098 209480 606556 209536
rect 600037 209478 606556 209480
rect 600037 209475 600103 209478
rect 38285 209400 38394 209405
rect 38285 209344 38290 209400
rect 38346 209344 38394 209400
rect 38285 209342 38394 209344
rect 38285 209339 38351 209342
rect 666553 209266 666619 209269
rect 666356 209264 666619 209266
rect 38150 208997 38210 209236
rect 666356 209208 666558 209264
rect 666614 209208 666619 209264
rect 666356 209206 666619 209208
rect 666553 209203 666619 209206
rect 38150 208992 38259 208997
rect 38150 208936 38198 208992
rect 38254 208936 38259 208992
rect 38150 208934 38259 208936
rect 38193 208931 38259 208934
rect 38150 208589 38210 208828
rect 581453 208722 581519 208725
rect 576380 208720 581519 208722
rect 576380 208664 581458 208720
rect 581514 208664 581519 208720
rect 576380 208662 581519 208664
rect 581453 208659 581519 208662
rect 38101 208584 38210 208589
rect 38101 208528 38106 208584
rect 38162 208528 38210 208584
rect 38101 208526 38210 208528
rect 599945 208586 600011 208589
rect 599945 208584 606556 208586
rect 599945 208528 599950 208584
rect 600006 208528 606556 208584
rect 599945 208526 606556 208528
rect 38101 208523 38167 208526
rect 599945 208523 600011 208526
rect 38518 208181 38578 208420
rect 38518 208176 38627 208181
rect 38518 208120 38566 208176
rect 38622 208120 38627 208176
rect 38518 208118 38627 208120
rect 38561 208115 38627 208118
rect 38334 207773 38394 208012
rect 38334 207768 38443 207773
rect 38334 207712 38382 207768
rect 38438 207712 38443 207768
rect 38334 207710 38443 207712
rect 38377 207707 38443 207710
rect 38518 207365 38578 207604
rect 599853 207498 599919 207501
rect 599853 207496 606556 207498
rect 599853 207440 599858 207496
rect 599914 207440 606556 207496
rect 599853 207438 606556 207440
rect 599853 207435 599919 207438
rect 38469 207360 38578 207365
rect 38469 207304 38474 207360
rect 38530 207304 38578 207360
rect 38469 207302 38578 207304
rect 38469 207299 38535 207302
rect 37966 206957 38026 207196
rect 582281 207090 582347 207093
rect 576380 207088 582347 207090
rect 576380 207032 582286 207088
rect 582342 207032 582347 207088
rect 576380 207030 582347 207032
rect 582281 207027 582347 207030
rect 37917 206952 38026 206957
rect 37917 206896 37922 206952
rect 37978 206896 38026 206952
rect 37917 206894 38026 206896
rect 37917 206891 37983 206894
rect 42701 206818 42767 206821
rect 41492 206816 42767 206818
rect 41492 206760 42706 206816
rect 42762 206760 42767 206816
rect 41492 206758 42767 206760
rect 42701 206755 42767 206758
rect 600773 206546 600839 206549
rect 600773 206544 606556 206546
rect 600773 206488 600778 206544
rect 600834 206488 606556 206544
rect 600773 206486 606556 206488
rect 600773 206483 600839 206486
rect 43253 206410 43319 206413
rect 41492 206408 43319 206410
rect 41492 206352 43258 206408
rect 43314 206352 43319 206408
rect 41492 206350 43319 206352
rect 43253 206347 43319 206350
rect 675569 206274 675635 206277
rect 675526 206272 675635 206274
rect 675526 206216 675574 206272
rect 675630 206216 675635 206272
rect 675526 206211 675635 206216
rect 43437 206002 43503 206005
rect 41492 206000 43503 206002
rect 41492 205944 43442 206000
rect 43498 205944 43503 206000
rect 41492 205942 43503 205944
rect 43437 205939 43503 205942
rect 667105 206002 667171 206005
rect 675385 206002 675451 206005
rect 667105 206000 675451 206002
rect 667105 205944 667110 206000
rect 667166 205944 675390 206000
rect 675446 205944 675451 206000
rect 667105 205942 675451 205944
rect 667105 205939 667171 205942
rect 675385 205939 675451 205942
rect 666553 205866 666619 205869
rect 666356 205864 666619 205866
rect 666356 205808 666558 205864
rect 666614 205808 666619 205864
rect 666356 205806 666619 205808
rect 666553 205803 666619 205806
rect 43069 205594 43135 205597
rect 582281 205594 582347 205597
rect 41492 205592 43135 205594
rect 41492 205536 43074 205592
rect 43130 205536 43135 205592
rect 41492 205534 43135 205536
rect 576380 205592 582347 205594
rect 576380 205536 582286 205592
rect 582342 205536 582347 205592
rect 576380 205534 582347 205536
rect 43069 205531 43135 205534
rect 582281 205531 582347 205534
rect 601141 205458 601207 205461
rect 601141 205456 606556 205458
rect 601141 205400 601146 205456
rect 601202 205400 606556 205456
rect 601141 205398 606556 205400
rect 601141 205395 601207 205398
rect 42333 205186 42399 205189
rect 41492 205184 42399 205186
rect 41492 205128 42338 205184
rect 42394 205128 42399 205184
rect 41492 205126 42399 205128
rect 42333 205123 42399 205126
rect 38377 204914 38443 204917
rect 41638 204914 41644 204916
rect 38377 204912 41644 204914
rect 38377 204856 38382 204912
rect 38438 204856 41644 204912
rect 38377 204854 41644 204856
rect 38377 204851 38443 204854
rect 41638 204852 41644 204854
rect 41708 204852 41714 204916
rect 674833 204914 674899 204917
rect 675526 204914 675586 206211
rect 674833 204912 675586 204914
rect 674833 204856 674838 204912
rect 674894 204856 675586 204912
rect 674833 204854 675586 204856
rect 674833 204851 674899 204854
rect 48221 204778 48287 204781
rect 41492 204776 48287 204778
rect 41492 204720 48226 204776
rect 48282 204720 48287 204776
rect 41492 204718 48287 204720
rect 48221 204715 48287 204718
rect 38285 204506 38351 204509
rect 41454 204506 41460 204508
rect 38285 204504 41460 204506
rect 38285 204448 38290 204504
rect 38346 204448 41460 204504
rect 38285 204446 41460 204448
rect 38285 204443 38351 204446
rect 41454 204444 41460 204446
rect 41524 204444 41530 204508
rect 601601 204506 601667 204509
rect 601601 204504 606556 204506
rect 601601 204448 601606 204504
rect 601662 204448 606556 204504
rect 601601 204446 606556 204448
rect 601601 204443 601667 204446
rect 30054 204101 30114 204340
rect 666553 204234 666619 204237
rect 666356 204232 666619 204234
rect 666356 204176 666558 204232
rect 666614 204176 666619 204232
rect 666356 204174 666619 204176
rect 666553 204171 666619 204174
rect 30054 204096 30163 204101
rect 580717 204098 580783 204101
rect 30054 204040 30102 204096
rect 30158 204040 30163 204096
rect 30054 204038 30163 204040
rect 576380 204096 580783 204098
rect 576380 204040 580722 204096
rect 580778 204040 580783 204096
rect 576380 204038 580783 204040
rect 30097 204035 30163 204038
rect 580717 204035 580783 204038
rect 31661 203690 31727 203693
rect 31661 203688 31770 203690
rect 31661 203632 31666 203688
rect 31722 203632 31770 203688
rect 31661 203627 31770 203632
rect 31710 203524 31770 203627
rect 599669 203418 599735 203421
rect 599669 203416 606556 203418
rect 599669 203360 599674 203416
rect 599730 203360 606556 203416
rect 599669 203358 606556 203360
rect 599669 203355 599735 203358
rect 581085 202602 581151 202605
rect 576380 202600 581151 202602
rect 576380 202544 581090 202600
rect 581146 202544 581151 202600
rect 576380 202542 581151 202544
rect 581085 202539 581151 202542
rect 8201 202466 8267 202469
rect 30097 202466 30163 202469
rect 8201 202464 30163 202466
rect 8201 202408 8206 202464
rect 8262 202408 30102 202464
rect 30158 202408 30163 202464
rect 8201 202406 30163 202408
rect 8201 202403 8267 202406
rect 30097 202403 30163 202406
rect 599945 202466 600011 202469
rect 599945 202464 606556 202466
rect 599945 202408 599950 202464
rect 600006 202408 606556 202464
rect 599945 202406 606556 202408
rect 599945 202403 600011 202406
rect 598933 201378 598999 201381
rect 598933 201376 606556 201378
rect 598933 201320 598938 201376
rect 598994 201320 606556 201376
rect 598933 201318 606556 201320
rect 598933 201315 598999 201318
rect 581085 201106 581151 201109
rect 576380 201104 581151 201106
rect 576380 201048 581090 201104
rect 581146 201048 581151 201104
rect 576380 201046 581151 201048
rect 581085 201043 581151 201046
rect 666553 200834 666619 200837
rect 666356 200832 666619 200834
rect 666356 200776 666558 200832
rect 666614 200776 666619 200832
rect 666356 200774 666619 200776
rect 666553 200771 666619 200774
rect 599945 200426 600011 200429
rect 599945 200424 606556 200426
rect 599945 200368 599950 200424
rect 600006 200368 606556 200424
rect 599945 200366 606556 200368
rect 599945 200363 600011 200366
rect 582281 199610 582347 199613
rect 576380 199608 582347 199610
rect 576380 199552 582286 199608
rect 582342 199552 582347 199608
rect 576380 199550 582347 199552
rect 582281 199547 582347 199550
rect 599945 199338 600011 199341
rect 599945 199336 606556 199338
rect 599945 199280 599950 199336
rect 600006 199280 606556 199336
rect 599945 199278 606556 199280
rect 599945 199275 600011 199278
rect 666553 199066 666619 199069
rect 666356 199064 666619 199066
rect 666356 199008 666558 199064
rect 666614 199008 666619 199064
rect 666356 199006 666619 199008
rect 666553 199003 666619 199006
rect 37825 198794 37891 198797
rect 41822 198794 41828 198796
rect 37825 198792 41828 198794
rect 37825 198736 37830 198792
rect 37886 198736 41828 198792
rect 37825 198734 41828 198736
rect 37825 198731 37891 198734
rect 41822 198732 41828 198734
rect 41892 198732 41898 198796
rect 599945 198386 600011 198389
rect 599945 198384 606556 198386
rect 599945 198328 599950 198384
rect 600006 198328 606556 198384
rect 599945 198326 606556 198328
rect 599945 198323 600011 198326
rect 582281 197978 582347 197981
rect 576380 197976 582347 197978
rect 576380 197920 582286 197976
rect 582342 197920 582347 197976
rect 576380 197918 582347 197920
rect 582281 197915 582347 197918
rect 599945 197298 600011 197301
rect 599945 197296 606556 197298
rect 599945 197240 599950 197296
rect 600006 197240 606556 197296
rect 599945 197238 606556 197240
rect 599945 197235 600011 197238
rect 580717 196482 580783 196485
rect 576380 196480 580783 196482
rect 576380 196424 580722 196480
rect 580778 196424 580783 196480
rect 576380 196422 580783 196424
rect 580717 196419 580783 196422
rect 599393 196346 599459 196349
rect 599393 196344 606556 196346
rect 599393 196288 599398 196344
rect 599454 196288 606556 196344
rect 599393 196286 606556 196288
rect 599393 196283 599459 196286
rect 666553 195666 666619 195669
rect 666356 195664 666619 195666
rect 666356 195608 666558 195664
rect 666614 195608 666619 195664
rect 666356 195606 666619 195608
rect 666553 195603 666619 195606
rect 599853 195258 599919 195261
rect 599853 195256 606556 195258
rect 599853 195200 599858 195256
rect 599914 195200 606556 195256
rect 599853 195198 606556 195200
rect 599853 195195 599919 195198
rect 582281 194986 582347 194989
rect 576380 194984 582347 194986
rect 576380 194928 582286 194984
rect 582342 194928 582347 194984
rect 576380 194926 582347 194928
rect 582281 194923 582347 194926
rect 599945 194306 600011 194309
rect 599945 194304 606556 194306
rect 599945 194248 599950 194304
rect 600006 194248 606556 194304
rect 599945 194246 606556 194248
rect 599945 194243 600011 194246
rect 670693 194034 670759 194037
rect 666356 194032 670759 194034
rect 666356 193976 670698 194032
rect 670754 193976 670759 194032
rect 666356 193974 670759 193976
rect 670693 193971 670759 193974
rect 582189 193490 582255 193493
rect 576380 193488 582255 193490
rect 576380 193432 582194 193488
rect 582250 193432 582255 193488
rect 576380 193430 582255 193432
rect 582189 193427 582255 193430
rect 599485 193218 599551 193221
rect 599485 193216 606556 193218
rect 599485 193160 599490 193216
rect 599546 193160 606556 193216
rect 599485 193158 606556 193160
rect 599485 193155 599551 193158
rect 599945 192266 600011 192269
rect 599945 192264 606556 192266
rect 599945 192208 599950 192264
rect 600006 192208 606556 192264
rect 599945 192206 606556 192208
rect 599945 192203 600011 192206
rect 582281 191994 582347 191997
rect 576380 191992 582347 191994
rect 576380 191936 582286 191992
rect 582342 191936 582347 191992
rect 576380 191934 582347 191936
rect 582281 191931 582347 191934
rect 599945 191178 600011 191181
rect 599945 191176 606556 191178
rect 599945 191120 599950 191176
rect 600006 191120 606556 191176
rect 599945 191118 606556 191120
rect 599945 191115 600011 191118
rect 670693 190634 670759 190637
rect 666356 190632 670759 190634
rect 666356 190576 670698 190632
rect 670754 190576 670759 190632
rect 666356 190574 670759 190576
rect 670693 190571 670759 190574
rect 581269 190498 581335 190501
rect 576380 190496 581335 190498
rect 576380 190440 581274 190496
rect 581330 190440 581335 190496
rect 576380 190438 581335 190440
rect 581269 190435 581335 190438
rect 601509 190226 601575 190229
rect 601509 190224 606556 190226
rect 601509 190168 601514 190224
rect 601570 190168 606556 190224
rect 601509 190166 606556 190168
rect 601509 190163 601575 190166
rect 601601 189138 601667 189141
rect 601601 189136 606556 189138
rect 601601 189080 601606 189136
rect 601662 189080 606556 189136
rect 601601 189078 606556 189080
rect 601601 189075 601667 189078
rect 666553 189002 666619 189005
rect 666356 189000 666619 189002
rect 666356 188944 666558 189000
rect 666614 188944 666619 189000
rect 666356 188942 666619 188944
rect 666553 188939 666619 188942
rect 579705 188866 579771 188869
rect 576380 188864 579771 188866
rect 576380 188808 579710 188864
rect 579766 188808 579771 188864
rect 576380 188806 579771 188808
rect 579705 188803 579771 188806
rect 599117 188186 599183 188189
rect 599117 188184 606556 188186
rect 599117 188128 599122 188184
rect 599178 188128 606556 188184
rect 599117 188126 606556 188128
rect 599117 188123 599183 188126
rect 582281 187370 582347 187373
rect 576380 187368 582347 187370
rect 576380 187312 582286 187368
rect 582342 187312 582347 187368
rect 576380 187310 582347 187312
rect 582281 187307 582347 187310
rect 599945 187098 600011 187101
rect 599945 187096 606556 187098
rect 599945 187040 599950 187096
rect 600006 187040 606556 187096
rect 599945 187038 606556 187040
rect 599945 187035 600011 187038
rect 600037 186146 600103 186149
rect 600037 186144 606556 186146
rect 600037 186088 600042 186144
rect 600098 186088 606556 186144
rect 600037 186086 606556 186088
rect 600037 186083 600103 186086
rect 579889 185874 579955 185877
rect 576380 185872 579955 185874
rect 576380 185816 579894 185872
rect 579950 185816 579955 185872
rect 576380 185814 579955 185816
rect 579889 185811 579955 185814
rect 666553 185602 666619 185605
rect 666356 185600 666619 185602
rect 666356 185544 666558 185600
rect 666614 185544 666619 185600
rect 666356 185542 666619 185544
rect 666553 185539 666619 185542
rect 599853 185058 599919 185061
rect 599853 185056 606556 185058
rect 599853 185000 599858 185056
rect 599914 185000 606556 185056
rect 599853 184998 606556 185000
rect 599853 184995 599919 184998
rect 580901 184378 580967 184381
rect 576380 184376 580967 184378
rect 576380 184320 580906 184376
rect 580962 184320 580967 184376
rect 576380 184318 580967 184320
rect 580901 184315 580967 184318
rect 41873 184244 41939 184245
rect 41822 184242 41828 184244
rect 41782 184182 41828 184242
rect 41892 184240 41939 184244
rect 41934 184184 41939 184240
rect 41822 184180 41828 184182
rect 41892 184180 41939 184184
rect 41873 184179 41939 184180
rect 599945 184106 600011 184109
rect 599945 184104 606556 184106
rect 599945 184048 599950 184104
rect 600006 184048 606556 184104
rect 599945 184046 606556 184048
rect 599945 184043 600011 184046
rect 666553 183834 666619 183837
rect 666356 183832 666619 183834
rect 666356 183776 666558 183832
rect 666614 183776 666619 183832
rect 666356 183774 666619 183776
rect 666553 183771 666619 183774
rect 41638 183364 41644 183428
rect 41708 183426 41714 183428
rect 41781 183426 41847 183429
rect 41708 183424 41847 183426
rect 41708 183368 41786 183424
rect 41842 183368 41847 183424
rect 41708 183366 41847 183368
rect 41708 183364 41714 183366
rect 41781 183363 41847 183366
rect 598933 183018 598999 183021
rect 598933 183016 606556 183018
rect 598933 182960 598938 183016
rect 598994 182960 606556 183016
rect 598933 182958 606556 182960
rect 598933 182955 598999 182958
rect 580257 182882 580323 182885
rect 576380 182880 580323 182882
rect 576380 182824 580262 182880
rect 580318 182824 580323 182880
rect 576380 182822 580323 182824
rect 580257 182819 580323 182822
rect 41454 182684 41460 182748
rect 41524 182746 41530 182748
rect 41781 182746 41847 182749
rect 41524 182744 41847 182746
rect 41524 182688 41786 182744
rect 41842 182688 41847 182744
rect 41524 182686 41847 182688
rect 41524 182684 41530 182686
rect 41781 182683 41847 182686
rect 600037 182066 600103 182069
rect 600037 182064 606556 182066
rect 600037 182008 600042 182064
rect 600098 182008 606556 182064
rect 600037 182006 606556 182008
rect 600037 182003 600103 182006
rect 580625 181386 580691 181389
rect 576380 181384 580691 181386
rect 576380 181328 580630 181384
rect 580686 181328 580691 181384
rect 576380 181326 580691 181328
rect 580625 181323 580691 181326
rect 600129 180978 600195 180981
rect 600129 180976 606556 180978
rect 600129 180920 600134 180976
rect 600190 180920 606556 180976
rect 600129 180918 606556 180920
rect 600129 180915 600195 180918
rect 666553 180434 666619 180437
rect 666356 180432 666619 180434
rect 666356 180376 666558 180432
rect 666614 180376 666619 180432
rect 666356 180374 666619 180376
rect 666553 180371 666619 180374
rect 599853 180026 599919 180029
rect 599853 180024 606556 180026
rect 599853 179968 599858 180024
rect 599914 179968 606556 180024
rect 599853 179966 606556 179968
rect 599853 179963 599919 179966
rect 580533 179754 580599 179757
rect 576380 179752 580599 179754
rect 576380 179696 580538 179752
rect 580594 179696 580599 179752
rect 576380 179694 580599 179696
rect 580533 179691 580599 179694
rect 599669 178938 599735 178941
rect 599669 178936 606556 178938
rect 599669 178880 599674 178936
rect 599730 178880 606556 178936
rect 599669 178878 606556 178880
rect 599669 178875 599735 178878
rect 670693 178802 670759 178805
rect 671981 178802 672047 178805
rect 666356 178800 672047 178802
rect 666356 178744 670698 178800
rect 670754 178744 671986 178800
rect 672042 178744 672047 178800
rect 666356 178742 672047 178744
rect 670693 178739 670759 178742
rect 671981 178739 672047 178742
rect 675845 178530 675911 178533
rect 675845 178528 676292 178530
rect 675845 178472 675850 178528
rect 675906 178472 676292 178528
rect 675845 178470 676292 178472
rect 675845 178467 675911 178470
rect 581085 178258 581151 178261
rect 576380 178256 581151 178258
rect 576380 178200 581090 178256
rect 581146 178200 581151 178256
rect 576380 178198 581151 178200
rect 581085 178195 581151 178198
rect 675937 178122 676003 178125
rect 675937 178120 676292 178122
rect 675937 178064 675942 178120
rect 675998 178064 676292 178120
rect 675937 178062 676292 178064
rect 675937 178059 676003 178062
rect 599761 177986 599827 177989
rect 599761 177984 606556 177986
rect 599761 177928 599766 177984
rect 599822 177928 606556 177984
rect 599761 177926 606556 177928
rect 599761 177923 599827 177926
rect 676029 177714 676095 177717
rect 676029 177712 676292 177714
rect 676029 177656 676034 177712
rect 676090 177656 676292 177712
rect 676029 177654 676292 177656
rect 676029 177651 676095 177654
rect 675293 177306 675359 177309
rect 675293 177304 676292 177306
rect 675293 177248 675298 177304
rect 675354 177248 676292 177304
rect 675293 177246 676292 177248
rect 675293 177243 675359 177246
rect 599945 176898 600011 176901
rect 674925 176898 674991 176901
rect 599945 176896 606556 176898
rect 599945 176840 599950 176896
rect 600006 176840 606556 176896
rect 599945 176838 606556 176840
rect 674906 176896 676292 176898
rect 674906 176840 674930 176896
rect 674986 176840 676292 176896
rect 674906 176838 676292 176840
rect 599945 176835 600011 176838
rect 674925 176835 674991 176838
rect 580717 176762 580783 176765
rect 576380 176760 580783 176762
rect 576380 176704 580722 176760
rect 580778 176704 580783 176760
rect 576380 176702 580783 176704
rect 580717 176699 580783 176702
rect 676029 176490 676095 176493
rect 676029 176488 676292 176490
rect 676029 176432 676034 176488
rect 676090 176432 676292 176488
rect 676029 176430 676292 176432
rect 676029 176427 676095 176430
rect 675937 176082 676003 176085
rect 675937 176080 676292 176082
rect 675937 176024 675942 176080
rect 675998 176024 676292 176080
rect 675937 176022 676292 176024
rect 675937 176019 676003 176022
rect 600405 175946 600471 175949
rect 600405 175944 606556 175946
rect 600405 175888 600410 175944
rect 600466 175888 606556 175944
rect 600405 175886 606556 175888
rect 600405 175883 600471 175886
rect 676029 175674 676095 175677
rect 676029 175672 676292 175674
rect 676029 175616 676034 175672
rect 676090 175616 676292 175672
rect 676029 175614 676292 175616
rect 676029 175611 676095 175614
rect 670693 175402 670759 175405
rect 666356 175400 670759 175402
rect 666356 175344 670698 175400
rect 670754 175344 670759 175400
rect 666356 175342 670759 175344
rect 670693 175339 670759 175342
rect 581453 175266 581519 175269
rect 576380 175264 581519 175266
rect 576380 175208 581458 175264
rect 581514 175208 581519 175264
rect 576380 175206 581519 175208
rect 581453 175203 581519 175206
rect 675385 175266 675451 175269
rect 675385 175264 676292 175266
rect 675385 175208 675390 175264
rect 675446 175208 676292 175264
rect 675385 175206 676292 175208
rect 675385 175203 675451 175206
rect 599945 174858 600011 174861
rect 676029 174858 676095 174861
rect 599945 174856 606556 174858
rect 599945 174800 599950 174856
rect 600006 174800 606556 174856
rect 599945 174798 606556 174800
rect 676029 174856 676292 174858
rect 676029 174800 676034 174856
rect 676090 174800 676292 174856
rect 676029 174798 676292 174800
rect 599945 174795 600011 174798
rect 676029 174795 676095 174798
rect 675753 174450 675819 174453
rect 675734 174448 676292 174450
rect 675734 174392 675758 174448
rect 675814 174392 676292 174448
rect 675734 174390 676292 174392
rect 675753 174387 675819 174390
rect 676029 174042 676095 174045
rect 676029 174040 676292 174042
rect 676029 173984 676034 174040
rect 676090 173984 676292 174040
rect 676029 173982 676292 173984
rect 676029 173979 676095 173982
rect 601325 173906 601391 173909
rect 601325 173904 606556 173906
rect 601325 173848 601330 173904
rect 601386 173848 606556 173904
rect 601325 173846 606556 173848
rect 601325 173843 601391 173846
rect 582281 173770 582347 173773
rect 576380 173768 582347 173770
rect 576380 173712 582286 173768
rect 582342 173712 582347 173768
rect 576380 173710 582347 173712
rect 582281 173707 582347 173710
rect 666553 173634 666619 173637
rect 672073 173634 672139 173637
rect 666356 173632 672139 173634
rect 666356 173576 666558 173632
rect 666614 173576 672078 173632
rect 672134 173576 672139 173632
rect 666356 173574 672139 173576
rect 666553 173571 666619 173574
rect 672073 173571 672139 173574
rect 676029 173634 676095 173637
rect 676029 173632 676292 173634
rect 676029 173576 676034 173632
rect 676090 173576 676292 173632
rect 676029 173574 676292 173576
rect 676029 173571 676095 173574
rect 675569 173226 675635 173229
rect 675569 173224 676292 173226
rect 675569 173168 675574 173224
rect 675630 173168 676292 173224
rect 675569 173166 676292 173168
rect 675569 173163 675635 173166
rect 599485 172818 599551 172821
rect 676029 172818 676095 172821
rect 599485 172816 606556 172818
rect 599485 172760 599490 172816
rect 599546 172760 606556 172816
rect 599485 172758 606556 172760
rect 676029 172816 676292 172818
rect 676029 172760 676034 172816
rect 676090 172760 676292 172816
rect 676029 172758 676292 172760
rect 599485 172755 599551 172758
rect 676029 172755 676095 172758
rect 675937 172410 676003 172413
rect 675937 172408 676292 172410
rect 675937 172352 675942 172408
rect 675998 172352 676292 172408
rect 675937 172350 676292 172352
rect 675937 172347 676003 172350
rect 579705 172274 579771 172277
rect 576380 172272 579771 172274
rect 576380 172216 579710 172272
rect 579766 172216 579771 172272
rect 576380 172214 579771 172216
rect 579705 172211 579771 172214
rect 675937 172002 676003 172005
rect 675937 172000 676292 172002
rect 675937 171944 675942 172000
rect 675998 171944 676292 172000
rect 675937 171942 676292 171944
rect 675937 171939 676003 171942
rect 599945 171866 600011 171869
rect 599945 171864 606556 171866
rect 599945 171808 599950 171864
rect 600006 171808 606556 171864
rect 599945 171806 606556 171808
rect 599945 171803 600011 171806
rect 675661 171594 675727 171597
rect 675661 171592 676292 171594
rect 675661 171536 675666 171592
rect 675722 171536 676292 171592
rect 675661 171534 676292 171536
rect 675661 171531 675727 171534
rect 676029 171186 676095 171189
rect 676029 171184 676292 171186
rect 676029 171128 676034 171184
rect 676090 171128 676292 171184
rect 676029 171126 676292 171128
rect 676029 171123 676095 171126
rect 599853 170778 599919 170781
rect 676029 170778 676095 170781
rect 599853 170776 606556 170778
rect 599853 170720 599858 170776
rect 599914 170720 606556 170776
rect 599853 170718 606556 170720
rect 676029 170776 676292 170778
rect 676029 170720 676034 170776
rect 676090 170720 676292 170776
rect 676029 170718 676292 170720
rect 599853 170715 599919 170718
rect 676029 170715 676095 170718
rect 580533 170642 580599 170645
rect 576380 170640 580599 170642
rect 576380 170584 580538 170640
rect 580594 170584 580599 170640
rect 576380 170582 580599 170584
rect 580533 170579 580599 170582
rect 675937 170370 676003 170373
rect 675937 170368 676292 170370
rect 675937 170312 675942 170368
rect 675998 170312 676292 170368
rect 675937 170310 676292 170312
rect 675937 170307 676003 170310
rect 666553 170234 666619 170237
rect 666356 170232 666619 170234
rect 666356 170176 666558 170232
rect 666614 170176 666619 170232
rect 666356 170174 666619 170176
rect 666553 170171 666619 170174
rect 675937 169962 676003 169965
rect 675937 169960 676292 169962
rect 675937 169904 675942 169960
rect 675998 169904 676292 169960
rect 675937 169902 676292 169904
rect 675937 169899 676003 169902
rect 599945 169826 600011 169829
rect 599945 169824 606556 169826
rect 599945 169768 599950 169824
rect 600006 169768 606556 169824
rect 599945 169766 606556 169768
rect 599945 169763 600011 169766
rect 676029 169554 676095 169557
rect 676029 169552 676292 169554
rect 676029 169496 676034 169552
rect 676090 169496 676292 169552
rect 676029 169494 676292 169496
rect 676029 169491 676095 169494
rect 582005 169146 582071 169149
rect 576380 169144 582071 169146
rect 576380 169088 582010 169144
rect 582066 169088 582071 169144
rect 576380 169086 582071 169088
rect 582005 169083 582071 169086
rect 675937 169146 676003 169149
rect 675937 169144 676292 169146
rect 675937 169088 675942 169144
rect 675998 169088 676292 169144
rect 675937 169086 676292 169088
rect 675937 169083 676003 169086
rect 599485 168738 599551 168741
rect 676029 168738 676095 168741
rect 599485 168736 606556 168738
rect 599485 168680 599490 168736
rect 599546 168680 606556 168736
rect 599485 168678 606556 168680
rect 676029 168736 676292 168738
rect 676029 168680 676034 168736
rect 676090 168680 676292 168736
rect 676029 168678 676292 168680
rect 599485 168675 599551 168678
rect 676029 168675 676095 168678
rect 666737 168602 666803 168605
rect 672165 168602 672231 168605
rect 666356 168600 672231 168602
rect 666356 168544 666742 168600
rect 666798 168544 672170 168600
rect 672226 168544 672231 168600
rect 666356 168542 672231 168544
rect 666737 168539 666803 168542
rect 672165 168539 672231 168542
rect 599485 167786 599551 167789
rect 599485 167784 606556 167786
rect 599485 167728 599490 167784
rect 599546 167728 606556 167784
rect 599485 167726 606556 167728
rect 599485 167723 599551 167726
rect 581085 167650 581151 167653
rect 576380 167648 581151 167650
rect 576380 167592 581090 167648
rect 581146 167592 581151 167648
rect 576380 167590 581151 167592
rect 581085 167587 581151 167590
rect 676029 167106 676095 167109
rect 676029 167104 676292 167106
rect 676029 167048 676034 167104
rect 676090 167048 676292 167104
rect 676029 167046 676292 167048
rect 676029 167043 676095 167046
rect 600037 166698 600103 166701
rect 600037 166696 606556 166698
rect 600037 166640 600042 166696
rect 600098 166640 606556 166696
rect 600037 166638 606556 166640
rect 600037 166635 600103 166638
rect 580165 166154 580231 166157
rect 576380 166152 580231 166154
rect 576380 166096 580170 166152
rect 580226 166096 580231 166152
rect 576380 166094 580231 166096
rect 580165 166091 580231 166094
rect 599945 165746 600011 165749
rect 599945 165744 606556 165746
rect 599945 165688 599950 165744
rect 600006 165688 606556 165744
rect 599945 165686 606556 165688
rect 599945 165683 600011 165686
rect 666737 165202 666803 165205
rect 666356 165200 666803 165202
rect 666356 165144 666742 165200
rect 666798 165144 666803 165200
rect 666356 165142 666803 165144
rect 666737 165139 666803 165142
rect 581637 164658 581703 164661
rect 576380 164656 581703 164658
rect 576380 164600 581642 164656
rect 581698 164600 581703 164656
rect 576380 164598 581703 164600
rect 581637 164595 581703 164598
rect 600037 164658 600103 164661
rect 600037 164656 606556 164658
rect 600037 164600 600042 164656
rect 600098 164600 606556 164656
rect 600037 164598 606556 164600
rect 600037 164595 600103 164598
rect 599945 163706 600011 163709
rect 599945 163704 606556 163706
rect 599945 163648 599950 163704
rect 600006 163648 606556 163704
rect 599945 163646 606556 163648
rect 599945 163643 600011 163646
rect 666737 163570 666803 163573
rect 672257 163570 672323 163573
rect 666356 163568 672323 163570
rect 666356 163512 666742 163568
rect 666798 163512 672262 163568
rect 672318 163512 672323 163568
rect 666356 163510 672323 163512
rect 666737 163507 666803 163510
rect 672257 163507 672323 163510
rect 581821 163162 581887 163165
rect 576380 163160 581887 163162
rect 576380 163104 581826 163160
rect 581882 163104 581887 163160
rect 576380 163102 581887 163104
rect 581821 163099 581887 163102
rect 600037 162618 600103 162621
rect 600037 162616 606556 162618
rect 600037 162560 600042 162616
rect 600098 162560 606556 162616
rect 600037 162558 606556 162560
rect 600037 162555 600103 162558
rect 599853 161666 599919 161669
rect 599853 161664 606556 161666
rect 599853 161608 599858 161664
rect 599914 161608 606556 161664
rect 599853 161606 606556 161608
rect 599853 161603 599919 161606
rect 579889 161530 579955 161533
rect 576380 161528 579955 161530
rect 576380 161472 579894 161528
rect 579950 161472 579955 161528
rect 576380 161470 579955 161472
rect 579889 161467 579955 161470
rect 599945 160578 600011 160581
rect 599945 160576 606556 160578
rect 599945 160520 599950 160576
rect 600006 160520 606556 160576
rect 599945 160518 606556 160520
rect 599945 160515 600011 160518
rect 666737 160170 666803 160173
rect 666356 160168 666803 160170
rect 666356 160112 666742 160168
rect 666798 160112 666803 160168
rect 666356 160110 666803 160112
rect 666737 160107 666803 160110
rect 582005 160034 582071 160037
rect 576380 160032 582071 160034
rect 576380 159976 582010 160032
rect 582066 159976 582071 160032
rect 576380 159974 582071 159976
rect 582005 159971 582071 159974
rect 599853 159626 599919 159629
rect 599853 159624 606556 159626
rect 599853 159568 599858 159624
rect 599914 159568 606556 159624
rect 599853 159566 606556 159568
rect 599853 159563 599919 159566
rect 579797 158538 579863 158541
rect 576380 158536 579863 158538
rect 576380 158480 579802 158536
rect 579858 158480 579863 158536
rect 576380 158478 579863 158480
rect 579797 158475 579863 158478
rect 600037 158538 600103 158541
rect 600037 158536 606556 158538
rect 600037 158480 600042 158536
rect 600098 158480 606556 158536
rect 600037 158478 606556 158480
rect 600037 158475 600103 158478
rect 666737 158402 666803 158405
rect 672349 158402 672415 158405
rect 666356 158400 672415 158402
rect 666356 158344 666742 158400
rect 666798 158344 672354 158400
rect 672410 158344 672415 158400
rect 666356 158342 672415 158344
rect 666737 158339 666803 158342
rect 672349 158339 672415 158342
rect 599945 157586 600011 157589
rect 599945 157584 606556 157586
rect 599945 157528 599950 157584
rect 600006 157528 606556 157584
rect 599945 157526 606556 157528
rect 599945 157523 600011 157526
rect 580441 157042 580507 157045
rect 576380 157040 580507 157042
rect 576380 156984 580446 157040
rect 580502 156984 580507 157040
rect 576380 156982 580507 156984
rect 580441 156979 580507 156982
rect 599853 156498 599919 156501
rect 599853 156496 606556 156498
rect 599853 156440 599858 156496
rect 599914 156440 606556 156496
rect 599853 156438 606556 156440
rect 599853 156435 599919 156438
rect 580257 155546 580323 155549
rect 576380 155544 580323 155546
rect 576380 155488 580262 155544
rect 580318 155488 580323 155544
rect 576380 155486 580323 155488
rect 580257 155483 580323 155486
rect 599945 155546 600011 155549
rect 599945 155544 606556 155546
rect 599945 155488 599950 155544
rect 600006 155488 606556 155544
rect 599945 155486 606556 155488
rect 599945 155483 600011 155486
rect 666737 155002 666803 155005
rect 666356 155000 666803 155002
rect 666356 154944 666742 155000
rect 666798 154944 666803 155000
rect 666356 154942 666803 154944
rect 666737 154939 666803 154942
rect 599853 154458 599919 154461
rect 599853 154456 606556 154458
rect 599853 154400 599858 154456
rect 599914 154400 606556 154456
rect 599853 154398 606556 154400
rect 599853 154395 599919 154398
rect 581269 154050 581335 154053
rect 576380 154048 581335 154050
rect 576380 153992 581274 154048
rect 581330 153992 581335 154048
rect 576380 153990 581335 153992
rect 581269 153987 581335 153990
rect 600037 153506 600103 153509
rect 600037 153504 606556 153506
rect 600037 153448 600042 153504
rect 600098 153448 606556 153504
rect 600037 153446 606556 153448
rect 600037 153443 600103 153446
rect 666737 153370 666803 153373
rect 672441 153370 672507 153373
rect 666356 153368 672507 153370
rect 666356 153312 666742 153368
rect 666798 153312 672446 153368
rect 672502 153312 672507 153368
rect 666356 153310 672507 153312
rect 666737 153307 666803 153310
rect 672441 153307 672507 153310
rect 582281 152418 582347 152421
rect 576380 152416 582347 152418
rect 576380 152360 582286 152416
rect 582342 152360 582347 152416
rect 576380 152358 582347 152360
rect 582281 152355 582347 152358
rect 599945 152418 600011 152421
rect 599945 152416 606556 152418
rect 599945 152360 599950 152416
rect 600006 152360 606556 152416
rect 599945 152358 606556 152360
rect 599945 152355 600011 152358
rect 600037 151466 600103 151469
rect 600037 151464 606556 151466
rect 600037 151408 600042 151464
rect 600098 151408 606556 151464
rect 600037 151406 606556 151408
rect 600037 151403 600103 151406
rect 582189 150922 582255 150925
rect 576380 150920 582255 150922
rect 576380 150864 582194 150920
rect 582250 150864 582255 150920
rect 576380 150862 582255 150864
rect 582189 150859 582255 150862
rect 599853 150378 599919 150381
rect 599853 150376 606556 150378
rect 599853 150320 599858 150376
rect 599914 150320 606556 150376
rect 599853 150318 606556 150320
rect 599853 150315 599919 150318
rect 666737 149970 666803 149973
rect 666356 149968 666803 149970
rect 666356 149912 666742 149968
rect 666798 149912 666803 149968
rect 666356 149910 666803 149912
rect 666737 149907 666803 149910
rect 580073 149426 580139 149429
rect 576380 149424 580139 149426
rect 576380 149368 580078 149424
rect 580134 149368 580139 149424
rect 576380 149366 580139 149368
rect 580073 149363 580139 149366
rect 599945 149426 600011 149429
rect 599945 149424 606556 149426
rect 599945 149368 599950 149424
rect 600006 149368 606556 149424
rect 599945 149366 606556 149368
rect 599945 149363 600011 149366
rect 599853 148338 599919 148341
rect 599853 148336 606556 148338
rect 599853 148280 599858 148336
rect 599914 148280 606556 148336
rect 599853 148278 606556 148280
rect 599853 148275 599919 148278
rect 666737 148202 666803 148205
rect 672533 148202 672599 148205
rect 666356 148200 672599 148202
rect 666356 148144 666742 148200
rect 666798 148144 672538 148200
rect 672594 148144 672599 148200
rect 666356 148142 672599 148144
rect 666737 148139 666803 148142
rect 672533 148139 672599 148142
rect 581177 147930 581243 147933
rect 576380 147928 581243 147930
rect 576380 147872 581182 147928
rect 581238 147872 581243 147928
rect 576380 147870 581243 147872
rect 581177 147867 581243 147870
rect 599945 147386 600011 147389
rect 599945 147384 606556 147386
rect 599945 147328 599950 147384
rect 600006 147328 606556 147384
rect 599945 147326 606556 147328
rect 599945 147323 600011 147326
rect 581729 146434 581795 146437
rect 576380 146432 581795 146434
rect 576380 146376 581734 146432
rect 581790 146376 581795 146432
rect 576380 146374 581795 146376
rect 581729 146371 581795 146374
rect 599853 146298 599919 146301
rect 599853 146296 606556 146298
rect 599853 146240 599858 146296
rect 599914 146240 606556 146296
rect 599853 146238 606556 146240
rect 599853 146235 599919 146238
rect 600037 145346 600103 145349
rect 600037 145344 606556 145346
rect 600037 145288 600042 145344
rect 600098 145288 606556 145344
rect 600037 145286 606556 145288
rect 600037 145283 600103 145286
rect 581637 144938 581703 144941
rect 666737 144938 666803 144941
rect 576380 144936 581703 144938
rect 576380 144880 581642 144936
rect 581698 144880 581703 144936
rect 576380 144878 581703 144880
rect 666356 144936 666803 144938
rect 666356 144880 666742 144936
rect 666798 144880 666803 144936
rect 666356 144878 666803 144880
rect 581637 144875 581703 144878
rect 666737 144875 666803 144878
rect 599945 144258 600011 144261
rect 599945 144256 606556 144258
rect 599945 144200 599950 144256
rect 600006 144200 606556 144256
rect 599945 144198 606556 144200
rect 599945 144195 600011 144198
rect 580625 143306 580691 143309
rect 576380 143304 580691 143306
rect 576380 143248 580630 143304
rect 580686 143248 580691 143304
rect 576380 143246 580691 143248
rect 580625 143243 580691 143246
rect 600037 143306 600103 143309
rect 600037 143304 606556 143306
rect 600037 143248 600042 143304
rect 600098 143248 606556 143304
rect 600037 143246 606556 143248
rect 600037 143243 600103 143246
rect 666737 143170 666803 143173
rect 672809 143170 672875 143173
rect 666356 143168 672875 143170
rect 666356 143112 666742 143168
rect 666798 143112 672814 143168
rect 672870 143112 672875 143168
rect 666356 143110 672875 143112
rect 666737 143107 666803 143110
rect 672809 143107 672875 143110
rect 599945 142218 600011 142221
rect 599945 142216 606556 142218
rect 599945 142160 599950 142216
rect 600006 142160 606556 142216
rect 599945 142158 606556 142160
rect 599945 142155 600011 142158
rect 581085 141810 581151 141813
rect 576380 141808 581151 141810
rect 576380 141752 581090 141808
rect 581146 141752 581151 141808
rect 576380 141750 581151 141752
rect 581085 141747 581151 141750
rect 599853 141266 599919 141269
rect 599853 141264 606556 141266
rect 599853 141208 599858 141264
rect 599914 141208 606556 141264
rect 599853 141206 606556 141208
rect 599853 141203 599919 141206
rect 582097 140314 582163 140317
rect 576380 140312 582163 140314
rect 576380 140256 582102 140312
rect 582158 140256 582163 140312
rect 576380 140254 582163 140256
rect 582097 140251 582163 140254
rect 600037 140178 600103 140181
rect 600037 140176 606556 140178
rect 600037 140120 600042 140176
rect 600098 140120 606556 140176
rect 600037 140118 606556 140120
rect 600037 140115 600103 140118
rect 666737 139770 666803 139773
rect 666356 139768 666803 139770
rect 666356 139712 666742 139768
rect 666798 139712 666803 139768
rect 666356 139710 666803 139712
rect 666737 139707 666803 139710
rect 599853 139226 599919 139229
rect 599853 139224 606556 139226
rect 599853 139168 599858 139224
rect 599914 139168 606556 139224
rect 599853 139166 606556 139168
rect 599853 139163 599919 139166
rect 580533 138818 580599 138821
rect 576380 138816 580599 138818
rect 576380 138760 580538 138816
rect 580594 138760 580599 138816
rect 576380 138758 580599 138760
rect 580533 138755 580599 138758
rect 672901 138458 672967 138461
rect 671316 138456 672967 138458
rect 671316 138400 672906 138456
rect 672962 138400 672967 138456
rect 671316 138398 672967 138400
rect 599945 138138 600011 138141
rect 670693 138138 670759 138141
rect 671316 138138 671376 138398
rect 672901 138395 672967 138398
rect 599945 138136 606556 138138
rect 599945 138080 599950 138136
rect 600006 138080 606556 138136
rect 599945 138078 606556 138080
rect 666356 138136 671376 138138
rect 666356 138080 670698 138136
rect 670754 138080 671376 138136
rect 666356 138078 671376 138080
rect 599945 138075 600011 138078
rect 670693 138075 670759 138078
rect 580901 137322 580967 137325
rect 576380 137320 580967 137322
rect 576380 137264 580906 137320
rect 580962 137264 580967 137320
rect 576380 137262 580967 137264
rect 580901 137259 580967 137262
rect 599853 137186 599919 137189
rect 599853 137184 606556 137186
rect 599853 137128 599858 137184
rect 599914 137128 606556 137184
rect 599853 137126 606556 137128
rect 599853 137123 599919 137126
rect 599945 136098 600011 136101
rect 599945 136096 606556 136098
rect 599945 136040 599950 136096
rect 600006 136040 606556 136096
rect 599945 136038 606556 136040
rect 599945 136035 600011 136038
rect 580717 135826 580783 135829
rect 576380 135824 580783 135826
rect 576380 135768 580722 135824
rect 580778 135768 580783 135824
rect 576380 135766 580783 135768
rect 580717 135763 580783 135766
rect 600037 135146 600103 135149
rect 600037 135144 606556 135146
rect 600037 135088 600042 135144
rect 600098 135088 606556 135144
rect 600037 135086 606556 135088
rect 600037 135083 600103 135086
rect 670693 134738 670759 134741
rect 666356 134736 670759 134738
rect 666356 134680 670698 134736
rect 670754 134680 670759 134736
rect 666356 134678 670759 134680
rect 670693 134675 670759 134678
rect 582281 134194 582347 134197
rect 576380 134192 582347 134194
rect 576380 134136 582286 134192
rect 582342 134136 582347 134192
rect 576380 134134 582347 134136
rect 582281 134131 582347 134134
rect 599853 134058 599919 134061
rect 599853 134056 606556 134058
rect 599853 134000 599858 134056
rect 599914 134000 606556 134056
rect 599853 133998 606556 134000
rect 599853 133995 599919 133998
rect 599945 133106 600011 133109
rect 676121 133106 676187 133109
rect 676262 133106 676322 133348
rect 599945 133104 606556 133106
rect 599945 133048 599950 133104
rect 600006 133048 606556 133104
rect 599945 133046 606556 133048
rect 676121 133104 676322 133106
rect 676121 133048 676126 133104
rect 676182 133048 676322 133104
rect 676121 133046 676322 133048
rect 599945 133043 600011 133046
rect 676121 133043 676187 133046
rect 666737 132970 666803 132973
rect 672993 132970 673059 132973
rect 666356 132968 673059 132970
rect 666356 132912 666742 132968
rect 666798 132912 672998 132968
rect 673054 132912 673059 132968
rect 666356 132910 673059 132912
rect 666737 132907 666803 132910
rect 672993 132907 673059 132910
rect 676029 132970 676095 132973
rect 676029 132968 676292 132970
rect 676029 132912 676034 132968
rect 676090 132912 676292 132968
rect 676029 132910 676292 132912
rect 676029 132907 676095 132910
rect 580809 132698 580875 132701
rect 576380 132696 580875 132698
rect 576380 132640 580814 132696
rect 580870 132640 580875 132696
rect 576380 132638 580875 132640
rect 580809 132635 580875 132638
rect 676213 132698 676279 132701
rect 676213 132696 676322 132698
rect 676213 132640 676218 132696
rect 676274 132640 676322 132696
rect 676213 132635 676322 132640
rect 676262 132532 676322 132635
rect 676029 132154 676095 132157
rect 676029 132152 676292 132154
rect 676029 132096 676034 132152
rect 676090 132096 676292 132152
rect 676029 132094 676292 132096
rect 676029 132091 676095 132094
rect 600037 132018 600103 132021
rect 600037 132016 606556 132018
rect 600037 131960 600042 132016
rect 600098 131960 606556 132016
rect 600037 131958 606556 131960
rect 600037 131955 600103 131958
rect 676029 131746 676095 131749
rect 676029 131744 676292 131746
rect 676029 131688 676034 131744
rect 676090 131688 676292 131744
rect 676029 131686 676292 131688
rect 676029 131683 676095 131686
rect 676213 131474 676279 131477
rect 676213 131472 676322 131474
rect 676213 131416 676218 131472
rect 676274 131416 676322 131472
rect 676213 131411 676322 131416
rect 676262 131308 676322 131411
rect 581821 131202 581887 131205
rect 576380 131200 581887 131202
rect 576380 131144 581826 131200
rect 581882 131144 581887 131200
rect 576380 131142 581887 131144
rect 581821 131139 581887 131142
rect 599853 131066 599919 131069
rect 599853 131064 606556 131066
rect 599853 131008 599858 131064
rect 599914 131008 606556 131064
rect 599853 131006 606556 131008
rect 599853 131003 599919 131006
rect 676029 130930 676095 130933
rect 676029 130928 676292 130930
rect 676029 130872 676034 130928
rect 676090 130872 676292 130928
rect 676029 130870 676292 130872
rect 676029 130867 676095 130870
rect 675293 130522 675359 130525
rect 675293 130520 676292 130522
rect 675293 130464 675298 130520
rect 675354 130464 676292 130520
rect 675293 130462 676292 130464
rect 675293 130459 675359 130462
rect 676029 130114 676095 130117
rect 676029 130112 676292 130114
rect 676029 130056 676034 130112
rect 676090 130056 676292 130112
rect 676029 130054 676292 130056
rect 676029 130051 676095 130054
rect 599945 129978 600011 129981
rect 599945 129976 606556 129978
rect 599945 129920 599950 129976
rect 600006 129920 606556 129976
rect 599945 129918 606556 129920
rect 599945 129915 600011 129918
rect 582005 129706 582071 129709
rect 576380 129704 582071 129706
rect 576380 129648 582010 129704
rect 582066 129648 582071 129704
rect 576380 129646 582071 129648
rect 582005 129643 582071 129646
rect 675753 129706 675819 129709
rect 675753 129704 676292 129706
rect 675753 129648 675758 129704
rect 675814 129648 676292 129704
rect 675753 129646 676292 129648
rect 675753 129643 675819 129646
rect 666737 129570 666803 129573
rect 666356 129568 666803 129570
rect 666356 129512 666742 129568
rect 666798 129512 666803 129568
rect 666356 129510 666803 129512
rect 666737 129507 666803 129510
rect 676213 129434 676279 129437
rect 676213 129432 676322 129434
rect 676213 129376 676218 129432
rect 676274 129376 676322 129432
rect 676213 129371 676322 129376
rect 676262 129268 676322 129371
rect 599853 129026 599919 129029
rect 599853 129024 606556 129026
rect 599853 128968 599858 129024
rect 599914 128968 606556 129024
rect 599853 128966 606556 128968
rect 599853 128963 599919 128966
rect 676029 128890 676095 128893
rect 676029 128888 676292 128890
rect 676029 128832 676034 128888
rect 676090 128832 676292 128888
rect 676029 128830 676292 128832
rect 676029 128827 676095 128830
rect 675937 128482 676003 128485
rect 675937 128480 676292 128482
rect 675937 128424 675942 128480
rect 675998 128424 676292 128480
rect 675937 128422 676292 128424
rect 675937 128419 676003 128422
rect 582189 128210 582255 128213
rect 576380 128208 582255 128210
rect 576380 128152 582194 128208
rect 582250 128152 582255 128208
rect 576380 128150 582255 128152
rect 582189 128147 582255 128150
rect 675569 128074 675635 128077
rect 675569 128072 676292 128074
rect 675569 128016 675574 128072
rect 675630 128016 676292 128072
rect 675569 128014 676292 128016
rect 675569 128011 675635 128014
rect 599945 127938 600011 127941
rect 666645 127938 666711 127941
rect 672625 127938 672691 127941
rect 599945 127936 606556 127938
rect 599945 127880 599950 127936
rect 600006 127880 606556 127936
rect 599945 127878 606556 127880
rect 666356 127936 672691 127938
rect 666356 127880 666650 127936
rect 666706 127880 672630 127936
rect 672686 127880 672691 127936
rect 666356 127878 672691 127880
rect 599945 127875 600011 127878
rect 666645 127875 666711 127878
rect 672625 127875 672691 127878
rect 676029 127666 676095 127669
rect 676029 127664 676292 127666
rect 676029 127608 676034 127664
rect 676090 127608 676292 127664
rect 676029 127606 676292 127608
rect 676029 127603 676095 127606
rect 675937 127258 676003 127261
rect 675937 127256 676292 127258
rect 675937 127200 675942 127256
rect 675998 127200 676292 127256
rect 675937 127198 676292 127200
rect 675937 127195 676003 127198
rect 599853 126986 599919 126989
rect 599853 126984 606556 126986
rect 599853 126928 599858 126984
rect 599914 126928 606556 126984
rect 599853 126926 606556 126928
rect 599853 126923 599919 126926
rect 676029 126850 676095 126853
rect 676029 126848 676292 126850
rect 676029 126792 676034 126848
rect 676090 126792 676292 126848
rect 676029 126790 676292 126792
rect 676029 126787 676095 126790
rect 581361 126714 581427 126717
rect 576380 126712 581427 126714
rect 576380 126656 581366 126712
rect 581422 126656 581427 126712
rect 576380 126654 581427 126656
rect 581361 126651 581427 126654
rect 676029 126442 676095 126445
rect 676029 126440 676292 126442
rect 676029 126384 676034 126440
rect 676090 126384 676292 126440
rect 676029 126382 676292 126384
rect 676029 126379 676095 126382
rect 675293 126034 675359 126037
rect 675293 126032 676292 126034
rect 675293 125976 675298 126032
rect 675354 125976 676292 126032
rect 675293 125974 676292 125976
rect 675293 125971 675359 125974
rect 599945 125898 600011 125901
rect 599945 125896 606556 125898
rect 599945 125840 599950 125896
rect 600006 125840 606556 125896
rect 599945 125838 606556 125840
rect 599945 125835 600011 125838
rect 675201 125626 675267 125629
rect 675201 125624 676292 125626
rect 675201 125568 675206 125624
rect 675262 125568 676292 125624
rect 675201 125566 676292 125568
rect 675201 125563 675267 125566
rect 675937 125218 676003 125221
rect 675937 125216 676292 125218
rect 675937 125160 675942 125216
rect 675998 125160 676292 125216
rect 675937 125158 676292 125160
rect 675937 125155 676003 125158
rect 581545 125082 581611 125085
rect 576380 125080 581611 125082
rect 576380 125024 581550 125080
rect 581606 125024 581611 125080
rect 576380 125022 581611 125024
rect 581545 125019 581611 125022
rect 599761 124946 599827 124949
rect 599761 124944 606556 124946
rect 599761 124888 599766 124944
rect 599822 124888 606556 124944
rect 599761 124886 606556 124888
rect 599761 124883 599827 124886
rect 675937 124810 676003 124813
rect 675937 124808 676292 124810
rect 675937 124752 675942 124808
rect 675998 124752 676292 124808
rect 675937 124750 676292 124752
rect 675937 124747 676003 124750
rect 666645 124538 666711 124541
rect 666356 124536 666711 124538
rect 666356 124480 666650 124536
rect 666706 124480 666711 124536
rect 666356 124478 666711 124480
rect 666645 124475 666711 124478
rect 675937 124402 676003 124405
rect 675937 124400 676292 124402
rect 675937 124344 675942 124400
rect 675998 124344 676292 124400
rect 675937 124342 676292 124344
rect 675937 124339 676003 124342
rect 676029 123994 676095 123997
rect 676029 123992 676292 123994
rect 676029 123936 676034 123992
rect 676090 123936 676292 123992
rect 676029 123934 676292 123936
rect 676029 123931 676095 123934
rect 600037 123858 600103 123861
rect 600037 123856 606556 123858
rect 600037 123800 600042 123856
rect 600098 123800 606556 123856
rect 600037 123798 606556 123800
rect 600037 123795 600103 123798
rect 581453 123586 581519 123589
rect 576380 123584 581519 123586
rect 576380 123528 581458 123584
rect 581514 123528 581519 123584
rect 576380 123526 581519 123528
rect 581453 123523 581519 123526
rect 675937 123586 676003 123589
rect 675937 123584 676292 123586
rect 675937 123528 675942 123584
rect 675998 123528 676292 123584
rect 675937 123526 676292 123528
rect 675937 123523 676003 123526
rect 599853 122906 599919 122909
rect 666645 122906 666711 122909
rect 672717 122906 672783 122909
rect 599853 122904 606556 122906
rect 599853 122848 599858 122904
rect 599914 122848 606556 122904
rect 599853 122846 606556 122848
rect 666356 122904 672783 122906
rect 666356 122848 666650 122904
rect 666706 122848 672722 122904
rect 672778 122848 672783 122904
rect 666356 122846 672783 122848
rect 599853 122843 599919 122846
rect 666645 122843 666711 122846
rect 672717 122843 672783 122846
rect 581913 122090 581979 122093
rect 576380 122088 581979 122090
rect 576380 122032 581918 122088
rect 581974 122032 581979 122088
rect 576380 122030 581979 122032
rect 581913 122027 581979 122030
rect 599945 121818 600011 121821
rect 599945 121816 606556 121818
rect 599945 121760 599950 121816
rect 600006 121760 606556 121816
rect 599945 121758 606556 121760
rect 599945 121755 600011 121758
rect 676262 121685 676322 121924
rect 676213 121680 676322 121685
rect 676213 121624 676218 121680
rect 676274 121624 676322 121680
rect 676213 121622 676322 121624
rect 676213 121619 676279 121622
rect 600037 120866 600103 120869
rect 600037 120864 606556 120866
rect 600037 120808 600042 120864
rect 600098 120808 606556 120864
rect 600037 120806 606556 120808
rect 600037 120803 600103 120806
rect 581269 120594 581335 120597
rect 576380 120592 581335 120594
rect 576380 120536 581274 120592
rect 581330 120536 581335 120592
rect 576380 120534 581335 120536
rect 581269 120531 581335 120534
rect 599945 119778 600011 119781
rect 599945 119776 606556 119778
rect 599945 119720 599950 119776
rect 600006 119720 606556 119776
rect 599945 119718 606556 119720
rect 599945 119715 600011 119718
rect 666645 119506 666711 119509
rect 666356 119504 666711 119506
rect 666356 119448 666650 119504
rect 666706 119448 666711 119504
rect 666356 119446 666711 119448
rect 666645 119443 666711 119446
rect 581729 119098 581795 119101
rect 576380 119096 581795 119098
rect 576380 119040 581734 119096
rect 581790 119040 581795 119096
rect 576380 119038 581795 119040
rect 581729 119035 581795 119038
rect 599853 118826 599919 118829
rect 599853 118824 606556 118826
rect 599853 118768 599858 118824
rect 599914 118768 606556 118824
rect 599853 118766 606556 118768
rect 599853 118763 599919 118766
rect 600037 117738 600103 117741
rect 600037 117736 606556 117738
rect 600037 117680 600042 117736
rect 600098 117680 606556 117736
rect 600037 117678 606556 117680
rect 600037 117675 600103 117678
rect 580993 117602 581059 117605
rect 576380 117600 581059 117602
rect 576380 117544 580998 117600
rect 581054 117544 581059 117600
rect 576380 117542 581059 117544
rect 580993 117539 581059 117542
rect 599945 116786 600011 116789
rect 599945 116784 606556 116786
rect 599945 116728 599950 116784
rect 600006 116728 606556 116784
rect 599945 116726 606556 116728
rect 599945 116723 600011 116726
rect 581637 115970 581703 115973
rect 576380 115968 581703 115970
rect 576380 115912 581642 115968
rect 581698 115912 581703 115968
rect 576380 115910 581703 115912
rect 581637 115907 581703 115910
rect 599853 115698 599919 115701
rect 599853 115696 606556 115698
rect 599853 115640 599858 115696
rect 599914 115640 606556 115696
rect 599853 115638 606556 115640
rect 599853 115635 599919 115638
rect 599945 114746 600011 114749
rect 599945 114744 606556 114746
rect 599945 114688 599950 114744
rect 600006 114688 606556 114744
rect 599945 114686 606556 114688
rect 599945 114683 600011 114686
rect 581177 114474 581243 114477
rect 576380 114472 581243 114474
rect 576380 114416 581182 114472
rect 581238 114416 581243 114472
rect 576380 114414 581243 114416
rect 581177 114411 581243 114414
rect 671981 114338 672047 114341
rect 666356 114336 672047 114338
rect 666356 114280 671986 114336
rect 672042 114280 672047 114336
rect 666356 114278 672047 114280
rect 671981 114275 672047 114278
rect 580942 113188 580948 113252
rect 581012 113250 581018 113252
rect 606526 113250 606586 113628
rect 581012 113190 606586 113250
rect 581012 113188 581018 113190
rect 579705 112978 579771 112981
rect 576380 112976 579771 112978
rect 576380 112920 579710 112976
rect 579766 112920 579771 112976
rect 576380 112918 579771 112920
rect 579705 112915 579771 112918
rect 599853 112706 599919 112709
rect 599853 112704 606556 112706
rect 599853 112648 599858 112704
rect 599914 112648 606556 112704
rect 599853 112646 606556 112648
rect 599853 112643 599919 112646
rect 599945 111618 600011 111621
rect 599945 111616 606556 111618
rect 599945 111560 599950 111616
rect 600006 111560 606556 111616
rect 599945 111558 606556 111560
rect 599945 111555 600011 111558
rect 579889 111482 579955 111485
rect 576380 111480 579955 111482
rect 576380 111424 579894 111480
rect 579950 111424 579955 111480
rect 576380 111422 579955 111424
rect 579889 111419 579955 111422
rect 600221 110666 600287 110669
rect 600221 110664 606556 110666
rect 600221 110608 600226 110664
rect 600282 110608 606556 110664
rect 600221 110606 606556 110608
rect 600221 110603 600287 110606
rect 581085 109986 581151 109989
rect 576380 109984 581151 109986
rect 576380 109928 581090 109984
rect 581146 109928 581151 109984
rect 576380 109926 581151 109928
rect 581085 109923 581151 109926
rect 599301 109578 599367 109581
rect 599301 109576 606556 109578
rect 599301 109520 599306 109576
rect 599362 109520 606556 109576
rect 599301 109518 606556 109520
rect 599301 109515 599367 109518
rect 672441 109306 672507 109309
rect 666356 109304 672507 109306
rect 666356 109248 672446 109304
rect 672502 109248 672507 109304
rect 666356 109246 672507 109248
rect 672441 109243 672507 109246
rect 600313 108626 600379 108629
rect 600313 108624 606556 108626
rect 600313 108568 600318 108624
rect 600374 108568 606556 108624
rect 600313 108566 606556 108568
rect 600313 108563 600379 108566
rect 580073 108490 580139 108493
rect 576380 108488 580139 108490
rect 576380 108432 580078 108488
rect 580134 108432 580139 108488
rect 576380 108430 580139 108432
rect 580073 108427 580139 108430
rect 599945 107538 600011 107541
rect 666921 107538 666987 107541
rect 599945 107536 606556 107538
rect 599945 107480 599950 107536
rect 600006 107480 606556 107536
rect 599945 107478 606556 107480
rect 666356 107536 666987 107538
rect 666356 107480 666926 107536
rect 666982 107480 666987 107536
rect 666356 107478 666987 107480
rect 599945 107475 600011 107478
rect 666921 107475 666987 107478
rect 580165 106858 580231 106861
rect 576380 106856 580231 106858
rect 576380 106800 580170 106856
rect 580226 106800 580231 106856
rect 576380 106798 580231 106800
rect 580165 106795 580231 106798
rect 600589 106586 600655 106589
rect 600589 106584 606556 106586
rect 600589 106528 600594 106584
rect 600650 106528 606556 106584
rect 600589 106526 606556 106528
rect 600589 106523 600655 106526
rect 672257 105906 672323 105909
rect 666356 105904 672323 105906
rect 666356 105848 672262 105904
rect 672318 105848 672323 105904
rect 666356 105846 672323 105848
rect 672257 105843 672323 105846
rect 600405 105498 600471 105501
rect 600405 105496 606556 105498
rect 600405 105440 600410 105496
rect 600466 105440 606556 105496
rect 600405 105438 606556 105440
rect 600405 105435 600471 105438
rect 579981 105362 580047 105365
rect 576380 105360 580047 105362
rect 576380 105304 579986 105360
rect 580042 105304 580047 105360
rect 576380 105302 580047 105304
rect 579981 105299 580047 105302
rect 600865 104546 600931 104549
rect 600865 104544 606556 104546
rect 600865 104488 600870 104544
rect 600926 104488 606556 104544
rect 600865 104486 606556 104488
rect 600865 104483 600931 104486
rect 672165 104138 672231 104141
rect 666356 104136 672231 104138
rect 666356 104080 672170 104136
rect 672226 104080 672231 104136
rect 666356 104078 672231 104080
rect 672165 104075 672231 104078
rect 580257 103866 580323 103869
rect 576380 103864 580323 103866
rect 576380 103808 580262 103864
rect 580318 103808 580323 103864
rect 576380 103806 580323 103808
rect 580257 103803 580323 103806
rect 600681 103458 600747 103461
rect 600681 103456 606556 103458
rect 600681 103400 600686 103456
rect 600742 103400 606556 103456
rect 600681 103398 606556 103400
rect 600681 103395 600747 103398
rect 600497 102506 600563 102509
rect 672349 102506 672415 102509
rect 600497 102504 606556 102506
rect 600497 102448 600502 102504
rect 600558 102448 606556 102504
rect 600497 102446 606556 102448
rect 666356 102504 672415 102506
rect 666356 102448 672354 102504
rect 672410 102448 672415 102504
rect 666356 102446 672415 102448
rect 600497 102443 600563 102446
rect 672349 102443 672415 102446
rect 580901 102370 580967 102373
rect 576380 102368 580967 102370
rect 576380 102312 580906 102368
rect 580962 102312 580967 102368
rect 576380 102310 580967 102312
rect 580901 102307 580967 102310
rect 600773 101418 600839 101421
rect 600773 101416 606556 101418
rect 600773 101360 600778 101416
rect 600834 101360 606556 101416
rect 600773 101358 606556 101360
rect 600773 101355 600839 101358
rect 580349 100874 580415 100877
rect 672073 100874 672139 100877
rect 576380 100872 580415 100874
rect 576380 100816 580354 100872
rect 580410 100816 580415 100872
rect 576380 100814 580415 100816
rect 666356 100872 672139 100874
rect 666356 100816 672078 100872
rect 672134 100816 672139 100872
rect 666356 100814 672139 100816
rect 580349 100811 580415 100814
rect 672073 100811 672139 100814
rect 599945 100466 600011 100469
rect 599945 100464 606556 100466
rect 599945 100408 599950 100464
rect 600006 100408 606556 100464
rect 599945 100406 606556 100408
rect 599945 100403 600011 100406
rect 580625 99378 580691 99381
rect 576380 99376 580691 99378
rect 576380 99320 580630 99376
rect 580686 99320 580691 99376
rect 576380 99318 580691 99320
rect 580625 99315 580691 99318
rect 580441 97746 580507 97749
rect 576380 97744 580507 97746
rect 576380 97688 580446 97744
rect 580502 97688 580507 97744
rect 576380 97686 580507 97688
rect 580441 97683 580507 97686
rect 580717 96250 580783 96253
rect 576380 96248 580783 96250
rect 576380 96192 580722 96248
rect 580778 96192 580783 96248
rect 576380 96190 580783 96192
rect 580717 96187 580783 96190
rect 628281 95978 628347 95981
rect 628238 95976 628347 95978
rect 628238 95920 628286 95976
rect 628342 95920 628347 95976
rect 628238 95915 628347 95920
rect 628238 95404 628298 95915
rect 640517 95706 640583 95709
rect 640517 95704 642466 95706
rect 640517 95648 640522 95704
rect 640578 95648 642466 95704
rect 640517 95646 642466 95648
rect 640517 95643 640583 95646
rect 580533 94754 580599 94757
rect 576380 94752 580599 94754
rect 576380 94696 580538 94752
rect 580594 94696 580599 94752
rect 576380 94694 580599 94696
rect 580533 94691 580599 94694
rect 642406 94588 642466 95646
rect 662086 95508 662092 95572
rect 662156 95570 662162 95572
rect 662229 95570 662295 95573
rect 662156 95568 662295 95570
rect 662156 95512 662234 95568
rect 662290 95512 662295 95568
rect 662156 95510 662295 95512
rect 662156 95508 662162 95510
rect 662229 95507 662295 95510
rect 657353 94754 657419 94757
rect 657310 94752 657419 94754
rect 657310 94696 657358 94752
rect 657414 94696 657419 94752
rect 657310 94691 657419 94696
rect 627913 94482 627979 94485
rect 627913 94480 628268 94482
rect 627913 94424 627918 94480
rect 627974 94424 628268 94480
rect 627913 94422 628268 94424
rect 627913 94419 627979 94422
rect 657310 94180 657370 94691
rect 663241 93802 663307 93805
rect 663198 93800 663307 93802
rect 663198 93744 663246 93800
rect 663302 93744 663307 93800
rect 663198 93739 663307 93744
rect 627269 93530 627335 93533
rect 627269 93528 628268 93530
rect 627269 93472 627274 93528
rect 627330 93472 628268 93528
rect 627269 93470 628268 93472
rect 627269 93467 627335 93470
rect 655329 93394 655395 93397
rect 655329 93392 656788 93394
rect 655329 93336 655334 93392
rect 655390 93336 656788 93392
rect 663198 93364 663258 93739
rect 655329 93334 656788 93336
rect 655329 93331 655395 93334
rect 582281 93258 582347 93261
rect 576380 93256 582347 93258
rect 576380 93200 582286 93256
rect 582342 93200 582347 93256
rect 576380 93198 582347 93200
rect 582281 93195 582347 93198
rect 663425 93122 663491 93125
rect 663382 93120 663491 93122
rect 663382 93064 663430 93120
rect 663486 93064 663491 93120
rect 663382 93059 663491 93064
rect 642725 92714 642791 92717
rect 642725 92712 642834 92714
rect 642725 92656 642730 92712
rect 642786 92656 642834 92712
rect 642725 92651 642834 92656
rect 626441 92578 626507 92581
rect 626441 92576 628268 92578
rect 626441 92520 626446 92576
rect 626502 92520 628268 92576
rect 626441 92518 628268 92520
rect 626441 92515 626507 92518
rect 642774 92140 642834 92651
rect 653949 92578 654015 92581
rect 653949 92576 656788 92578
rect 653949 92520 653954 92576
rect 654010 92520 656788 92576
rect 663382 92548 663442 93059
rect 653949 92518 656788 92520
rect 653949 92515 654015 92518
rect 663517 92306 663583 92309
rect 663517 92304 663626 92306
rect 663517 92248 663522 92304
rect 663578 92248 663626 92304
rect 663517 92243 663626 92248
rect 580809 91762 580875 91765
rect 576380 91760 580875 91762
rect 576380 91704 580814 91760
rect 580870 91704 580875 91760
rect 663566 91732 663626 92243
rect 576380 91702 580875 91704
rect 580809 91699 580875 91702
rect 625889 91626 625955 91629
rect 625889 91624 628268 91626
rect 625889 91568 625894 91624
rect 625950 91568 628268 91624
rect 625889 91566 628268 91568
rect 625889 91563 625955 91566
rect 654041 91490 654107 91493
rect 654041 91488 656788 91490
rect 654041 91432 654046 91488
rect 654102 91432 656788 91488
rect 654041 91430 656788 91432
rect 654041 91427 654107 91430
rect 663517 91082 663583 91085
rect 663517 91080 663626 91082
rect 663517 91024 663522 91080
rect 663578 91024 663626 91080
rect 663517 91019 663626 91024
rect 623957 90674 624023 90677
rect 653121 90674 653187 90677
rect 623957 90672 628268 90674
rect 623957 90616 623962 90672
rect 624018 90616 628268 90672
rect 623957 90614 628268 90616
rect 653121 90672 656788 90674
rect 653121 90616 653126 90672
rect 653182 90616 656788 90672
rect 663566 90644 663626 91019
rect 653121 90614 656788 90616
rect 623957 90611 624023 90614
rect 653121 90611 653187 90614
rect 656985 90402 657051 90405
rect 663609 90402 663675 90405
rect 656942 90400 657051 90402
rect 656942 90344 656990 90400
rect 657046 90344 657051 90400
rect 656942 90339 657051 90344
rect 663566 90400 663675 90402
rect 663566 90344 663614 90400
rect 663670 90344 663675 90400
rect 663566 90339 663675 90344
rect 581821 90266 581887 90269
rect 576380 90264 581887 90266
rect 576380 90208 581826 90264
rect 581882 90208 581887 90264
rect 576380 90206 581887 90208
rect 581821 90203 581887 90206
rect 656942 89828 657002 90339
rect 663566 89828 663626 90339
rect 623773 89722 623839 89725
rect 645853 89722 645919 89725
rect 623773 89720 628268 89722
rect 623773 89664 623778 89720
rect 623834 89664 628268 89720
rect 623773 89662 628268 89664
rect 642988 89720 645919 89722
rect 642988 89664 645858 89720
rect 645914 89664 645919 89720
rect 642988 89662 645919 89664
rect 623773 89659 623839 89662
rect 645853 89659 645919 89662
rect 663425 89586 663491 89589
rect 663382 89584 663491 89586
rect 663382 89528 663430 89584
rect 663486 89528 663491 89584
rect 663382 89523 663491 89528
rect 663382 89012 663442 89523
rect 623221 88906 623287 88909
rect 623221 88904 628268 88906
rect 623221 88848 623226 88904
rect 623282 88848 628268 88904
rect 623221 88846 628268 88848
rect 623221 88843 623287 88846
rect 662137 88772 662203 88773
rect 662086 88708 662092 88772
rect 662156 88770 662203 88772
rect 662156 88768 662248 88770
rect 662198 88712 662248 88768
rect 662156 88710 662248 88712
rect 662156 88708 662203 88710
rect 662137 88707 662203 88708
rect 582097 88634 582163 88637
rect 576380 88632 582163 88634
rect 576380 88576 582102 88632
rect 582158 88576 582163 88632
rect 576380 88574 582163 88576
rect 582097 88571 582163 88574
rect 622485 87954 622551 87957
rect 622485 87952 628268 87954
rect 622485 87896 622490 87952
rect 622546 87896 628268 87952
rect 622485 87894 628268 87896
rect 622485 87891 622551 87894
rect 582005 87138 582071 87141
rect 646037 87138 646103 87141
rect 576380 87136 582071 87138
rect 576380 87080 582010 87136
rect 582066 87080 582071 87136
rect 576380 87078 582071 87080
rect 642988 87136 646103 87138
rect 642988 87080 646042 87136
rect 646098 87080 646103 87136
rect 642988 87078 646103 87080
rect 582005 87075 582071 87078
rect 646037 87075 646103 87078
rect 623405 87002 623471 87005
rect 623405 87000 628268 87002
rect 623405 86944 623410 87000
rect 623466 86944 628268 87000
rect 623405 86942 628268 86944
rect 623405 86939 623471 86942
rect 623497 86050 623563 86053
rect 623497 86048 628268 86050
rect 623497 85992 623502 86048
rect 623558 85992 628268 86048
rect 623497 85990 628268 85992
rect 623497 85987 623563 85990
rect 582189 85642 582255 85645
rect 576380 85640 582255 85642
rect 576380 85584 582194 85640
rect 582250 85584 582255 85640
rect 576380 85582 582255 85584
rect 582189 85579 582255 85582
rect 623313 85098 623379 85101
rect 623313 85096 628268 85098
rect 623313 85040 623318 85096
rect 623374 85040 628268 85096
rect 623313 85038 628268 85040
rect 623313 85035 623379 85038
rect 646129 84690 646195 84693
rect 642988 84688 646195 84690
rect 642988 84632 646134 84688
rect 646190 84632 646195 84688
rect 642988 84630 646195 84632
rect 646129 84627 646195 84630
rect 581913 84146 581979 84149
rect 576380 84144 581979 84146
rect 576380 84088 581918 84144
rect 581974 84088 581979 84144
rect 576380 84086 581979 84088
rect 581913 84083 581979 84086
rect 623129 84146 623195 84149
rect 623129 84144 628268 84146
rect 623129 84088 623134 84144
rect 623190 84088 628268 84144
rect 623129 84086 628268 84088
rect 623129 84083 623195 84086
rect 622117 83194 622183 83197
rect 622117 83192 628268 83194
rect 622117 83136 622122 83192
rect 622178 83136 628268 83192
rect 622117 83134 628268 83136
rect 622117 83131 622183 83134
rect 579613 82650 579679 82653
rect 576380 82648 579679 82650
rect 576380 82592 579618 82648
rect 579674 82592 579679 82648
rect 576380 82590 579679 82592
rect 579613 82587 579679 82590
rect 622301 82242 622367 82245
rect 645945 82242 646011 82245
rect 622301 82240 628268 82242
rect 622301 82184 622306 82240
rect 622362 82184 628268 82240
rect 622301 82182 628268 82184
rect 642988 82240 646011 82242
rect 642988 82184 645950 82240
rect 646006 82184 646011 82240
rect 642988 82182 646011 82184
rect 622301 82179 622367 82182
rect 645945 82179 646011 82182
rect 622485 81426 622551 81429
rect 622485 81424 628268 81426
rect 622485 81368 622490 81424
rect 622546 81368 628268 81424
rect 622485 81366 628268 81368
rect 622485 81363 622551 81366
rect 581453 81154 581519 81157
rect 576380 81152 581519 81154
rect 576380 81096 581458 81152
rect 581514 81096 581519 81152
rect 576380 81094 581519 81096
rect 581453 81091 581519 81094
rect 581269 79522 581335 79525
rect 576380 79520 581335 79522
rect 576380 79464 581274 79520
rect 581330 79464 581335 79520
rect 576380 79462 581335 79464
rect 581269 79459 581335 79462
rect 581729 78026 581795 78029
rect 576380 78024 581795 78026
rect 576380 77968 581734 78024
rect 581790 77968 581795 78024
rect 576380 77966 581795 77968
rect 581729 77963 581795 77966
rect 581361 76530 581427 76533
rect 576380 76528 581427 76530
rect 576380 76472 581366 76528
rect 581422 76472 581427 76528
rect 576380 76470 581427 76472
rect 581361 76467 581427 76470
rect 581637 75034 581703 75037
rect 576380 75032 581703 75034
rect 576380 74976 581642 75032
rect 581698 74976 581703 75032
rect 576380 74974 581703 74976
rect 581637 74971 581703 74974
rect 580942 73538 580948 73540
rect 576380 73478 580948 73538
rect 580942 73476 580948 73478
rect 581012 73476 581018 73540
rect 581545 72042 581611 72045
rect 576380 72040 581611 72042
rect 576380 71984 581550 72040
rect 581606 71984 581611 72040
rect 576380 71982 581611 71984
rect 581545 71979 581611 71982
rect 580993 70410 581059 70413
rect 576380 70408 581059 70410
rect 576380 70352 580998 70408
rect 581054 70352 581059 70408
rect 576380 70350 581059 70352
rect 580993 70347 581059 70350
rect 580717 68914 580783 68917
rect 576380 68912 580783 68914
rect 576380 68856 580722 68912
rect 580778 68856 580783 68912
rect 576380 68854 580783 68856
rect 580717 68851 580783 68854
rect 581177 67418 581243 67421
rect 576380 67416 581243 67418
rect 576380 67360 581182 67416
rect 581238 67360 581243 67416
rect 576380 67358 581243 67360
rect 581177 67355 581243 67358
rect 579613 65922 579679 65925
rect 576380 65920 579679 65922
rect 576380 65864 579618 65920
rect 579674 65864 579679 65920
rect 576380 65862 579679 65864
rect 579613 65859 579679 65862
rect 581085 64426 581151 64429
rect 576380 64424 581151 64426
rect 576380 64368 581090 64424
rect 581146 64368 581151 64424
rect 576380 64366 581151 64368
rect 581085 64363 581151 64366
rect 580809 62930 580875 62933
rect 576380 62928 580875 62930
rect 576380 62872 580814 62928
rect 580870 62872 580875 62928
rect 576380 62870 580875 62872
rect 580809 62867 580875 62870
rect 582189 61298 582255 61301
rect 576380 61296 582255 61298
rect 576380 61240 582194 61296
rect 582250 61240 582255 61296
rect 576380 61238 582255 61240
rect 582189 61235 582255 61238
rect 582097 59802 582163 59805
rect 576380 59800 582163 59802
rect 576380 59744 582102 59800
rect 582158 59744 582163 59800
rect 576380 59742 582163 59744
rect 582097 59739 582163 59742
rect 582281 58306 582347 58309
rect 576380 58304 582347 58306
rect 576380 58248 582286 58304
rect 582342 58248 582347 58304
rect 576380 58246 582347 58248
rect 582281 58243 582347 58246
rect 581821 56810 581887 56813
rect 576380 56808 581887 56810
rect 576380 56752 581826 56808
rect 581882 56752 581887 56808
rect 576380 56750 581887 56752
rect 581821 56747 581887 56750
rect 582005 55314 582071 55317
rect 576380 55312 582071 55314
rect 576380 55256 582010 55312
rect 582066 55256 582071 55312
rect 576380 55254 582071 55256
rect 582005 55251 582071 55254
rect 580901 53818 580967 53821
rect 576380 53816 580967 53818
rect 576380 53760 580906 53816
rect 580962 53760 580967 53816
rect 576380 53758 580967 53760
rect 580901 53755 580967 53758
rect 666553 48514 666619 48517
rect 662094 48512 666619 48514
rect 661480 48456 666558 48512
rect 666614 48456 666619 48512
rect 661480 48454 666619 48456
rect 661480 48452 662154 48454
rect 666553 48451 666619 48454
rect 216121 48242 216187 48245
rect 521694 48242 521700 48244
rect 216121 48240 521700 48242
rect 216121 48184 216126 48240
rect 216182 48184 521700 48240
rect 216121 48182 521700 48184
rect 216121 48179 216187 48182
rect 521694 48180 521700 48182
rect 521764 48180 521770 48244
rect 661174 47565 661234 47761
rect 661125 47560 661234 47565
rect 661125 47504 661130 47560
rect 661186 47504 661234 47560
rect 661125 47502 661234 47504
rect 661125 47499 661191 47502
rect 665173 47426 665239 47429
rect 661388 47424 665239 47426
rect 661388 47368 665178 47424
rect 665234 47368 665239 47424
rect 661388 47366 665239 47368
rect 665173 47363 665239 47366
rect 470133 43618 470199 43621
rect 575841 43618 575907 43621
rect 470133 43616 575907 43618
rect 470133 43560 470138 43616
rect 470194 43560 575846 43616
rect 575902 43560 575907 43616
rect 470133 43558 575907 43560
rect 470133 43555 470199 43558
rect 575841 43555 575907 43558
rect 416589 43482 416655 43485
rect 577957 43482 578023 43485
rect 416589 43480 578023 43482
rect 416589 43424 416594 43480
rect 416650 43424 577962 43480
rect 578018 43424 578023 43480
rect 416589 43422 578023 43424
rect 416589 43419 416655 43422
rect 577957 43419 578023 43422
rect 415393 43346 415459 43349
rect 586421 43346 586487 43349
rect 415393 43344 586487 43346
rect 415393 43288 415398 43344
rect 415454 43288 586426 43344
rect 586482 43288 586487 43344
rect 415393 43286 586487 43288
rect 415393 43283 415459 43286
rect 586421 43283 586487 43286
rect 307293 43210 307359 43213
rect 575657 43210 575723 43213
rect 307293 43208 575723 43210
rect 307293 43152 307298 43208
rect 307354 43152 575662 43208
rect 575718 43152 575723 43208
rect 307293 43150 575723 43152
rect 307293 43147 307359 43150
rect 575657 43147 575723 43150
rect 521745 42124 521811 42125
rect 521694 42060 521700 42124
rect 521764 42122 521811 42124
rect 521764 42120 521856 42122
rect 521806 42064 521856 42120
rect 521764 42062 521856 42064
rect 521764 42060 521811 42062
rect 521745 42059 521811 42060
rect 187601 41850 187667 41853
rect 361941 41850 362007 41853
rect 419993 41850 420059 41853
rect 427905 41850 427971 41853
rect 187601 41848 187710 41850
rect 187601 41792 187606 41848
rect 187662 41792 187710 41848
rect 187601 41787 187710 41792
rect 361941 41848 362050 41850
rect 361941 41792 361946 41848
rect 362002 41792 362050 41848
rect 361941 41787 362050 41792
rect 419993 41848 427971 41850
rect 419993 41792 419998 41848
rect 420054 41792 427910 41848
rect 427966 41792 427971 41848
rect 419993 41790 427971 41792
rect 419993 41787 420059 41790
rect 427905 41787 427971 41790
rect 471697 41850 471763 41853
rect 513281 41850 513347 41853
rect 518525 41850 518591 41853
rect 471697 41848 477510 41850
rect 471697 41792 471702 41848
rect 471758 41792 477510 41848
rect 471697 41790 477510 41792
rect 471697 41787 471763 41790
rect 187650 41306 187710 41787
rect 209773 41306 209839 41309
rect 212441 41306 212507 41309
rect 187650 41304 212507 41306
rect 187650 41248 209778 41304
rect 209834 41248 212446 41304
rect 212502 41248 212507 41304
rect 187650 41246 212507 41248
rect 361990 41306 362050 41787
rect 477450 41442 477510 41790
rect 513281 41848 518591 41850
rect 513281 41792 513286 41848
rect 513342 41792 518530 41848
rect 518586 41792 518591 41848
rect 513281 41790 518591 41792
rect 513281 41787 513347 41790
rect 518525 41787 518591 41790
rect 568573 41442 568639 41445
rect 477450 41440 568639 41442
rect 477450 41384 568578 41440
rect 568634 41384 568639 41440
rect 477450 41382 568639 41384
rect 568573 41379 568639 41382
rect 530301 41306 530367 41309
rect 361990 41304 530367 41306
rect 361990 41248 530306 41304
rect 530362 41248 530367 41304
rect 361990 41246 530367 41248
rect 209773 41243 209839 41246
rect 212441 41243 212507 41246
rect 530301 41243 530367 41246
rect 427905 41170 427971 41173
rect 530393 41170 530459 41173
rect 427905 41168 530459 41170
rect 427905 41112 427910 41168
rect 427966 41112 530398 41168
rect 530454 41112 530459 41168
rect 427905 41110 530459 41112
rect 427905 41107 427971 41110
rect 530393 41107 530459 41110
rect 475469 41034 475535 41037
rect 549253 41034 549319 41037
rect 475469 41032 549319 41034
rect 475469 40976 475474 41032
rect 475530 40976 549258 41032
rect 549314 40976 549319 41032
rect 475469 40974 549319 40976
rect 475469 40971 475535 40974
rect 549253 40971 549319 40974
rect 230933 16690 230999 16693
rect 225676 16688 230999 16690
rect 225676 16632 230938 16688
rect 230994 16632 230999 16688
rect 225676 16630 230999 16632
rect 230933 16627 230999 16630
rect 230749 15194 230815 15197
rect 225676 15192 230815 15194
rect 225676 15136 230754 15192
rect 230810 15136 230815 15192
rect 225676 15134 230815 15136
rect 230749 15131 230815 15134
rect 230657 13698 230723 13701
rect 225676 13696 230723 13698
rect 225676 13640 230662 13696
rect 230718 13640 230723 13696
rect 225676 13638 230723 13640
rect 230657 13635 230723 13638
rect 230841 12202 230907 12205
rect 225676 12200 230907 12202
rect 225676 12144 230846 12200
rect 230902 12144 230907 12200
rect 225676 12142 230907 12144
rect 230841 12139 230907 12142
rect 230381 10706 230447 10709
rect 225676 10704 230447 10706
rect 225676 10648 230386 10704
rect 230442 10648 230447 10704
rect 225676 10646 230447 10648
rect 230381 10643 230447 10646
rect 230565 9210 230631 9213
rect 225676 9208 230631 9210
rect 225676 9152 230570 9208
rect 230626 9152 230631 9208
rect 225676 9150 230631 9152
rect 230565 9147 230631 9150
rect 230473 7714 230539 7717
rect 225676 7712 230539 7714
rect 225676 7656 230478 7712
rect 230534 7656 230539 7712
rect 225676 7654 230539 7656
rect 230473 7651 230539 7654
rect 229369 6218 229435 6221
rect 225676 6216 229435 6218
rect 225676 6160 229374 6216
rect 229430 6160 229435 6216
rect 225676 6158 229435 6160
rect 229369 6155 229435 6158
<< via3 >>
rect 221400 993820 234879 995620
rect 240878 993820 254357 995620
rect 274000 993820 287479 995620
rect 293478 993820 306957 995620
rect 375800 993820 389279 995620
rect 395278 993820 408757 995620
rect 679204 886620 679268 886684
rect 679204 885804 679268 885868
rect 679204 884988 679268 885052
rect 41828 807876 41892 807940
rect 41828 795016 41892 795020
rect 41828 794960 41878 795016
rect 41878 794960 41892 795016
rect 41828 794956 41892 794960
rect 674972 788292 675036 788356
rect 674604 787204 674668 787268
rect 674788 786660 674852 786724
rect 676812 745316 676876 745380
rect 676628 745180 676692 745244
rect 674052 742868 674116 742932
rect 673868 742460 673932 742524
rect 674236 741644 674300 741708
rect 675156 739740 675220 739804
rect 673684 739060 673748 739124
rect 674420 738652 674484 738716
rect 675340 738032 675404 738036
rect 675340 737976 675390 738032
rect 675390 737976 675404 738032
rect 675340 737972 675404 737976
rect 673500 730764 673564 730828
rect 674604 730764 674668 730828
rect 674604 711996 674668 712060
rect 674788 711180 674852 711244
rect 673500 709548 673564 709612
rect 676076 707236 676140 707300
rect 676076 706828 676140 706892
rect 676996 699348 677060 699412
rect 676812 699212 676876 699276
rect 673500 698260 673564 698324
rect 676076 697172 676140 697236
rect 674972 695540 675036 695604
rect 674604 694724 674668 694788
rect 674788 694588 674852 694652
rect 677180 692956 677244 693020
rect 676628 690100 676692 690164
rect 673868 687108 673932 687172
rect 674052 685748 674116 685812
rect 674236 680308 674300 680372
rect 674972 680308 675036 680372
rect 676628 680308 676692 680372
rect 677364 680308 677428 680372
rect 30604 678948 30668 679012
rect 674052 678812 674116 678876
rect 676076 677968 676140 677972
rect 676076 677912 676126 677968
rect 676126 677912 676140 677968
rect 676076 677908 676140 677912
rect 60780 676500 60844 676564
rect 676076 676472 676140 676476
rect 676076 676416 676126 676472
rect 676126 676416 676140 676472
rect 676076 676412 676140 676416
rect 30604 676016 30668 676020
rect 30604 675960 30618 676016
rect 30618 675960 30668 676016
rect 30604 675956 30668 675960
rect 674236 674052 674300 674116
rect 674972 674052 675036 674116
rect 42564 670652 42628 670716
rect 676628 668612 676692 668676
rect 675156 665620 675220 665684
rect 42564 665076 42628 665140
rect 673684 663988 673748 664052
rect 674420 663580 674484 663644
rect 675708 662356 675772 662420
rect 676996 662084 677060 662148
rect 676812 661676 676876 661740
rect 673868 652836 673932 652900
rect 674052 652156 674116 652220
rect 674236 651612 674300 651676
rect 675156 649164 675220 649228
rect 674972 633056 675036 633120
rect 676076 633056 676140 633120
rect 42380 627464 42444 627468
rect 42380 627408 42430 627464
rect 42430 627408 42444 627464
rect 42380 627404 42444 627408
rect 43484 626996 43548 627060
rect 676628 624412 676692 624476
rect 43484 622100 43548 622164
rect 674788 621828 674852 621892
rect 673500 621012 673564 621076
rect 42380 620936 42444 620940
rect 42380 620880 42394 620936
rect 42394 620880 42444 620936
rect 42380 620876 42444 620880
rect 674420 620604 674484 620668
rect 674972 619380 675036 619444
rect 674604 618972 674668 619036
rect 677180 617476 677244 617540
rect 677364 617068 677428 617132
rect 677180 610132 677244 610196
rect 677364 609996 677428 610060
rect 673684 608092 673748 608156
rect 673500 607276 673564 607340
rect 674788 605100 674852 605164
rect 674972 604964 675036 605028
rect 674604 604420 674668 604484
rect 674420 601836 674484 601900
rect 43116 585304 43180 585308
rect 43116 585248 43130 585304
rect 43130 585248 43180 585304
rect 43116 585244 43180 585248
rect 43116 581360 43180 581364
rect 43116 581304 43130 581360
rect 43130 581304 43180 581360
rect 43116 581300 43180 581304
rect 676076 579260 676140 579324
rect 676628 577628 676692 577692
rect 676812 576812 676876 576876
rect 674236 576540 674300 576604
rect 673868 575724 673932 575788
rect 674052 574092 674116 574156
rect 675156 573684 675220 573748
rect 677180 571916 677244 571980
rect 676996 571508 677060 571572
rect 677364 571508 677428 571572
rect 674052 562668 674116 562732
rect 675156 562260 675220 562324
rect 674236 561172 674300 561236
rect 42564 556004 42628 556068
rect 675340 554976 675404 554980
rect 675340 554920 675354 554976
rect 675354 554920 675404 554976
rect 675340 554916 675404 554920
rect 675340 554644 675404 554708
rect 41644 553828 41708 553892
rect 42932 553148 42996 553212
rect 42196 552740 42260 552804
rect 42380 552332 42444 552396
rect 42012 551516 42076 551580
rect 41460 550972 41524 551036
rect 41828 550700 41892 550764
rect 674420 546484 674484 546548
rect 39988 546348 40052 546412
rect 674604 543628 674668 543692
rect 673500 543492 673564 543556
rect 676076 543288 676140 543352
rect 675892 539616 675956 539620
rect 675892 539560 675942 539616
rect 675942 539560 675956 539616
rect 675892 539556 675956 539560
rect 42380 538732 42444 538796
rect 41828 535740 41892 535804
rect 675892 534924 675956 534988
rect 673684 533836 673748 533900
rect 676628 533428 676692 533492
rect 42196 533020 42260 533084
rect 674972 533020 675036 533084
rect 41644 532884 41708 532948
rect 41460 532748 41524 532812
rect 674788 532748 674852 532812
rect 676812 532612 676876 532676
rect 42932 530708 42996 530772
rect 42012 530164 42076 530228
rect 676996 526900 677060 526964
rect 674052 491404 674116 491468
rect 674236 491268 674300 491332
rect 675156 485148 675220 485212
rect 42564 455908 42628 455972
rect 42380 450800 42444 450804
rect 42380 450744 42430 450800
rect 42430 450744 42444 450800
rect 42380 450740 42444 450744
rect 42380 445904 42444 445908
rect 42380 445848 42430 445904
rect 42430 445848 42444 445904
rect 42380 445844 42444 445848
rect 42380 440736 42444 440740
rect 42380 440680 42430 440736
rect 42430 440680 42444 440736
rect 42380 440676 42444 440680
rect 42380 428844 42444 428908
rect 675156 402188 675220 402252
rect 674972 400556 675036 400620
rect 674788 399740 674852 399804
rect 675156 357444 675220 357508
rect 674972 355812 675036 355876
rect 674788 354996 674852 355060
rect 41644 338948 41708 339012
rect 42012 338812 42076 338876
rect 41828 337588 41892 337652
rect 42196 329700 42260 329764
rect 42012 315616 42076 315620
rect 42012 315560 42026 315616
rect 42026 315560 42076 315616
rect 42012 315556 42076 315560
rect 42196 313848 42260 313852
rect 42196 313792 42210 313848
rect 42210 313792 42260 313848
rect 42196 313788 42260 313792
rect 41828 313168 41892 313172
rect 41828 313112 41842 313168
rect 41842 313112 41892 313168
rect 41828 313108 41892 313112
rect 41644 312292 41708 312356
rect 41828 296788 41892 296852
rect 60780 275980 60844 276044
rect 41644 270404 41708 270468
rect 675156 264556 675220 264620
rect 41644 252588 41708 252652
rect 41644 225932 41708 225996
rect 675156 219812 675220 219876
rect 41644 204852 41708 204916
rect 41460 204444 41524 204508
rect 41828 198732 41892 198796
rect 41828 184240 41892 184244
rect 41828 184184 41878 184240
rect 41878 184184 41892 184240
rect 41828 184180 41892 184184
rect 41644 183364 41708 183428
rect 41460 182684 41524 182748
rect 580948 113188 581012 113252
rect 662092 95508 662156 95572
rect 662092 88768 662156 88772
rect 662092 88712 662142 88768
rect 662142 88712 662156 88768
rect 662092 88708 662156 88712
rect 580948 73476 581012 73540
rect 521700 48180 521764 48244
rect 521700 42120 521764 42124
rect 521700 42064 521750 42120
rect 521750 42064 521764 42120
rect 521700 42060 521764 42064
<< metal4 >>
rect 221000 995620 235279 996020
rect 221000 993820 221400 995620
rect 234879 993820 235279 995620
rect 221000 993420 235279 993820
tri 221000 983518 230902 993420 ne
rect 230902 983518 235279 993420
rect 240478 995620 254757 996020
rect 240478 993820 240878 995620
rect 254357 993820 254757 995620
rect 273600 995620 287879 996020
rect 273600 993820 274000 995620
rect 287479 993820 287879 995620
rect 240478 992116 254800 993820
rect 240478 984242 246202 992116
tri 240478 983518 241202 984242 ne
rect 230902 982718 235902 983518
rect 241202 982718 246202 984242
tri 246202 983518 254800 992116 nw
rect 273600 992520 287879 993820
tri 273600 983518 282602 992520 ne
rect 282602 983795 287879 992520
rect 282602 982718 287602 983795
tri 287602 983518 287879 983795 nw
rect 293078 995620 307357 996020
rect 293078 993820 293478 995620
rect 306957 993820 307357 995620
rect 375400 995620 389679 996020
rect 375400 993820 375800 995620
rect 389279 993820 389679 995620
rect 293078 993016 307400 993820
rect 293078 983518 297902 993016
tri 297902 983518 307400 993016 nw
rect 375400 992420 389679 993820
tri 375400 983518 384302 992420 ne
rect 384302 983895 389679 992420
rect 292902 982718 297902 983518
rect 384302 982718 389302 983895
tri 389302 983518 389679 983895 nw
rect 394878 995620 409157 996020
rect 394878 993820 395278 995620
rect 408757 993820 409157 995620
rect 394878 993116 409200 993820
rect 394878 983518 399602 993116
tri 399602 983518 409200 993116 nw
rect 394602 982718 399602 983518
rect 679203 886684 679269 886685
rect 679203 886620 679204 886684
rect 679268 886620 679269 886684
rect 679203 886619 679269 886620
rect 679206 885869 679266 886619
rect 679203 885868 679269 885869
rect 679203 885804 679204 885868
rect 679268 885804 679269 885868
rect 679203 885803 679269 885804
rect 679206 885053 679266 885803
rect 679203 885052 679269 885053
rect 679203 884988 679204 885052
rect 679268 884988 679269 885052
rect 679203 884987 679269 884988
rect 41827 807940 41893 807941
rect 41827 807876 41828 807940
rect 41892 807876 41893 807940
rect 41827 807875 41893 807876
rect 41830 795021 41890 807875
rect 41827 795020 41893 795021
rect 41827 794956 41828 795020
rect 41892 794956 41893 795020
rect 41827 794955 41893 794956
rect 674971 788356 675037 788357
rect 674971 788292 674972 788356
rect 675036 788292 675037 788356
rect 674971 788291 675037 788292
rect 674603 787268 674669 787269
rect 674603 787204 674604 787268
rect 674668 787204 674669 787268
rect 674603 787203 674669 787204
rect 674051 742932 674117 742933
rect 674051 742868 674052 742932
rect 674116 742868 674117 742932
rect 674051 742867 674117 742868
rect 673867 742524 673933 742525
rect 673867 742460 673868 742524
rect 673932 742460 673933 742524
rect 673867 742459 673933 742460
rect 673683 739124 673749 739125
rect 673683 739060 673684 739124
rect 673748 739060 673749 739124
rect 673683 739059 673749 739060
rect 673499 730828 673565 730829
rect 673499 730764 673500 730828
rect 673564 730764 673565 730828
rect 673499 730763 673565 730764
rect 673502 709613 673562 730763
rect 673499 709612 673565 709613
rect 673499 709548 673500 709612
rect 673564 709548 673565 709612
rect 673499 709547 673565 709548
rect 673499 698324 673565 698325
rect 673499 698260 673500 698324
rect 673564 698260 673565 698324
rect 673499 698259 673565 698260
rect 30603 679012 30669 679013
rect 30603 678948 30604 679012
rect 30668 678948 30669 679012
rect 30603 678947 30669 678948
rect 30606 676021 30666 678947
rect 60779 676564 60845 676565
rect 60779 676500 60780 676564
rect 60844 676500 60845 676564
rect 60779 676499 60845 676500
rect 30603 676020 30669 676021
rect 30603 675956 30604 676020
rect 30668 675956 30669 676020
rect 30603 675955 30669 675956
rect 42563 670716 42629 670717
rect 42563 670652 42564 670716
rect 42628 670652 42629 670716
rect 42563 670651 42629 670652
rect 42566 665141 42626 670651
rect 42563 665140 42629 665141
rect 42563 665076 42564 665140
rect 42628 665076 42629 665140
rect 42563 665075 42629 665076
rect 42379 627468 42445 627469
rect 42379 627404 42380 627468
rect 42444 627404 42445 627468
rect 42379 627403 42445 627404
rect 42382 620941 42442 627403
rect 43483 627060 43549 627061
rect 43483 626996 43484 627060
rect 43548 626996 43549 627060
rect 43483 626995 43549 626996
rect 43486 622165 43546 626995
rect 43483 622164 43549 622165
rect 43483 622100 43484 622164
rect 43548 622100 43549 622164
rect 43483 622099 43549 622100
rect 42379 620940 42445 620941
rect 42379 620876 42380 620940
rect 42444 620876 42445 620940
rect 42379 620875 42445 620876
rect 43115 585308 43181 585309
rect 43115 585244 43116 585308
rect 43180 585244 43181 585308
rect 43115 585243 43181 585244
rect 43118 581365 43178 585243
rect 43115 581364 43181 581365
rect 43115 581300 43116 581364
rect 43180 581300 43181 581364
rect 43115 581299 43181 581300
rect 42563 556068 42629 556069
rect 42563 556004 42564 556068
rect 42628 556004 42629 556068
rect 42563 556003 42629 556004
rect 41643 553892 41709 553893
rect 41643 553828 41644 553892
rect 41708 553828 41709 553892
rect 41643 553827 41709 553828
rect 41459 551036 41525 551037
rect 41459 550972 41460 551036
rect 41524 550972 41525 551036
rect 41459 550971 41525 550972
rect 39987 546412 40053 546413
rect 39987 546348 39988 546412
rect 40052 546348 40053 546412
rect 39987 546347 40053 546348
rect 39990 462329 40050 546347
rect 41462 532813 41522 550971
rect 41646 532949 41706 553827
rect 42195 552804 42261 552805
rect 42195 552740 42196 552804
rect 42260 552740 42261 552804
rect 42195 552739 42261 552740
rect 42011 551580 42077 551581
rect 42011 551516 42012 551580
rect 42076 551516 42077 551580
rect 42011 551515 42077 551516
rect 41827 550764 41893 550765
rect 41827 550700 41828 550764
rect 41892 550700 41893 550764
rect 41827 550699 41893 550700
rect 41830 535805 41890 550699
rect 41827 535804 41893 535805
rect 41827 535740 41828 535804
rect 41892 535740 41893 535804
rect 41827 535739 41893 535740
rect 41643 532948 41709 532949
rect 41643 532884 41644 532948
rect 41708 532884 41709 532948
rect 41643 532883 41709 532884
rect 41459 532812 41525 532813
rect 41459 532748 41460 532812
rect 41524 532748 41525 532812
rect 41459 532747 41525 532748
rect 42014 530229 42074 551515
rect 42198 533085 42258 552739
rect 42379 552396 42445 552397
rect 42379 552332 42380 552396
rect 42444 552332 42445 552396
rect 42379 552331 42445 552332
rect 42382 538797 42442 552331
rect 42379 538796 42445 538797
rect 42379 538732 42380 538796
rect 42444 538732 42445 538796
rect 42379 538731 42445 538732
rect 42195 533084 42261 533085
rect 42195 533020 42196 533084
rect 42260 533020 42261 533084
rect 42195 533019 42261 533020
rect 42011 530228 42077 530229
rect 42011 530164 42012 530228
rect 42076 530164 42077 530228
rect 42011 530163 42077 530164
rect 42566 455973 42626 556003
rect 42931 553212 42997 553213
rect 42931 553148 42932 553212
rect 42996 553148 42997 553212
rect 42931 553147 42997 553148
rect 42934 530773 42994 553147
rect 42931 530772 42997 530773
rect 42931 530708 42932 530772
rect 42996 530708 42997 530772
rect 42931 530707 42997 530708
rect 42563 455972 42629 455973
rect 42563 455908 42564 455972
rect 42628 455908 42629 455972
rect 42563 455907 42629 455908
rect 42379 450804 42445 450805
rect 42379 450740 42380 450804
rect 42444 450740 42445 450804
rect 42379 450739 42445 450740
rect 42382 445909 42442 450739
rect 42379 445908 42445 445909
rect 42379 445844 42380 445908
rect 42444 445844 42445 445908
rect 42379 445843 42445 445844
rect 42379 440740 42445 440741
rect 42379 440676 42380 440740
rect 42444 440676 42445 440740
rect 42379 440675 42445 440676
rect 42382 428909 42442 440675
rect 42379 428908 42445 428909
rect 42379 428844 42380 428908
rect 42444 428844 42445 428908
rect 42379 428843 42445 428844
rect 41643 339012 41709 339013
rect 41643 338948 41644 339012
rect 41708 338948 41709 339012
rect 41643 338947 41709 338948
rect 41646 312357 41706 338947
rect 42011 338876 42077 338877
rect 42011 338812 42012 338876
rect 42076 338812 42077 338876
rect 42011 338811 42077 338812
rect 41827 337652 41893 337653
rect 41827 337588 41828 337652
rect 41892 337588 41893 337652
rect 41827 337587 41893 337588
rect 41830 313173 41890 337587
rect 42014 315621 42074 338811
rect 42195 329764 42261 329765
rect 42195 329700 42196 329764
rect 42260 329700 42261 329764
rect 42195 329699 42261 329700
rect 42011 315620 42077 315621
rect 42011 315556 42012 315620
rect 42076 315556 42077 315620
rect 42011 315555 42077 315556
rect 42198 313853 42258 329699
rect 42195 313852 42261 313853
rect 42195 313788 42196 313852
rect 42260 313788 42261 313852
rect 42195 313787 42261 313788
rect 41827 313172 41893 313173
rect 41827 313108 41828 313172
rect 41892 313108 41893 313172
rect 41827 313107 41893 313108
rect 41643 312356 41709 312357
rect 41643 312292 41644 312356
rect 41708 312292 41709 312356
rect 41643 312291 41709 312292
rect 41827 296852 41893 296853
rect 41827 296850 41828 296852
rect 41646 296790 41828 296850
rect 41646 270469 41706 296790
rect 41827 296788 41828 296790
rect 41892 296788 41893 296852
rect 41827 296787 41893 296788
rect 60782 276045 60842 676499
rect 673502 621077 673562 698259
rect 673686 664053 673746 739059
rect 673870 687173 673930 742459
rect 673867 687172 673933 687173
rect 673867 687108 673868 687172
rect 673932 687108 673933 687172
rect 673867 687107 673933 687108
rect 674054 685813 674114 742867
rect 674235 741708 674301 741709
rect 674235 741644 674236 741708
rect 674300 741644 674301 741708
rect 674235 741643 674301 741644
rect 674051 685812 674117 685813
rect 674051 685748 674052 685812
rect 674116 685748 674117 685812
rect 674051 685747 674117 685748
rect 674238 681050 674298 741643
rect 674419 738716 674485 738717
rect 674419 738652 674420 738716
rect 674484 738652 674485 738716
rect 674419 738651 674485 738652
rect 674054 680990 674298 681050
rect 674054 678877 674114 680990
rect 674235 680372 674301 680373
rect 674235 680308 674236 680372
rect 674300 680308 674301 680372
rect 674235 680307 674301 680308
rect 674051 678876 674117 678877
rect 674051 678812 674052 678876
rect 674116 678812 674117 678876
rect 674051 678811 674117 678812
rect 674238 674117 674298 680307
rect 674235 674116 674301 674117
rect 674235 674052 674236 674116
rect 674300 674052 674301 674116
rect 674235 674051 674301 674052
rect 673683 664052 673749 664053
rect 673683 663988 673684 664052
rect 673748 663988 673749 664052
rect 673683 663987 673749 663988
rect 674422 663645 674482 738651
rect 674606 730829 674666 787203
rect 674787 786724 674853 786725
rect 674787 786660 674788 786724
rect 674852 786660 674853 786724
rect 674787 786659 674853 786660
rect 674603 730828 674669 730829
rect 674603 730764 674604 730828
rect 674668 730764 674669 730828
rect 674603 730763 674669 730764
rect 674790 730690 674850 786659
rect 674606 730630 674850 730690
rect 674606 712061 674666 730630
rect 674974 730010 675034 788291
rect 676811 745380 676877 745381
rect 676811 745316 676812 745380
rect 676876 745316 676877 745380
rect 676811 745315 676877 745316
rect 676627 745244 676693 745245
rect 676627 745180 676628 745244
rect 676692 745180 676693 745244
rect 676627 745179 676693 745180
rect 675155 739804 675221 739805
rect 675155 739740 675156 739804
rect 675220 739740 675221 739804
rect 675155 739739 675221 739740
rect 674790 729950 675034 730010
rect 674603 712060 674669 712061
rect 674603 711996 674604 712060
rect 674668 711996 674669 712060
rect 674603 711995 674669 711996
rect 674790 711245 674850 729950
rect 675158 729330 675218 739739
rect 675339 738036 675405 738037
rect 675339 737972 675340 738036
rect 675404 737972 675405 738036
rect 675339 737971 675405 737972
rect 674974 729270 675218 729330
rect 674787 711244 674853 711245
rect 674787 711180 674788 711244
rect 674852 711180 674853 711244
rect 674787 711179 674853 711180
rect 674974 709350 675034 729270
rect 675342 728650 675402 737971
rect 675158 728590 675402 728650
rect 675158 719130 675218 728590
rect 676630 723227 676690 745179
rect 676630 723151 676720 723227
rect 676660 721626 676720 723151
rect 676630 721549 676720 721626
rect 675158 719070 675770 719130
rect 674974 709290 675218 709350
rect 674971 695604 675037 695605
rect 674971 695540 674972 695604
rect 675036 695540 675037 695604
rect 674971 695539 675037 695540
rect 674603 694788 674669 694789
rect 674603 694724 674604 694788
rect 674668 694724 674669 694788
rect 674603 694723 674669 694724
rect 674419 663644 674485 663645
rect 674419 663580 674420 663644
rect 674484 663580 674485 663644
rect 674419 663579 674485 663580
rect 673867 652900 673933 652901
rect 673867 652836 673868 652900
rect 673932 652836 673933 652900
rect 673867 652835 673933 652836
rect 673499 621076 673565 621077
rect 673499 621012 673500 621076
rect 673564 621012 673565 621076
rect 673499 621011 673565 621012
rect 673683 608156 673749 608157
rect 673683 608092 673684 608156
rect 673748 608092 673749 608156
rect 673683 608091 673749 608092
rect 673499 607340 673565 607341
rect 673499 607276 673500 607340
rect 673564 607276 673565 607340
rect 673499 607275 673565 607276
rect 673502 543557 673562 607275
rect 673499 543556 673565 543557
rect 673499 543492 673500 543556
rect 673564 543492 673565 543556
rect 673499 543491 673565 543492
rect 673686 533901 673746 608091
rect 673870 575789 673930 652835
rect 674051 652220 674117 652221
rect 674051 652156 674052 652220
rect 674116 652156 674117 652220
rect 674051 652155 674117 652156
rect 673867 575788 673933 575789
rect 673867 575724 673868 575788
rect 673932 575724 673933 575788
rect 673867 575723 673933 575724
rect 674054 574157 674114 652155
rect 674235 651676 674301 651677
rect 674235 651612 674236 651676
rect 674300 651612 674301 651676
rect 674235 651611 674301 651612
rect 674238 576605 674298 651611
rect 674606 651390 674666 694723
rect 674787 694652 674853 694653
rect 674787 694588 674788 694652
rect 674852 694588 674853 694652
rect 674787 694587 674853 694588
rect 674422 651330 674666 651390
rect 674422 620669 674482 651330
rect 674790 641610 674850 694587
rect 674974 680373 675034 695539
rect 674971 680372 675037 680373
rect 674971 680308 674972 680372
rect 675036 680308 675037 680372
rect 674971 680307 675037 680308
rect 675158 678650 675218 709290
rect 675710 681750 675770 719070
rect 676630 707570 676690 721549
rect 676078 707510 676690 707570
rect 676078 707301 676138 707510
rect 676075 707300 676141 707301
rect 676075 707236 676076 707300
rect 676140 707236 676141 707300
rect 676075 707235 676141 707236
rect 676075 706892 676141 706893
rect 676075 706828 676076 706892
rect 676140 706890 676141 706892
rect 676814 706890 676874 745315
rect 676140 706830 676874 706890
rect 676140 706828 676141 706830
rect 676075 706827 676141 706828
rect 676995 699412 677061 699413
rect 676995 699348 676996 699412
rect 677060 699348 677061 699412
rect 676995 699347 677061 699348
rect 676811 699276 676877 699277
rect 676811 699212 676812 699276
rect 676876 699212 676877 699276
rect 676811 699211 676877 699212
rect 676075 697236 676141 697237
rect 676075 697172 676076 697236
rect 676140 697172 676141 697236
rect 676075 697171 676141 697172
rect 674974 678590 675218 678650
rect 675342 681690 675770 681750
rect 674974 675250 675034 678590
rect 675342 677970 675402 681690
rect 676078 677973 676138 697171
rect 676627 690164 676693 690165
rect 676627 690100 676628 690164
rect 676692 690100 676693 690164
rect 676627 690099 676693 690100
rect 676630 680373 676690 690099
rect 676627 680372 676693 680373
rect 676627 680308 676628 680372
rect 676692 680308 676693 680372
rect 676627 680307 676693 680308
rect 675158 677910 675402 677970
rect 676075 677972 676141 677973
rect 675158 675930 675218 677910
rect 676075 677908 676076 677972
rect 676140 677908 676141 677972
rect 676075 677907 676141 677908
rect 676075 676476 676141 676477
rect 676075 676412 676076 676476
rect 676140 676412 676141 676476
rect 676075 676411 676141 676412
rect 675158 675870 675770 675930
rect 674974 675190 675218 675250
rect 674971 674116 675037 674117
rect 674971 674052 674972 674116
rect 675036 674052 675037 674116
rect 674971 674051 675037 674052
rect 674606 641550 674850 641610
rect 674419 620668 674485 620669
rect 674419 620604 674420 620668
rect 674484 620604 674485 620668
rect 674419 620603 674485 620604
rect 674606 619037 674666 641550
rect 674974 633770 675034 674051
rect 675158 665685 675218 675190
rect 675155 665684 675221 665685
rect 675155 665620 675156 665684
rect 675220 665620 675221 665684
rect 675155 665619 675221 665620
rect 675710 662421 675770 675870
rect 675707 662420 675773 662421
rect 675707 662356 675708 662420
rect 675772 662356 675773 662420
rect 675707 662355 675773 662356
rect 675155 649228 675221 649229
rect 675155 649164 675156 649228
rect 675220 649164 675221 649228
rect 675155 649163 675221 649164
rect 674790 633710 675034 633770
rect 674790 621893 674850 633710
rect 674971 633120 675037 633121
rect 674971 633056 674972 633120
rect 675036 633056 675037 633120
rect 674971 633055 675037 633056
rect 674787 621892 674853 621893
rect 674787 621828 674788 621892
rect 674852 621828 674853 621892
rect 674787 621827 674853 621828
rect 674974 619445 675034 633055
rect 674971 619444 675037 619445
rect 674971 619380 674972 619444
rect 675036 619380 675037 619444
rect 674971 619379 675037 619380
rect 674603 619036 674669 619037
rect 674603 618972 674604 619036
rect 674668 618972 674669 619036
rect 674603 618971 674669 618972
rect 674787 605164 674853 605165
rect 674787 605100 674788 605164
rect 674852 605100 674853 605164
rect 674787 605099 674853 605100
rect 674603 604484 674669 604485
rect 674603 604420 674604 604484
rect 674668 604420 674669 604484
rect 674603 604419 674669 604420
rect 674419 601900 674485 601901
rect 674419 601836 674420 601900
rect 674484 601836 674485 601900
rect 674419 601835 674485 601836
rect 674235 576604 674301 576605
rect 674235 576540 674236 576604
rect 674300 576540 674301 576604
rect 674235 576539 674301 576540
rect 674051 574156 674117 574157
rect 674051 574092 674052 574156
rect 674116 574092 674117 574156
rect 674051 574091 674117 574092
rect 674051 562732 674117 562733
rect 674051 562668 674052 562732
rect 674116 562668 674117 562732
rect 674051 562667 674117 562668
rect 673683 533900 673749 533901
rect 673683 533836 673684 533900
rect 673748 533836 673749 533900
rect 673683 533835 673749 533836
rect 674054 491469 674114 562667
rect 674235 561236 674301 561237
rect 674235 561172 674236 561236
rect 674300 561172 674301 561236
rect 674235 561171 674301 561172
rect 674051 491468 674117 491469
rect 674051 491404 674052 491468
rect 674116 491404 674117 491468
rect 674051 491403 674117 491404
rect 674238 491333 674298 561171
rect 674422 546549 674482 601835
rect 674419 546548 674485 546549
rect 674419 546484 674420 546548
rect 674484 546484 674485 546548
rect 674419 546483 674485 546484
rect 674606 543693 674666 604419
rect 674603 543692 674669 543693
rect 674603 543628 674604 543692
rect 674668 543628 674669 543692
rect 674603 543627 674669 543628
rect 674790 532813 674850 605099
rect 674971 605028 675037 605029
rect 674971 604964 674972 605028
rect 675036 604964 675037 605028
rect 674971 604963 675037 604964
rect 674974 533085 675034 604963
rect 675158 573749 675218 649163
rect 676078 633121 676138 676411
rect 676627 668676 676693 668677
rect 676627 668612 676628 668676
rect 676692 668612 676693 668676
rect 676627 668611 676693 668612
rect 676630 633131 676690 668611
rect 676814 661741 676874 699211
rect 676998 662149 677058 699347
rect 677179 693020 677245 693021
rect 677179 692956 677180 693020
rect 677244 692956 677245 693020
rect 677179 692955 677245 692956
rect 676995 662148 677061 662149
rect 676995 662084 676996 662148
rect 677060 662084 677061 662148
rect 676995 662083 677061 662084
rect 676811 661740 676877 661741
rect 676811 661676 676812 661740
rect 676876 661676 676877 661740
rect 676811 661675 676877 661676
rect 676075 633120 676141 633121
rect 676075 633056 676076 633120
rect 676140 633056 676141 633120
rect 676630 633056 676730 633131
rect 676075 633055 676141 633056
rect 676670 631304 676730 633056
rect 676630 631227 676730 631304
rect 676630 624477 676690 631227
rect 676627 624476 676693 624477
rect 676627 624412 676628 624476
rect 676692 624412 676693 624476
rect 676627 624411 676693 624412
rect 677182 617541 677242 692955
rect 677363 680372 677429 680373
rect 677363 680308 677364 680372
rect 677428 680308 677429 680372
rect 677363 680307 677429 680308
rect 677179 617540 677245 617541
rect 677179 617476 677180 617540
rect 677244 617476 677245 617540
rect 677179 617475 677245 617476
rect 677366 617133 677426 680307
rect 677363 617132 677429 617133
rect 677363 617068 677364 617132
rect 677428 617068 677429 617132
rect 677363 617067 677429 617068
rect 677179 610196 677245 610197
rect 677179 610132 677180 610196
rect 677244 610132 677245 610196
rect 677179 610131 677245 610132
rect 676075 579324 676141 579325
rect 676075 579260 676076 579324
rect 676140 579260 676141 579324
rect 676075 579259 676141 579260
rect 675155 573748 675221 573749
rect 675155 573684 675156 573748
rect 675220 573684 675221 573748
rect 675155 573683 675221 573684
rect 675155 562324 675221 562325
rect 675155 562260 675156 562324
rect 675220 562260 675221 562324
rect 675155 562259 675221 562260
rect 674971 533084 675037 533085
rect 674971 533020 674972 533084
rect 675036 533020 675037 533084
rect 674971 533019 675037 533020
rect 674787 532812 674853 532813
rect 674787 532748 674788 532812
rect 674852 532748 674853 532812
rect 674787 532747 674853 532748
rect 674235 491332 674301 491333
rect 674235 491268 674236 491332
rect 674300 491268 674301 491332
rect 674235 491267 674301 491268
rect 675158 485213 675218 562259
rect 675339 554980 675405 554981
rect 675339 554916 675340 554980
rect 675404 554916 675405 554980
rect 675339 554915 675405 554916
rect 675342 554709 675402 554915
rect 675339 554708 675405 554709
rect 675339 554644 675340 554708
rect 675404 554644 675405 554708
rect 675339 554643 675405 554644
rect 676078 543353 676138 579259
rect 676627 577692 676693 577693
rect 676627 577628 676628 577692
rect 676692 577628 676693 577692
rect 676627 577627 676693 577628
rect 676075 543352 676141 543353
rect 676075 543288 676076 543352
rect 676140 543288 676141 543352
rect 676075 543287 676141 543288
rect 676630 542911 676690 577627
rect 676811 576876 676877 576877
rect 676811 576812 676812 576876
rect 676876 576812 676877 576876
rect 676811 576811 676877 576812
rect 676630 542822 676710 542911
rect 676650 541027 676710 542822
rect 676630 540938 676710 541027
rect 675891 539620 675957 539621
rect 675891 539556 675892 539620
rect 675956 539556 675957 539620
rect 675891 539555 675957 539556
rect 675894 534989 675954 539555
rect 675891 534988 675957 534989
rect 675891 534924 675892 534988
rect 675956 534924 675957 534988
rect 675891 534923 675957 534924
rect 676630 533493 676690 540938
rect 676627 533492 676693 533493
rect 676627 533428 676628 533492
rect 676692 533428 676693 533492
rect 676627 533427 676693 533428
rect 676814 532677 676874 576811
rect 677182 571981 677242 610131
rect 677363 610060 677429 610061
rect 677363 609996 677364 610060
rect 677428 609996 677429 610060
rect 677363 609995 677429 609996
rect 677179 571980 677245 571981
rect 677179 571916 677180 571980
rect 677244 571916 677245 571980
rect 677179 571915 677245 571916
rect 677366 571573 677426 609995
rect 676995 571572 677061 571573
rect 676995 571508 676996 571572
rect 677060 571508 677061 571572
rect 676995 571507 677061 571508
rect 677363 571572 677429 571573
rect 677363 571508 677364 571572
rect 677428 571508 677429 571572
rect 677363 571507 677429 571508
rect 676811 532676 676877 532677
rect 676811 532612 676812 532676
rect 676876 532612 676877 532676
rect 676811 532611 676877 532612
rect 676998 526965 677058 571507
rect 676995 526964 677061 526965
rect 676995 526900 676996 526964
rect 677060 526900 677061 526964
rect 676995 526899 677061 526900
rect 675155 485212 675221 485213
rect 675155 485148 675156 485212
rect 675220 485148 675221 485212
rect 675155 485147 675221 485148
rect 675155 402252 675221 402253
rect 675155 402188 675156 402252
rect 675220 402188 675221 402252
rect 675155 402187 675221 402188
rect 674971 400620 675037 400621
rect 674971 400556 674972 400620
rect 675036 400556 675037 400620
rect 674971 400555 675037 400556
rect 674787 399804 674853 399805
rect 674787 399740 674788 399804
rect 674852 399740 674853 399804
rect 674787 399739 674853 399740
rect 674790 355061 674850 399739
rect 674974 355877 675034 400555
rect 675158 357509 675218 402187
rect 675155 357508 675221 357509
rect 675155 357444 675156 357508
rect 675220 357444 675221 357508
rect 675155 357443 675221 357444
rect 674971 355876 675037 355877
rect 674971 355812 674972 355876
rect 675036 355812 675037 355876
rect 674971 355811 675037 355812
rect 674974 355798 675034 355811
rect 674787 355060 674853 355061
rect 674787 354996 674788 355060
rect 674852 354996 674853 355060
rect 674787 354995 674853 354996
rect 674790 354980 674850 354995
rect 60779 276044 60845 276045
rect 60779 275980 60780 276044
rect 60844 275980 60845 276044
rect 60779 275979 60845 275980
rect 41643 270468 41709 270469
rect 41643 270404 41644 270468
rect 41708 270404 41709 270468
rect 41643 270403 41709 270404
rect 675155 264620 675221 264621
rect 675155 264556 675156 264620
rect 675220 264556 675221 264620
rect 675155 264555 675221 264556
rect 41643 252652 41709 252653
rect 41643 252588 41644 252652
rect 41708 252588 41709 252652
rect 41643 252587 41709 252588
rect 41646 246010 41706 252587
rect 675158 251038 675218 264555
rect 675158 250978 677018 251038
rect 40346 245950 41706 246010
rect 40346 237622 40406 245950
rect 676958 244786 677018 250978
rect 675158 244726 677018 244786
rect 40346 237562 41706 237622
rect 41646 225997 41706 237562
rect 41643 225996 41709 225997
rect 41643 225932 41644 225996
rect 41708 225932 41709 225996
rect 41643 225931 41709 225932
rect 675158 219877 675218 244726
rect 675155 219876 675221 219877
rect 675155 219812 675156 219876
rect 675220 219812 675221 219876
rect 675155 219811 675221 219812
rect 41643 204916 41709 204917
rect 41643 204852 41644 204916
rect 41708 204852 41709 204916
rect 41643 204851 41709 204852
rect 41459 204508 41525 204509
rect 41459 204444 41460 204508
rect 41524 204444 41525 204508
rect 41459 204443 41525 204444
rect 41462 182749 41522 204443
rect 41646 183429 41706 204851
rect 41827 198796 41893 198797
rect 41827 198732 41828 198796
rect 41892 198732 41893 198796
rect 41827 198731 41893 198732
rect 41830 184245 41890 198731
rect 41827 184244 41893 184245
rect 41827 184180 41828 184244
rect 41892 184180 41893 184244
rect 41827 184179 41893 184180
rect 41643 183428 41709 183429
rect 41643 183364 41644 183428
rect 41708 183364 41709 183428
rect 41643 183363 41709 183364
rect 41459 182748 41525 182749
rect 41459 182684 41460 182748
rect 41524 182684 41525 182748
rect 41459 182683 41525 182684
rect 580947 113252 581013 113253
rect 580947 113188 580948 113252
rect 581012 113188 581013 113252
rect 580947 113187 581013 113188
rect 580950 73541 581010 113187
rect 662091 95572 662157 95573
rect 662091 95508 662092 95572
rect 662156 95508 662157 95572
rect 662091 95507 662157 95508
rect 662094 88773 662154 95507
rect 662091 88772 662157 88773
rect 662091 88708 662092 88772
rect 662156 88708 662157 88772
rect 662091 88707 662157 88708
rect 580947 73540 581013 73541
rect 580947 73476 580948 73540
rect 581012 73476 581013 73540
rect 580947 73475 581013 73476
rect 521699 48244 521765 48245
rect 521699 48180 521700 48244
rect 521764 48180 521765 48244
rect 521699 48179 521765 48180
rect 521702 42125 521762 48179
rect 521699 42124 521765 42125
rect 521699 42060 521700 42124
rect 521764 42060 521765 42124
rect 521699 42059 521765 42060
<< via4 >>
rect 221400 993820 234879 995620
rect 240878 993820 254357 995620
rect 274000 993820 287479 995620
rect 293478 993820 306957 995620
rect 375800 993820 389279 995620
rect 395278 993820 408757 995620
<< metal5 >>
rect 78610 1018624 90778 1030788
rect 130010 1018624 142178 1030788
rect 181410 1018624 193578 1030788
rect 231810 1018624 243978 1030788
rect 284410 1018624 296578 1030788
rect 334810 1018624 346978 1030788
rect 386210 1018624 398378 1030788
rect 475210 1018624 487378 1030788
rect 526610 1018624 538778 1030788
rect 577010 1018624 589178 1030788
rect 628410 1018624 640578 1030788
rect 221000 995620 235279 996020
rect 221000 993820 221400 995620
rect 234879 993820 235279 995620
rect 221000 993420 235279 993820
tri 221000 983518 230902 993420 ne
rect 230902 983518 235279 993420
rect 240478 995620 254757 996020
rect 240478 993820 240878 995620
rect 254357 993820 254757 995620
rect 273600 995620 287879 996020
rect 273600 993820 274000 995620
rect 287479 993820 287879 995620
rect 240478 992116 254800 993820
rect 240478 984242 246202 992116
tri 240478 983518 241202 984242 ne
rect 230902 982718 235902 983518
rect 241202 982718 246202 984242
tri 246202 983518 254800 992116 nw
rect 273600 992520 287879 993820
tri 273600 983518 282602 992520 ne
rect 282602 983795 287879 992520
rect 282602 982718 287602 983795
tri 287602 983518 287879 983795 nw
rect 293078 995620 307357 996020
rect 293078 993820 293478 995620
rect 306957 993820 307357 995620
rect 375400 995620 389679 996020
rect 375400 993820 375800 995620
rect 389279 993820 389679 995620
rect 293078 993016 307400 993820
rect 293078 983518 297902 993016
tri 297902 983518 307400 993016 nw
rect 375400 992420 389679 993820
tri 375400 983518 384302 992420 ne
rect 384302 983895 389679 992420
rect 292902 982718 297902 983518
rect 384302 982718 389302 983895
tri 389302 983518 389679 983895 nw
rect 394878 995620 409157 996020
rect 394878 993820 395278 995620
rect 408757 993820 409157 995620
rect 394878 993116 409200 993820
rect 394878 983518 399602 993116
tri 399602 983518 409200 993116 nw
rect 394602 982718 399602 983518
rect 6811 956610 18975 968778
rect 6167 914054 19619 924934
rect 697980 909666 711432 920546
rect 6811 871210 18975 883378
rect 698512 863640 711002 876160
rect 6811 829010 18975 841178
rect 698624 819822 710788 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710788 517390
rect 6811 484410 18975 496578
rect 697980 461866 711432 472746
rect 6167 443228 7258 453734
rect 8732 443228 19619 453734
rect 6167 442854 6970 443228
rect 9444 442854 19619 443228
rect 698624 417022 710788 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 621364 266578 630312 269344
rect 621454 262586 630402 265352
rect 621420 258566 630368 261332
rect 621518 254554 630436 257262
rect 621850 250624 630856 253288
rect 621912 246680 630918 249344
rect 621702 242714 630708 245378
rect 6598 227040 19088 239560
rect 621626 238638 630632 241302
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18975 123778
rect 698512 101240 711002 113760
rect 6167 70054 19619 80934
rect 80222 6811 92390 18975
rect 136713 7143 144149 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19619
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18975
rect 624222 6811 636390 18975
use caravel_clocking  clocking
timestamp 1637790566
transform 1 0 205746 0 1 5488
box -38 -48 20000 12000
use copyright_block_a  copyright_block_a_0
timestamp 1636248774
transform 1 0 149582 0 1 16298
box -262 -9464 35048 2764
use caravan_logo  caravan_logo_0
timestamp 1636751500
transform 1 0 310698 0 1 5742
box 2240 2560 37000 11520
use xres_buf  rstb_level
timestamp 1637551221
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use open_source  open_source_0 hexdigits
timestamp 1635801696
transform 1 0 260430 0 1 2174
box 752 5164 29030 16242
use user_id_textblock  user_id_textblock_0
timestamp 1608324878
transform 1 0 96272 0 1 6890
box -656 1508 33720 10344
use housekeeping  housekeeping
timestamp 1637790566
transform 1 0 606434 0 1 100002
box 0 0 60046 110190
use digital_pll  pll
timestamp 1637790566
transform 1 0 628146 0 1 80944
box 0 0 15000 15000
use user_id_programming  user_id_value
timestamp 1637790566
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use gpio_defaults_block  gpio_01_defaults\[0\]
timestamp 1637790566
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1637790566
transform -1 0 710203 0 1 121000
box 882 167 34000 13000
use caravan_motto  caravan_motto_0
timestamp 1637698689
transform 1 0 886 0 1 288
box 367960 10204 399802 14768
use simple_por  por
timestamp 1637617477
transform 1 0 650146 0 -1 55282
box -52 -62 11344 8684
use mgmt_core_wrapper  soc
timestamp 1637416673
transform 1 0 52034 0 1 53002
box 382 -400 524400 164400
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1637790566
transform 1 0 7631 0 1 202600
box 882 167 34000 13000
use gpio_defaults_block  gpio_01_defaults\[1\]
timestamp 1637790566
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1637790566
transform -1 0 710203 0 1 166200
box 882 167 34000 13000
use gpio_defaults_block  gpio_37_defaults
timestamp 1637790566
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1637790566
transform 1 0 7631 0 1 245800
box 882 167 34000 13000
use mgmt_protect  mgmt_buffers
timestamp 1637790566
transform 1 0 192180 0 1 232036
box -400 -400 220400 32400
use spare_logic_block  spare_logic_block_3
timestamp 1637790566
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic_block_1
timestamp 1637790566
transform 1 0 168632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic_block_2
timestamp 1637790566
transform 1 0 428632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic_block_0
timestamp 1637790566
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use gpio_defaults_block  gpio_234_defaults\[0\]
timestamp 1637790566
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1637790566
transform -1 0 710203 0 1 211200
box 882 167 34000 13000
use gpio_defaults_block  gpio_36_defaults
timestamp 1637790566
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_defaults_block  gpio_234_defaults\[1\]
timestamp 1637790566
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1637790566
transform -1 0 710203 0 1 256400
box 882 167 34000 13000
use gpio_defaults_block  gpio_35_defaults
timestamp 1637790566
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1637790566
transform 1 0 7631 0 1 289000
box 882 167 34000 13000
use gpio_defaults_block  gpio_234_defaults\[2\]
timestamp 1637790566
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1637790566
transform -1 0 710203 0 1 301400
box 882 167 34000 13000
use gpio_defaults_block  gpio_32_defaults
timestamp 1637790566
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_33_defaults
timestamp 1637790566
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_34_defaults
timestamp 1637790566
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1637790566
transform 1 0 7631 0 1 418600
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1637790566
transform 1 0 7631 0 1 375400
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1637790566
transform 1 0 7631 0 1 332200
box 882 167 34000 13000
use gpio_defaults_block  gpio_5_defaults
timestamp 1637790566
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_6_defaults
timestamp 1637790566
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_7_defaults
timestamp 1637790566
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1637790566
transform -1 0 710203 0 1 346400
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1637790566
transform -1 0 710203 0 1 391600
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1637790566
transform -1 0 710203 0 1 479800
box 882 167 34000 13000
use gpio_defaults_block  gpio_31_defaults
timestamp 1637790566
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_30_defaults
timestamp 1637790566
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1637790566
transform 1 0 7631 0 1 546200
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1637790566
transform 1 0 7631 0 1 589400
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1637790566
transform 1 0 7631 0 1 632600
box 882 167 34000 13000
use gpio_defaults_block  gpio_9_defaults
timestamp 1637790566
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_8_defaults
timestamp 1637790566
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_10_defaults
timestamp 1637790566
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1637790566
transform -1 0 710203 0 1 614000
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1637790566
transform -1 0 710203 0 1 568800
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1637790566
transform -1 0 710203 0 1 523800
box 882 167 34000 13000
use gpio_defaults_block  gpio_29_defaults
timestamp 1637790566
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_28_defaults
timestamp 1637790566
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_defaults_block  gpio_27_defaults
timestamp 1637790566
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1637790566
transform 1 0 7631 0 1 675800
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1637790566
transform 1 0 7631 0 1 719000
box 882 167 34000 13000
use gpio_defaults_block  gpio_12_defaults
timestamp 1637790566
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_11_defaults
timestamp 1637790566
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1637790566
transform -1 0 710203 0 1 704200
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1637790566
transform -1 0 710203 0 1 659000
box 882 167 34000 13000
use gpio_defaults_block  gpio_26_defaults
timestamp 1637790566
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_defaults_block  gpio_14_defaults
timestamp 1637790566
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1637790566
transform 1 0 7631 0 1 762200
box 882 167 34000 13000
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1637790566
transform 1 0 7631 0 1 805400
box 882 167 34000 13000
use gpio_defaults_block  gpio_13_defaults
timestamp 1637790566
transform -1 0 709467 0 1 897800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1637790566
transform -1 0 710203 0 1 884800
box 882 167 34000 13000
use caravan_power_routing  caravan_power_routing_0
timestamp 1637791793
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use user_analog_project_wrapper  mprj
timestamp 1632839657
transform 1 0 65308 0 1 278718
box -800 -800 584800 704800
use chip_io_alt  padframe
timestamp 1637691079
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< labels >>
flabel metal5 s 187640 6598 200160 19088 0 FreeSans 24000 0 0 0 clock
port 0 nsew signal input
flabel metal5 s 351040 6598 363560 19088 0 FreeSans 24000 0 0 0 flash_clk
port 1 nsew signal tristate
flabel metal5 s 296240 6598 308760 19088 0 FreeSans 24000 0 0 0 flash_csb
port 2 nsew signal tristate
flabel metal5 s 405840 6598 418360 19088 0 FreeSans 24000 0 0 0 flash_io0
port 3 nsew signal tristate
flabel metal5 s 460640 6598 473160 19088 0 FreeSans 24000 0 0 0 flash_io1
port 4 nsew signal tristate
flabel metal5 s 515440 6598 527960 19088 0 FreeSans 24000 0 0 0 gpio
port 5 nsew signal bidirectional
flabel metal5 s 698512 101240 711002 113760 0 FreeSans 24000 0 0 0 mprj_io[0]
port 6 nsew signal bidirectional
flabel metal5 s 698512 684440 711002 696960 0 FreeSans 24000 0 0 0 mprj_io[10]
port 7 nsew signal bidirectional
flabel metal5 s 698512 729440 711002 741960 0 FreeSans 24000 0 0 0 mprj_io[11]
port 8 nsew signal bidirectional
flabel metal5 s 698512 774440 711002 786960 0 FreeSans 24000 0 0 0 mprj_io[12]
port 9 nsew signal bidirectional
flabel metal5 s 698512 863640 711002 876160 0 FreeSans 24000 0 0 0 mprj_io[13]
port 10 nsew signal bidirectional
flabel metal5 s 698512 952840 711002 965360 0 FreeSans 24000 0 0 0 mprj_io[14]
port 11 nsew signal bidirectional
flabel metal5 s 628240 1018512 640760 1031002 0 FreeSans 24000 0 0 0 mprj_io[15]
port 12 nsew signal bidirectional
flabel metal5 s 526440 1018512 538960 1031002 0 FreeSans 24000 0 0 0 mprj_io[16]
port 13 nsew signal bidirectional
flabel metal5 s 475040 1018512 487560 1031002 0 FreeSans 24000 0 0 0 mprj_io[17]
port 14 nsew signal bidirectional
flabel metal5 s 386040 1018512 398560 1031002 0 FreeSans 24000 0 0 0 mprj_io[18]
port 15 nsew signal bidirectional
flabel metal5 s 284240 1018512 296760 1031002 0 FreeSans 24000 0 0 0 mprj_io[19]
port 16 nsew signal bidirectional
flabel metal5 s 698512 146440 711002 158960 0 FreeSans 24000 0 0 0 mprj_io[1]
port 17 nsew signal bidirectional
flabel metal5 s 232640 1018512 245160 1031002 0 FreeSans 24000 0 0 0 mprj_io[20]
port 18 nsew signal bidirectional
flabel metal5 s 181240 1018512 193760 1031002 0 FreeSans 24000 0 0 0 mprj_io[21]
port 19 nsew signal bidirectional
flabel metal5 s 129840 1018512 142360 1031002 0 FreeSans 24000 0 0 0 mprj_io[22]
port 20 nsew signal bidirectional
flabel metal5 s 78440 1018512 90960 1031002 0 FreeSans 24000 0 0 0 mprj_io[23]
port 21 nsew signal bidirectional
flabel metal5 s 6598 956440 19088 968960 0 FreeSans 24000 0 0 0 mprj_io[24]
port 22 nsew signal bidirectional
flabel metal5 s 6598 786640 19088 799160 0 FreeSans 24000 0 0 0 mprj_io[25]
port 23 nsew signal bidirectional
flabel metal5 s 6598 743440 19088 755960 0 FreeSans 24000 0 0 0 mprj_io[26]
port 24 nsew signal bidirectional
flabel metal5 s 6598 700240 19088 712760 0 FreeSans 24000 0 0 0 mprj_io[27]
port 25 nsew signal bidirectional
flabel metal5 s 6598 657040 19088 669560 0 FreeSans 24000 0 0 0 mprj_io[28]
port 26 nsew signal bidirectional
flabel metal5 s 6598 613840 19088 626360 0 FreeSans 24000 0 0 0 mprj_io[29]
port 27 nsew signal bidirectional
flabel metal5 s 698512 191440 711002 203960 0 FreeSans 24000 0 0 0 mprj_io[2]
port 28 nsew signal bidirectional
flabel metal5 s 6598 570640 19088 583160 0 FreeSans 24000 0 0 0 mprj_io[30]
port 29 nsew signal bidirectional
flabel metal5 s 6598 527440 19088 539960 0 FreeSans 24000 0 0 0 mprj_io[31]
port 30 nsew signal bidirectional
flabel metal5 s 6598 399840 19088 412360 0 FreeSans 24000 0 0 0 mprj_io[32]
port 31 nsew signal bidirectional
flabel metal5 s 6598 356640 19088 369160 0 FreeSans 24000 0 0 0 mprj_io[33]
port 32 nsew signal bidirectional
flabel metal5 s 6598 313440 19088 325960 0 FreeSans 24000 0 0 0 mprj_io[34]
port 33 nsew signal bidirectional
flabel metal5 s 6598 270240 19088 282760 0 FreeSans 24000 0 0 0 mprj_io[35]
port 34 nsew signal bidirectional
flabel metal5 s 6598 227040 19088 239560 0 FreeSans 24000 0 0 0 mprj_io[36]
port 35 nsew signal bidirectional
flabel metal5 s 6598 183840 19088 196360 0 FreeSans 24000 0 0 0 mprj_io[37]
port 36 nsew signal bidirectional
flabel metal5 s 698512 236640 711002 249160 0 FreeSans 24000 0 0 0 mprj_io[3]
port 37 nsew signal bidirectional
flabel metal5 s 698512 281640 711002 294160 0 FreeSans 24000 0 0 0 mprj_io[4]
port 38 nsew signal bidirectional
flabel metal5 s 698512 326640 711002 339160 0 FreeSans 24000 0 0 0 mprj_io[5]
port 39 nsew signal bidirectional
flabel metal5 s 698512 371840 711002 384360 0 FreeSans 24000 0 0 0 mprj_io[6]
port 40 nsew signal bidirectional
flabel metal5 s 698512 549040 711002 561560 0 FreeSans 24000 0 0 0 mprj_io[7]
port 41 nsew signal bidirectional
flabel metal5 s 698512 594240 711002 606760 0 FreeSans 24000 0 0 0 mprj_io[8]
port 42 nsew signal bidirectional
flabel metal5 s 698512 639240 711002 651760 0 FreeSans 24000 0 0 0 mprj_io[9]
port 43 nsew signal bidirectional
flabel metal5 s 136713 7143 144150 18309 0 FreeSans 24000 0 0 0 resetb
port 44 nsew signal input
flabel metal5 s 6167 70054 19619 80934 0 FreeSans 24000 0 0 0 vccd
port 45 nsew signal bidirectional
flabel metal5 s 697980 909666 711432 920546 0 FreeSans 24000 0 0 0 vccd1
port 46 nsew signal bidirectional
flabel metal5 s 6167 914054 19619 924934 0 FreeSans 24000 0 0 0 vccd2
port 47 nsew signal bidirectional
flabel metal5 s 624222 6811 636390 18975 0 FreeSans 24000 0 0 0 vdda
port 48 nsew signal bidirectional
flabel metal5 s 698624 819822 710788 831990 0 FreeSans 24000 0 0 0 vdda1
port 49 nsew signal bidirectional
flabel metal5 s 698624 505222 710788 517390 0 FreeSans 24000 0 0 0 vdda1_2
port 50 nsew signal bidirectional
flabel metal5 s 6811 484410 18975 496578 0 FreeSans 24000 0 0 0 vdda2
port 51 nsew signal bidirectional
flabel metal5 s 6811 111610 18975 123778 0 FreeSans 24000 0 0 0 vddio
port 52 nsew signal bidirectional
flabel metal5 s 6811 871210 18975 883378 0 FreeSans 24000 0 0 0 vddio_2
port 53 nsew signal bidirectional
flabel metal5 s 80222 6811 92390 18975 0 FreeSans 24000 0 0 0 vssa
port 54 nsew signal bidirectional
flabel metal5 s 577010 1018624 589178 1030788 0 FreeSans 24000 0 0 0 vssa1
port 55 nsew signal bidirectional
flabel metal5 s 698624 417022 710788 429190 0 FreeSans 24000 0 0 0 vssa1_2
port 56 nsew signal bidirectional
flabel metal5 s 6811 829010 18975 841178 0 FreeSans 24000 0 0 0 vssa2
port 57 nsew signal bidirectional
flabel metal5 s 243266 6167 254146 19619 0 FreeSans 24000 0 0 0 vssd
port 58 nsew signal bidirectional
flabel metal5 s 697980 461866 711432 472746 0 FreeSans 24000 0 0 0 vssd1
port 59 nsew signal bidirectional
flabel metal5 s 6167 442854 19619 453734 0 FreeSans 24000 0 0 0 vssd2
port 60 nsew signal bidirectional
flabel metal5 s 570422 6811 582590 18975 0 FreeSans 24000 0 0 0 vssio
port 61 nsew signal bidirectional
flabel metal5 s 334810 1018624 346978 1030788 0 FreeSans 24000 0 0 0 vssio_2
port 62 nsew signal bidirectional
flabel metal5 621960 246802 629984 249230 0 FreeSans 16000 0 0 0 vccd1_core
flabel metal5 621948 250708 629990 253036 0 FreeSans 16000 0 0 0 vssd1_core
flabel metal5 621550 262640 629508 265144 0 FreeSans 16000 0 0 0 vdda1_core
flabel metal5 621514 266692 629472 269196 0 FreeSans 16000 0 0 0 vssa1_core
flabel metal5 590480 230750 595228 233134 0 FreeSans 16000 0 0 0 vccd_core
flabel metal5 590522 234770 595540 236910 0 FreeSans 16000 0 0 0 vssd_core
flabel metal5 621512 258708 630212 261250 0 FreeSans 16000 0 0 0 vssa2_core
flabel metal5 621598 254668 630298 257210 0 FreeSans 16000 0 0 0 vdda2_core
flabel metal5 621936 242776 630636 245318 0 FreeSans 16000 0 0 0 vssd2_core
flabel metal5 621794 238736 630494 241278 0 FreeSans 16000 0 0 0 vccd2_core
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
