magic
tech sky130A
magscale 1 2
timestamp 1665142205
<< isosubstrate >>
rect 926 1576 2738 4794
<< viali >>
rect 8769 11781 8803 11815
rect 9781 11781 9815 11815
rect 1317 11713 1351 11747
rect 8217 11713 8251 11747
rect 1225 11645 1259 11679
rect 3433 11645 3467 11679
rect 3617 11645 3651 11679
rect 3801 11645 3835 11679
rect 3985 11645 4019 11679
rect 4261 11645 4295 11679
rect 6193 11645 6227 11679
rect 6377 11645 6411 11679
rect 6653 11645 6687 11679
rect 9321 11645 9355 11679
rect 9597 11645 9631 11679
rect 10057 11645 10091 11679
rect 6561 11577 6595 11611
rect 2513 11509 2547 11543
rect 5181 11509 5215 11543
rect 1685 11305 1719 11339
rect 6193 11237 6227 11271
rect 1501 11169 1535 11203
rect 3893 11169 3927 11203
rect 5365 11169 5399 11203
rect 7021 11169 7055 11203
rect 7297 11169 7331 11203
rect 7573 11169 7607 11203
rect 9413 11169 9447 11203
rect 3433 11101 3467 11135
rect 3525 11101 3559 11135
rect 5929 11101 5963 11135
rect 6745 11101 6779 11135
rect 7941 11101 7975 11135
rect 1317 11033 1351 11067
rect 7205 11033 7239 11067
rect 9973 11033 10007 11067
rect 3175 10965 3209 10999
rect 1317 10761 1351 10795
rect 8769 10761 8803 10795
rect 1409 10625 1443 10659
rect 3433 10625 3467 10659
rect 5825 10625 5859 10659
rect 8493 10625 8527 10659
rect 9321 10625 9355 10659
rect 3801 10557 3835 10591
rect 5917 10557 5951 10591
rect 6285 10557 6319 10591
rect 7757 10557 7791 10591
rect 8321 10557 8355 10591
rect 9597 10557 9631 10591
rect 9965 10557 9999 10591
rect 1685 10489 1719 10523
rect 4077 10489 4111 10523
rect 9781 10489 9815 10523
rect 3709 10421 3743 10455
rect 1685 10149 1719 10183
rect 5929 10149 5963 10183
rect 1409 10081 1443 10115
rect 3433 10081 3467 10115
rect 5365 10081 5399 10115
rect 7021 10081 7055 10115
rect 8861 10081 8895 10115
rect 3525 10013 3559 10047
rect 3893 10013 3927 10047
rect 6285 10013 6319 10047
rect 6929 10013 6963 10047
rect 7389 10013 7423 10047
rect 9597 10013 9631 10047
rect 9781 10013 9815 10047
rect 9965 10013 9999 10047
rect 1317 9877 1351 9911
rect 9421 9877 9455 9911
rect 6285 9605 6319 9639
rect 8769 9605 8803 9639
rect 3617 9537 3651 9571
rect 6017 9537 6051 9571
rect 8585 9537 8619 9571
rect 9321 9537 9355 9571
rect 9597 9537 9631 9571
rect 9965 9537 9999 9571
rect 3433 9469 3467 9503
rect 3985 9469 4019 9503
rect 5457 9469 5491 9503
rect 6462 9469 6496 9503
rect 6561 9469 6595 9503
rect 9873 9469 9907 9503
rect 1409 9401 1443 9435
rect 3157 9401 3191 9435
rect 6837 9401 6871 9435
rect 9505 9401 9539 9435
rect 1225 9333 1259 9367
rect 6193 9061 6227 9095
rect 7941 9061 7975 9095
rect 8309 9061 8343 9095
rect 1317 8993 1351 9027
rect 1869 8993 1903 9027
rect 2697 8993 2731 9027
rect 5641 8993 5675 9027
rect 1961 8925 1995 8959
rect 2973 8925 3007 8959
rect 4721 8925 4755 8959
rect 5365 8925 5399 8959
rect 5825 8925 5859 8959
rect 8217 8925 8251 8959
rect 9597 8857 9631 8891
rect 2605 8789 2639 8823
rect 4813 8789 4847 8823
rect 6009 8789 6043 8823
rect 2145 8585 2179 8619
rect 9873 8585 9907 8619
rect 8769 8517 8803 8551
rect 1409 8449 1443 8483
rect 5457 8449 5491 8483
rect 6285 8449 6319 8483
rect 9689 8449 9723 8483
rect 1593 8381 1627 8415
rect 3433 8381 3467 8415
rect 3617 8381 3651 8415
rect 4077 8381 4111 8415
rect 6193 8381 6227 8415
rect 8401 8381 8435 8415
rect 9321 8381 9355 8415
rect 9965 8381 9999 8415
rect 1225 8313 1259 8347
rect 3893 8313 3927 8347
rect 6561 8313 6595 8347
rect 8309 8313 8343 8347
rect 8493 8245 8527 8279
rect 1317 8041 1351 8075
rect 9973 8041 10007 8075
rect 1409 7905 1443 7939
rect 3341 7905 3375 7939
rect 5365 7905 5399 7939
rect 7021 7905 7055 7939
rect 7297 7905 7331 7939
rect 7573 7905 7607 7939
rect 9413 7905 9447 7939
rect 3525 7837 3559 7871
rect 3893 7837 3927 7871
rect 6193 7837 6227 7871
rect 7941 7837 7975 7871
rect 2513 7769 2547 7803
rect 6837 7769 6871 7803
rect 7389 7769 7423 7803
rect 5929 7701 5963 7735
rect 3801 7497 3835 7531
rect 8861 7497 8895 7531
rect 6185 7429 6219 7463
rect 1409 7361 1443 7395
rect 3157 7361 3191 7395
rect 3985 7361 4019 7395
rect 6009 7361 6043 7395
rect 8217 7361 8251 7395
rect 8585 7361 8619 7395
rect 3433 7293 3467 7327
rect 3617 7293 3651 7327
rect 6745 7293 6779 7327
rect 8769 7293 8803 7327
rect 9505 7293 9539 7327
rect 9689 7293 9723 7327
rect 9781 7293 9815 7327
rect 5733 7225 5767 7259
rect 9045 7225 9079 7259
rect 1317 7157 1351 7191
rect 8585 6885 8619 6919
rect 3893 6817 3927 6851
rect 5365 6817 5399 6851
rect 6653 6817 6687 6851
rect 8861 6817 8895 6851
rect 9229 6817 9263 6851
rect 9505 6817 9539 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 3433 6749 3467 6783
rect 3525 6749 3559 6783
rect 6285 6749 6319 6783
rect 6377 6749 6411 6783
rect 6837 6749 6871 6783
rect 9873 6749 9907 6783
rect 9137 6681 9171 6715
rect 1317 6613 1351 6647
rect 5929 6613 5963 6647
rect 1225 6409 1259 6443
rect 8493 6409 8527 6443
rect 9321 6409 9355 6443
rect 9505 6409 9539 6443
rect 10057 6409 10091 6443
rect 3709 6341 3743 6375
rect 4905 6341 4939 6375
rect 8769 6341 8803 6375
rect 3893 6273 3927 6307
rect 5273 6273 5307 6307
rect 5641 6273 5675 6307
rect 7849 6273 7883 6307
rect 9137 6273 9171 6307
rect 1409 6205 1443 6239
rect 1593 6205 1627 6239
rect 3433 6205 3467 6239
rect 3801 6199 3835 6233
rect 4629 6205 4663 6239
rect 5089 6205 5123 6239
rect 7113 6205 7147 6239
rect 8953 6205 8987 6239
rect 9873 6205 9907 6239
rect 9459 6137 9493 6171
rect 2145 6069 2179 6103
rect 4537 6069 4571 6103
rect 7677 6069 7711 6103
rect 3709 5865 3743 5899
rect 1777 5797 1811 5831
rect 3433 5797 3467 5831
rect 4261 5797 4295 5831
rect 6561 5797 6595 5831
rect 9689 5797 9723 5831
rect 1225 5729 1259 5763
rect 3893 5729 3927 5763
rect 8585 5729 8619 5763
rect 9229 5729 9263 5763
rect 9505 5729 9539 5763
rect 9965 5729 9999 5763
rect 1409 5661 1443 5695
rect 3985 5661 4019 5695
rect 6009 5661 6043 5695
rect 6193 5661 6227 5695
rect 6377 5661 6411 5695
rect 7941 5661 7975 5695
rect 8953 5661 8987 5695
rect 1593 5593 1627 5627
rect 8861 5525 8895 5559
rect 3709 5321 3743 5355
rect 5733 5321 5767 5355
rect 9421 5253 9455 5287
rect 3341 5185 3375 5219
rect 3525 5185 3559 5219
rect 5549 5185 5583 5219
rect 9781 5185 9815 5219
rect 3801 5117 3835 5151
rect 6285 5117 6319 5151
rect 6469 5117 6503 5151
rect 6653 5117 6687 5151
rect 7021 5117 7055 5151
rect 7389 5117 7423 5151
rect 8861 5117 8895 5151
rect 9597 5117 9631 5151
rect 9965 5117 9999 5151
rect 6837 5049 6871 5083
rect 9045 4981 9079 5015
rect 7389 4777 7423 4811
rect 9597 4777 9631 4811
rect 3433 4641 3467 4675
rect 3893 4641 3927 4675
rect 4445 4641 4479 4675
rect 5917 4641 5951 4675
rect 6745 4641 6779 4675
rect 7021 4641 7055 4675
rect 7481 4641 7515 4675
rect 7665 4641 7699 4675
rect 8309 4641 8343 4675
rect 4077 4573 4111 4607
rect 7941 4573 7975 4607
rect 8033 4573 8067 4607
rect 6929 4505 6963 4539
rect 3801 4437 3835 4471
rect 6477 4437 6511 4471
rect 5089 4097 5123 4131
rect 9413 4097 9447 4131
rect 3341 4029 3375 4063
rect 5181 4029 5215 4063
rect 5365 4029 5399 4063
rect 5549 4029 5583 4063
rect 5733 4029 5767 4063
rect 6285 4029 6319 4063
rect 8493 4029 8527 4063
rect 8033 3961 8067 3995
rect 5917 3893 5951 3927
rect 8953 3689 8987 3723
rect 9597 3689 9631 3723
rect 9137 3621 9171 3655
rect 3525 3553 3559 3587
rect 3985 3553 4019 3587
rect 6101 3553 6135 3587
rect 6377 3553 6411 3587
rect 8769 3553 8803 3587
rect 9781 3553 9815 3587
rect 3893 3485 3927 3519
rect 5089 3485 5123 3519
rect 8585 3485 8619 3519
rect 8125 3417 8159 3451
rect 9413 3417 9447 3451
rect 8401 3349 8435 3383
rect 9965 3349 9999 3383
rect 5273 3145 5307 3179
rect 6009 3145 6043 3179
rect 4629 3077 4663 3111
rect 5549 3077 5583 3111
rect 5733 3009 5767 3043
rect 6837 3009 6871 3043
rect 3341 2941 3375 2975
rect 5365 2941 5399 2975
rect 8033 2941 8067 2975
rect 8125 2941 8159 2975
rect 10057 2873 10091 2907
rect 3801 2601 3835 2635
rect 4169 2601 4203 2635
rect 5181 2601 5215 2635
rect 5365 2601 5399 2635
rect 6009 2601 6043 2635
rect 8953 2601 8987 2635
rect 9873 2601 9907 2635
rect 9505 2533 9539 2567
rect 3617 2465 3651 2499
rect 3985 2465 4019 2499
rect 4077 2465 4111 2499
rect 4445 2465 4479 2499
rect 4537 2465 4571 2499
rect 4813 2465 4847 2499
rect 4997 2465 5031 2499
rect 8125 2465 8159 2499
rect 8585 2465 8619 2499
rect 8769 2465 8803 2499
rect 9321 2465 9355 2499
rect 10057 2465 10091 2499
rect 4721 2397 4755 2431
rect 7481 2397 7515 2431
rect 9137 2397 9171 2431
rect 8401 2329 8435 2363
rect 3433 2261 3467 2295
rect 5641 2261 5675 2295
rect 5917 2261 5951 2295
rect 9689 2261 9723 2295
rect 3341 2057 3375 2091
rect 3525 2057 3559 2091
rect 3985 2057 4019 2091
rect 4169 2057 4203 2091
rect 4445 2057 4479 2091
rect 6009 2057 6043 2091
rect 3709 1989 3743 2023
rect 6837 1921 6871 1955
rect 4629 1853 4663 1887
rect 8033 1853 8067 1887
rect 8125 1853 8159 1887
rect 9873 1853 9907 1887
rect 5825 1717 5859 1751
rect 3341 1513 3375 1547
rect 3617 1513 3651 1547
rect 8125 1513 8159 1547
rect 9045 1513 9079 1547
rect 9689 1513 9723 1547
rect 6009 1377 6043 1411
rect 6193 1377 6227 1411
rect 8861 1377 8895 1411
rect 9505 1377 9539 1411
rect 9873 1377 9907 1411
rect 9965 1377 9999 1411
rect 5457 1309 5491 1343
rect 8493 1309 8527 1343
rect 8309 1173 8343 1207
rect 8677 1173 8711 1207
rect 9321 1173 9355 1207
rect 1317 969 1351 1003
rect 1869 969 1903 1003
rect 2973 969 3007 1003
rect 3157 969 3191 1003
rect 3341 969 3375 1003
rect 3709 969 3743 1003
rect 3893 969 3927 1003
rect 8769 969 8803 1003
rect 9045 969 9079 1003
rect 9689 969 9723 1003
rect 9873 969 9907 1003
rect 1593 901 1627 935
rect 2145 833 2179 867
rect 1225 765 1259 799
rect 1501 765 1535 799
rect 1777 765 1811 799
rect 2053 765 2087 799
rect 2421 697 2455 731
rect 2513 629 2547 663
rect 2789 629 2823 663
rect 7665 901 7699 935
rect 9137 833 9171 867
rect 9505 833 9539 867
rect 6009 765 6043 799
rect 8585 765 8619 799
rect 10057 765 10091 799
rect 6285 697 6319 731
rect 6561 697 6595 731
rect 5089 629 5123 663
rect 9321 629 9355 663
<< obsli1 >>
rect 0 12986 853 13014
rect 0 12969 9963 12986
rect 0 11815 33962 12969
rect 0 11781 8769 11815
rect 8803 11781 9781 11815
rect 9815 11781 33962 11815
rect 0 11747 33962 11781
rect 0 11713 1317 11747
rect 1351 11713 8217 11747
rect 8251 11713 33962 11747
rect 0 11679 33962 11713
rect 0 11645 1225 11679
rect 1259 11645 3433 11679
rect 3467 11645 3617 11679
rect 3651 11645 3801 11679
rect 3835 11645 3985 11679
rect 4019 11645 4261 11679
rect 4295 11645 6193 11679
rect 6227 11645 6377 11679
rect 6411 11645 6653 11679
rect 6687 11645 9321 11679
rect 9355 11645 9597 11679
rect 9631 11645 10057 11679
rect 10091 11645 33962 11679
rect 0 11611 33962 11645
rect 0 11577 6561 11611
rect 6595 11577 33962 11611
rect 0 11543 33962 11577
rect 0 11509 2513 11543
rect 2547 11509 5181 11543
rect 5215 11509 33962 11543
rect 0 11481 33962 11509
rect 0 6005 853 11481
rect 9800 11067 33962 11481
rect 9800 11033 9973 11067
rect 10007 11033 33962 11067
rect 9800 10591 33962 11033
rect 9800 10557 9965 10591
rect 9999 10557 33962 10591
rect 9800 10523 33962 10557
rect 9815 10489 33962 10523
rect 9800 10047 33962 10489
rect 9815 10013 9965 10047
rect 9999 10013 33962 10047
rect 9800 9571 33962 10013
rect 9800 9537 9965 9571
rect 9999 9537 33962 9571
rect 9800 9503 33962 9537
rect 9800 9469 9873 9503
rect 9907 9469 33962 9503
rect 9800 8619 33962 9469
rect 9800 8585 9873 8619
rect 9907 8585 33962 8619
rect 9800 8415 33962 8585
rect 9800 8381 9965 8415
rect 9999 8381 33962 8415
rect 9800 8075 33962 8381
rect 9800 8041 9973 8075
rect 10007 8041 33962 8075
rect 9800 7327 33962 8041
rect 9815 7293 33962 7327
rect 9800 6783 33962 7293
rect 9800 6749 9873 6783
rect 9907 6749 33962 6783
rect 9800 6443 33962 6749
rect 9800 6409 10057 6443
rect 10091 6409 33962 6443
rect 9800 6239 33962 6409
rect 9800 6205 9873 6239
rect 9907 6205 33962 6239
rect 0 5831 3359 6005
rect 0 5797 1777 5831
rect 1811 5797 3359 5831
rect 0 5763 3359 5797
rect 9800 5763 33962 6205
rect 0 5729 1225 5763
rect 1259 5729 3359 5763
rect 9800 5729 9965 5763
rect 9999 5729 33962 5763
rect 0 5695 3359 5729
rect 0 5661 1409 5695
rect 1443 5661 3359 5695
rect 0 5627 3359 5661
rect 0 5593 1593 5627
rect 1627 5593 3359 5627
rect 0 5219 3359 5593
rect 9800 5219 33962 5729
rect 0 5185 3341 5219
rect 9815 5185 33962 5219
rect 0 4063 3359 5185
rect 9800 5151 33962 5185
rect 9800 5117 9965 5151
rect 9999 5117 33962 5151
rect 0 4029 3341 4063
rect 0 2975 3359 4029
rect 9800 3587 33962 5117
rect 9815 3553 33962 3587
rect 9800 3383 33962 3553
rect 9800 3349 9965 3383
rect 9999 3349 33962 3383
rect 0 2941 3341 2975
rect 0 2091 3359 2941
rect 9800 2907 33962 3349
rect 9800 2873 10057 2907
rect 10091 2873 33962 2907
rect 9800 2635 33962 2873
rect 9800 2601 9873 2635
rect 9907 2601 33962 2635
rect 9800 2499 33962 2601
rect 9800 2465 10057 2499
rect 10091 2465 33962 2499
rect 0 2057 3341 2091
rect 0 1547 3359 2057
rect 9800 1887 33962 2465
rect 9800 1853 9873 1887
rect 9907 1853 33962 1887
rect 0 1513 3341 1547
rect 0 1003 3359 1513
rect 9800 1411 33962 1853
rect 9800 1377 9873 1411
rect 9907 1377 9965 1411
rect 9999 1377 33962 1411
rect 9800 1048 33962 1377
rect 3366 1003 33962 1048
rect 0 969 1317 1003
rect 1351 969 1869 1003
rect 1903 969 2973 1003
rect 3007 969 3157 1003
rect 3191 969 3341 1003
rect 3375 969 3709 1003
rect 3743 969 3893 1003
rect 3927 969 8769 1003
rect 8803 969 9045 1003
rect 9079 969 9689 1003
rect 9723 969 9873 1003
rect 9907 969 33962 1003
rect 0 935 3359 969
rect 0 901 1593 935
rect 1627 901 3359 935
rect 0 867 3359 901
rect 0 833 2145 867
rect 2179 833 3359 867
rect 0 799 3359 833
rect 0 765 1225 799
rect 1259 765 1501 799
rect 1535 765 1777 799
rect 1811 765 2053 799
rect 2087 765 3359 799
rect 0 731 3359 765
rect 0 697 2421 731
rect 2455 697 3359 731
rect 0 663 3359 697
rect 0 629 2513 663
rect 2547 629 2789 663
rect 2823 629 3359 663
rect 0 0 3359 629
rect 3366 935 33962 969
rect 3366 901 7665 935
rect 7699 901 33962 935
rect 3366 867 33962 901
rect 3366 833 9137 867
rect 9171 833 9505 867
rect 9539 833 33962 867
rect 3366 799 33962 833
rect 3366 765 6009 799
rect 6043 765 8585 799
rect 8619 765 10057 799
rect 10091 765 33962 799
rect 3366 731 33962 765
rect 3366 697 6285 731
rect 6319 697 6561 731
rect 6595 697 33962 731
rect 3366 663 33962 697
rect 3366 629 5089 663
rect 5123 629 9321 663
rect 9355 629 33962 663
rect 3366 0 33962 629
<< metal1 >>
rect 1210 12180 1216 12232
rect 1268 12220 1274 12232
rect 6086 12220 6092 12232
rect 1268 12192 6092 12220
rect 1268 12180 1274 12192
rect 6086 12180 6092 12192
rect 6144 12180 6150 12232
rect 2682 12044 2688 12096
rect 2740 12084 2746 12096
rect 3602 12084 3608 12096
rect 2740 12056 3608 12084
rect 2740 12044 2746 12056
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 920 11994 10396 12016
rect 920 11942 2566 11994
rect 2618 11942 2630 11994
rect 2682 11942 2694 11994
rect 2746 11942 2758 11994
rect 2810 11942 2822 11994
rect 2874 11942 7566 11994
rect 7618 11942 7630 11994
rect 7682 11942 7694 11994
rect 7746 11942 7758 11994
rect 7810 11942 7822 11994
rect 7874 11942 10396 11994
rect 920 11920 10396 11942
rect 6362 11880 6368 11892
rect 2746 11852 6368 11880
rect 2746 11824 2774 11852
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 6454 11840 6460 11892
rect 6512 11880 6518 11892
rect 7282 11880 7288 11892
rect 6512 11852 7288 11880
rect 6512 11840 6518 11852
rect 7282 11840 7288 11852
rect 7340 11880 7346 11892
rect 7340 11852 9628 11880
rect 7340 11840 7346 11852
rect 2682 11772 2688 11824
rect 2740 11784 2774 11824
rect 2740 11772 2746 11784
rect 3694 11772 3700 11824
rect 3752 11812 3758 11824
rect 8757 11815 8815 11821
rect 8757 11812 8769 11815
rect 3752 11784 8769 11812
rect 3752 11772 3758 11784
rect 8757 11781 8769 11784
rect 8803 11781 8815 11815
rect 8757 11775 8815 11781
rect 1305 11747 1363 11753
rect 1305 11713 1317 11747
rect 1351 11744 1363 11747
rect 7006 11744 7012 11756
rect 1351 11716 7012 11744
rect 1351 11713 1363 11716
rect 1305 11707 1363 11713
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 8202 11744 8208 11756
rect 8163 11716 8208 11744
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 1213 11679 1271 11685
rect 1213 11645 1225 11679
rect 1259 11645 1271 11679
rect 1213 11639 1271 11645
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11645 3479 11679
rect 3602 11676 3608 11688
rect 3563 11648 3608 11676
rect 3421 11639 3479 11645
rect 1228 11608 1256 11639
rect 3436 11608 3464 11639
rect 3602 11636 3608 11648
rect 3660 11636 3666 11688
rect 3786 11676 3792 11688
rect 3747 11648 3792 11676
rect 3786 11636 3792 11648
rect 3844 11636 3850 11688
rect 3973 11679 4031 11685
rect 3973 11645 3985 11679
rect 4019 11676 4031 11679
rect 4062 11676 4068 11688
rect 4019 11648 4068 11676
rect 4019 11645 4031 11648
rect 3973 11639 4031 11645
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4246 11636 4252 11688
rect 4304 11676 4310 11688
rect 4304 11648 4349 11676
rect 4304 11636 4310 11648
rect 6086 11636 6092 11688
rect 6144 11676 6150 11688
rect 6181 11679 6239 11685
rect 6181 11676 6193 11679
rect 6144 11648 6193 11676
rect 6144 11636 6150 11648
rect 6181 11645 6193 11648
rect 6227 11645 6239 11679
rect 6181 11639 6239 11645
rect 6365 11679 6423 11685
rect 6365 11645 6377 11679
rect 6411 11676 6423 11679
rect 6454 11676 6460 11688
rect 6411 11648 6460 11676
rect 6411 11645 6423 11648
rect 6365 11639 6423 11645
rect 6454 11636 6460 11648
rect 6512 11636 6518 11688
rect 6638 11676 6644 11688
rect 6599 11648 6644 11676
rect 6638 11636 6644 11648
rect 6696 11636 6702 11688
rect 6914 11636 6920 11688
rect 6972 11676 6978 11688
rect 9600 11685 9628 11852
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 17954 11880 17960 11892
rect 13872 11852 17960 11880
rect 13872 11840 13878 11852
rect 17954 11840 17960 11852
rect 18012 11840 18018 11892
rect 9769 11815 9827 11821
rect 9769 11781 9781 11815
rect 9815 11781 9827 11815
rect 9769 11775 9827 11781
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 6972 11648 9321 11676
rect 6972 11636 6978 11648
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 6549 11611 6607 11617
rect 1228 11580 2774 11608
rect 3436 11580 6500 11608
rect 2498 11540 2504 11552
rect 2459 11512 2504 11540
rect 2498 11500 2504 11512
rect 2556 11500 2562 11552
rect 2746 11540 2774 11580
rect 4154 11540 4160 11552
rect 2746 11512 4160 11540
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 5169 11543 5227 11549
rect 5169 11509 5181 11543
rect 5215 11540 5227 11543
rect 5442 11540 5448 11552
rect 5215 11512 5448 11540
rect 5215 11509 5227 11512
rect 5169 11503 5227 11509
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 6472 11540 6500 11580
rect 6549 11577 6561 11611
rect 6595 11608 6607 11611
rect 7466 11608 7472 11620
rect 6595 11580 7472 11608
rect 6595 11577 6607 11580
rect 6549 11571 6607 11577
rect 7466 11568 7472 11580
rect 7524 11568 7530 11620
rect 8478 11568 8484 11620
rect 8536 11608 8542 11620
rect 9784 11608 9812 11775
rect 10045 11679 10103 11685
rect 10045 11645 10057 11679
rect 10091 11645 10103 11679
rect 10045 11639 10103 11645
rect 8536 11580 9812 11608
rect 8536 11568 8542 11580
rect 6822 11540 6828 11552
rect 6472 11512 6828 11540
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 10060 11540 10088 11639
rect 8904 11512 10088 11540
rect 8904 11500 8910 11512
rect 920 11450 10396 11472
rect 920 11398 5066 11450
rect 5118 11398 5130 11450
rect 5182 11398 5194 11450
rect 5246 11398 5258 11450
rect 5310 11398 5322 11450
rect 5374 11398 10396 11450
rect 920 11376 10396 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 3878 11336 3884 11348
rect 1719 11308 3884 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 3970 11296 3976 11348
rect 4028 11336 4034 11348
rect 4028 11308 4200 11336
rect 4028 11296 4034 11308
rect 2682 11228 2688 11280
rect 2740 11228 2746 11280
rect 3142 11228 3148 11280
rect 3200 11268 3206 11280
rect 4172 11268 4200 11308
rect 4338 11296 4344 11348
rect 4396 11336 4402 11348
rect 4396 11308 7328 11336
rect 4396 11296 4402 11308
rect 6181 11271 6239 11277
rect 3200 11240 3464 11268
rect 4172 11240 4278 11268
rect 3200 11228 3206 11240
rect 1489 11203 1547 11209
rect 1489 11169 1501 11203
rect 1535 11169 1547 11203
rect 3436 11200 3464 11240
rect 6181 11237 6193 11271
rect 6227 11268 6239 11271
rect 6270 11268 6276 11280
rect 6227 11240 6276 11268
rect 6227 11237 6239 11240
rect 6181 11231 6239 11237
rect 6270 11228 6276 11240
rect 6328 11228 6334 11280
rect 3694 11200 3700 11212
rect 3436 11172 3700 11200
rect 1489 11163 1547 11169
rect 1504 11132 1532 11163
rect 3694 11160 3700 11172
rect 3752 11200 3758 11212
rect 3881 11203 3939 11209
rect 3881 11200 3893 11203
rect 3752 11172 3893 11200
rect 3752 11160 3758 11172
rect 3881 11169 3893 11172
rect 3927 11169 3939 11203
rect 3881 11163 3939 11169
rect 4798 11160 4804 11212
rect 4856 11200 4862 11212
rect 7300 11209 7328 11308
rect 8386 11228 8392 11280
rect 8444 11228 8450 11280
rect 5353 11203 5411 11209
rect 5353 11200 5365 11203
rect 4856 11172 5365 11200
rect 4856 11160 4862 11172
rect 5353 11169 5365 11172
rect 5399 11169 5411 11203
rect 7009 11203 7067 11209
rect 7009 11200 7021 11203
rect 5353 11163 5411 11169
rect 5460 11172 7021 11200
rect 2130 11132 2136 11144
rect 1504 11104 2136 11132
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 3418 11132 3424 11144
rect 3379 11104 3424 11132
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 3513 11135 3571 11141
rect 3513 11101 3525 11135
rect 3559 11132 3571 11135
rect 3602 11132 3608 11144
rect 3559 11104 3608 11132
rect 3559 11101 3571 11104
rect 3513 11095 3571 11101
rect 3602 11092 3608 11104
rect 3660 11092 3666 11144
rect 1305 11067 1363 11073
rect 1305 11033 1317 11067
rect 1351 11064 1363 11067
rect 5460 11064 5488 11172
rect 7009 11169 7021 11172
rect 7055 11169 7067 11203
rect 7009 11163 7067 11169
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11169 7343 11203
rect 7285 11163 7343 11169
rect 7561 11203 7619 11209
rect 7561 11169 7573 11203
rect 7607 11200 7619 11203
rect 7607 11172 8064 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 5917 11135 5975 11141
rect 5917 11101 5929 11135
rect 5963 11132 5975 11135
rect 6362 11132 6368 11144
rect 5963 11104 6368 11132
rect 5963 11101 5975 11104
rect 5917 11095 5975 11101
rect 6362 11092 6368 11104
rect 6420 11092 6426 11144
rect 6730 11132 6736 11144
rect 6691 11104 6736 11132
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 7926 11132 7932 11144
rect 7887 11104 7932 11132
rect 7926 11092 7932 11104
rect 7984 11092 7990 11144
rect 8036 11132 8064 11172
rect 8938 11160 8944 11212
rect 8996 11200 9002 11212
rect 9401 11203 9459 11209
rect 9401 11200 9413 11203
rect 8996 11172 9413 11200
rect 8996 11160 9002 11172
rect 9401 11169 9413 11172
rect 9447 11169 9459 11203
rect 9401 11163 9459 11169
rect 8570 11132 8576 11144
rect 8036 11104 8576 11132
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 1351 11036 2176 11064
rect 1351 11033 1363 11036
rect 1305 11027 1363 11033
rect 2148 10996 2176 11036
rect 4816 11036 5488 11064
rect 2682 10996 2688 11008
rect 2148 10968 2688 10996
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 3163 10999 3221 11005
rect 3163 10965 3175 10999
rect 3209 10996 3221 10999
rect 3326 10996 3332 11008
rect 3209 10968 3332 10996
rect 3209 10965 3221 10968
rect 3163 10959 3221 10965
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 3510 10956 3516 11008
rect 3568 10996 3574 11008
rect 3786 10996 3792 11008
rect 3568 10968 3792 10996
rect 3568 10956 3574 10968
rect 3786 10956 3792 10968
rect 3844 10996 3850 11008
rect 4816 10996 4844 11036
rect 5626 11024 5632 11076
rect 5684 11064 5690 11076
rect 7193 11067 7251 11073
rect 7193 11064 7205 11067
rect 5684 11036 7205 11064
rect 5684 11024 5690 11036
rect 7193 11033 7205 11036
rect 7239 11033 7251 11067
rect 7193 11027 7251 11033
rect 9858 11024 9864 11076
rect 9916 11064 9922 11076
rect 9961 11067 10019 11073
rect 9961 11064 9973 11067
rect 9916 11036 9973 11064
rect 9916 11024 9922 11036
rect 9961 11033 9973 11036
rect 10007 11033 10019 11067
rect 9961 11027 10019 11033
rect 3844 10968 4844 10996
rect 3844 10956 3850 10968
rect 920 10906 10396 10928
rect 920 10854 2566 10906
rect 2618 10854 2630 10906
rect 2682 10854 2694 10906
rect 2746 10854 2758 10906
rect 2810 10854 2822 10906
rect 2874 10854 7566 10906
rect 7618 10854 7630 10906
rect 7682 10854 7694 10906
rect 7746 10854 7758 10906
rect 7810 10854 7822 10906
rect 7874 10854 10396 10906
rect 920 10832 10396 10854
rect 1302 10792 1308 10804
rect 1263 10764 1308 10792
rect 1302 10752 1308 10764
rect 1360 10752 1366 10804
rect 6914 10792 6920 10804
rect 2746 10764 3280 10792
rect 1394 10656 1400 10668
rect 1307 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10656 1458 10668
rect 2746 10656 2774 10764
rect 1452 10628 2774 10656
rect 1452 10616 1458 10628
rect 3252 10600 3280 10764
rect 5368 10764 6920 10792
rect 3421 10659 3479 10665
rect 3421 10625 3433 10659
rect 3467 10656 3479 10659
rect 5368 10656 5396 10764
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7248 10764 7880 10792
rect 7248 10752 7254 10764
rect 7374 10684 7380 10736
rect 7432 10724 7438 10736
rect 7852 10724 7880 10764
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 8757 10795 8815 10801
rect 8757 10792 8769 10795
rect 7984 10764 8769 10792
rect 7984 10752 7990 10764
rect 8757 10761 8769 10764
rect 8803 10761 8815 10795
rect 8757 10755 8815 10761
rect 8294 10724 8300 10736
rect 7432 10696 7788 10724
rect 7852 10696 8300 10724
rect 7432 10684 7438 10696
rect 3467 10628 5396 10656
rect 5813 10659 5871 10665
rect 3467 10625 3479 10628
rect 3421 10619 3479 10625
rect 5813 10625 5825 10659
rect 5859 10656 5871 10659
rect 6730 10656 6736 10668
rect 5859 10628 6736 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 7760 10656 7788 10696
rect 8294 10684 8300 10696
rect 8352 10724 8358 10736
rect 8352 10696 9352 10724
rect 8352 10684 8358 10696
rect 9324 10665 9352 10696
rect 8481 10659 8539 10665
rect 8481 10656 8493 10659
rect 7760 10628 8493 10656
rect 8481 10625 8493 10628
rect 8527 10625 8539 10659
rect 8481 10619 8539 10625
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10625 9367 10659
rect 9309 10619 9367 10625
rect 2774 10548 2780 10600
rect 2832 10548 2838 10600
rect 3234 10548 3240 10600
rect 3292 10588 3298 10600
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 3292 10560 3801 10588
rect 3292 10548 3298 10560
rect 3789 10557 3801 10560
rect 3835 10557 3847 10591
rect 5902 10588 5908 10600
rect 5863 10560 5908 10588
rect 3789 10551 3847 10557
rect 5902 10548 5908 10560
rect 5960 10548 5966 10600
rect 6270 10588 6276 10600
rect 6231 10560 6276 10588
rect 6270 10548 6276 10560
rect 6328 10548 6334 10600
rect 7466 10548 7472 10600
rect 7524 10588 7530 10600
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7524 10560 7757 10588
rect 7524 10548 7530 10560
rect 7745 10557 7757 10560
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 8309 10591 8367 10597
rect 8309 10557 8321 10591
rect 8355 10588 8367 10591
rect 9122 10588 9128 10600
rect 8355 10560 9128 10588
rect 8355 10557 8367 10560
rect 8309 10551 8367 10557
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9582 10588 9588 10600
rect 9543 10560 9588 10588
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 1673 10523 1731 10529
rect 1673 10489 1685 10523
rect 1719 10489 1731 10523
rect 4065 10523 4123 10529
rect 4065 10520 4077 10523
rect 1673 10483 1731 10489
rect 3528 10492 4077 10520
rect 1688 10452 1716 10483
rect 2958 10452 2964 10464
rect 1688 10424 2964 10452
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 3050 10412 3056 10464
rect 3108 10452 3114 10464
rect 3528 10452 3556 10492
rect 4065 10489 4077 10492
rect 4111 10489 4123 10523
rect 5350 10520 5356 10532
rect 5290 10492 5356 10520
rect 4065 10483 4123 10489
rect 5350 10480 5356 10492
rect 5408 10480 5414 10532
rect 9769 10523 9827 10529
rect 9769 10520 9781 10523
rect 7406 10492 9781 10520
rect 9769 10489 9781 10492
rect 9815 10489 9827 10523
rect 9769 10483 9827 10489
rect 3108 10424 3556 10452
rect 3697 10455 3755 10461
rect 3108 10412 3114 10424
rect 3697 10421 3709 10455
rect 3743 10452 3755 10455
rect 4706 10452 4712 10464
rect 3743 10424 4712 10452
rect 3743 10421 3755 10424
rect 3697 10415 3755 10421
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 8662 10412 8668 10464
rect 8720 10452 8726 10464
rect 9968 10452 9996 10551
rect 8720 10424 9996 10452
rect 8720 10412 8726 10424
rect 920 10362 10396 10384
rect 920 10310 5066 10362
rect 5118 10310 5130 10362
rect 5182 10310 5194 10362
rect 5246 10310 5258 10362
rect 5310 10310 5322 10362
rect 5374 10310 10396 10362
rect 920 10288 10396 10310
rect 6270 10248 6276 10260
rect 1688 10220 6276 10248
rect 1688 10189 1716 10220
rect 6270 10208 6276 10220
rect 6328 10208 6334 10260
rect 8110 10248 8116 10260
rect 7024 10220 8116 10248
rect 1673 10183 1731 10189
rect 1673 10149 1685 10183
rect 1719 10149 1731 10183
rect 3510 10180 3516 10192
rect 2898 10166 3516 10180
rect 1673 10143 1731 10149
rect 2884 10152 3516 10166
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 2130 10004 2136 10056
rect 2188 10044 2194 10056
rect 2884 10044 2912 10152
rect 3510 10140 3516 10152
rect 3568 10140 3574 10192
rect 5626 10180 5632 10192
rect 5014 10152 5632 10180
rect 5626 10140 5632 10152
rect 5684 10140 5690 10192
rect 5917 10183 5975 10189
rect 5917 10149 5929 10183
rect 5963 10180 5975 10183
rect 7024 10180 7052 10220
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 5963 10152 7052 10180
rect 8484 10192 8536 10198
rect 5963 10149 5975 10152
rect 5917 10143 5975 10149
rect 8484 10134 8536 10140
rect 3421 10115 3479 10121
rect 3421 10081 3433 10115
rect 3467 10112 3479 10115
rect 3694 10112 3700 10124
rect 3467 10084 3700 10112
rect 3467 10081 3479 10084
rect 3421 10075 3479 10081
rect 3694 10072 3700 10084
rect 3752 10072 3758 10124
rect 5353 10115 5411 10121
rect 5353 10081 5365 10115
rect 5399 10112 5411 10115
rect 7006 10112 7012 10124
rect 5399 10084 5580 10112
rect 6967 10084 7012 10112
rect 5399 10081 5411 10084
rect 5353 10075 5411 10081
rect 5552 10056 5580 10084
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 8662 10072 8668 10124
rect 8720 10112 8726 10124
rect 8849 10115 8907 10121
rect 8849 10112 8861 10115
rect 8720 10084 8861 10112
rect 8720 10072 8726 10084
rect 8849 10081 8861 10084
rect 8895 10081 8907 10115
rect 8849 10075 8907 10081
rect 3510 10044 3516 10056
rect 2188 10016 2912 10044
rect 3471 10016 3516 10044
rect 2188 10004 2194 10016
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 3878 10044 3884 10056
rect 3620 10016 3884 10044
rect 2958 9936 2964 9988
rect 3016 9976 3022 9988
rect 3620 9976 3648 10016
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 5534 10004 5540 10056
rect 5592 10004 5598 10056
rect 6270 10044 6276 10056
rect 6231 10016 6276 10044
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10044 6975 10047
rect 7098 10044 7104 10056
rect 6963 10016 7104 10044
rect 6963 10013 6975 10016
rect 6917 10007 6975 10013
rect 7098 10004 7104 10016
rect 7156 10044 7162 10056
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 7156 10016 7389 10044
rect 7156 10004 7162 10016
rect 7377 10013 7389 10016
rect 7423 10013 7435 10047
rect 7377 10007 7435 10013
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 9585 10047 9643 10053
rect 9585 10044 9597 10047
rect 9456 10016 9597 10044
rect 9456 10004 9462 10016
rect 9585 10013 9597 10016
rect 9631 10013 9643 10047
rect 9766 10044 9772 10056
rect 9727 10016 9772 10044
rect 9585 10007 9643 10013
rect 9766 10004 9772 10016
rect 9824 10004 9830 10056
rect 9953 10047 10011 10053
rect 9953 10013 9965 10047
rect 9999 10044 10011 10047
rect 10226 10044 10232 10056
rect 9999 10016 10232 10044
rect 9999 10013 10011 10016
rect 9953 10007 10011 10013
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 3016 9948 3648 9976
rect 4816 9948 6040 9976
rect 3016 9936 3022 9948
rect 1305 9911 1363 9917
rect 1305 9877 1317 9911
rect 1351 9908 1363 9911
rect 3786 9908 3792 9920
rect 1351 9880 3792 9908
rect 1351 9877 1363 9880
rect 1305 9871 1363 9877
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 3878 9868 3884 9920
rect 3936 9908 3942 9920
rect 4816 9908 4844 9948
rect 3936 9880 4844 9908
rect 6012 9908 6040 9948
rect 7926 9908 7932 9920
rect 6012 9880 7932 9908
rect 3936 9868 3942 9880
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 8754 9868 8760 9920
rect 8812 9908 8818 9920
rect 9409 9911 9467 9917
rect 9409 9908 9421 9911
rect 8812 9880 9421 9908
rect 8812 9868 8818 9880
rect 9409 9877 9421 9880
rect 9455 9877 9467 9911
rect 9409 9871 9467 9877
rect 920 9818 10396 9840
rect 920 9766 2566 9818
rect 2618 9766 2630 9818
rect 2682 9766 2694 9818
rect 2746 9766 2758 9818
rect 2810 9766 2822 9818
rect 2874 9766 7566 9818
rect 7618 9766 7630 9818
rect 7682 9766 7694 9818
rect 7746 9766 7758 9818
rect 7810 9766 7822 9818
rect 7874 9766 10396 9818
rect 920 9744 10396 9766
rect 3694 9664 3700 9716
rect 3752 9704 3758 9716
rect 3752 9676 9352 9704
rect 3752 9664 3758 9676
rect 4982 9596 4988 9648
rect 5040 9636 5046 9648
rect 6273 9639 6331 9645
rect 6273 9636 6285 9639
rect 5040 9608 6285 9636
rect 5040 9596 5046 9608
rect 6273 9605 6285 9608
rect 6319 9605 6331 9639
rect 6273 9599 6331 9605
rect 7926 9596 7932 9648
rect 7984 9636 7990 9648
rect 8757 9639 8815 9645
rect 8757 9636 8769 9639
rect 7984 9608 8769 9636
rect 7984 9596 7990 9608
rect 8757 9605 8769 9608
rect 8803 9605 8815 9639
rect 8757 9599 8815 9605
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 3605 9571 3663 9577
rect 3605 9568 3617 9571
rect 2464 9540 3617 9568
rect 2464 9528 2470 9540
rect 3605 9537 3617 9540
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 5718 9528 5724 9580
rect 5776 9568 5782 9580
rect 6005 9571 6063 9577
rect 6005 9568 6017 9571
rect 5776 9540 6017 9568
rect 5776 9528 5782 9540
rect 6005 9537 6017 9540
rect 6051 9537 6063 9571
rect 6005 9531 6063 9537
rect 7282 9528 7288 9580
rect 7340 9568 7346 9580
rect 7466 9568 7472 9580
rect 7340 9540 7472 9568
rect 7340 9528 7346 9540
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 7558 9528 7564 9580
rect 7616 9568 7622 9580
rect 7616 9540 8064 9568
rect 7616 9528 7622 9540
rect 2038 9460 2044 9512
rect 2096 9460 2102 9512
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9469 3479 9503
rect 3973 9503 4031 9509
rect 3973 9500 3985 9503
rect 3421 9463 3479 9469
rect 3528 9472 3985 9500
rect 1302 9392 1308 9444
rect 1360 9432 1366 9444
rect 1397 9435 1455 9441
rect 1397 9432 1409 9435
rect 1360 9404 1409 9432
rect 1360 9392 1366 9404
rect 1397 9401 1409 9404
rect 1443 9401 1455 9435
rect 3142 9432 3148 9444
rect 3103 9404 3148 9432
rect 1397 9395 1455 9401
rect 3142 9392 3148 9404
rect 3200 9392 3206 9444
rect 3234 9392 3240 9444
rect 3292 9432 3298 9444
rect 3436 9432 3464 9463
rect 3292 9404 3464 9432
rect 3292 9392 3298 9404
rect 1213 9367 1271 9373
rect 1213 9333 1225 9367
rect 1259 9364 1271 9367
rect 2774 9364 2780 9376
rect 1259 9336 2780 9364
rect 1259 9333 1271 9336
rect 1213 9327 1271 9333
rect 2774 9324 2780 9336
rect 2832 9324 2838 9376
rect 2958 9324 2964 9376
rect 3016 9364 3022 9376
rect 3528 9364 3556 9472
rect 3973 9469 3985 9472
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 5166 9460 5172 9512
rect 5224 9500 5230 9512
rect 5445 9503 5503 9509
rect 5445 9500 5457 9503
rect 5224 9472 5457 9500
rect 5224 9460 5230 9472
rect 5445 9469 5457 9472
rect 5491 9469 5503 9503
rect 5445 9463 5503 9469
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 6450 9503 6508 9509
rect 6450 9500 6462 9503
rect 5868 9472 6462 9500
rect 5868 9460 5874 9472
rect 6450 9469 6462 9472
rect 6496 9469 6508 9503
rect 6450 9463 6508 9469
rect 6549 9503 6607 9509
rect 6549 9469 6561 9503
rect 6595 9469 6607 9503
rect 8036 9500 8064 9540
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 9324 9577 9352 9676
rect 8573 9571 8631 9577
rect 8573 9568 8585 9571
rect 8352 9540 8585 9568
rect 8352 9528 8358 9540
rect 8573 9537 8585 9540
rect 8619 9537 8631 9571
rect 8573 9531 8631 9537
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 9490 9528 9496 9580
rect 9548 9568 9554 9580
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 9548 9540 9597 9568
rect 9548 9528 9554 9540
rect 9585 9537 9597 9540
rect 9631 9537 9643 9571
rect 9950 9568 9956 9580
rect 9911 9540 9956 9568
rect 9585 9531 9643 9537
rect 9950 9528 9956 9540
rect 10008 9528 10014 9580
rect 8036 9472 9076 9500
rect 6549 9463 6607 9469
rect 4522 9392 4528 9444
rect 4580 9392 4586 9444
rect 6564 9432 6592 9463
rect 6730 9432 6736 9444
rect 6564 9404 6736 9432
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 6825 9435 6883 9441
rect 6825 9401 6837 9435
rect 6871 9432 6883 9435
rect 7098 9432 7104 9444
rect 6871 9404 7104 9432
rect 6871 9401 6883 9404
rect 6825 9395 6883 9401
rect 7098 9392 7104 9404
rect 7156 9392 7162 9444
rect 7282 9392 7288 9444
rect 7340 9392 7346 9444
rect 3016 9336 3556 9364
rect 3016 9324 3022 9336
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 5166 9364 5172 9376
rect 4120 9336 5172 9364
rect 4120 9324 4126 9336
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 5994 9364 6000 9376
rect 5684 9336 6000 9364
rect 5684 9324 5690 9336
rect 5994 9324 6000 9336
rect 6052 9364 6058 9376
rect 8846 9364 8852 9376
rect 6052 9336 8852 9364
rect 6052 9324 6058 9336
rect 8846 9324 8852 9336
rect 8904 9324 8910 9376
rect 9048 9364 9076 9472
rect 9214 9460 9220 9512
rect 9272 9500 9278 9512
rect 9861 9503 9919 9509
rect 9861 9500 9873 9503
rect 9272 9472 9873 9500
rect 9272 9460 9278 9472
rect 9861 9469 9873 9472
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 9122 9392 9128 9444
rect 9180 9432 9186 9444
rect 9493 9435 9551 9441
rect 9493 9432 9505 9435
rect 9180 9404 9505 9432
rect 9180 9392 9186 9404
rect 9493 9401 9505 9404
rect 9539 9401 9551 9435
rect 9493 9395 9551 9401
rect 10226 9364 10232 9376
rect 9048 9336 10232 9364
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 920 9274 10396 9296
rect 920 9222 5066 9274
rect 5118 9222 5130 9274
rect 5182 9222 5194 9274
rect 5246 9222 5258 9274
rect 5310 9222 5322 9274
rect 5374 9222 10396 9274
rect 920 9200 10396 9222
rect 3970 9120 3976 9172
rect 4028 9160 4034 9172
rect 4028 9132 8340 9160
rect 4028 9120 4034 9132
rect 3234 9092 3240 9104
rect 2700 9064 3240 9092
rect 1302 9024 1308 9036
rect 1263 8996 1308 9024
rect 1302 8984 1308 8996
rect 1360 8984 1366 9036
rect 2700 9033 2728 9064
rect 3234 9052 3240 9064
rect 3292 9052 3298 9104
rect 6181 9095 6239 9101
rect 6181 9061 6193 9095
rect 6227 9092 6239 9095
rect 6270 9092 6276 9104
rect 6227 9064 6276 9092
rect 6227 9061 6239 9064
rect 6181 9055 6239 9061
rect 6270 9052 6276 9064
rect 6328 9052 6334 9104
rect 7466 9052 7472 9104
rect 7524 9052 7530 9104
rect 7929 9095 7987 9101
rect 7929 9061 7941 9095
rect 7975 9092 7987 9095
rect 8018 9092 8024 9104
rect 7975 9064 8024 9092
rect 7975 9061 7987 9064
rect 7929 9055 7987 9061
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 8312 9101 8340 9132
rect 8297 9095 8355 9101
rect 8297 9061 8309 9095
rect 8343 9061 8355 9095
rect 8297 9055 8355 9061
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 2685 9027 2743 9033
rect 1903 8996 2636 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 1946 8956 1952 8968
rect 1907 8928 1952 8956
rect 1946 8916 1952 8928
rect 2004 8916 2010 8968
rect 2608 8956 2636 8996
rect 2685 8993 2697 9027
rect 2731 8993 2743 9027
rect 2685 8987 2743 8993
rect 4062 8984 4068 9036
rect 4120 8984 4126 9036
rect 4614 8984 4620 9036
rect 4672 9024 4678 9036
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 4672 8996 5641 9024
rect 4672 8984 4678 8996
rect 5629 8993 5641 8996
rect 5675 9024 5687 9027
rect 5675 8996 6776 9024
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 2958 8956 2964 8968
rect 2608 8928 2964 8956
rect 2958 8916 2964 8928
rect 3016 8916 3022 8968
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 4755 8928 5365 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 5353 8925 5365 8928
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 5813 8959 5871 8965
rect 5813 8925 5825 8959
rect 5859 8956 5871 8959
rect 6270 8956 6276 8968
rect 5859 8928 6276 8956
rect 5859 8925 5871 8928
rect 5813 8919 5871 8925
rect 6270 8916 6276 8928
rect 6328 8916 6334 8968
rect 6748 8956 6776 8996
rect 7282 8956 7288 8968
rect 6748 8928 7288 8956
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 4430 8848 4436 8900
rect 4488 8888 4494 8900
rect 6086 8888 6092 8900
rect 4488 8860 6092 8888
rect 4488 8848 4494 8860
rect 6086 8848 6092 8860
rect 6144 8848 6150 8900
rect 6178 8848 6184 8900
rect 6236 8888 6242 8900
rect 8220 8888 8248 8919
rect 8846 8888 8852 8900
rect 6236 8860 6960 8888
rect 8220 8860 8852 8888
rect 6236 8848 6242 8860
rect 2314 8780 2320 8832
rect 2372 8820 2378 8832
rect 2593 8823 2651 8829
rect 2593 8820 2605 8823
rect 2372 8792 2605 8820
rect 2372 8780 2378 8792
rect 2593 8789 2605 8792
rect 2639 8789 2651 8823
rect 2593 8783 2651 8789
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 4246 8820 4252 8832
rect 3200 8792 4252 8820
rect 3200 8780 3206 8792
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4798 8820 4804 8832
rect 4759 8792 4804 8820
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 5997 8823 6055 8829
rect 5997 8789 6009 8823
rect 6043 8820 6055 8823
rect 6730 8820 6736 8832
rect 6043 8792 6736 8820
rect 6043 8789 6055 8792
rect 5997 8783 6055 8789
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 6932 8820 6960 8860
rect 8846 8848 8852 8860
rect 8904 8888 8910 8900
rect 9585 8891 9643 8897
rect 9585 8888 9597 8891
rect 8904 8860 9597 8888
rect 8904 8848 8910 8860
rect 9585 8857 9597 8860
rect 9631 8857 9643 8891
rect 9585 8851 9643 8857
rect 7374 8820 7380 8832
rect 6932 8792 7380 8820
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 7466 8780 7472 8832
rect 7524 8820 7530 8832
rect 9766 8820 9772 8832
rect 7524 8792 9772 8820
rect 7524 8780 7530 8792
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 920 8730 10396 8752
rect 920 8678 2566 8730
rect 2618 8678 2630 8730
rect 2682 8678 2694 8730
rect 2746 8678 2758 8730
rect 2810 8678 2822 8730
rect 2874 8678 7566 8730
rect 7618 8678 7630 8730
rect 7682 8678 7694 8730
rect 7746 8678 7758 8730
rect 7810 8678 7822 8730
rect 7874 8678 10396 8730
rect 920 8656 10396 8678
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8616 2191 8619
rect 3970 8616 3976 8628
rect 2179 8588 3976 8616
rect 2179 8585 2191 8588
rect 2133 8579 2191 8585
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4522 8576 4528 8628
rect 4580 8616 4586 8628
rect 5718 8616 5724 8628
rect 4580 8588 5724 8616
rect 4580 8576 4586 8588
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 8662 8616 8668 8628
rect 5828 8588 8668 8616
rect 3786 8548 3792 8560
rect 3620 8520 3792 8548
rect 1397 8483 1455 8489
rect 1397 8449 1409 8483
rect 1443 8480 1455 8483
rect 3142 8480 3148 8492
rect 1443 8452 3148 8480
rect 1443 8449 1455 8452
rect 1397 8443 1455 8449
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3620 8480 3648 8520
rect 3786 8508 3792 8520
rect 3844 8508 3850 8560
rect 4430 8508 4436 8560
rect 4488 8548 4494 8560
rect 5828 8548 5856 8588
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 9861 8619 9919 8625
rect 9861 8616 9873 8619
rect 9732 8588 9873 8616
rect 9732 8576 9738 8588
rect 9861 8585 9873 8588
rect 9907 8585 9919 8619
rect 9861 8579 9919 8585
rect 4488 8520 5856 8548
rect 4488 8508 4494 8520
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 8757 8551 8815 8557
rect 8757 8548 8769 8551
rect 8352 8520 8769 8548
rect 8352 8508 8358 8520
rect 8757 8517 8769 8520
rect 8803 8517 8815 8551
rect 10226 8548 10232 8560
rect 8757 8511 8815 8517
rect 9692 8520 10232 8548
rect 5442 8480 5448 8492
rect 3436 8452 3648 8480
rect 5403 8452 5448 8480
rect 1581 8415 1639 8421
rect 1581 8381 1593 8415
rect 1627 8412 1639 8415
rect 2130 8412 2136 8424
rect 1627 8384 2136 8412
rect 1627 8381 1639 8384
rect 1581 8375 1639 8381
rect 2130 8372 2136 8384
rect 2188 8372 2194 8424
rect 3436 8421 3464 8452
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 5994 8440 6000 8492
rect 6052 8480 6058 8492
rect 6273 8483 6331 8489
rect 6273 8480 6285 8483
rect 6052 8452 6285 8480
rect 6052 8440 6058 8452
rect 6273 8449 6285 8452
rect 6319 8480 6331 8483
rect 6546 8480 6552 8492
rect 6319 8452 6552 8480
rect 6319 8449 6331 8452
rect 6273 8443 6331 8449
rect 6546 8440 6552 8452
rect 6604 8480 6610 8492
rect 8846 8480 8852 8492
rect 6604 8452 8852 8480
rect 6604 8440 6610 8452
rect 8846 8440 8852 8452
rect 8904 8440 8910 8492
rect 9692 8489 9720 8520
rect 10226 8508 10232 8520
rect 10284 8508 10290 8560
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8449 9735 8483
rect 9677 8443 9735 8449
rect 3421 8415 3479 8421
rect 3421 8381 3433 8415
rect 3467 8381 3479 8415
rect 3605 8415 3663 8421
rect 3605 8412 3617 8415
rect 3421 8375 3479 8381
rect 3528 8384 3617 8412
rect 1213 8347 1271 8353
rect 1213 8313 1225 8347
rect 1259 8344 1271 8347
rect 1302 8344 1308 8356
rect 1259 8316 1308 8344
rect 1259 8313 1271 8316
rect 1213 8307 1271 8313
rect 1302 8304 1308 8316
rect 1360 8304 1366 8356
rect 1486 8304 1492 8356
rect 1544 8344 1550 8356
rect 3528 8344 3556 8384
rect 3605 8381 3617 8384
rect 3651 8381 3663 8415
rect 3605 8375 3663 8381
rect 3786 8372 3792 8424
rect 3844 8412 3850 8424
rect 4065 8415 4123 8421
rect 4065 8412 4077 8415
rect 3844 8384 4077 8412
rect 3844 8372 3850 8384
rect 4065 8381 4077 8384
rect 4111 8381 4123 8415
rect 6178 8412 6184 8424
rect 6139 8384 6184 8412
rect 4065 8375 4123 8381
rect 6178 8372 6184 8384
rect 6236 8372 6242 8424
rect 7926 8372 7932 8424
rect 7984 8412 7990 8424
rect 8389 8415 8447 8421
rect 8389 8412 8401 8415
rect 7984 8384 8401 8412
rect 7984 8372 7990 8384
rect 8389 8381 8401 8384
rect 8435 8381 8447 8415
rect 8389 8375 8447 8381
rect 8478 8372 8484 8424
rect 8536 8412 8542 8424
rect 8754 8412 8760 8424
rect 8536 8384 8760 8412
rect 8536 8372 8542 8384
rect 8754 8372 8760 8384
rect 8812 8372 8818 8424
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 1544 8316 3556 8344
rect 3881 8347 3939 8353
rect 1544 8304 1550 8316
rect 3881 8313 3893 8347
rect 3927 8344 3939 8347
rect 4246 8344 4252 8356
rect 3927 8316 4252 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 4246 8304 4252 8316
rect 4304 8304 4310 8356
rect 6546 8344 6552 8356
rect 5184 8316 5396 8344
rect 6507 8316 6552 8344
rect 3326 8236 3332 8288
rect 3384 8276 3390 8288
rect 5184 8276 5212 8316
rect 3384 8248 5212 8276
rect 5368 8276 5396 8316
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 7558 8304 7564 8356
rect 7616 8304 7622 8356
rect 8297 8347 8355 8353
rect 8297 8313 8309 8347
rect 8343 8344 8355 8347
rect 9324 8344 9352 8375
rect 9766 8372 9772 8424
rect 9824 8412 9830 8424
rect 9953 8415 10011 8421
rect 9953 8412 9965 8415
rect 9824 8384 9965 8412
rect 9824 8372 9830 8384
rect 9953 8381 9965 8384
rect 9999 8381 10011 8415
rect 9953 8375 10011 8381
rect 8343 8316 9352 8344
rect 8343 8313 8355 8316
rect 8297 8307 8355 8313
rect 7834 8276 7840 8288
rect 5368 8248 7840 8276
rect 3384 8236 3390 8248
rect 7834 8236 7840 8248
rect 7892 8236 7898 8288
rect 8478 8276 8484 8288
rect 8439 8248 8484 8276
rect 8478 8236 8484 8248
rect 8536 8236 8542 8288
rect 920 8186 10396 8208
rect 920 8134 5066 8186
rect 5118 8134 5130 8186
rect 5182 8134 5194 8186
rect 5246 8134 5258 8186
rect 5310 8134 5322 8186
rect 5374 8134 10396 8186
rect 920 8112 10396 8134
rect 1305 8075 1363 8081
rect 1305 8041 1317 8075
rect 1351 8072 1363 8075
rect 1351 8044 7604 8072
rect 1351 8041 1363 8044
rect 1305 8035 1363 8041
rect 2222 7964 2228 8016
rect 2280 8004 2286 8016
rect 2280 7976 3556 8004
rect 2280 7964 2286 7976
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1762 7936 1768 7948
rect 1443 7908 1768 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1762 7896 1768 7908
rect 1820 7896 1826 7948
rect 3326 7936 3332 7948
rect 3287 7908 3332 7936
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 3528 7936 3556 7976
rect 4614 7964 4620 8016
rect 4672 7964 4678 8016
rect 6270 7964 6276 8016
rect 6328 8004 6334 8016
rect 7466 8004 7472 8016
rect 6328 7976 7472 8004
rect 6328 7964 6334 7976
rect 3528 7908 4016 7936
rect 1118 7828 1124 7880
rect 1176 7868 1182 7880
rect 3513 7871 3571 7877
rect 3513 7868 3525 7871
rect 1176 7840 3525 7868
rect 1176 7828 1182 7840
rect 3513 7837 3525 7840
rect 3559 7837 3571 7871
rect 3881 7871 3939 7877
rect 3881 7868 3893 7871
rect 3513 7831 3571 7837
rect 3620 7840 3893 7868
rect 2498 7800 2504 7812
rect 2459 7772 2504 7800
rect 2498 7760 2504 7772
rect 2556 7760 2562 7812
rect 3142 7692 3148 7744
rect 3200 7732 3206 7744
rect 3620 7732 3648 7840
rect 3881 7837 3893 7840
rect 3927 7837 3939 7871
rect 3988 7868 4016 7908
rect 4890 7896 4896 7948
rect 4948 7936 4954 7948
rect 7024 7945 7052 7976
rect 7466 7964 7472 7976
rect 7524 7964 7530 8016
rect 5353 7939 5411 7945
rect 5353 7936 5365 7939
rect 4948 7908 5365 7936
rect 4948 7896 4954 7908
rect 5353 7905 5365 7908
rect 5399 7905 5411 7939
rect 5353 7899 5411 7905
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7905 7067 7939
rect 7282 7936 7288 7948
rect 7243 7908 7288 7936
rect 7009 7899 7067 7905
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 7576 7945 7604 8044
rect 7834 8032 7840 8084
rect 7892 8072 7898 8084
rect 9961 8075 10019 8081
rect 9961 8072 9973 8075
rect 7892 8044 9973 8072
rect 7892 8032 7898 8044
rect 9961 8041 9973 8044
rect 10007 8041 10019 8075
rect 9961 8035 10019 8041
rect 9674 8004 9680 8016
rect 9062 7976 9680 8004
rect 9674 7964 9680 7976
rect 9732 7964 9738 8016
rect 7561 7939 7619 7945
rect 7561 7905 7573 7939
rect 7607 7905 7619 7939
rect 9398 7936 9404 7948
rect 9359 7908 9404 7936
rect 7561 7899 7619 7905
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 4246 7868 4252 7880
rect 3988 7840 4252 7868
rect 3881 7831 3939 7837
rect 4246 7828 4252 7840
rect 4304 7828 4310 7880
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 6181 7871 6239 7877
rect 6181 7868 6193 7871
rect 5684 7840 6193 7868
rect 5684 7828 5690 7840
rect 6181 7837 6193 7840
rect 6227 7837 6239 7871
rect 6181 7831 6239 7837
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7868 7987 7871
rect 8294 7868 8300 7880
rect 7975 7840 8300 7868
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 6546 7760 6552 7812
rect 6604 7800 6610 7812
rect 6825 7803 6883 7809
rect 6825 7800 6837 7803
rect 6604 7772 6837 7800
rect 6604 7760 6610 7772
rect 6825 7769 6837 7772
rect 6871 7800 6883 7803
rect 6871 7772 7236 7800
rect 6871 7769 6883 7772
rect 6825 7763 6883 7769
rect 4798 7732 4804 7744
rect 3200 7704 4804 7732
rect 3200 7692 3206 7704
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 5917 7735 5975 7741
rect 5917 7701 5929 7735
rect 5963 7732 5975 7735
rect 6270 7732 6276 7744
rect 5963 7704 6276 7732
rect 5963 7701 5975 7704
rect 5917 7695 5975 7701
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 7208 7732 7236 7772
rect 7282 7760 7288 7812
rect 7340 7800 7346 7812
rect 7377 7803 7435 7809
rect 7377 7800 7389 7803
rect 7340 7772 7389 7800
rect 7340 7760 7346 7772
rect 7377 7769 7389 7772
rect 7423 7769 7435 7803
rect 7377 7763 7435 7769
rect 8202 7732 8208 7744
rect 7208 7704 8208 7732
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 920 7642 10396 7664
rect 920 7590 2566 7642
rect 2618 7590 2630 7642
rect 2682 7590 2694 7642
rect 2746 7590 2758 7642
rect 2810 7590 2822 7642
rect 2874 7590 7566 7642
rect 7618 7590 7630 7642
rect 7682 7590 7694 7642
rect 7746 7590 7758 7642
rect 7810 7590 7822 7642
rect 7874 7590 10396 7642
rect 920 7568 10396 7590
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 3789 7531 3847 7537
rect 3789 7528 3801 7531
rect 2740 7500 3801 7528
rect 2740 7488 2746 7500
rect 3789 7497 3801 7500
rect 3835 7528 3847 7531
rect 4062 7528 4068 7540
rect 3835 7500 4068 7528
rect 3835 7497 3847 7500
rect 3789 7491 3847 7497
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4212 7500 8524 7528
rect 4212 7488 4218 7500
rect 3694 7420 3700 7472
rect 3752 7460 3758 7472
rect 4706 7460 4712 7472
rect 3752 7432 4712 7460
rect 3752 7420 3758 7432
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 6178 7469 6184 7472
rect 6173 7460 6184 7469
rect 6139 7432 6184 7460
rect 6173 7423 6184 7432
rect 6178 7420 6184 7423
rect 6236 7420 6242 7472
rect 8496 7460 8524 7500
rect 8570 7488 8576 7540
rect 8628 7528 8634 7540
rect 8849 7531 8907 7537
rect 8849 7528 8861 7531
rect 8628 7500 8861 7528
rect 8628 7488 8634 7500
rect 8849 7497 8861 7500
rect 8895 7497 8907 7531
rect 8849 7491 8907 7497
rect 8496 7432 8708 7460
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7392 1455 7395
rect 1946 7392 1952 7404
rect 1443 7364 1952 7392
rect 1443 7361 1455 7364
rect 1397 7355 1455 7361
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 3142 7392 3148 7404
rect 3103 7364 3148 7392
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7392 4031 7395
rect 5626 7392 5632 7404
rect 4019 7364 5632 7392
rect 4019 7361 4031 7364
rect 3973 7355 4031 7361
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5994 7392 6000 7404
rect 5955 7364 6000 7392
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 8202 7392 8208 7404
rect 8163 7364 8208 7392
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 8478 7352 8484 7404
rect 8536 7392 8542 7404
rect 8573 7395 8631 7401
rect 8573 7392 8585 7395
rect 8536 7364 8585 7392
rect 8536 7352 8542 7364
rect 8573 7361 8585 7364
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 3421 7327 3479 7333
rect 3421 7293 3433 7327
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7324 3663 7327
rect 4246 7324 4252 7336
rect 3651 7296 4252 7324
rect 3651 7293 3663 7296
rect 3605 7287 3663 7293
rect 2682 7216 2688 7268
rect 2740 7216 2746 7268
rect 3234 7216 3240 7268
rect 3292 7256 3298 7268
rect 3436 7256 3464 7287
rect 4246 7284 4252 7296
rect 4304 7284 4310 7336
rect 6730 7324 6736 7336
rect 6691 7296 6736 7324
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 8680 7324 8708 7432
rect 8757 7327 8815 7333
rect 8757 7324 8769 7327
rect 8680 7296 8769 7324
rect 8757 7293 8769 7296
rect 8803 7293 8815 7327
rect 8757 7287 8815 7293
rect 9122 7284 9128 7336
rect 9180 7324 9186 7336
rect 9493 7327 9551 7333
rect 9493 7324 9505 7327
rect 9180 7296 9505 7324
rect 9180 7284 9186 7296
rect 9493 7293 9505 7296
rect 9539 7293 9551 7327
rect 9674 7324 9680 7336
rect 9635 7296 9680 7324
rect 9493 7287 9551 7293
rect 9674 7284 9680 7296
rect 9732 7284 9738 7336
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7324 9827 7327
rect 9815 7296 16574 7324
rect 9815 7293 9827 7296
rect 9769 7287 9827 7293
rect 5442 7256 5448 7268
rect 3292 7228 3464 7256
rect 5290 7228 5448 7256
rect 3292 7216 3298 7228
rect 5442 7216 5448 7228
rect 5500 7216 5506 7268
rect 5626 7216 5632 7268
rect 5684 7256 5690 7268
rect 5721 7259 5779 7265
rect 5721 7256 5733 7259
rect 5684 7228 5733 7256
rect 5684 7216 5690 7228
rect 5721 7225 5733 7228
rect 5767 7225 5779 7259
rect 5721 7219 5779 7225
rect 7282 7216 7288 7268
rect 7340 7216 7346 7268
rect 8570 7216 8576 7268
rect 8628 7256 8634 7268
rect 9033 7259 9091 7265
rect 9033 7256 9045 7259
rect 8628 7228 9045 7256
rect 8628 7216 8634 7228
rect 9033 7225 9045 7228
rect 9079 7225 9091 7259
rect 9033 7219 9091 7225
rect 1305 7191 1363 7197
rect 1305 7157 1317 7191
rect 1351 7188 1363 7191
rect 9784 7188 9812 7287
rect 1351 7160 9812 7188
rect 16546 7188 16574 7296
rect 17954 7188 17960 7200
rect 16546 7160 17960 7188
rect 1351 7157 1363 7160
rect 1305 7151 1363 7157
rect 17954 7148 17960 7160
rect 18012 7148 18018 7200
rect 920 7098 10396 7120
rect 920 7046 5066 7098
rect 5118 7046 5130 7098
rect 5182 7046 5194 7098
rect 5246 7046 5258 7098
rect 5310 7046 5322 7098
rect 5374 7046 10396 7098
rect 920 7024 10396 7046
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 2038 6984 2044 6996
rect 1728 6956 2044 6984
rect 1728 6944 1734 6956
rect 2038 6944 2044 6956
rect 2096 6984 2102 6996
rect 3786 6984 3792 6996
rect 2096 6956 3792 6984
rect 2096 6944 2102 6956
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 4338 6944 4344 6996
rect 4396 6984 4402 6996
rect 5442 6984 5448 6996
rect 4396 6956 5448 6984
rect 4396 6944 4402 6956
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 8202 6984 8208 6996
rect 7616 6956 8208 6984
rect 7616 6944 7622 6956
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 4890 6876 4896 6928
rect 4948 6876 4954 6928
rect 8220 6916 8248 6944
rect 8142 6888 8248 6916
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 8573 6919 8631 6925
rect 8573 6916 8585 6919
rect 8352 6888 8585 6916
rect 8352 6876 8358 6888
rect 8573 6885 8585 6888
rect 8619 6885 8631 6919
rect 8573 6879 8631 6885
rect 3142 6848 3148 6860
rect 2806 6820 3148 6848
rect 3142 6808 3148 6820
rect 3200 6808 3206 6860
rect 3881 6851 3939 6857
rect 3881 6848 3893 6851
rect 3344 6820 3893 6848
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 2314 6780 2320 6792
rect 1719 6752 2320 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 2314 6740 2320 6752
rect 2372 6780 2378 6792
rect 2372 6752 2728 6780
rect 2372 6740 2378 6752
rect 2700 6712 2728 6752
rect 3344 6712 3372 6820
rect 3881 6817 3893 6820
rect 3927 6817 3939 6851
rect 3881 6811 3939 6817
rect 4798 6808 4804 6860
rect 4856 6848 4862 6860
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 4856 6820 5365 6848
rect 4856 6808 4862 6820
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 6641 6851 6699 6857
rect 6641 6848 6653 6851
rect 5353 6811 5411 6817
rect 5552 6820 6653 6848
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 2700 6684 3372 6712
rect 1302 6644 1308 6656
rect 1263 6616 1308 6644
rect 1302 6604 1308 6616
rect 1360 6604 1366 6656
rect 3436 6644 3464 6743
rect 3510 6740 3516 6792
rect 3568 6780 3574 6792
rect 3568 6752 3613 6780
rect 3568 6740 3574 6752
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 4522 6780 4528 6792
rect 3844 6752 4528 6780
rect 3844 6740 3850 6752
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 3878 6644 3884 6656
rect 3436 6616 3884 6644
rect 3878 6604 3884 6616
rect 3936 6604 3942 6656
rect 4522 6604 4528 6656
rect 4580 6644 4586 6656
rect 5552 6644 5580 6820
rect 6641 6817 6653 6820
rect 6687 6817 6699 6851
rect 6641 6811 6699 6817
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 9217 6851 9275 6857
rect 8904 6820 8949 6848
rect 8904 6808 8910 6820
rect 9217 6817 9229 6851
rect 9263 6848 9275 6851
rect 9306 6848 9312 6860
rect 9263 6820 9312 6848
rect 9263 6817 9275 6820
rect 9217 6811 9275 6817
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 9490 6848 9496 6860
rect 9451 6820 9496 6848
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 6273 6783 6331 6789
rect 6273 6780 6285 6783
rect 5776 6752 6285 6780
rect 5776 6740 5782 6752
rect 6273 6749 6285 6752
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6780 6423 6783
rect 6546 6780 6552 6792
rect 6411 6752 6552 6780
rect 6411 6749 6423 6752
rect 6365 6743 6423 6749
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6780 6883 6783
rect 7374 6780 7380 6792
rect 6871 6752 7380 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 7374 6740 7380 6752
rect 7432 6740 7438 6792
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 4580 6616 5580 6644
rect 5917 6647 5975 6653
rect 4580 6604 4586 6616
rect 5917 6613 5929 6647
rect 5963 6644 5975 6647
rect 6178 6644 6184 6656
rect 5963 6616 6184 6644
rect 5963 6613 5975 6616
rect 5917 6607 5975 6613
rect 6178 6604 6184 6616
rect 6236 6604 6242 6656
rect 6564 6644 6592 6740
rect 9122 6712 9128 6724
rect 9083 6684 9128 6712
rect 9122 6672 9128 6684
rect 9180 6672 9186 6724
rect 9490 6672 9496 6724
rect 9548 6712 9554 6724
rect 9876 6712 9904 6743
rect 9548 6684 9904 6712
rect 9548 6672 9554 6684
rect 6564 6616 10456 6644
rect 920 6554 10396 6576
rect 920 6502 2566 6554
rect 2618 6502 2630 6554
rect 2682 6502 2694 6554
rect 2746 6502 2758 6554
rect 2810 6502 2822 6554
rect 2874 6502 7566 6554
rect 7618 6502 7630 6554
rect 7682 6502 7694 6554
rect 7746 6502 7758 6554
rect 7810 6502 7822 6554
rect 7874 6502 10396 6554
rect 920 6480 10396 6502
rect 1210 6440 1216 6452
rect 1171 6412 1216 6440
rect 1210 6400 1216 6412
rect 1268 6400 1274 6452
rect 2866 6400 2872 6452
rect 2924 6440 2930 6452
rect 3142 6440 3148 6452
rect 2924 6412 3148 6440
rect 2924 6400 2930 6412
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 6914 6440 6920 6452
rect 3804 6412 6920 6440
rect 3510 6332 3516 6384
rect 3568 6372 3574 6384
rect 3697 6375 3755 6381
rect 3697 6372 3709 6375
rect 3568 6344 3709 6372
rect 3568 6332 3574 6344
rect 3697 6341 3709 6344
rect 3743 6341 3755 6375
rect 3697 6335 3755 6341
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 2774 6304 2780 6316
rect 1360 6276 2780 6304
rect 1360 6264 1366 6276
rect 2774 6264 2780 6276
rect 2832 6264 2838 6316
rect 3804 6304 3832 6412
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 8018 6440 8024 6452
rect 7524 6412 8024 6440
rect 7524 6400 7530 6412
rect 8018 6400 8024 6412
rect 8076 6440 8082 6452
rect 8481 6443 8539 6449
rect 8481 6440 8493 6443
rect 8076 6412 8493 6440
rect 8076 6400 8082 6412
rect 8481 6409 8493 6412
rect 8527 6409 8539 6443
rect 8481 6403 8539 6409
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 9309 6443 9367 6449
rect 9309 6440 9321 6443
rect 9272 6412 9321 6440
rect 9272 6400 9278 6412
rect 9309 6409 9321 6412
rect 9355 6409 9367 6443
rect 9309 6403 9367 6409
rect 9493 6443 9551 6449
rect 9493 6409 9505 6443
rect 9539 6409 9551 6443
rect 9493 6403 9551 6409
rect 10045 6443 10103 6449
rect 10045 6409 10057 6443
rect 10091 6440 10103 6443
rect 10428 6440 10456 6616
rect 10091 6412 10456 6440
rect 10091 6409 10103 6412
rect 10045 6403 10103 6409
rect 4890 6372 4896 6384
rect 4851 6344 4896 6372
rect 4890 6332 4896 6344
rect 4948 6332 4954 6384
rect 8110 6332 8116 6384
rect 8168 6372 8174 6384
rect 8757 6375 8815 6381
rect 8757 6372 8769 6375
rect 8168 6344 8769 6372
rect 8168 6332 8174 6344
rect 8757 6341 8769 6344
rect 8803 6341 8815 6375
rect 9508 6372 9536 6403
rect 8757 6335 8815 6341
rect 9048 6344 9536 6372
rect 3436 6276 3832 6304
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6205 1455 6239
rect 1397 6199 1455 6205
rect 1412 6168 1440 6199
rect 1486 6196 1492 6248
rect 1544 6236 1550 6248
rect 1581 6239 1639 6245
rect 1581 6236 1593 6239
rect 1544 6208 1593 6236
rect 1544 6196 1550 6208
rect 1581 6205 1593 6208
rect 1627 6236 1639 6239
rect 3050 6236 3056 6248
rect 1627 6208 3056 6236
rect 1627 6205 1639 6208
rect 1581 6199 1639 6205
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 3436 6245 3464 6276
rect 3878 6264 3884 6316
rect 3936 6304 3942 6316
rect 3936 6276 3981 6304
rect 3936 6264 3942 6276
rect 4246 6264 4252 6316
rect 4304 6304 4310 6316
rect 5261 6307 5319 6313
rect 5261 6304 5273 6307
rect 4304 6276 5273 6304
rect 4304 6264 4310 6276
rect 5261 6273 5273 6276
rect 5307 6273 5319 6307
rect 5626 6304 5632 6316
rect 5587 6276 5632 6304
rect 5261 6267 5319 6273
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7432 6276 7849 6304
rect 7432 6264 7438 6276
rect 7837 6273 7849 6276
rect 7883 6273 7895 6307
rect 7837 6267 7895 6273
rect 8662 6264 8668 6316
rect 8720 6304 8726 6316
rect 9048 6304 9076 6344
rect 8720 6276 9076 6304
rect 9125 6307 9183 6313
rect 8720 6264 8726 6276
rect 9125 6273 9137 6307
rect 9171 6304 9183 6307
rect 9674 6304 9680 6316
rect 9171 6276 9680 6304
rect 9171 6273 9183 6276
rect 9125 6267 9183 6273
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6236 3479 6239
rect 3510 6236 3516 6248
rect 3467 6208 3516 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 3789 6233 3847 6239
rect 3789 6230 3801 6233
rect 3712 6202 3801 6230
rect 1670 6168 1676 6180
rect 1412 6140 1676 6168
rect 1670 6128 1676 6140
rect 1728 6128 1734 6180
rect 1762 6128 1768 6180
rect 1820 6168 1826 6180
rect 3712 6168 3740 6202
rect 3789 6199 3801 6202
rect 3835 6230 3847 6233
rect 3835 6202 3924 6230
rect 3835 6199 3847 6202
rect 3789 6193 3847 6199
rect 1820 6140 3740 6168
rect 3896 6168 3924 6202
rect 4154 6196 4160 6248
rect 4212 6236 4218 6248
rect 4617 6239 4675 6245
rect 4617 6236 4629 6239
rect 4212 6208 4629 6236
rect 4212 6196 4218 6208
rect 4617 6205 4629 6208
rect 4663 6236 4675 6239
rect 4706 6236 4712 6248
rect 4663 6208 4712 6236
rect 4663 6205 4675 6208
rect 4617 6199 4675 6205
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 4982 6196 4988 6248
rect 5040 6236 5046 6248
rect 5077 6239 5135 6245
rect 5077 6236 5089 6239
rect 5040 6208 5089 6236
rect 5040 6196 5046 6208
rect 5077 6205 5089 6208
rect 5123 6205 5135 6239
rect 5077 6199 5135 6205
rect 6546 6196 6552 6248
rect 6604 6236 6610 6248
rect 7101 6239 7159 6245
rect 7101 6236 7113 6239
rect 6604 6208 7113 6236
rect 6604 6196 6610 6208
rect 7101 6205 7113 6208
rect 7147 6205 7159 6239
rect 8938 6236 8944 6248
rect 8899 6208 8944 6236
rect 7101 6199 7159 6205
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 9858 6236 9864 6248
rect 9819 6208 9864 6236
rect 9858 6196 9864 6208
rect 9916 6196 9922 6248
rect 4430 6168 4436 6180
rect 3896 6140 4436 6168
rect 1820 6128 1826 6140
rect 4430 6128 4436 6140
rect 4488 6128 4494 6180
rect 6914 6168 6920 6180
rect 6762 6140 6920 6168
rect 6914 6128 6920 6140
rect 6972 6128 6978 6180
rect 8956 6168 8984 6196
rect 9447 6171 9505 6177
rect 9447 6168 9459 6171
rect 8956 6140 9459 6168
rect 9447 6137 9459 6140
rect 9493 6137 9505 6171
rect 9447 6131 9505 6137
rect 2133 6103 2191 6109
rect 2133 6069 2145 6103
rect 2179 6100 2191 6103
rect 3786 6100 3792 6112
rect 2179 6072 3792 6100
rect 2179 6069 2191 6072
rect 2133 6063 2191 6069
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 4154 6100 4160 6112
rect 4028 6072 4160 6100
rect 4028 6060 4034 6072
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 4522 6100 4528 6112
rect 4483 6072 4528 6100
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 7665 6103 7723 6109
rect 7665 6069 7677 6103
rect 7711 6100 7723 6103
rect 8018 6100 8024 6112
rect 7711 6072 8024 6100
rect 7711 6069 7723 6072
rect 7665 6063 7723 6069
rect 8018 6060 8024 6072
rect 8076 6060 8082 6112
rect 8754 6060 8760 6112
rect 8812 6100 8818 6112
rect 9766 6100 9772 6112
rect 8812 6072 9772 6100
rect 8812 6060 8818 6072
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 920 6010 10396 6032
rect 920 5958 5066 6010
rect 5118 5958 5130 6010
rect 5182 5958 5194 6010
rect 5246 5958 5258 6010
rect 5310 5958 5322 6010
rect 5374 5958 10396 6010
rect 920 5936 10396 5958
rect 3142 5856 3148 5908
rect 3200 5896 3206 5908
rect 3697 5899 3755 5905
rect 3697 5896 3709 5899
rect 3200 5868 3709 5896
rect 3200 5856 3206 5868
rect 3697 5865 3709 5868
rect 3743 5865 3755 5899
rect 3697 5859 3755 5865
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4890 5896 4896 5908
rect 4028 5868 4896 5896
rect 4028 5856 4034 5868
rect 4890 5856 4896 5868
rect 4948 5896 4954 5908
rect 11054 5896 11060 5908
rect 4948 5868 11060 5896
rect 4948 5856 4954 5868
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 1394 5788 1400 5840
rect 1452 5828 1458 5840
rect 1765 5831 1823 5837
rect 1765 5828 1777 5831
rect 1452 5800 1777 5828
rect 1452 5788 1458 5800
rect 1765 5797 1777 5800
rect 1811 5797 1823 5831
rect 1765 5791 1823 5797
rect 3421 5831 3479 5837
rect 3421 5797 3433 5831
rect 3467 5828 3479 5831
rect 4154 5828 4160 5840
rect 3467 5800 4160 5828
rect 3467 5797 3479 5800
rect 3421 5791 3479 5797
rect 1213 5763 1271 5769
rect 1213 5729 1225 5763
rect 1259 5760 1271 5763
rect 1302 5760 1308 5772
rect 1259 5732 1308 5760
rect 1259 5729 1271 5732
rect 1213 5723 1271 5729
rect 1302 5720 1308 5732
rect 1360 5720 1366 5772
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5692 1455 5695
rect 1780 5692 1808 5791
rect 4154 5788 4160 5800
rect 4212 5788 4218 5840
rect 4249 5831 4307 5837
rect 4249 5797 4261 5831
rect 4295 5828 4307 5831
rect 4522 5828 4528 5840
rect 4295 5800 4528 5828
rect 4295 5797 4307 5800
rect 4249 5791 4307 5797
rect 4522 5788 4528 5800
rect 4580 5788 4586 5840
rect 4982 5788 4988 5840
rect 5040 5788 5046 5840
rect 6546 5828 6552 5840
rect 6507 5800 6552 5828
rect 6546 5788 6552 5800
rect 6604 5788 6610 5840
rect 8202 5788 8208 5840
rect 8260 5828 8266 5840
rect 8260 5800 9260 5828
rect 8260 5788 8266 5800
rect 3878 5720 3884 5772
rect 3936 5760 3942 5772
rect 3936 5732 3981 5760
rect 3936 5720 3942 5732
rect 5810 5720 5816 5772
rect 5868 5760 5874 5772
rect 8573 5763 8631 5769
rect 5868 5732 6408 5760
rect 5868 5720 5874 5732
rect 3234 5692 3240 5704
rect 1443 5664 1532 5692
rect 1780 5664 3240 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 1504 5556 1532 5664
rect 3234 5652 3240 5664
rect 3292 5692 3298 5704
rect 3970 5692 3976 5704
rect 3292 5664 3976 5692
rect 3292 5652 3298 5664
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 4798 5692 4804 5704
rect 4080 5664 4804 5692
rect 1581 5627 1639 5633
rect 1581 5593 1593 5627
rect 1627 5624 1639 5627
rect 4080 5624 4108 5664
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 5994 5692 6000 5704
rect 5955 5664 6000 5692
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 6086 5652 6092 5704
rect 6144 5692 6150 5704
rect 6380 5701 6408 5732
rect 8573 5729 8585 5763
rect 8619 5760 8631 5763
rect 9122 5760 9128 5772
rect 8619 5732 9128 5760
rect 8619 5729 8631 5732
rect 8573 5723 8631 5729
rect 9122 5720 9128 5732
rect 9180 5720 9186 5772
rect 9232 5769 9260 5800
rect 9306 5788 9312 5840
rect 9364 5828 9370 5840
rect 9677 5831 9735 5837
rect 9677 5828 9689 5831
rect 9364 5800 9689 5828
rect 9364 5788 9370 5800
rect 9677 5797 9689 5800
rect 9723 5797 9735 5831
rect 9677 5791 9735 5797
rect 9217 5763 9275 5769
rect 9217 5729 9229 5763
rect 9263 5729 9275 5763
rect 9217 5723 9275 5729
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5729 9551 5763
rect 9953 5763 10011 5769
rect 9953 5760 9965 5763
rect 9493 5723 9551 5729
rect 9692 5732 9965 5760
rect 6181 5695 6239 5701
rect 6181 5692 6193 5695
rect 6144 5664 6193 5692
rect 6144 5652 6150 5664
rect 6181 5661 6193 5664
rect 6227 5661 6239 5695
rect 6181 5655 6239 5661
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 6546 5692 6552 5704
rect 6411 5664 6552 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 1627 5596 4108 5624
rect 6196 5624 6224 5655
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5692 7987 5695
rect 8110 5692 8116 5704
rect 7975 5664 8116 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8812 5664 8953 5692
rect 8812 5652 8818 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 6822 5624 6828 5636
rect 6196 5596 6828 5624
rect 1627 5593 1639 5596
rect 1581 5587 1639 5593
rect 6822 5584 6828 5596
rect 6880 5584 6886 5636
rect 2866 5556 2872 5568
rect 1504 5528 2872 5556
rect 2866 5516 2872 5528
rect 2924 5556 2930 5568
rect 3878 5556 3884 5568
rect 2924 5528 3884 5556
rect 2924 5516 2930 5528
rect 3878 5516 3884 5528
rect 3936 5556 3942 5568
rect 4982 5556 4988 5568
rect 3936 5528 4988 5556
rect 3936 5516 3942 5528
rect 4982 5516 4988 5528
rect 5040 5516 5046 5568
rect 8478 5516 8484 5568
rect 8536 5556 8542 5568
rect 8849 5559 8907 5565
rect 8849 5556 8861 5559
rect 8536 5528 8861 5556
rect 8536 5516 8542 5528
rect 8849 5525 8861 5528
rect 8895 5525 8907 5559
rect 8849 5519 8907 5525
rect 9122 5516 9128 5568
rect 9180 5556 9186 5568
rect 9232 5556 9260 5723
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 9508 5692 9536 5723
rect 9692 5704 9720 5732
rect 9953 5729 9965 5732
rect 9999 5760 10011 5763
rect 10042 5760 10048 5772
rect 9999 5732 10048 5760
rect 9999 5729 10011 5732
rect 9953 5723 10011 5729
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 9364 5664 9536 5692
rect 9364 5652 9370 5664
rect 9674 5652 9680 5704
rect 9732 5652 9738 5704
rect 9646 5596 16574 5624
rect 9180 5528 9260 5556
rect 9180 5516 9186 5528
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 9646 5556 9674 5596
rect 9364 5528 9674 5556
rect 16546 5568 16574 5596
rect 16546 5528 16580 5568
rect 9364 5516 9370 5528
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 920 5466 10396 5488
rect 920 5414 2566 5466
rect 2618 5414 2630 5466
rect 2682 5414 2694 5466
rect 2746 5414 2758 5466
rect 2810 5414 2822 5466
rect 2874 5414 7566 5466
rect 7618 5414 7630 5466
rect 7682 5414 7694 5466
rect 7746 5414 7758 5466
rect 7810 5414 7822 5466
rect 7874 5414 10396 5466
rect 920 5392 10396 5414
rect 1670 5312 1676 5364
rect 1728 5352 1734 5364
rect 2774 5352 2780 5364
rect 1728 5324 2780 5352
rect 1728 5312 1734 5324
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 3694 5352 3700 5364
rect 3655 5324 3700 5352
rect 3694 5312 3700 5324
rect 3752 5312 3758 5364
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 5721 5355 5779 5361
rect 5721 5352 5733 5355
rect 5684 5324 5733 5352
rect 5684 5312 5690 5324
rect 5721 5321 5733 5324
rect 5767 5321 5779 5355
rect 5721 5315 5779 5321
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 7650 5352 7656 5364
rect 7064 5324 7656 5352
rect 7064 5312 7070 5324
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 9306 5352 9312 5364
rect 8168 5324 9312 5352
rect 8168 5312 8174 5324
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 5810 5244 5816 5296
rect 5868 5284 5874 5296
rect 6454 5284 6460 5296
rect 5868 5256 6460 5284
rect 5868 5244 5874 5256
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 8294 5244 8300 5296
rect 8352 5284 8358 5296
rect 9409 5287 9467 5293
rect 9409 5284 9421 5287
rect 8352 5256 9421 5284
rect 8352 5244 8358 5256
rect 9409 5253 9421 5256
rect 9455 5253 9467 5287
rect 9409 5247 9467 5253
rect 2958 5176 2964 5228
rect 3016 5216 3022 5228
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 3016 5188 3341 5216
rect 3016 5176 3022 5188
rect 3329 5185 3341 5188
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 3513 5219 3571 5225
rect 3513 5185 3525 5219
rect 3559 5216 3571 5219
rect 3878 5216 3884 5228
rect 3559 5188 3884 5216
rect 3559 5185 3571 5188
rect 3513 5179 3571 5185
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 5537 5219 5595 5225
rect 5537 5216 5549 5219
rect 4488 5188 5549 5216
rect 4488 5176 4494 5188
rect 5537 5185 5549 5188
rect 5583 5216 5595 5219
rect 7926 5216 7932 5228
rect 5583 5188 7932 5216
rect 5583 5185 5595 5188
rect 5537 5179 5595 5185
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 9769 5219 9827 5225
rect 9769 5185 9781 5219
rect 9815 5216 9827 5219
rect 10318 5216 10324 5228
rect 9815 5188 10324 5216
rect 9815 5185 9827 5188
rect 9769 5179 9827 5185
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 3786 5148 3792 5160
rect 2924 5120 3792 5148
rect 2924 5108 2930 5120
rect 3786 5108 3792 5120
rect 3844 5108 3850 5160
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 6273 5151 6331 5157
rect 6273 5148 6285 5151
rect 6052 5120 6285 5148
rect 6052 5108 6058 5120
rect 6273 5117 6285 5120
rect 6319 5117 6331 5151
rect 6454 5148 6460 5160
rect 6415 5120 6460 5148
rect 6273 5111 6331 5117
rect 6454 5108 6460 5120
rect 6512 5108 6518 5160
rect 6546 5108 6552 5160
rect 6604 5148 6610 5160
rect 6641 5151 6699 5157
rect 6641 5148 6653 5151
rect 6604 5120 6653 5148
rect 6604 5108 6610 5120
rect 6641 5117 6653 5120
rect 6687 5117 6699 5151
rect 7006 5148 7012 5160
rect 6967 5120 7012 5148
rect 6641 5111 6699 5117
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 7466 5148 7472 5160
rect 7423 5120 7472 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5148 8907 5151
rect 9585 5151 9643 5157
rect 9585 5148 9597 5151
rect 8895 5120 9597 5148
rect 8895 5117 8907 5120
rect 8849 5111 8907 5117
rect 9585 5117 9597 5120
rect 9631 5117 9643 5151
rect 9585 5111 9643 5117
rect 9953 5151 10011 5157
rect 9953 5117 9965 5151
rect 9999 5117 10011 5151
rect 9953 5111 10011 5117
rect 8484 5092 8536 5098
rect 6086 5040 6092 5092
rect 6144 5080 6150 5092
rect 6825 5083 6883 5089
rect 6825 5080 6837 5083
rect 6144 5052 6837 5080
rect 6144 5040 6150 5052
rect 6825 5049 6837 5052
rect 6871 5049 6883 5083
rect 6825 5043 6883 5049
rect 9766 5040 9772 5092
rect 9824 5080 9830 5092
rect 9968 5080 9996 5111
rect 10134 5080 10140 5092
rect 9824 5052 10140 5080
rect 9824 5040 9830 5052
rect 10134 5040 10140 5052
rect 10192 5040 10198 5092
rect 8484 5034 8536 5040
rect 9030 5012 9036 5024
rect 8991 4984 9036 5012
rect 9030 4972 9036 4984
rect 9088 4972 9094 5024
rect 3036 4922 10396 4944
rect 3036 4870 5066 4922
rect 5118 4870 5130 4922
rect 5182 4870 5194 4922
rect 5246 4870 5258 4922
rect 5310 4870 5322 4922
rect 5374 4870 10396 4922
rect 3036 4848 10396 4870
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 4028 4780 6224 4808
rect 4028 4768 4034 4780
rect 4798 4700 4804 4752
rect 4856 4700 4862 4752
rect 2958 4632 2964 4684
rect 3016 4672 3022 4684
rect 3234 4672 3240 4684
rect 3016 4644 3240 4672
rect 3016 4632 3022 4644
rect 3234 4632 3240 4644
rect 3292 4672 3298 4684
rect 3421 4675 3479 4681
rect 3421 4672 3433 4675
rect 3292 4644 3433 4672
rect 3292 4632 3298 4644
rect 3421 4641 3433 4644
rect 3467 4641 3479 4675
rect 3878 4672 3884 4684
rect 3839 4644 3884 4672
rect 3421 4635 3479 4641
rect 3878 4632 3884 4644
rect 3936 4632 3942 4684
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 4522 4672 4528 4684
rect 4479 4644 4528 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 5905 4675 5963 4681
rect 5905 4641 5917 4675
rect 5951 4672 5963 4675
rect 6086 4672 6092 4684
rect 5951 4644 6092 4672
rect 5951 4641 5963 4644
rect 5905 4635 5963 4641
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4604 4123 4607
rect 4154 4604 4160 4616
rect 4111 4576 4160 4604
rect 4111 4573 4123 4576
rect 4065 4567 4123 4573
rect 4154 4564 4160 4576
rect 4212 4564 4218 4616
rect 6196 4604 6224 4780
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7377 4811 7435 4817
rect 7377 4808 7389 4811
rect 7064 4780 7389 4808
rect 7064 4768 7070 4780
rect 7377 4777 7389 4780
rect 7423 4777 7435 4811
rect 9582 4808 9588 4820
rect 9543 4780 9588 4808
rect 7377 4771 7435 4777
rect 9582 4768 9588 4780
rect 9640 4768 9646 4820
rect 7926 4740 7932 4752
rect 7484 4712 7932 4740
rect 6546 4632 6552 4684
rect 6604 4672 6610 4684
rect 6733 4675 6791 4681
rect 6733 4672 6745 4675
rect 6604 4644 6745 4672
rect 6604 4632 6610 4644
rect 6733 4641 6745 4644
rect 6779 4641 6791 4675
rect 6733 4635 6791 4641
rect 6822 4632 6828 4684
rect 6880 4672 6886 4684
rect 7484 4681 7512 4712
rect 7926 4700 7932 4712
rect 7984 4700 7990 4752
rect 7009 4675 7067 4681
rect 7009 4672 7021 4675
rect 6880 4644 7021 4672
rect 6880 4632 6886 4644
rect 7009 4641 7021 4644
rect 7055 4641 7067 4675
rect 7009 4635 7067 4641
rect 7469 4675 7527 4681
rect 7469 4641 7481 4675
rect 7515 4641 7527 4675
rect 7650 4672 7656 4684
rect 7611 4644 7656 4672
rect 7469 4635 7527 4641
rect 7650 4632 7656 4644
rect 7708 4632 7714 4684
rect 8297 4675 8355 4681
rect 8297 4672 8309 4675
rect 7760 4644 8309 4672
rect 7760 4604 7788 4644
rect 8297 4641 8309 4644
rect 8343 4641 8355 4675
rect 8297 4635 8355 4641
rect 6196 4576 7788 4604
rect 7929 4607 7987 4613
rect 7929 4573 7941 4607
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 8021 4607 8079 4613
rect 8021 4573 8033 4607
rect 8067 4604 8079 4607
rect 8386 4604 8392 4616
rect 8067 4576 8392 4604
rect 8067 4573 8079 4576
rect 8021 4567 8079 4573
rect 5994 4496 6000 4548
rect 6052 4536 6058 4548
rect 6638 4536 6644 4548
rect 6052 4508 6644 4536
rect 6052 4496 6058 4508
rect 6638 4496 6644 4508
rect 6696 4496 6702 4548
rect 6914 4536 6920 4548
rect 6875 4508 6920 4536
rect 6914 4496 6920 4508
rect 6972 4496 6978 4548
rect 7282 4496 7288 4548
rect 7340 4536 7346 4548
rect 7944 4536 7972 4567
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 7340 4508 7972 4536
rect 7340 4496 7346 4508
rect 3789 4471 3847 4477
rect 3789 4437 3801 4471
rect 3835 4468 3847 4471
rect 4614 4468 4620 4480
rect 3835 4440 4620 4468
rect 3835 4437 3847 4440
rect 3789 4431 3847 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 6086 4428 6092 4480
rect 6144 4468 6150 4480
rect 6465 4471 6523 4477
rect 6465 4468 6477 4471
rect 6144 4440 6477 4468
rect 6144 4428 6150 4440
rect 6465 4437 6477 4440
rect 6511 4437 6523 4471
rect 6465 4431 6523 4437
rect 3036 4378 10396 4400
rect 3036 4326 7566 4378
rect 7618 4326 7630 4378
rect 7682 4326 7694 4378
rect 7746 4326 7758 4378
rect 7810 4326 7822 4378
rect 7874 4326 10396 4378
rect 3036 4304 10396 4326
rect 3786 4088 3792 4140
rect 3844 4128 3850 4140
rect 4890 4128 4896 4140
rect 3844 4100 4896 4128
rect 3844 4088 3850 4100
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 9398 4128 9404 4140
rect 5123 4100 7972 4128
rect 9359 4100 9404 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 3329 4063 3387 4069
rect 3329 4029 3341 4063
rect 3375 4060 3387 4063
rect 4338 4060 4344 4072
rect 3375 4032 4344 4060
rect 3375 4029 3387 4032
rect 3329 4023 3387 4029
rect 4338 4020 4344 4032
rect 4396 4020 4402 4072
rect 5169 4063 5227 4069
rect 5169 4029 5181 4063
rect 5215 4029 5227 4063
rect 5350 4060 5356 4072
rect 5311 4032 5356 4060
rect 5169 4023 5227 4029
rect 4890 3952 4896 4004
rect 4948 3992 4954 4004
rect 5184 3992 5212 4023
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 5534 4060 5540 4072
rect 5495 4032 5540 4060
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5626 4020 5632 4072
rect 5684 4060 5690 4072
rect 5721 4063 5779 4069
rect 5721 4060 5733 4063
rect 5684 4032 5733 4060
rect 5684 4020 5690 4032
rect 5721 4029 5733 4032
rect 5767 4060 5779 4063
rect 5810 4060 5816 4072
rect 5767 4032 5816 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 5810 4020 5816 4032
rect 5868 4020 5874 4072
rect 6270 4060 6276 4072
rect 6231 4032 6276 4060
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 5442 3992 5448 4004
rect 4948 3964 5448 3992
rect 4948 3952 4954 3964
rect 5442 3952 5448 3964
rect 5500 3952 5506 4004
rect 5905 3927 5963 3933
rect 5905 3893 5917 3927
rect 5951 3924 5963 3927
rect 5994 3924 6000 3936
rect 5951 3896 6000 3924
rect 5951 3893 5963 3896
rect 5905 3887 5963 3893
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 7944 3924 7972 4100
rect 9398 4088 9404 4100
rect 9456 4088 9462 4140
rect 8481 4063 8539 4069
rect 8481 4029 8493 4063
rect 8527 4060 8539 4063
rect 8570 4060 8576 4072
rect 8527 4032 8576 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 12406 4032 16574 4060
rect 8021 3995 8079 4001
rect 8021 3961 8033 3995
rect 8067 3992 8079 3995
rect 12406 3992 12434 4032
rect 8067 3964 12434 3992
rect 16546 4004 16574 4032
rect 16546 3964 16580 4004
rect 8067 3961 8079 3964
rect 8021 3955 8079 3961
rect 16574 3952 16580 3964
rect 16632 3952 16638 4004
rect 22094 3924 22100 3936
rect 7944 3896 22100 3924
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 3036 3834 10396 3856
rect 3036 3782 5066 3834
rect 5118 3782 5130 3834
rect 5182 3782 5194 3834
rect 5246 3782 5258 3834
rect 5310 3782 5322 3834
rect 5374 3782 10396 3834
rect 3036 3760 10396 3782
rect 6638 3680 6644 3732
rect 6696 3720 6702 3732
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 6696 3692 8953 3720
rect 6696 3680 6702 3692
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 8941 3683 8999 3689
rect 9490 3680 9496 3732
rect 9548 3720 9554 3732
rect 9585 3723 9643 3729
rect 9585 3720 9597 3723
rect 9548 3692 9597 3720
rect 9548 3680 9554 3692
rect 9585 3689 9597 3692
rect 9631 3689 9643 3723
rect 9585 3683 9643 3689
rect 3878 3612 3884 3664
rect 3936 3612 3942 3664
rect 9030 3612 9036 3664
rect 9088 3652 9094 3664
rect 9125 3655 9183 3661
rect 9125 3652 9137 3655
rect 9088 3624 9137 3652
rect 9088 3612 9094 3624
rect 9125 3621 9137 3624
rect 9171 3621 9183 3655
rect 9125 3615 9183 3621
rect 3513 3587 3571 3593
rect 3513 3553 3525 3587
rect 3559 3584 3571 3587
rect 3896 3584 3924 3612
rect 3559 3556 3924 3584
rect 3973 3587 4031 3593
rect 3559 3553 3571 3556
rect 3513 3547 3571 3553
rect 3973 3553 3985 3587
rect 4019 3584 4031 3587
rect 4062 3584 4068 3596
rect 4019 3556 4068 3584
rect 4019 3553 4031 3556
rect 3973 3547 4031 3553
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 6086 3584 6092 3596
rect 6047 3556 6092 3584
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6362 3584 6368 3596
rect 6323 3556 6368 3584
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 8757 3587 8815 3593
rect 8757 3553 8769 3587
rect 8803 3584 8815 3587
rect 9582 3584 9588 3596
rect 8803 3556 9588 3584
rect 8803 3553 8815 3556
rect 8757 3547 8815 3553
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 9766 3584 9772 3596
rect 9727 3556 9772 3584
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 3881 3519 3939 3525
rect 3881 3485 3893 3519
rect 3927 3516 3939 3519
rect 4798 3516 4804 3528
rect 3927 3488 4804 3516
rect 3927 3485 3939 3488
rect 3881 3479 3939 3485
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5074 3516 5080 3528
rect 5035 3488 5080 3516
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 8573 3519 8631 3525
rect 8573 3516 8585 3519
rect 5184 3488 8585 3516
rect 2682 3408 2688 3460
rect 2740 3448 2746 3460
rect 5184 3448 5212 3488
rect 8573 3485 8585 3488
rect 8619 3485 8631 3519
rect 16666 3516 16672 3528
rect 8573 3479 8631 3485
rect 9324 3488 16672 3516
rect 2740 3420 5212 3448
rect 8113 3451 8171 3457
rect 2740 3408 2746 3420
rect 8113 3417 8125 3451
rect 8159 3448 8171 3451
rect 9324 3448 9352 3488
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 8159 3420 9352 3448
rect 9401 3451 9459 3457
rect 8159 3417 8171 3420
rect 8113 3411 8171 3417
rect 9401 3417 9413 3451
rect 9447 3417 9459 3451
rect 9401 3411 9459 3417
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 8389 3383 8447 3389
rect 8389 3380 8401 3383
rect 5040 3352 8401 3380
rect 5040 3340 5046 3352
rect 8389 3349 8401 3352
rect 8435 3349 8447 3383
rect 8389 3343 8447 3349
rect 9214 3340 9220 3392
rect 9272 3380 9278 3392
rect 9416 3380 9444 3411
rect 9272 3352 9444 3380
rect 9272 3340 9278 3352
rect 9490 3340 9496 3392
rect 9548 3380 9554 3392
rect 9953 3383 10011 3389
rect 9953 3380 9965 3383
rect 9548 3352 9965 3380
rect 9548 3340 9554 3352
rect 9953 3349 9965 3352
rect 9999 3349 10011 3383
rect 9953 3343 10011 3349
rect 3036 3290 10396 3312
rect 3036 3238 7566 3290
rect 7618 3238 7630 3290
rect 7682 3238 7694 3290
rect 7746 3238 7758 3290
rect 7810 3238 7822 3290
rect 7874 3238 10396 3290
rect 3036 3216 10396 3238
rect 3602 3136 3608 3188
rect 3660 3176 3666 3188
rect 5261 3179 5319 3185
rect 5261 3176 5273 3179
rect 3660 3148 5273 3176
rect 3660 3136 3666 3148
rect 5261 3145 5273 3148
rect 5307 3145 5319 3179
rect 5994 3176 6000 3188
rect 5907 3148 6000 3176
rect 5261 3139 5319 3145
rect 5994 3136 6000 3148
rect 6052 3176 6058 3188
rect 6730 3176 6736 3188
rect 6052 3148 6736 3176
rect 6052 3136 6058 3148
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 4338 3068 4344 3120
rect 4396 3108 4402 3120
rect 4617 3111 4675 3117
rect 4617 3108 4629 3111
rect 4396 3080 4629 3108
rect 4396 3068 4402 3080
rect 4617 3077 4629 3080
rect 4663 3108 4675 3111
rect 4982 3108 4988 3120
rect 4663 3080 4988 3108
rect 4663 3077 4675 3080
rect 4617 3071 4675 3077
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 5537 3111 5595 3117
rect 5537 3077 5549 3111
rect 5583 3108 5595 3111
rect 7282 3108 7288 3120
rect 5583 3080 7288 3108
rect 5583 3077 5595 3080
rect 5537 3071 5595 3077
rect 7282 3068 7288 3080
rect 7340 3108 7346 3120
rect 9214 3108 9220 3120
rect 7340 3080 9220 3108
rect 7340 3068 7346 3080
rect 9214 3068 9220 3080
rect 9272 3068 9278 3120
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 5721 3043 5779 3049
rect 5721 3040 5733 3043
rect 4120 3012 5733 3040
rect 4120 3000 4126 3012
rect 5721 3009 5733 3012
rect 5767 3040 5779 3043
rect 6454 3040 6460 3052
rect 5767 3012 6460 3040
rect 5767 3009 5779 3012
rect 5721 3003 5779 3009
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 6822 3040 6828 3052
rect 6783 3012 6828 3040
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 7248 3012 8156 3040
rect 7248 3000 7254 3012
rect 2866 2932 2872 2984
rect 2924 2972 2930 2984
rect 3329 2975 3387 2981
rect 3329 2972 3341 2975
rect 2924 2944 3341 2972
rect 2924 2932 2930 2944
rect 3329 2941 3341 2944
rect 3375 2941 3387 2975
rect 3329 2935 3387 2941
rect 4982 2932 4988 2984
rect 5040 2972 5046 2984
rect 8128 2981 8156 3012
rect 5353 2975 5411 2981
rect 5353 2972 5365 2975
rect 5040 2944 5365 2972
rect 5040 2932 5046 2944
rect 5353 2941 5365 2944
rect 5399 2941 5411 2975
rect 5353 2935 5411 2941
rect 8021 2975 8079 2981
rect 8021 2941 8033 2975
rect 8067 2941 8079 2975
rect 8021 2935 8079 2941
rect 8113 2975 8171 2981
rect 8113 2941 8125 2975
rect 8159 2941 8171 2975
rect 8113 2935 8171 2941
rect 8036 2904 8064 2935
rect 8662 2904 8668 2916
rect 8036 2876 8668 2904
rect 8662 2864 8668 2876
rect 8720 2864 8726 2916
rect 10045 2907 10103 2913
rect 10045 2873 10057 2907
rect 10091 2904 10103 2907
rect 16850 2904 16856 2916
rect 10091 2876 16856 2904
rect 10091 2873 10103 2876
rect 10045 2867 10103 2873
rect 16850 2864 16856 2876
rect 16908 2864 16914 2916
rect 3036 2746 10396 2768
rect 3036 2694 5066 2746
rect 5118 2694 5130 2746
rect 5182 2694 5194 2746
rect 5246 2694 5258 2746
rect 5310 2694 5322 2746
rect 5374 2694 10396 2746
rect 3036 2672 10396 2694
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 3789 2635 3847 2641
rect 3789 2632 3801 2635
rect 2832 2604 3801 2632
rect 2832 2592 2838 2604
rect 3789 2601 3801 2604
rect 3835 2601 3847 2635
rect 3789 2595 3847 2601
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 4246 2632 4252 2644
rect 4203 2604 4252 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4430 2592 4436 2644
rect 4488 2592 4494 2644
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 5169 2635 5227 2641
rect 5169 2632 5181 2635
rect 5040 2604 5181 2632
rect 5040 2592 5046 2604
rect 5169 2601 5181 2604
rect 5215 2632 5227 2635
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 5215 2604 5365 2632
rect 5215 2601 5227 2604
rect 5169 2595 5227 2601
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 5994 2632 6000 2644
rect 5955 2604 6000 2632
rect 5353 2595 5411 2601
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 7282 2592 7288 2644
rect 7340 2632 7346 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 7340 2604 8953 2632
rect 7340 2592 7346 2604
rect 4448 2564 4476 2592
rect 4080 2536 4568 2564
rect 3602 2496 3608 2508
rect 3563 2468 3608 2496
rect 3602 2456 3608 2468
rect 3660 2456 3666 2508
rect 3786 2456 3792 2508
rect 3844 2496 3850 2508
rect 4080 2505 4108 2536
rect 3973 2499 4031 2505
rect 3973 2496 3985 2499
rect 3844 2468 3985 2496
rect 3844 2456 3850 2468
rect 3973 2465 3985 2468
rect 4019 2465 4031 2499
rect 3973 2459 4031 2465
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 4154 2456 4160 2508
rect 4212 2496 4218 2508
rect 4540 2505 4568 2536
rect 4433 2499 4491 2505
rect 4433 2496 4445 2499
rect 4212 2468 4445 2496
rect 4212 2456 4218 2468
rect 4433 2465 4445 2468
rect 4479 2465 4491 2499
rect 4433 2459 4491 2465
rect 4525 2499 4583 2505
rect 4525 2465 4537 2499
rect 4571 2465 4583 2499
rect 4525 2459 4583 2465
rect 4801 2499 4859 2505
rect 4801 2465 4813 2499
rect 4847 2465 4859 2499
rect 4801 2459 4859 2465
rect 3326 2388 3332 2440
rect 3384 2428 3390 2440
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 3384 2400 4721 2428
rect 3384 2388 3390 2400
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 3970 2320 3976 2372
rect 4028 2360 4034 2372
rect 4816 2360 4844 2459
rect 4890 2456 4896 2508
rect 4948 2496 4954 2508
rect 4985 2499 5043 2505
rect 4985 2496 4997 2499
rect 4948 2468 4997 2496
rect 4948 2456 4954 2468
rect 4985 2465 4997 2468
rect 5031 2465 5043 2499
rect 4985 2459 5043 2465
rect 8113 2499 8171 2505
rect 8113 2465 8125 2499
rect 8159 2496 8171 2499
rect 8294 2496 8300 2508
rect 8159 2468 8300 2496
rect 8159 2465 8171 2468
rect 8113 2459 8171 2465
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 8386 2456 8392 2508
rect 8444 2494 8450 2508
rect 8573 2499 8631 2505
rect 8573 2494 8585 2499
rect 8444 2466 8585 2494
rect 8444 2456 8450 2466
rect 8573 2465 8585 2466
rect 8619 2465 8631 2499
rect 8573 2459 8631 2465
rect 7469 2431 7527 2437
rect 4028 2332 4844 2360
rect 5368 2400 6592 2428
rect 4028 2320 4034 2332
rect 3421 2295 3479 2301
rect 3421 2261 3433 2295
rect 3467 2292 3479 2295
rect 5368 2292 5396 2400
rect 5626 2292 5632 2304
rect 3467 2264 5396 2292
rect 5587 2264 5632 2292
rect 3467 2261 3479 2264
rect 3421 2255 3479 2261
rect 5626 2252 5632 2264
rect 5684 2252 5690 2304
rect 5810 2252 5816 2304
rect 5868 2292 5874 2304
rect 5905 2295 5963 2301
rect 5905 2292 5917 2295
rect 5868 2264 5917 2292
rect 5868 2252 5874 2264
rect 5905 2261 5917 2264
rect 5951 2292 5963 2295
rect 6086 2292 6092 2304
rect 5951 2264 6092 2292
rect 5951 2261 5963 2264
rect 5905 2255 5963 2261
rect 6086 2252 6092 2264
rect 6144 2252 6150 2304
rect 6564 2292 6592 2400
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 8680 2428 8708 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 9861 2635 9919 2641
rect 9861 2632 9873 2635
rect 9640 2604 9873 2632
rect 9640 2592 9646 2604
rect 9861 2601 9873 2604
rect 9907 2601 9919 2635
rect 9861 2595 9919 2601
rect 10042 2592 10048 2644
rect 10100 2592 10106 2644
rect 8846 2524 8852 2576
rect 8904 2564 8910 2576
rect 9493 2567 9551 2573
rect 9493 2564 9505 2567
rect 8904 2536 9505 2564
rect 8904 2524 8910 2536
rect 9493 2533 9505 2536
rect 9539 2533 9551 2567
rect 10060 2564 10088 2592
rect 9493 2527 9551 2533
rect 9600 2536 10088 2564
rect 8754 2456 8760 2508
rect 8812 2496 8818 2508
rect 9309 2499 9367 2505
rect 9309 2496 9321 2499
rect 8812 2468 8857 2496
rect 8956 2468 9321 2496
rect 8812 2456 8818 2468
rect 8956 2428 8984 2468
rect 9309 2465 9321 2468
rect 9355 2465 9367 2499
rect 9309 2459 9367 2465
rect 7515 2400 8524 2428
rect 8680 2400 8984 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 8110 2320 8116 2372
rect 8168 2360 8174 2372
rect 8389 2363 8447 2369
rect 8389 2360 8401 2363
rect 8168 2332 8401 2360
rect 8168 2320 8174 2332
rect 8389 2329 8401 2332
rect 8435 2329 8447 2363
rect 8496 2360 8524 2400
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 9088 2400 9137 2428
rect 9088 2388 9094 2400
rect 9125 2397 9137 2400
rect 9171 2428 9183 2431
rect 9214 2428 9220 2440
rect 9171 2400 9220 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 9600 2428 9628 2536
rect 10042 2496 10048 2508
rect 10003 2468 10048 2496
rect 10042 2456 10048 2468
rect 10100 2496 10106 2508
rect 16942 2496 16948 2508
rect 10100 2468 16948 2496
rect 10100 2456 10106 2468
rect 16942 2456 16948 2468
rect 17000 2456 17006 2508
rect 9324 2400 9628 2428
rect 9324 2360 9352 2400
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 9784 2360 9812 2388
rect 8496 2332 9352 2360
rect 9600 2332 9812 2360
rect 8389 2323 8447 2329
rect 9600 2292 9628 2332
rect 6564 2264 9628 2292
rect 9677 2295 9735 2301
rect 9677 2261 9689 2295
rect 9723 2292 9735 2295
rect 9766 2292 9772 2304
rect 9723 2264 9772 2292
rect 9723 2261 9735 2264
rect 9677 2255 9735 2261
rect 9766 2252 9772 2264
rect 9824 2292 9830 2304
rect 10134 2292 10140 2304
rect 9824 2264 10140 2292
rect 9824 2252 9830 2264
rect 10134 2252 10140 2264
rect 10192 2252 10198 2304
rect 3036 2202 10396 2224
rect 3036 2150 7566 2202
rect 7618 2150 7630 2202
rect 7682 2150 7694 2202
rect 7746 2150 7758 2202
rect 7810 2150 7822 2202
rect 7874 2150 10396 2202
rect 3036 2128 10396 2150
rect 3234 2048 3240 2100
rect 3292 2088 3298 2100
rect 3329 2091 3387 2097
rect 3329 2088 3341 2091
rect 3292 2060 3341 2088
rect 3292 2048 3298 2060
rect 3329 2057 3341 2060
rect 3375 2057 3387 2091
rect 3510 2088 3516 2100
rect 3471 2060 3516 2088
rect 3329 2051 3387 2057
rect 3510 2048 3516 2060
rect 3568 2048 3574 2100
rect 3878 2048 3884 2100
rect 3936 2088 3942 2100
rect 3973 2091 4031 2097
rect 3973 2088 3985 2091
rect 3936 2060 3985 2088
rect 3936 2048 3942 2060
rect 3973 2057 3985 2060
rect 4019 2057 4031 2091
rect 3973 2051 4031 2057
rect 4062 2048 4068 2100
rect 4120 2088 4126 2100
rect 4157 2091 4215 2097
rect 4157 2088 4169 2091
rect 4120 2060 4169 2088
rect 4120 2048 4126 2060
rect 4157 2057 4169 2060
rect 4203 2057 4215 2091
rect 4157 2051 4215 2057
rect 4433 2091 4491 2097
rect 4433 2057 4445 2091
rect 4479 2088 4491 2091
rect 4614 2088 4620 2100
rect 4479 2060 4620 2088
rect 4479 2057 4491 2060
rect 4433 2051 4491 2057
rect 4614 2048 4620 2060
rect 4672 2048 4678 2100
rect 5997 2091 6055 2097
rect 5997 2057 6009 2091
rect 6043 2088 6055 2091
rect 10042 2088 10048 2100
rect 6043 2060 10048 2088
rect 6043 2057 6055 2060
rect 5997 2051 6055 2057
rect 10042 2048 10048 2060
rect 10100 2048 10106 2100
rect 3050 1980 3056 2032
rect 3108 2020 3114 2032
rect 3697 2023 3755 2029
rect 3697 2020 3709 2023
rect 3108 1992 3709 2020
rect 3108 1980 3114 1992
rect 3697 1989 3709 1992
rect 3743 1989 3755 2023
rect 3697 1983 3755 1989
rect 8110 1980 8116 2032
rect 8168 2020 8174 2032
rect 16574 2020 16580 2032
rect 8168 1992 16580 2020
rect 8168 1980 8174 1992
rect 16574 1980 16580 1992
rect 16632 1980 16638 2032
rect 6822 1952 6828 1964
rect 6783 1924 6828 1952
rect 6822 1912 6828 1924
rect 6880 1912 6886 1964
rect 22278 1952 22284 1964
rect 6932 1924 22284 1952
rect 3602 1844 3608 1896
rect 3660 1884 3666 1896
rect 4617 1887 4675 1893
rect 4617 1884 4629 1887
rect 3660 1856 4629 1884
rect 3660 1844 3666 1856
rect 4617 1853 4629 1856
rect 4663 1884 4675 1887
rect 6932 1884 6960 1924
rect 22278 1912 22284 1924
rect 22336 1912 22342 1964
rect 8018 1884 8024 1896
rect 4663 1856 6960 1884
rect 7979 1856 8024 1884
rect 4663 1853 4675 1856
rect 4617 1847 4675 1853
rect 8018 1844 8024 1856
rect 8076 1844 8082 1896
rect 8113 1887 8171 1893
rect 8113 1853 8125 1887
rect 8159 1884 8171 1887
rect 9858 1884 9864 1896
rect 8159 1856 9720 1884
rect 9819 1856 9864 1884
rect 8159 1853 8171 1856
rect 8113 1847 8171 1853
rect 8570 1776 8576 1828
rect 8628 1816 8634 1828
rect 9306 1816 9312 1828
rect 8628 1788 9312 1816
rect 8628 1776 8634 1788
rect 9306 1776 9312 1788
rect 9364 1776 9370 1828
rect 9692 1816 9720 1856
rect 9858 1844 9864 1856
rect 9916 1844 9922 1896
rect 16758 1816 16764 1828
rect 9692 1788 16764 1816
rect 16758 1776 16764 1788
rect 16816 1776 16822 1828
rect 5813 1751 5871 1757
rect 5813 1717 5825 1751
rect 5859 1748 5871 1751
rect 10042 1748 10048 1760
rect 5859 1720 10048 1748
rect 5859 1717 5871 1720
rect 5813 1711 5871 1717
rect 10042 1708 10048 1720
rect 10100 1708 10106 1760
rect 3036 1658 10396 1680
rect 3036 1606 5066 1658
rect 5118 1606 5130 1658
rect 5182 1606 5194 1658
rect 5246 1606 5258 1658
rect 5310 1606 5322 1658
rect 5374 1606 10396 1658
rect 3036 1584 10396 1606
rect 3234 1504 3240 1556
rect 3292 1544 3298 1556
rect 3329 1547 3387 1553
rect 3329 1544 3341 1547
rect 3292 1516 3341 1544
rect 3292 1504 3298 1516
rect 3329 1513 3341 1516
rect 3375 1513 3387 1547
rect 3329 1507 3387 1513
rect 3605 1547 3663 1553
rect 3605 1513 3617 1547
rect 3651 1544 3663 1547
rect 5534 1544 5540 1556
rect 3651 1516 5540 1544
rect 3651 1513 3663 1516
rect 3605 1507 3663 1513
rect 5534 1504 5540 1516
rect 5592 1504 5598 1556
rect 8110 1544 8116 1556
rect 8071 1516 8116 1544
rect 8110 1504 8116 1516
rect 8168 1504 8174 1556
rect 8938 1504 8944 1556
rect 8996 1544 9002 1556
rect 9033 1547 9091 1553
rect 9033 1544 9045 1547
rect 8996 1516 9045 1544
rect 8996 1504 9002 1516
rect 9033 1513 9045 1516
rect 9079 1513 9091 1547
rect 9033 1507 9091 1513
rect 9122 1504 9128 1556
rect 9180 1544 9186 1556
rect 9677 1547 9735 1553
rect 9677 1544 9689 1547
rect 9180 1516 9689 1544
rect 9180 1504 9186 1516
rect 9677 1513 9689 1516
rect 9723 1513 9735 1547
rect 9677 1507 9735 1513
rect 9214 1476 9220 1488
rect 6012 1448 9220 1476
rect 6012 1417 6040 1448
rect 9214 1436 9220 1448
rect 9272 1436 9278 1488
rect 5997 1411 6055 1417
rect 5997 1377 6009 1411
rect 6043 1377 6055 1411
rect 6178 1408 6184 1420
rect 6139 1380 6184 1408
rect 5997 1371 6055 1377
rect 6178 1368 6184 1380
rect 6236 1368 6242 1420
rect 8846 1408 8852 1420
rect 8807 1380 8852 1408
rect 8846 1368 8852 1380
rect 8904 1368 8910 1420
rect 9493 1411 9551 1417
rect 9493 1377 9505 1411
rect 9539 1408 9551 1411
rect 9582 1408 9588 1420
rect 9539 1380 9588 1408
rect 9539 1377 9551 1380
rect 9493 1371 9551 1377
rect 9582 1368 9588 1380
rect 9640 1368 9646 1420
rect 9861 1411 9919 1417
rect 9861 1377 9873 1411
rect 9907 1408 9919 1411
rect 9953 1411 10011 1417
rect 9953 1408 9965 1411
rect 9907 1380 9965 1408
rect 9907 1377 9919 1380
rect 9861 1371 9919 1377
rect 9953 1377 9965 1380
rect 9999 1408 10011 1411
rect 10318 1408 10324 1420
rect 9999 1380 10324 1408
rect 9999 1377 10011 1380
rect 9953 1371 10011 1377
rect 5442 1340 5448 1352
rect 5403 1312 5448 1340
rect 5442 1300 5448 1312
rect 5500 1300 5506 1352
rect 6086 1300 6092 1352
rect 6144 1340 6150 1352
rect 8481 1343 8539 1349
rect 8481 1340 8493 1343
rect 6144 1312 8493 1340
rect 6144 1300 6150 1312
rect 8481 1309 8493 1312
rect 8527 1309 8539 1343
rect 8481 1303 8539 1309
rect 9306 1300 9312 1352
rect 9364 1340 9370 1352
rect 9876 1340 9904 1371
rect 10318 1368 10324 1380
rect 10376 1368 10382 1420
rect 9364 1312 9904 1340
rect 9364 1300 9370 1312
rect 8754 1272 8760 1284
rect 2746 1244 8760 1272
rect 2314 1164 2320 1216
rect 2372 1204 2378 1216
rect 2746 1204 2774 1244
rect 8754 1232 8760 1244
rect 8812 1232 8818 1284
rect 10226 1272 10232 1284
rect 9140 1244 10232 1272
rect 2372 1176 2774 1204
rect 2372 1164 2378 1176
rect 5626 1164 5632 1216
rect 5684 1204 5690 1216
rect 8297 1207 8355 1213
rect 8297 1204 8309 1207
rect 5684 1176 8309 1204
rect 5684 1164 5690 1176
rect 8297 1173 8309 1176
rect 8343 1204 8355 1207
rect 8570 1204 8576 1216
rect 8343 1176 8576 1204
rect 8343 1173 8355 1176
rect 8297 1167 8355 1173
rect 8570 1164 8576 1176
rect 8628 1164 8634 1216
rect 8665 1207 8723 1213
rect 8665 1173 8677 1207
rect 8711 1204 8723 1207
rect 9140 1204 9168 1244
rect 10226 1232 10232 1244
rect 10284 1232 10290 1284
rect 9306 1204 9312 1216
rect 8711 1176 9168 1204
rect 9267 1176 9312 1204
rect 8711 1173 8723 1176
rect 8665 1167 8723 1173
rect 9306 1164 9312 1176
rect 9364 1164 9370 1216
rect 920 1114 10396 1136
rect 920 1062 2566 1114
rect 2618 1062 2630 1114
rect 2682 1062 2694 1114
rect 2746 1062 2758 1114
rect 2810 1062 2822 1114
rect 2874 1062 7566 1114
rect 7618 1062 7630 1114
rect 7682 1062 7694 1114
rect 7746 1062 7758 1114
rect 7810 1062 7822 1114
rect 7874 1062 10396 1114
rect 920 1040 10396 1062
rect 1118 960 1124 1012
rect 1176 1000 1182 1012
rect 1305 1003 1363 1009
rect 1305 1000 1317 1003
rect 1176 972 1317 1000
rect 1176 960 1182 972
rect 1305 969 1317 972
rect 1351 969 1363 1003
rect 1305 963 1363 969
rect 1857 1003 1915 1009
rect 1857 969 1869 1003
rect 1903 1000 1915 1003
rect 2406 1000 2412 1012
rect 1903 972 2412 1000
rect 1903 969 1915 972
rect 1857 963 1915 969
rect 2406 960 2412 972
rect 2464 960 2470 1012
rect 2958 1000 2964 1012
rect 2871 972 2964 1000
rect 2958 960 2964 972
rect 3016 1000 3022 1012
rect 3145 1003 3203 1009
rect 3145 1000 3157 1003
rect 3016 972 3157 1000
rect 3016 960 3022 972
rect 3145 969 3157 972
rect 3191 1000 3203 1003
rect 3329 1003 3387 1009
rect 3329 1000 3341 1003
rect 3191 972 3341 1000
rect 3191 969 3203 972
rect 3145 963 3203 969
rect 3329 969 3341 972
rect 3375 1000 3387 1003
rect 3697 1003 3755 1009
rect 3697 1000 3709 1003
rect 3375 972 3709 1000
rect 3375 969 3387 972
rect 3329 963 3387 969
rect 3697 969 3709 972
rect 3743 1000 3755 1003
rect 3881 1003 3939 1009
rect 3881 1000 3893 1003
rect 3743 972 3893 1000
rect 3743 969 3755 972
rect 3697 963 3755 969
rect 3881 969 3893 972
rect 3927 1000 3939 1003
rect 4982 1000 4988 1012
rect 3927 972 4988 1000
rect 3927 969 3939 972
rect 3881 963 3939 969
rect 4982 960 4988 972
rect 5040 960 5046 1012
rect 8754 1000 8760 1012
rect 8715 972 8760 1000
rect 8754 960 8760 972
rect 8812 960 8818 1012
rect 9030 1000 9036 1012
rect 8991 972 9036 1000
rect 9030 960 9036 972
rect 9088 960 9094 1012
rect 9674 1000 9680 1012
rect 9635 972 9680 1000
rect 9674 960 9680 972
rect 9732 960 9738 1012
rect 9861 1003 9919 1009
rect 9861 969 9873 1003
rect 9907 1000 9919 1003
rect 9950 1000 9956 1012
rect 9907 972 9956 1000
rect 9907 969 9919 972
rect 9861 963 9919 969
rect 9950 960 9956 972
rect 10008 960 10014 1012
rect 1581 935 1639 941
rect 1581 901 1593 935
rect 1627 932 1639 935
rect 3418 932 3424 944
rect 1627 904 3424 932
rect 1627 901 1639 904
rect 1581 895 1639 901
rect 3418 892 3424 904
rect 3476 892 3482 944
rect 7653 935 7711 941
rect 7653 901 7665 935
rect 7699 932 7711 935
rect 13814 932 13820 944
rect 7699 904 13820 932
rect 7699 901 7711 904
rect 7653 895 7711 901
rect 13814 892 13820 904
rect 13872 892 13878 944
rect 2133 867 2191 873
rect 2133 833 2145 867
rect 2179 864 2191 867
rect 5902 864 5908 876
rect 2179 836 5908 864
rect 2179 833 2191 836
rect 2133 827 2191 833
rect 5902 824 5908 836
rect 5960 824 5966 876
rect 9125 867 9183 873
rect 9125 864 9137 867
rect 6012 836 9137 864
rect 1213 799 1271 805
rect 1213 765 1225 799
rect 1259 796 1271 799
rect 1489 799 1547 805
rect 1489 796 1501 799
rect 1259 768 1501 796
rect 1259 765 1271 768
rect 1213 759 1271 765
rect 1489 765 1501 768
rect 1535 796 1547 799
rect 1765 799 1823 805
rect 1765 796 1777 799
rect 1535 768 1777 796
rect 1535 765 1547 768
rect 1489 759 1547 765
rect 1765 765 1777 768
rect 1811 796 1823 799
rect 2041 799 2099 805
rect 2041 796 2053 799
rect 1811 768 2053 796
rect 1811 765 1823 768
rect 1765 759 1823 765
rect 2041 765 2053 768
rect 2087 796 2099 799
rect 2958 796 2964 808
rect 2087 768 2964 796
rect 2087 765 2099 768
rect 2041 759 2099 765
rect 2958 756 2964 768
rect 3016 756 3022 808
rect 6012 805 6040 836
rect 9125 833 9137 836
rect 9171 833 9183 867
rect 9125 827 9183 833
rect 9493 867 9551 873
rect 9493 833 9505 867
rect 9539 864 9551 867
rect 9766 864 9772 876
rect 9539 836 9772 864
rect 9539 833 9551 836
rect 9493 827 9551 833
rect 9766 824 9772 836
rect 9824 824 9830 876
rect 5997 799 6055 805
rect 5997 765 6009 799
rect 6043 765 6055 799
rect 5997 759 6055 765
rect 8573 799 8631 805
rect 8573 765 8585 799
rect 8619 796 8631 799
rect 9306 796 9312 808
rect 8619 768 9312 796
rect 8619 765 8631 768
rect 8573 759 8631 765
rect 9306 756 9312 768
rect 9364 756 9370 808
rect 10042 796 10048 808
rect 10003 768 10048 796
rect 10042 756 10048 768
rect 10100 756 10106 808
rect 2409 731 2467 737
rect 2409 697 2421 731
rect 2455 728 2467 731
rect 3050 728 3056 740
rect 2455 700 3056 728
rect 2455 697 2467 700
rect 2409 691 2467 697
rect 3050 688 3056 700
rect 3108 688 3114 740
rect 5626 728 5632 740
rect 5000 700 5632 728
rect 2314 620 2320 672
rect 2372 660 2378 672
rect 2501 663 2559 669
rect 2501 660 2513 663
rect 2372 632 2513 660
rect 2372 620 2378 632
rect 2501 629 2513 632
rect 2547 629 2559 663
rect 2501 623 2559 629
rect 2777 663 2835 669
rect 2777 629 2789 663
rect 2823 660 2835 663
rect 5000 660 5028 700
rect 5626 688 5632 700
rect 5684 728 5690 740
rect 6273 731 6331 737
rect 6273 728 6285 731
rect 5684 700 6285 728
rect 5684 688 5690 700
rect 6273 697 6285 700
rect 6319 697 6331 731
rect 6273 691 6331 697
rect 6549 731 6607 737
rect 6549 697 6561 731
rect 6595 728 6607 731
rect 8846 728 8852 740
rect 6595 700 8852 728
rect 6595 697 6607 700
rect 6549 691 6607 697
rect 8846 688 8852 700
rect 8904 688 8910 740
rect 2823 632 5028 660
rect 5077 663 5135 669
rect 2823 629 2835 632
rect 2777 623 2835 629
rect 5077 629 5089 663
rect 5123 660 5135 663
rect 5442 660 5448 672
rect 5123 632 5448 660
rect 5123 629 5135 632
rect 5077 623 5135 629
rect 5442 620 5448 632
rect 5500 620 5506 672
rect 9214 620 9220 672
rect 9272 660 9278 672
rect 9309 663 9367 669
rect 9309 660 9321 663
rect 9272 632 9321 660
rect 9272 620 9278 632
rect 9309 629 9321 632
rect 9355 629 9367 663
rect 9309 623 9367 629
rect 920 570 10396 592
rect 920 518 5066 570
rect 5118 518 5130 570
rect 5182 518 5194 570
rect 5246 518 5258 570
rect 5310 518 5322 570
rect 5374 518 10396 570
rect 920 496 10396 518
<< via1 >>
rect 1216 12180 1268 12232
rect 6092 12180 6144 12232
rect 2688 12044 2740 12096
rect 3608 12044 3660 12096
rect 2566 11942 2618 11994
rect 2630 11942 2682 11994
rect 2694 11942 2746 11994
rect 2758 11942 2810 11994
rect 2822 11942 2874 11994
rect 7566 11942 7618 11994
rect 7630 11942 7682 11994
rect 7694 11942 7746 11994
rect 7758 11942 7810 11994
rect 7822 11942 7874 11994
rect 6368 11840 6420 11892
rect 6460 11840 6512 11892
rect 7288 11840 7340 11892
rect 2688 11772 2740 11824
rect 3700 11772 3752 11824
rect 7012 11704 7064 11756
rect 8208 11747 8260 11756
rect 8208 11713 8217 11747
rect 8217 11713 8251 11747
rect 8251 11713 8260 11747
rect 8208 11704 8260 11713
rect 3608 11679 3660 11688
rect 3608 11645 3617 11679
rect 3617 11645 3651 11679
rect 3651 11645 3660 11679
rect 3608 11636 3660 11645
rect 3792 11679 3844 11688
rect 3792 11645 3801 11679
rect 3801 11645 3835 11679
rect 3835 11645 3844 11679
rect 3792 11636 3844 11645
rect 4068 11636 4120 11688
rect 4252 11679 4304 11688
rect 4252 11645 4261 11679
rect 4261 11645 4295 11679
rect 4295 11645 4304 11679
rect 4252 11636 4304 11645
rect 6092 11636 6144 11688
rect 6460 11636 6512 11688
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 6920 11636 6972 11688
rect 13820 11840 13872 11892
rect 17960 11840 18012 11892
rect 2504 11543 2556 11552
rect 2504 11509 2513 11543
rect 2513 11509 2547 11543
rect 2547 11509 2556 11543
rect 2504 11500 2556 11509
rect 4160 11500 4212 11552
rect 5448 11500 5500 11552
rect 7472 11568 7524 11620
rect 8484 11568 8536 11620
rect 6828 11500 6880 11552
rect 8852 11500 8904 11552
rect 5066 11398 5118 11450
rect 5130 11398 5182 11450
rect 5194 11398 5246 11450
rect 5258 11398 5310 11450
rect 5322 11398 5374 11450
rect 3884 11296 3936 11348
rect 3976 11296 4028 11348
rect 2688 11228 2740 11280
rect 3148 11228 3200 11280
rect 4344 11296 4396 11348
rect 6276 11228 6328 11280
rect 3700 11160 3752 11212
rect 4804 11160 4856 11212
rect 8392 11228 8444 11280
rect 2136 11092 2188 11144
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 3608 11092 3660 11144
rect 6368 11092 6420 11144
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 8944 11160 8996 11212
rect 8576 11092 8628 11144
rect 2688 10956 2740 11008
rect 3332 10956 3384 11008
rect 3516 10956 3568 11008
rect 3792 10956 3844 11008
rect 5632 11024 5684 11076
rect 9864 11024 9916 11076
rect 2566 10854 2618 10906
rect 2630 10854 2682 10906
rect 2694 10854 2746 10906
rect 2758 10854 2810 10906
rect 2822 10854 2874 10906
rect 7566 10854 7618 10906
rect 7630 10854 7682 10906
rect 7694 10854 7746 10906
rect 7758 10854 7810 10906
rect 7822 10854 7874 10906
rect 1308 10795 1360 10804
rect 1308 10761 1317 10795
rect 1317 10761 1351 10795
rect 1351 10761 1360 10795
rect 1308 10752 1360 10761
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 6920 10752 6972 10804
rect 7196 10752 7248 10804
rect 7380 10684 7432 10736
rect 7932 10752 7984 10804
rect 6736 10616 6788 10668
rect 8300 10684 8352 10736
rect 2780 10548 2832 10600
rect 3240 10548 3292 10600
rect 5908 10591 5960 10600
rect 5908 10557 5917 10591
rect 5917 10557 5951 10591
rect 5951 10557 5960 10591
rect 5908 10548 5960 10557
rect 6276 10591 6328 10600
rect 6276 10557 6285 10591
rect 6285 10557 6319 10591
rect 6319 10557 6328 10591
rect 6276 10548 6328 10557
rect 7472 10548 7524 10600
rect 9128 10548 9180 10600
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 2964 10412 3016 10464
rect 3056 10412 3108 10464
rect 5356 10480 5408 10532
rect 4712 10412 4764 10464
rect 8668 10412 8720 10464
rect 5066 10310 5118 10362
rect 5130 10310 5182 10362
rect 5194 10310 5246 10362
rect 5258 10310 5310 10362
rect 5322 10310 5374 10362
rect 6276 10208 6328 10260
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 2136 10004 2188 10056
rect 3516 10140 3568 10192
rect 5632 10140 5684 10192
rect 8116 10208 8168 10260
rect 8484 10140 8536 10192
rect 3700 10072 3752 10124
rect 7012 10115 7064 10124
rect 7012 10081 7021 10115
rect 7021 10081 7055 10115
rect 7055 10081 7064 10115
rect 7012 10072 7064 10081
rect 8668 10072 8720 10124
rect 3516 10047 3568 10056
rect 3516 10013 3525 10047
rect 3525 10013 3559 10047
rect 3559 10013 3568 10047
rect 3516 10004 3568 10013
rect 3884 10047 3936 10056
rect 2964 9936 3016 9988
rect 3884 10013 3893 10047
rect 3893 10013 3927 10047
rect 3927 10013 3936 10047
rect 3884 10004 3936 10013
rect 5540 10004 5592 10056
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 7104 10004 7156 10056
rect 9404 10004 9456 10056
rect 9772 10047 9824 10056
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 10232 10004 10284 10056
rect 3792 9868 3844 9920
rect 3884 9868 3936 9920
rect 7932 9868 7984 9920
rect 8760 9868 8812 9920
rect 2566 9766 2618 9818
rect 2630 9766 2682 9818
rect 2694 9766 2746 9818
rect 2758 9766 2810 9818
rect 2822 9766 2874 9818
rect 7566 9766 7618 9818
rect 7630 9766 7682 9818
rect 7694 9766 7746 9818
rect 7758 9766 7810 9818
rect 7822 9766 7874 9818
rect 3700 9664 3752 9716
rect 4988 9596 5040 9648
rect 7932 9596 7984 9648
rect 2412 9528 2464 9580
rect 5724 9528 5776 9580
rect 7288 9528 7340 9580
rect 7472 9528 7524 9580
rect 7564 9528 7616 9580
rect 2044 9460 2096 9512
rect 1308 9392 1360 9444
rect 3148 9435 3200 9444
rect 3148 9401 3157 9435
rect 3157 9401 3191 9435
rect 3191 9401 3200 9435
rect 3148 9392 3200 9401
rect 3240 9392 3292 9444
rect 2780 9324 2832 9376
rect 2964 9324 3016 9376
rect 5172 9460 5224 9512
rect 5816 9460 5868 9512
rect 8300 9528 8352 9580
rect 9496 9528 9548 9580
rect 9956 9571 10008 9580
rect 9956 9537 9965 9571
rect 9965 9537 9999 9571
rect 9999 9537 10008 9571
rect 9956 9528 10008 9537
rect 4528 9392 4580 9444
rect 6736 9392 6788 9444
rect 7104 9392 7156 9444
rect 7288 9392 7340 9444
rect 4068 9324 4120 9376
rect 5172 9324 5224 9376
rect 5632 9324 5684 9376
rect 6000 9324 6052 9376
rect 8852 9324 8904 9376
rect 9220 9460 9272 9512
rect 9128 9392 9180 9444
rect 10232 9324 10284 9376
rect 5066 9222 5118 9274
rect 5130 9222 5182 9274
rect 5194 9222 5246 9274
rect 5258 9222 5310 9274
rect 5322 9222 5374 9274
rect 3976 9120 4028 9172
rect 1308 9027 1360 9036
rect 1308 8993 1317 9027
rect 1317 8993 1351 9027
rect 1351 8993 1360 9027
rect 1308 8984 1360 8993
rect 3240 9052 3292 9104
rect 6276 9052 6328 9104
rect 7472 9052 7524 9104
rect 8024 9052 8076 9104
rect 1952 8959 2004 8968
rect 1952 8925 1961 8959
rect 1961 8925 1995 8959
rect 1995 8925 2004 8959
rect 1952 8916 2004 8925
rect 4068 8984 4120 9036
rect 4620 8984 4672 9036
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 6276 8916 6328 8968
rect 7288 8916 7340 8968
rect 4436 8848 4488 8900
rect 6092 8848 6144 8900
rect 6184 8848 6236 8900
rect 2320 8780 2372 8832
rect 3148 8780 3200 8832
rect 4252 8780 4304 8832
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 6736 8780 6788 8832
rect 8852 8848 8904 8900
rect 7380 8780 7432 8832
rect 7472 8780 7524 8832
rect 9772 8780 9824 8832
rect 2566 8678 2618 8730
rect 2630 8678 2682 8730
rect 2694 8678 2746 8730
rect 2758 8678 2810 8730
rect 2822 8678 2874 8730
rect 7566 8678 7618 8730
rect 7630 8678 7682 8730
rect 7694 8678 7746 8730
rect 7758 8678 7810 8730
rect 7822 8678 7874 8730
rect 3976 8576 4028 8628
rect 4528 8576 4580 8628
rect 5724 8576 5776 8628
rect 3148 8440 3200 8492
rect 3792 8508 3844 8560
rect 4436 8508 4488 8560
rect 8668 8576 8720 8628
rect 9680 8576 9732 8628
rect 8300 8508 8352 8560
rect 5448 8483 5500 8492
rect 2136 8372 2188 8424
rect 5448 8449 5457 8483
rect 5457 8449 5491 8483
rect 5491 8449 5500 8483
rect 5448 8440 5500 8449
rect 6000 8440 6052 8492
rect 6552 8440 6604 8492
rect 8852 8440 8904 8492
rect 10232 8508 10284 8560
rect 1308 8304 1360 8356
rect 1492 8304 1544 8356
rect 3792 8372 3844 8424
rect 6184 8415 6236 8424
rect 6184 8381 6193 8415
rect 6193 8381 6227 8415
rect 6227 8381 6236 8415
rect 6184 8372 6236 8381
rect 7932 8372 7984 8424
rect 8484 8372 8536 8424
rect 8760 8372 8812 8424
rect 4252 8304 4304 8356
rect 6552 8347 6604 8356
rect 3332 8236 3384 8288
rect 6552 8313 6561 8347
rect 6561 8313 6595 8347
rect 6595 8313 6604 8347
rect 6552 8304 6604 8313
rect 7564 8304 7616 8356
rect 9772 8372 9824 8424
rect 7840 8236 7892 8288
rect 8484 8279 8536 8288
rect 8484 8245 8493 8279
rect 8493 8245 8527 8279
rect 8527 8245 8536 8279
rect 8484 8236 8536 8245
rect 5066 8134 5118 8186
rect 5130 8134 5182 8186
rect 5194 8134 5246 8186
rect 5258 8134 5310 8186
rect 5322 8134 5374 8186
rect 2228 7964 2280 8016
rect 1768 7896 1820 7948
rect 3332 7939 3384 7948
rect 3332 7905 3341 7939
rect 3341 7905 3375 7939
rect 3375 7905 3384 7939
rect 3332 7896 3384 7905
rect 4620 7964 4672 8016
rect 6276 7964 6328 8016
rect 1124 7828 1176 7880
rect 2504 7803 2556 7812
rect 2504 7769 2513 7803
rect 2513 7769 2547 7803
rect 2547 7769 2556 7803
rect 2504 7760 2556 7769
rect 3148 7692 3200 7744
rect 4896 7896 4948 7948
rect 7472 7964 7524 8016
rect 7288 7939 7340 7948
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 7840 8032 7892 8084
rect 9680 7964 9732 8016
rect 9404 7939 9456 7948
rect 9404 7905 9413 7939
rect 9413 7905 9447 7939
rect 9447 7905 9456 7939
rect 9404 7896 9456 7905
rect 4252 7828 4304 7880
rect 5632 7828 5684 7880
rect 8300 7828 8352 7880
rect 6552 7760 6604 7812
rect 4804 7692 4856 7744
rect 6276 7692 6328 7744
rect 7288 7760 7340 7812
rect 8208 7692 8260 7744
rect 2566 7590 2618 7642
rect 2630 7590 2682 7642
rect 2694 7590 2746 7642
rect 2758 7590 2810 7642
rect 2822 7590 2874 7642
rect 7566 7590 7618 7642
rect 7630 7590 7682 7642
rect 7694 7590 7746 7642
rect 7758 7590 7810 7642
rect 7822 7590 7874 7642
rect 2688 7488 2740 7540
rect 4068 7488 4120 7540
rect 4160 7488 4212 7540
rect 3700 7420 3752 7472
rect 4712 7420 4764 7472
rect 6184 7463 6236 7472
rect 6184 7429 6185 7463
rect 6185 7429 6219 7463
rect 6219 7429 6236 7463
rect 6184 7420 6236 7429
rect 8576 7488 8628 7540
rect 1952 7352 2004 7404
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 5632 7352 5684 7404
rect 6000 7395 6052 7404
rect 6000 7361 6009 7395
rect 6009 7361 6043 7395
rect 6043 7361 6052 7395
rect 6000 7352 6052 7361
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 8484 7352 8536 7404
rect 2688 7216 2740 7268
rect 3240 7216 3292 7268
rect 4252 7284 4304 7336
rect 6736 7327 6788 7336
rect 6736 7293 6745 7327
rect 6745 7293 6779 7327
rect 6779 7293 6788 7327
rect 6736 7284 6788 7293
rect 9128 7284 9180 7336
rect 9680 7327 9732 7336
rect 9680 7293 9689 7327
rect 9689 7293 9723 7327
rect 9723 7293 9732 7327
rect 9680 7284 9732 7293
rect 5448 7216 5500 7268
rect 5632 7216 5684 7268
rect 7288 7216 7340 7268
rect 8576 7216 8628 7268
rect 17960 7148 18012 7200
rect 5066 7046 5118 7098
rect 5130 7046 5182 7098
rect 5194 7046 5246 7098
rect 5258 7046 5310 7098
rect 5322 7046 5374 7098
rect 1676 6944 1728 6996
rect 2044 6944 2096 6996
rect 3792 6944 3844 6996
rect 4344 6944 4396 6996
rect 5448 6944 5500 6996
rect 7564 6944 7616 6996
rect 8208 6944 8260 6996
rect 4896 6876 4948 6928
rect 8300 6876 8352 6928
rect 3148 6808 3200 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 2320 6740 2372 6792
rect 4804 6808 4856 6860
rect 1308 6647 1360 6656
rect 1308 6613 1317 6647
rect 1317 6613 1351 6647
rect 1351 6613 1360 6647
rect 1308 6604 1360 6613
rect 3516 6783 3568 6792
rect 3516 6749 3525 6783
rect 3525 6749 3559 6783
rect 3559 6749 3568 6783
rect 3516 6740 3568 6749
rect 3792 6740 3844 6792
rect 4528 6740 4580 6792
rect 3884 6604 3936 6656
rect 4528 6604 4580 6656
rect 8852 6851 8904 6860
rect 8852 6817 8861 6851
rect 8861 6817 8895 6851
rect 8895 6817 8904 6851
rect 8852 6808 8904 6817
rect 9312 6808 9364 6860
rect 9496 6851 9548 6860
rect 9496 6817 9505 6851
rect 9505 6817 9539 6851
rect 9539 6817 9548 6851
rect 9496 6808 9548 6817
rect 5724 6740 5776 6792
rect 6552 6740 6604 6792
rect 7380 6740 7432 6792
rect 6184 6604 6236 6656
rect 9128 6715 9180 6724
rect 9128 6681 9137 6715
rect 9137 6681 9171 6715
rect 9171 6681 9180 6715
rect 9128 6672 9180 6681
rect 9496 6672 9548 6724
rect 2566 6502 2618 6554
rect 2630 6502 2682 6554
rect 2694 6502 2746 6554
rect 2758 6502 2810 6554
rect 2822 6502 2874 6554
rect 7566 6502 7618 6554
rect 7630 6502 7682 6554
rect 7694 6502 7746 6554
rect 7758 6502 7810 6554
rect 7822 6502 7874 6554
rect 1216 6443 1268 6452
rect 1216 6409 1225 6443
rect 1225 6409 1259 6443
rect 1259 6409 1268 6443
rect 1216 6400 1268 6409
rect 2872 6400 2924 6452
rect 3148 6400 3200 6452
rect 3516 6332 3568 6384
rect 1308 6264 1360 6316
rect 2780 6264 2832 6316
rect 6920 6400 6972 6452
rect 7472 6400 7524 6452
rect 8024 6400 8076 6452
rect 9220 6400 9272 6452
rect 4896 6375 4948 6384
rect 4896 6341 4905 6375
rect 4905 6341 4939 6375
rect 4939 6341 4948 6375
rect 4896 6332 4948 6341
rect 8116 6332 8168 6384
rect 1492 6196 1544 6248
rect 3056 6196 3108 6248
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 4252 6264 4304 6316
rect 5632 6307 5684 6316
rect 5632 6273 5641 6307
rect 5641 6273 5675 6307
rect 5675 6273 5684 6307
rect 5632 6264 5684 6273
rect 7380 6264 7432 6316
rect 8668 6264 8720 6316
rect 9680 6264 9732 6316
rect 3516 6196 3568 6248
rect 1676 6128 1728 6180
rect 1768 6128 1820 6180
rect 4160 6196 4212 6248
rect 4712 6196 4764 6248
rect 4988 6196 5040 6248
rect 6552 6196 6604 6248
rect 8944 6239 8996 6248
rect 8944 6205 8953 6239
rect 8953 6205 8987 6239
rect 8987 6205 8996 6239
rect 8944 6196 8996 6205
rect 9864 6239 9916 6248
rect 9864 6205 9873 6239
rect 9873 6205 9907 6239
rect 9907 6205 9916 6239
rect 9864 6196 9916 6205
rect 4436 6128 4488 6180
rect 6920 6128 6972 6180
rect 3792 6060 3844 6112
rect 3976 6060 4028 6112
rect 4160 6060 4212 6112
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 8024 6060 8076 6112
rect 8760 6060 8812 6112
rect 9772 6060 9824 6112
rect 5066 5958 5118 6010
rect 5130 5958 5182 6010
rect 5194 5958 5246 6010
rect 5258 5958 5310 6010
rect 5322 5958 5374 6010
rect 3148 5856 3200 5908
rect 3976 5856 4028 5908
rect 4896 5856 4948 5908
rect 11060 5856 11112 5908
rect 1400 5788 1452 5840
rect 1308 5720 1360 5772
rect 4160 5788 4212 5840
rect 4528 5788 4580 5840
rect 4988 5788 5040 5840
rect 6552 5831 6604 5840
rect 6552 5797 6561 5831
rect 6561 5797 6595 5831
rect 6595 5797 6604 5831
rect 6552 5788 6604 5797
rect 8208 5788 8260 5840
rect 3884 5763 3936 5772
rect 3884 5729 3893 5763
rect 3893 5729 3927 5763
rect 3927 5729 3936 5763
rect 3884 5720 3936 5729
rect 5816 5720 5868 5772
rect 3240 5652 3292 5704
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 4804 5652 4856 5704
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 6092 5652 6144 5704
rect 9128 5720 9180 5772
rect 9312 5788 9364 5840
rect 6552 5652 6604 5704
rect 8116 5652 8168 5704
rect 8760 5652 8812 5704
rect 6828 5584 6880 5636
rect 2872 5516 2924 5568
rect 3884 5516 3936 5568
rect 4988 5516 5040 5568
rect 8484 5516 8536 5568
rect 9128 5516 9180 5568
rect 9312 5652 9364 5704
rect 10048 5720 10100 5772
rect 9680 5652 9732 5704
rect 9312 5516 9364 5568
rect 16580 5516 16632 5568
rect 2566 5414 2618 5466
rect 2630 5414 2682 5466
rect 2694 5414 2746 5466
rect 2758 5414 2810 5466
rect 2822 5414 2874 5466
rect 7566 5414 7618 5466
rect 7630 5414 7682 5466
rect 7694 5414 7746 5466
rect 7758 5414 7810 5466
rect 7822 5414 7874 5466
rect 1676 5312 1728 5364
rect 2780 5312 2832 5364
rect 3700 5355 3752 5364
rect 3700 5321 3709 5355
rect 3709 5321 3743 5355
rect 3743 5321 3752 5355
rect 3700 5312 3752 5321
rect 5632 5312 5684 5364
rect 7012 5312 7064 5364
rect 7656 5312 7708 5364
rect 8116 5312 8168 5364
rect 9312 5312 9364 5364
rect 5816 5244 5868 5296
rect 6460 5244 6512 5296
rect 8300 5244 8352 5296
rect 2964 5176 3016 5228
rect 3884 5176 3936 5228
rect 4436 5176 4488 5228
rect 7932 5176 7984 5228
rect 10324 5176 10376 5228
rect 2872 5108 2924 5160
rect 3792 5151 3844 5160
rect 3792 5117 3801 5151
rect 3801 5117 3835 5151
rect 3835 5117 3844 5151
rect 3792 5108 3844 5117
rect 6000 5108 6052 5160
rect 6460 5151 6512 5160
rect 6460 5117 6469 5151
rect 6469 5117 6503 5151
rect 6503 5117 6512 5151
rect 6460 5108 6512 5117
rect 6552 5108 6604 5160
rect 7012 5151 7064 5160
rect 7012 5117 7021 5151
rect 7021 5117 7055 5151
rect 7055 5117 7064 5151
rect 7012 5108 7064 5117
rect 7472 5108 7524 5160
rect 6092 5040 6144 5092
rect 8484 5040 8536 5092
rect 9772 5040 9824 5092
rect 10140 5040 10192 5092
rect 9036 5015 9088 5024
rect 9036 4981 9045 5015
rect 9045 4981 9079 5015
rect 9079 4981 9088 5015
rect 9036 4972 9088 4981
rect 5066 4870 5118 4922
rect 5130 4870 5182 4922
rect 5194 4870 5246 4922
rect 5258 4870 5310 4922
rect 5322 4870 5374 4922
rect 3976 4768 4028 4820
rect 4804 4700 4856 4752
rect 2964 4632 3016 4684
rect 3240 4632 3292 4684
rect 3884 4675 3936 4684
rect 3884 4641 3893 4675
rect 3893 4641 3927 4675
rect 3927 4641 3936 4675
rect 3884 4632 3936 4641
rect 4528 4632 4580 4684
rect 6092 4632 6144 4684
rect 4160 4564 4212 4616
rect 7012 4768 7064 4820
rect 9588 4811 9640 4820
rect 9588 4777 9597 4811
rect 9597 4777 9631 4811
rect 9631 4777 9640 4811
rect 9588 4768 9640 4777
rect 6552 4632 6604 4684
rect 6828 4632 6880 4684
rect 7932 4700 7984 4752
rect 7656 4675 7708 4684
rect 7656 4641 7665 4675
rect 7665 4641 7699 4675
rect 7699 4641 7708 4675
rect 7656 4632 7708 4641
rect 6000 4496 6052 4548
rect 6644 4496 6696 4548
rect 6920 4539 6972 4548
rect 6920 4505 6929 4539
rect 6929 4505 6963 4539
rect 6963 4505 6972 4539
rect 6920 4496 6972 4505
rect 7288 4496 7340 4548
rect 8392 4564 8444 4616
rect 4620 4428 4672 4480
rect 6092 4428 6144 4480
rect 7566 4326 7618 4378
rect 7630 4326 7682 4378
rect 7694 4326 7746 4378
rect 7758 4326 7810 4378
rect 7822 4326 7874 4378
rect 3792 4088 3844 4140
rect 4896 4088 4948 4140
rect 9404 4131 9456 4140
rect 4344 4020 4396 4072
rect 5356 4063 5408 4072
rect 4896 3952 4948 4004
rect 5356 4029 5365 4063
rect 5365 4029 5399 4063
rect 5399 4029 5408 4063
rect 5356 4020 5408 4029
rect 5540 4063 5592 4072
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 5632 4020 5684 4072
rect 5816 4020 5868 4072
rect 6276 4063 6328 4072
rect 6276 4029 6285 4063
rect 6285 4029 6319 4063
rect 6319 4029 6328 4063
rect 6276 4020 6328 4029
rect 5448 3952 5500 4004
rect 6000 3884 6052 3936
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 9404 4088 9456 4097
rect 8576 4020 8628 4072
rect 16580 3952 16632 4004
rect 22100 3884 22152 3936
rect 5066 3782 5118 3834
rect 5130 3782 5182 3834
rect 5194 3782 5246 3834
rect 5258 3782 5310 3834
rect 5322 3782 5374 3834
rect 6644 3680 6696 3732
rect 9496 3680 9548 3732
rect 3884 3612 3936 3664
rect 9036 3612 9088 3664
rect 4068 3544 4120 3596
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 9588 3544 9640 3596
rect 9772 3587 9824 3596
rect 9772 3553 9781 3587
rect 9781 3553 9815 3587
rect 9815 3553 9824 3587
rect 9772 3544 9824 3553
rect 4804 3476 4856 3528
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 2688 3408 2740 3460
rect 16672 3476 16724 3528
rect 4988 3340 5040 3392
rect 9220 3340 9272 3392
rect 9496 3340 9548 3392
rect 7566 3238 7618 3290
rect 7630 3238 7682 3290
rect 7694 3238 7746 3290
rect 7758 3238 7810 3290
rect 7822 3238 7874 3290
rect 3608 3136 3660 3188
rect 6000 3179 6052 3188
rect 6000 3145 6009 3179
rect 6009 3145 6043 3179
rect 6043 3145 6052 3179
rect 6000 3136 6052 3145
rect 6736 3136 6788 3188
rect 4344 3068 4396 3120
rect 4988 3068 5040 3120
rect 7288 3068 7340 3120
rect 9220 3068 9272 3120
rect 4068 3000 4120 3052
rect 6460 3000 6512 3052
rect 6828 3043 6880 3052
rect 6828 3009 6837 3043
rect 6837 3009 6871 3043
rect 6871 3009 6880 3043
rect 6828 3000 6880 3009
rect 7196 3000 7248 3052
rect 2872 2932 2924 2984
rect 4988 2932 5040 2984
rect 8668 2864 8720 2916
rect 16856 2864 16908 2916
rect 5066 2694 5118 2746
rect 5130 2694 5182 2746
rect 5194 2694 5246 2746
rect 5258 2694 5310 2746
rect 5322 2694 5374 2746
rect 2780 2592 2832 2644
rect 4252 2592 4304 2644
rect 4436 2592 4488 2644
rect 4988 2592 5040 2644
rect 6000 2635 6052 2644
rect 6000 2601 6009 2635
rect 6009 2601 6043 2635
rect 6043 2601 6052 2635
rect 6000 2592 6052 2601
rect 7288 2592 7340 2644
rect 3608 2499 3660 2508
rect 3608 2465 3617 2499
rect 3617 2465 3651 2499
rect 3651 2465 3660 2499
rect 3608 2456 3660 2465
rect 3792 2456 3844 2508
rect 4160 2456 4212 2508
rect 3332 2388 3384 2440
rect 3976 2320 4028 2372
rect 4896 2456 4948 2508
rect 8300 2456 8352 2508
rect 8392 2456 8444 2508
rect 5632 2295 5684 2304
rect 5632 2261 5641 2295
rect 5641 2261 5675 2295
rect 5675 2261 5684 2295
rect 5632 2252 5684 2261
rect 5816 2252 5868 2304
rect 6092 2252 6144 2304
rect 9588 2592 9640 2644
rect 10048 2592 10100 2644
rect 8852 2524 8904 2576
rect 8760 2499 8812 2508
rect 8760 2465 8769 2499
rect 8769 2465 8803 2499
rect 8803 2465 8812 2499
rect 8760 2456 8812 2465
rect 8116 2320 8168 2372
rect 9036 2388 9088 2440
rect 9220 2388 9272 2440
rect 10048 2499 10100 2508
rect 10048 2465 10057 2499
rect 10057 2465 10091 2499
rect 10091 2465 10100 2499
rect 10048 2456 10100 2465
rect 16948 2456 17000 2508
rect 9772 2388 9824 2440
rect 9772 2252 9824 2304
rect 10140 2252 10192 2304
rect 7566 2150 7618 2202
rect 7630 2150 7682 2202
rect 7694 2150 7746 2202
rect 7758 2150 7810 2202
rect 7822 2150 7874 2202
rect 3240 2048 3292 2100
rect 3516 2091 3568 2100
rect 3516 2057 3525 2091
rect 3525 2057 3559 2091
rect 3559 2057 3568 2091
rect 3516 2048 3568 2057
rect 3884 2048 3936 2100
rect 4068 2048 4120 2100
rect 4620 2048 4672 2100
rect 10048 2048 10100 2100
rect 3056 1980 3108 2032
rect 8116 1980 8168 2032
rect 16580 1980 16632 2032
rect 6828 1955 6880 1964
rect 6828 1921 6837 1955
rect 6837 1921 6871 1955
rect 6871 1921 6880 1955
rect 6828 1912 6880 1921
rect 3608 1844 3660 1896
rect 22284 1912 22336 1964
rect 8024 1887 8076 1896
rect 8024 1853 8033 1887
rect 8033 1853 8067 1887
rect 8067 1853 8076 1887
rect 8024 1844 8076 1853
rect 9864 1887 9916 1896
rect 8576 1776 8628 1828
rect 9312 1776 9364 1828
rect 9864 1853 9873 1887
rect 9873 1853 9907 1887
rect 9907 1853 9916 1887
rect 9864 1844 9916 1853
rect 16764 1776 16816 1828
rect 10048 1708 10100 1760
rect 5066 1606 5118 1658
rect 5130 1606 5182 1658
rect 5194 1606 5246 1658
rect 5258 1606 5310 1658
rect 5322 1606 5374 1658
rect 3240 1504 3292 1556
rect 5540 1504 5592 1556
rect 8116 1547 8168 1556
rect 8116 1513 8125 1547
rect 8125 1513 8159 1547
rect 8159 1513 8168 1547
rect 8116 1504 8168 1513
rect 8944 1504 8996 1556
rect 9128 1504 9180 1556
rect 9220 1436 9272 1488
rect 6184 1411 6236 1420
rect 6184 1377 6193 1411
rect 6193 1377 6227 1411
rect 6227 1377 6236 1411
rect 6184 1368 6236 1377
rect 8852 1411 8904 1420
rect 8852 1377 8861 1411
rect 8861 1377 8895 1411
rect 8895 1377 8904 1411
rect 8852 1368 8904 1377
rect 9588 1368 9640 1420
rect 5448 1343 5500 1352
rect 5448 1309 5457 1343
rect 5457 1309 5491 1343
rect 5491 1309 5500 1343
rect 5448 1300 5500 1309
rect 6092 1300 6144 1352
rect 9312 1300 9364 1352
rect 10324 1368 10376 1420
rect 2320 1164 2372 1216
rect 8760 1232 8812 1284
rect 5632 1164 5684 1216
rect 8576 1164 8628 1216
rect 10232 1232 10284 1284
rect 9312 1207 9364 1216
rect 9312 1173 9321 1207
rect 9321 1173 9355 1207
rect 9355 1173 9364 1207
rect 9312 1164 9364 1173
rect 2566 1062 2618 1114
rect 2630 1062 2682 1114
rect 2694 1062 2746 1114
rect 2758 1062 2810 1114
rect 2822 1062 2874 1114
rect 7566 1062 7618 1114
rect 7630 1062 7682 1114
rect 7694 1062 7746 1114
rect 7758 1062 7810 1114
rect 7822 1062 7874 1114
rect 1124 960 1176 1012
rect 2412 960 2464 1012
rect 2964 1003 3016 1012
rect 2964 969 2973 1003
rect 2973 969 3007 1003
rect 3007 969 3016 1003
rect 2964 960 3016 969
rect 4988 960 5040 1012
rect 8760 1003 8812 1012
rect 8760 969 8769 1003
rect 8769 969 8803 1003
rect 8803 969 8812 1003
rect 8760 960 8812 969
rect 9036 1003 9088 1012
rect 9036 969 9045 1003
rect 9045 969 9079 1003
rect 9079 969 9088 1003
rect 9036 960 9088 969
rect 9680 1003 9732 1012
rect 9680 969 9689 1003
rect 9689 969 9723 1003
rect 9723 969 9732 1003
rect 9680 960 9732 969
rect 9956 960 10008 1012
rect 3424 892 3476 944
rect 13820 892 13872 944
rect 5908 824 5960 876
rect 2964 756 3016 808
rect 9772 824 9824 876
rect 9312 756 9364 808
rect 10048 799 10100 808
rect 10048 765 10057 799
rect 10057 765 10091 799
rect 10091 765 10100 799
rect 10048 756 10100 765
rect 3056 688 3108 740
rect 2320 620 2372 672
rect 5632 688 5684 740
rect 8852 688 8904 740
rect 5448 620 5500 672
rect 9220 620 9272 672
rect 5066 518 5118 570
rect 5130 518 5182 570
rect 5194 518 5246 570
rect 5258 518 5310 570
rect 5322 518 5374 570
<< obsm1 >>
rect 24000 0 34000 13000
<< metal2 >>
rect 938 12322 994 13000
rect 938 12294 1256 12322
rect 938 12200 994 12294
rect 1228 12238 1256 12294
rect 1216 12232 1268 12238
rect 1398 12200 1454 13000
rect 1858 12322 1914 13000
rect 1504 12294 1914 12322
rect 1216 12174 1268 12180
rect 1412 11121 1440 12200
rect 1398 11112 1454 11121
rect 1398 11047 1454 11056
rect 1308 10804 1360 10810
rect 1412 10792 1440 11047
rect 1360 10764 1440 10792
rect 1308 10746 1360 10752
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 10130 1440 10610
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1308 9444 1360 9450
rect 1308 9386 1360 9392
rect 1214 9344 1270 9353
rect 1214 9279 1270 9288
rect 1124 7880 1176 7886
rect 1124 7822 1176 7828
rect 1136 1018 1164 7822
rect 1228 6458 1256 9279
rect 1320 9042 1348 9386
rect 1308 9036 1360 9042
rect 1308 8978 1360 8984
rect 1504 8362 1532 12294
rect 1858 12200 1914 12294
rect 2318 12322 2374 13000
rect 2778 12322 2834 13000
rect 3238 12322 3294 13000
rect 3698 12322 3754 13000
rect 2318 12294 2728 12322
rect 2318 12200 2374 12294
rect 2700 12102 2728 12294
rect 2778 12294 3004 12322
rect 2778 12200 2834 12294
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2566 11996 2874 12005
rect 2566 11994 2572 11996
rect 2628 11994 2652 11996
rect 2708 11994 2732 11996
rect 2788 11994 2812 11996
rect 2868 11994 2874 11996
rect 2628 11942 2630 11994
rect 2810 11942 2812 11994
rect 2566 11940 2572 11942
rect 2628 11940 2652 11942
rect 2708 11940 2732 11942
rect 2788 11940 2812 11942
rect 2868 11940 2874 11942
rect 2566 11931 2874 11940
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2502 11656 2558 11665
rect 2502 11591 2558 11600
rect 2516 11558 2544 11591
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2700 11286 2728 11766
rect 2688 11280 2740 11286
rect 2688 11222 2740 11228
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2148 10554 2176 11086
rect 2700 11014 2728 11222
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2566 10908 2874 10917
rect 2566 10906 2572 10908
rect 2628 10906 2652 10908
rect 2708 10906 2732 10908
rect 2788 10906 2812 10908
rect 2868 10906 2874 10908
rect 2628 10854 2630 10906
rect 2810 10854 2812 10906
rect 2566 10852 2572 10854
rect 2628 10852 2652 10854
rect 2708 10852 2732 10854
rect 2788 10852 2812 10854
rect 2868 10852 2874 10854
rect 2566 10843 2874 10852
rect 2778 10704 2834 10713
rect 2778 10639 2834 10648
rect 2792 10606 2820 10639
rect 2780 10600 2832 10606
rect 2148 10526 2268 10554
rect 2976 10554 3004 12294
rect 3068 12294 3294 12322
rect 3068 10577 3096 12294
rect 3238 12200 3294 12294
rect 3344 12294 3754 12322
rect 3148 11280 3200 11286
rect 3148 11222 3200 11228
rect 2780 10542 2832 10548
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2044 9512 2096 9518
rect 2148 9500 2176 9998
rect 2096 9472 2176 9500
rect 2044 9454 2096 9460
rect 1952 8968 2004 8974
rect 1952 8910 2004 8916
rect 1308 8356 1360 8362
rect 1308 8298 1360 8304
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1320 8265 1348 8298
rect 1306 8256 1362 8265
rect 1306 8191 1362 8200
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1308 6656 1360 6662
rect 1308 6598 1360 6604
rect 1216 6452 1268 6458
rect 1216 6394 1268 6400
rect 1320 6322 1348 6598
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1320 5778 1348 6258
rect 1412 5846 1440 6734
rect 1504 6254 1532 8298
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1492 6248 1544 6254
rect 1492 6190 1544 6196
rect 1688 6186 1716 6938
rect 1780 6186 1808 7890
rect 1964 7410 1992 8910
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 2056 7002 2084 9454
rect 2134 8528 2190 8537
rect 2134 8463 2190 8472
rect 2148 8430 2176 8463
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1768 6180 1820 6186
rect 1768 6122 1820 6128
rect 1400 5840 1452 5846
rect 1400 5782 1452 5788
rect 1308 5772 1360 5778
rect 1308 5714 1360 5720
rect 1688 5370 1716 6122
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 2148 4536 2176 8366
rect 2240 8022 2268 10526
rect 2884 10526 3004 10554
rect 3054 10568 3110 10577
rect 2884 10033 2912 10526
rect 3054 10503 3110 10512
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2870 10024 2926 10033
rect 2976 9994 3004 10406
rect 2870 9959 2926 9968
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2962 9888 3018 9897
rect 2566 9820 2874 9829
rect 2962 9823 3018 9832
rect 2566 9818 2572 9820
rect 2628 9818 2652 9820
rect 2708 9818 2732 9820
rect 2788 9818 2812 9820
rect 2868 9818 2874 9820
rect 2628 9766 2630 9818
rect 2810 9766 2812 9818
rect 2566 9764 2572 9766
rect 2628 9764 2652 9766
rect 2708 9764 2732 9766
rect 2788 9764 2812 9766
rect 2868 9764 2874 9766
rect 2566 9755 2874 9764
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2228 8016 2280 8022
rect 2228 7958 2280 7964
rect 2332 6798 2360 8774
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2148 4508 2360 4536
rect 2332 1222 2360 4508
rect 2320 1216 2372 1222
rect 2320 1158 2372 1164
rect 1124 1012 1176 1018
rect 1124 954 1176 960
rect 2332 678 2360 1158
rect 2424 1018 2452 9522
rect 2778 9480 2834 9489
rect 2976 9466 3004 9823
rect 2778 9415 2834 9424
rect 2884 9438 3004 9466
rect 2792 9382 2820 9415
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2884 8820 2912 9438
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 8974 3004 9318
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2884 8792 3004 8820
rect 2566 8732 2874 8741
rect 2566 8730 2572 8732
rect 2628 8730 2652 8732
rect 2708 8730 2732 8732
rect 2788 8730 2812 8732
rect 2868 8730 2874 8732
rect 2628 8678 2630 8730
rect 2810 8678 2812 8730
rect 2566 8676 2572 8678
rect 2628 8676 2652 8678
rect 2708 8676 2732 8678
rect 2788 8676 2812 8678
rect 2868 8676 2874 8678
rect 2566 8667 2874 8676
rect 2502 7848 2558 7857
rect 2502 7783 2504 7792
rect 2556 7783 2558 7792
rect 2504 7754 2556 7760
rect 2566 7644 2874 7653
rect 2566 7642 2572 7644
rect 2628 7642 2652 7644
rect 2708 7642 2732 7644
rect 2788 7642 2812 7644
rect 2868 7642 2874 7644
rect 2628 7590 2630 7642
rect 2810 7590 2812 7642
rect 2566 7588 2572 7590
rect 2628 7588 2652 7590
rect 2708 7588 2732 7590
rect 2788 7588 2812 7590
rect 2868 7588 2874 7590
rect 2566 7579 2874 7588
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2700 7274 2728 7482
rect 2688 7268 2740 7274
rect 2688 7210 2740 7216
rect 2566 6556 2874 6565
rect 2566 6554 2572 6556
rect 2628 6554 2652 6556
rect 2708 6554 2732 6556
rect 2788 6554 2812 6556
rect 2868 6554 2874 6556
rect 2628 6502 2630 6554
rect 2810 6502 2812 6554
rect 2566 6500 2572 6502
rect 2628 6500 2652 6502
rect 2708 6500 2732 6502
rect 2788 6500 2812 6502
rect 2868 6500 2874 6502
rect 2566 6491 2874 6500
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2778 6352 2834 6361
rect 2778 6287 2780 6296
rect 2832 6287 2834 6296
rect 2780 6258 2832 6264
rect 2884 5574 2912 6394
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2566 5468 2874 5477
rect 2566 5466 2572 5468
rect 2628 5466 2652 5468
rect 2708 5466 2732 5468
rect 2788 5466 2812 5468
rect 2868 5466 2874 5468
rect 2628 5414 2630 5466
rect 2810 5414 2812 5466
rect 2566 5412 2572 5414
rect 2628 5412 2652 5414
rect 2708 5412 2732 5414
rect 2788 5412 2812 5414
rect 2868 5412 2874 5414
rect 2566 5403 2874 5412
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2688 3460 2740 3466
rect 2686 3428 2688 3437
rect 2740 3428 2742 3437
rect 2686 3363 2742 3372
rect 2792 2650 2820 5306
rect 2976 5234 3004 8792
rect 3068 6338 3096 10406
rect 3160 9450 3188 11222
rect 3344 11098 3372 12294
rect 3698 12200 3754 12294
rect 4158 12458 4214 13000
rect 4158 12430 4476 12458
rect 4158 12200 4214 12430
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11694 3648 12038
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3620 11257 3648 11630
rect 3606 11248 3662 11257
rect 3712 11218 3740 11766
rect 3896 11750 4292 11778
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3606 11183 3662 11192
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3252 11070 3372 11098
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3252 10690 3280 11070
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3344 10849 3372 10950
rect 3330 10840 3386 10849
rect 3330 10775 3386 10784
rect 3252 10662 3372 10690
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3252 9450 3280 10542
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3252 9110 3280 9386
rect 3240 9104 3292 9110
rect 3240 9046 3292 9052
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3160 8498 3188 8774
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3148 7744 3200 7750
rect 3148 7686 3200 7692
rect 3160 7410 3188 7686
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3252 7274 3280 9046
rect 3344 8401 3372 10662
rect 3330 8392 3386 8401
rect 3330 8327 3386 8336
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3344 7954 3372 8230
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3160 6458 3188 6802
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3068 6310 3188 6338
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 2964 5228 3016 5234
rect 2964 5170 3016 5176
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2884 2990 2912 5102
rect 2976 4690 3004 5170
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 3068 2038 3096 6190
rect 3160 5914 3188 6310
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3252 5710 3280 7210
rect 3436 7018 3464 11086
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3528 10198 3556 10950
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3344 6990 3464 7018
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3252 2106 3280 4626
rect 3344 2446 3372 6990
rect 3528 6882 3556 9998
rect 3436 6854 3556 6882
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 3240 2100 3292 2106
rect 3240 2042 3292 2048
rect 3056 2032 3108 2038
rect 3056 1974 3108 1980
rect 2566 1116 2874 1125
rect 2566 1114 2572 1116
rect 2628 1114 2652 1116
rect 2708 1114 2732 1116
rect 2788 1114 2812 1116
rect 2868 1114 2874 1116
rect 2628 1062 2630 1114
rect 2810 1062 2812 1114
rect 2566 1060 2572 1062
rect 2628 1060 2652 1062
rect 2708 1060 2732 1062
rect 2788 1060 2812 1062
rect 2868 1060 2874 1062
rect 2566 1051 2874 1060
rect 2412 1012 2464 1018
rect 2412 954 2464 960
rect 2964 1012 3016 1018
rect 2964 954 3016 960
rect 2976 814 3004 954
rect 2964 808 3016 814
rect 2964 750 3016 756
rect 3068 746 3096 1974
rect 3252 1562 3280 2042
rect 3240 1556 3292 1562
rect 3240 1498 3292 1504
rect 3436 950 3464 6854
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3528 6390 3556 6734
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3528 2106 3556 6190
rect 3620 3194 3648 11086
rect 3804 11014 3832 11630
rect 3896 11354 3924 11750
rect 4264 11694 4292 11750
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3712 9722 3740 10066
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3896 9926 3924 9998
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3804 9081 3832 9862
rect 3988 9674 4016 11290
rect 3896 9646 4016 9674
rect 3790 9072 3846 9081
rect 3790 9007 3846 9016
rect 3804 8566 3832 9007
rect 3896 8673 3924 9646
rect 4080 9382 4108 11630
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3882 8664 3938 8673
rect 3988 8634 4016 9114
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 3882 8599 3938 8608
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3882 8392 3938 8401
rect 3700 7472 3752 7478
rect 3700 7414 3752 7420
rect 3712 5370 3740 7414
rect 3804 7002 3832 8366
rect 3882 8327 3938 8336
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3804 6798 3832 6938
rect 3792 6792 3844 6798
rect 3896 6769 3924 8327
rect 3792 6734 3844 6740
rect 3882 6760 3938 6769
rect 3882 6695 3938 6704
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3896 6322 3924 6598
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3988 6118 4016 8570
rect 4080 7546 4108 8978
rect 4172 7546 4200 11494
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4356 11121 4384 11290
rect 4342 11112 4398 11121
rect 4342 11047 4398 11056
rect 4250 8936 4306 8945
rect 4250 8871 4306 8880
rect 4264 8838 4292 8871
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4250 8664 4306 8673
rect 4250 8599 4306 8608
rect 4264 8362 4292 8599
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4080 7313 4108 7482
rect 4066 7304 4122 7313
rect 4066 7239 4122 7248
rect 4066 6760 4122 6769
rect 4066 6695 4122 6704
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3804 5166 3832 6054
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3988 5794 4016 5850
rect 3896 5778 4016 5794
rect 3884 5772 4016 5778
rect 3936 5766 4016 5772
rect 3884 5714 3936 5720
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3896 5234 3924 5510
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3896 4690 3924 5170
rect 3988 4826 4016 5646
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3804 3516 3832 4082
rect 3896 3670 3924 4626
rect 3884 3664 3936 3670
rect 3884 3606 3936 3612
rect 3804 3488 3924 3516
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3790 2544 3846 2553
rect 3608 2508 3660 2514
rect 3790 2479 3792 2488
rect 3608 2450 3660 2456
rect 3844 2479 3846 2488
rect 3792 2450 3844 2456
rect 3516 2100 3568 2106
rect 3516 2042 3568 2048
rect 3620 1902 3648 2450
rect 3896 2106 3924 3488
rect 3988 2378 4016 4762
rect 4080 3602 4108 6695
rect 4172 6474 4200 7482
rect 4264 7342 4292 7822
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4264 6905 4292 7278
rect 4356 7002 4384 11047
rect 4448 8906 4476 12430
rect 4618 12322 4674 13000
rect 4618 12294 4752 12322
rect 4618 12200 4674 12294
rect 4724 10470 4752 12294
rect 5078 12200 5134 13000
rect 5538 12322 5594 13000
rect 5538 12294 5856 12322
rect 5538 12200 5594 12294
rect 5092 11540 5120 12200
rect 4908 11512 5120 11540
rect 5448 11552 5500 11558
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4540 8634 4568 9386
rect 4724 9058 4752 10406
rect 4816 9353 4844 11154
rect 4908 9489 4936 11512
rect 5448 11494 5500 11500
rect 5066 11452 5374 11461
rect 5066 11450 5072 11452
rect 5128 11450 5152 11452
rect 5208 11450 5232 11452
rect 5288 11450 5312 11452
rect 5368 11450 5374 11452
rect 5128 11398 5130 11450
rect 5310 11398 5312 11450
rect 5066 11396 5072 11398
rect 5128 11396 5152 11398
rect 5208 11396 5232 11398
rect 5288 11396 5312 11398
rect 5368 11396 5374 11398
rect 5066 11387 5374 11396
rect 5354 10568 5410 10577
rect 5354 10503 5356 10512
rect 5408 10503 5410 10512
rect 5356 10474 5408 10480
rect 5066 10364 5374 10373
rect 5066 10362 5072 10364
rect 5128 10362 5152 10364
rect 5208 10362 5232 10364
rect 5288 10362 5312 10364
rect 5368 10362 5374 10364
rect 5128 10310 5130 10362
rect 5310 10310 5312 10362
rect 5066 10308 5072 10310
rect 5128 10308 5152 10310
rect 5208 10308 5232 10310
rect 5288 10308 5312 10310
rect 5368 10308 5374 10310
rect 5066 10299 5374 10308
rect 5460 10305 5488 11494
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5538 10568 5594 10577
rect 5538 10503 5594 10512
rect 5446 10296 5502 10305
rect 5446 10231 5502 10240
rect 5552 10180 5580 10503
rect 5644 10198 5672 11018
rect 5368 10152 5580 10180
rect 5632 10192 5684 10198
rect 4988 9648 5040 9654
rect 5368 9625 5396 10152
rect 5632 10134 5684 10140
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 4988 9590 5040 9596
rect 5354 9616 5410 9625
rect 4894 9480 4950 9489
rect 4894 9415 4950 9424
rect 4802 9344 4858 9353
rect 4802 9279 4858 9288
rect 4632 9042 4752 9058
rect 4620 9036 4752 9042
rect 4672 9030 4752 9036
rect 4620 8978 4672 8984
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4448 8265 4476 8502
rect 4434 8256 4490 8265
rect 4434 8191 4490 8200
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4344 6996 4396 7002
rect 4344 6938 4396 6944
rect 4250 6896 4306 6905
rect 4250 6831 4306 6840
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 6662 4568 6734
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4172 6446 4384 6474
rect 4158 6352 4214 6361
rect 4158 6287 4214 6296
rect 4252 6316 4304 6322
rect 4172 6254 4200 6287
rect 4252 6258 4304 6264
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4172 5846 4200 6054
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4068 3596 4120 3602
rect 4068 3538 4120 3544
rect 4080 3058 4108 3538
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 4080 2106 4108 2994
rect 4172 2514 4200 4558
rect 4264 2650 4292 6258
rect 4356 4078 4384 6446
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4448 5234 4476 6122
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4540 5846 4568 6054
rect 4528 5840 4580 5846
rect 4528 5782 4580 5788
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4356 3126 4384 4014
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4448 2650 4476 5170
rect 4540 4690 4568 5782
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4632 4486 4660 7958
rect 4816 7750 4844 8774
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4908 7562 4936 7890
rect 4724 7534 4936 7562
rect 4724 7478 4752 7534
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4724 2774 4752 6190
rect 4816 5710 4844 6802
rect 4908 6390 4936 6870
rect 4896 6384 4948 6390
rect 4896 6326 4948 6332
rect 5000 6254 5028 9590
rect 5354 9551 5410 9560
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5184 9382 5212 9454
rect 5172 9376 5224 9382
rect 5172 9318 5224 9324
rect 5066 9276 5374 9285
rect 5066 9274 5072 9276
rect 5128 9274 5152 9276
rect 5208 9274 5232 9276
rect 5288 9274 5312 9276
rect 5368 9274 5374 9276
rect 5128 9222 5130 9274
rect 5310 9222 5312 9274
rect 5066 9220 5072 9222
rect 5128 9220 5152 9222
rect 5208 9220 5232 9222
rect 5288 9220 5312 9222
rect 5368 9220 5374 9222
rect 5066 9211 5374 9220
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5066 8188 5374 8197
rect 5066 8186 5072 8188
rect 5128 8186 5152 8188
rect 5208 8186 5232 8188
rect 5288 8186 5312 8188
rect 5368 8186 5374 8188
rect 5128 8134 5130 8186
rect 5310 8134 5312 8186
rect 5066 8132 5072 8134
rect 5128 8132 5152 8134
rect 5208 8132 5232 8134
rect 5288 8132 5312 8134
rect 5368 8132 5374 8134
rect 5066 8123 5374 8132
rect 5460 7449 5488 8434
rect 5446 7440 5502 7449
rect 5446 7375 5502 7384
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5460 7177 5488 7210
rect 5446 7168 5502 7177
rect 5066 7100 5374 7109
rect 5446 7103 5502 7112
rect 5066 7098 5072 7100
rect 5128 7098 5152 7100
rect 5208 7098 5232 7100
rect 5288 7098 5312 7100
rect 5368 7098 5374 7100
rect 5128 7046 5130 7098
rect 5310 7046 5312 7098
rect 5066 7044 5072 7046
rect 5128 7044 5152 7046
rect 5208 7044 5232 7046
rect 5288 7044 5312 7046
rect 5368 7044 5374 7046
rect 5066 7035 5374 7044
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4816 3534 4844 4694
rect 4908 4146 4936 5850
rect 5000 5846 5028 6190
rect 5066 6012 5374 6021
rect 5066 6010 5072 6012
rect 5128 6010 5152 6012
rect 5208 6010 5232 6012
rect 5288 6010 5312 6012
rect 5368 6010 5374 6012
rect 5128 5958 5130 6010
rect 5310 5958 5312 6010
rect 5066 5956 5072 5958
rect 5128 5956 5152 5958
rect 5208 5956 5232 5958
rect 5288 5956 5312 5958
rect 5368 5956 5374 5958
rect 5066 5947 5374 5956
rect 4988 5840 5040 5846
rect 4988 5782 5040 5788
rect 5000 5574 5028 5782
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 5066 4924 5374 4933
rect 5066 4922 5072 4924
rect 5128 4922 5152 4924
rect 5208 4922 5232 4924
rect 5288 4922 5312 4924
rect 5368 4922 5374 4924
rect 5128 4870 5130 4922
rect 5310 4870 5312 4922
rect 5066 4868 5072 4870
rect 5128 4868 5152 4870
rect 5208 4868 5232 4870
rect 5288 4868 5312 4870
rect 5368 4868 5374 4870
rect 5066 4859 5374 4868
rect 5354 4176 5410 4185
rect 4896 4140 4948 4146
rect 5354 4111 5410 4120
rect 4896 4082 4948 4088
rect 5368 4078 5396 4111
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5460 4010 5488 6938
rect 5552 4078 5580 9998
rect 5828 9625 5856 12294
rect 5998 12200 6054 13000
rect 6458 12322 6514 13000
rect 10046 12336 10102 12345
rect 6458 12294 6592 12322
rect 6092 12232 6144 12238
rect 5908 10600 5960 10606
rect 5908 10542 5960 10548
rect 5814 9616 5870 9625
rect 5724 9580 5776 9586
rect 5814 9551 5870 9560
rect 5724 9522 5776 9528
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5644 8537 5672 9318
rect 5736 8809 5764 9522
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5722 8800 5778 8809
rect 5722 8735 5778 8744
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5630 8528 5686 8537
rect 5630 8463 5686 8472
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5644 7410 5672 7822
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5644 6322 5672 7210
rect 5736 6798 5764 8570
rect 5828 7177 5856 9454
rect 5814 7168 5870 7177
rect 5814 7103 5870 7112
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5722 6624 5778 6633
rect 5722 6559 5778 6568
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5644 5370 5672 6258
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4632 2746 4752 2774
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4632 2106 4660 2746
rect 4908 2514 4936 3946
rect 5538 3904 5594 3913
rect 5066 3836 5374 3845
rect 5538 3839 5594 3848
rect 5066 3834 5072 3836
rect 5128 3834 5152 3836
rect 5208 3834 5232 3836
rect 5288 3834 5312 3836
rect 5368 3834 5374 3836
rect 5128 3782 5130 3834
rect 5310 3782 5312 3834
rect 5066 3780 5072 3782
rect 5128 3780 5152 3782
rect 5208 3780 5232 3782
rect 5288 3780 5312 3782
rect 5368 3780 5374 3782
rect 5066 3771 5374 3780
rect 5080 3528 5132 3534
rect 5078 3496 5080 3505
rect 5132 3496 5134 3505
rect 5078 3431 5134 3440
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 5000 3126 5028 3334
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 5000 2990 5028 3062
rect 4988 2984 5040 2990
rect 4988 2926 5040 2932
rect 5000 2650 5028 2926
rect 5066 2748 5374 2757
rect 5066 2746 5072 2748
rect 5128 2746 5152 2748
rect 5208 2746 5232 2748
rect 5288 2746 5312 2748
rect 5368 2746 5374 2748
rect 5128 2694 5130 2746
rect 5310 2694 5312 2746
rect 5066 2692 5072 2694
rect 5128 2692 5152 2694
rect 5208 2692 5232 2694
rect 5288 2692 5312 2694
rect 5368 2692 5374 2694
rect 5066 2683 5374 2692
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 4896 2508 4948 2514
rect 4896 2450 4948 2456
rect 3884 2100 3936 2106
rect 3884 2042 3936 2048
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 4620 2100 4672 2106
rect 4620 2042 4672 2048
rect 3608 1896 3660 1902
rect 3608 1838 3660 1844
rect 5000 1018 5028 2586
rect 5066 1660 5374 1669
rect 5066 1658 5072 1660
rect 5128 1658 5152 1660
rect 5208 1658 5232 1660
rect 5288 1658 5312 1660
rect 5368 1658 5374 1660
rect 5128 1606 5130 1658
rect 5310 1606 5312 1658
rect 5066 1604 5072 1606
rect 5128 1604 5152 1606
rect 5208 1604 5232 1606
rect 5288 1604 5312 1606
rect 5368 1604 5374 1606
rect 5066 1595 5374 1604
rect 5552 1562 5580 3839
rect 5644 2310 5672 4014
rect 5736 2774 5764 6559
rect 5828 5778 5856 7103
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5828 4078 5856 5238
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5736 2746 5856 2774
rect 5828 2310 5856 2746
rect 5632 2304 5684 2310
rect 5632 2246 5684 2252
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5540 1556 5592 1562
rect 5540 1498 5592 1504
rect 5448 1352 5500 1358
rect 5446 1320 5448 1329
rect 5500 1320 5502 1329
rect 5446 1255 5502 1264
rect 5644 1222 5672 2246
rect 5632 1216 5684 1222
rect 5632 1158 5684 1164
rect 4988 1012 5040 1018
rect 4988 954 5040 960
rect 3424 944 3476 950
rect 3424 886 3476 892
rect 5644 746 5672 1158
rect 5920 882 5948 10542
rect 6012 9382 6040 12200
rect 6458 12200 6514 12294
rect 6092 12174 6144 12180
rect 6104 11694 6132 12174
rect 6564 12050 6592 12294
rect 10046 12271 10102 12280
rect 6196 12022 6592 12050
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6104 10441 6132 11630
rect 6090 10432 6146 10441
rect 6090 10367 6146 10376
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 6104 9194 6132 10367
rect 6012 9166 6132 9194
rect 6012 8673 6040 9166
rect 6196 8906 6224 12022
rect 7566 11996 7874 12005
rect 7566 11994 7572 11996
rect 7628 11994 7652 11996
rect 7708 11994 7732 11996
rect 7788 11994 7812 11996
rect 7868 11994 7874 11996
rect 7628 11942 7630 11994
rect 7810 11942 7812 11994
rect 7566 11940 7572 11942
rect 7628 11940 7652 11942
rect 7708 11940 7732 11942
rect 7788 11940 7812 11942
rect 7868 11940 7874 11942
rect 7566 11931 7874 11940
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6380 11234 6408 11834
rect 6472 11694 6500 11834
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6288 10606 6316 11222
rect 6380 11206 6500 11234
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6288 10266 6316 10542
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6288 9110 6316 9998
rect 6276 9104 6328 9110
rect 6276 9046 6328 9052
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 5998 8664 6054 8673
rect 5998 8599 6054 8608
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6012 7410 6040 8434
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6104 5710 6132 8842
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6196 7478 6224 8366
rect 6288 8022 6316 8910
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6012 5166 6040 5646
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 6104 4690 6132 5034
rect 6092 4684 6144 4690
rect 6092 4626 6144 4632
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 6012 3942 6040 4490
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6104 3602 6132 4422
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6012 2650 6040 3130
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 6104 1358 6132 2246
rect 6196 1426 6224 6598
rect 6288 4078 6316 7686
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6380 3602 6408 11086
rect 6472 5302 6500 11206
rect 6550 9344 6606 9353
rect 6550 9279 6606 9288
rect 6564 8498 6592 9279
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6564 7818 6592 8298
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6552 6792 6604 6798
rect 6550 6760 6552 6769
rect 6604 6760 6606 6769
rect 6550 6695 6606 6704
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6564 5846 6592 6190
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6564 5166 6592 5646
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6472 3058 6500 5102
rect 6564 4690 6592 5102
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6656 4554 6684 11630
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6748 10674 6776 11086
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6748 9353 6776 9386
rect 6734 9344 6790 9353
rect 6734 9279 6790 9288
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6748 7342 6776 8774
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6840 5794 6868 11494
rect 6932 10810 6960 11630
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6918 10704 6974 10713
rect 6918 10639 6974 10648
rect 6932 6458 6960 10639
rect 7024 10130 7052 11698
rect 7194 10840 7250 10849
rect 7194 10775 7196 10784
rect 7248 10775 7250 10784
rect 7196 10746 7248 10752
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 7116 9450 7144 9998
rect 7300 9586 7328 11834
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7300 9450 7328 9522
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7392 9330 7420 10678
rect 7484 10606 7512 11562
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 7566 10908 7874 10917
rect 7566 10906 7572 10908
rect 7628 10906 7652 10908
rect 7708 10906 7732 10908
rect 7788 10906 7812 10908
rect 7868 10906 7874 10908
rect 7628 10854 7630 10906
rect 7810 10854 7812 10906
rect 7566 10852 7572 10854
rect 7628 10852 7652 10854
rect 7708 10852 7732 10854
rect 7788 10852 7812 10854
rect 7868 10852 7874 10854
rect 7566 10843 7874 10852
rect 7944 10810 7972 11086
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7566 9820 7874 9829
rect 7566 9818 7572 9820
rect 7628 9818 7652 9820
rect 7708 9818 7732 9820
rect 7788 9818 7812 9820
rect 7868 9818 7874 9820
rect 7628 9766 7630 9818
rect 7810 9766 7812 9818
rect 7566 9764 7572 9766
rect 7628 9764 7652 9766
rect 7708 9764 7732 9766
rect 7788 9764 7812 9766
rect 7868 9764 7874 9766
rect 7566 9755 7874 9764
rect 7944 9654 7972 9862
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7300 9302 7420 9330
rect 7300 8974 7328 9302
rect 7484 9110 7512 9522
rect 7576 9489 7604 9522
rect 7562 9480 7618 9489
rect 7562 9415 7618 9424
rect 7472 9104 7524 9110
rect 7472 9046 7524 9052
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7288 8968 7340 8974
rect 7102 8936 7158 8945
rect 7484 8945 7512 9046
rect 7288 8910 7340 8916
rect 7470 8936 7526 8945
rect 7102 8871 7158 8880
rect 7116 7018 7144 8871
rect 7194 8800 7250 8809
rect 7194 8735 7250 8744
rect 7024 6990 7144 7018
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6748 5766 6868 5794
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6748 4434 6776 5766
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6840 4690 6868 5578
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6656 4406 6776 4434
rect 6656 3738 6684 4406
rect 6840 4298 6868 4626
rect 6932 4554 6960 6122
rect 7024 5370 7052 6990
rect 7102 6896 7158 6905
rect 7102 6831 7158 6840
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7024 4826 7052 5102
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6920 4548 6972 4554
rect 6920 4490 6972 4496
rect 6748 4270 6868 4298
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6748 3194 6776 4270
rect 6826 4176 6882 4185
rect 6826 4111 6882 4120
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6840 3058 6868 4111
rect 7116 3641 7144 6831
rect 7102 3632 7158 3641
rect 7102 3567 7158 3576
rect 7208 3058 7236 8735
rect 7300 7954 7328 8910
rect 7470 8871 7526 8880
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7300 7274 7328 7754
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7392 6882 7420 8774
rect 7484 8344 7512 8774
rect 7566 8732 7874 8741
rect 7566 8730 7572 8732
rect 7628 8730 7652 8732
rect 7708 8730 7732 8732
rect 7788 8730 7812 8732
rect 7868 8730 7874 8732
rect 7628 8678 7630 8730
rect 7810 8678 7812 8730
rect 7566 8676 7572 8678
rect 7628 8676 7652 8678
rect 7708 8676 7732 8678
rect 7788 8676 7812 8678
rect 7868 8676 7874 8678
rect 7566 8667 7874 8676
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7564 8356 7616 8362
rect 7484 8316 7564 8344
rect 7484 8022 7512 8316
rect 7564 8298 7616 8304
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7852 8090 7880 8230
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7484 6984 7512 7958
rect 7566 7644 7874 7653
rect 7566 7642 7572 7644
rect 7628 7642 7652 7644
rect 7708 7642 7732 7644
rect 7788 7642 7812 7644
rect 7868 7642 7874 7644
rect 7628 7590 7630 7642
rect 7810 7590 7812 7642
rect 7566 7588 7572 7590
rect 7628 7588 7652 7590
rect 7708 7588 7732 7590
rect 7788 7588 7812 7590
rect 7868 7588 7874 7590
rect 7566 7579 7874 7588
rect 7564 6996 7616 7002
rect 7484 6956 7564 6984
rect 7564 6938 7616 6944
rect 7300 6854 7420 6882
rect 7300 4554 7328 6854
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7392 6322 7420 6734
rect 7566 6556 7874 6565
rect 7566 6554 7572 6556
rect 7628 6554 7652 6556
rect 7708 6554 7732 6556
rect 7788 6554 7812 6556
rect 7868 6554 7874 6556
rect 7628 6502 7630 6554
rect 7810 6502 7812 6554
rect 7566 6500 7572 6502
rect 7628 6500 7652 6502
rect 7708 6500 7732 6502
rect 7788 6500 7812 6502
rect 7868 6500 7874 6502
rect 7566 6491 7874 6500
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7484 5166 7512 6394
rect 7566 5468 7874 5477
rect 7566 5466 7572 5468
rect 7628 5466 7652 5468
rect 7708 5466 7732 5468
rect 7788 5466 7812 5468
rect 7868 5466 7874 5468
rect 7628 5414 7630 5466
rect 7810 5414 7812 5466
rect 7566 5412 7572 5414
rect 7628 5412 7652 5414
rect 7708 5412 7732 5414
rect 7788 5412 7812 5414
rect 7868 5412 7874 5414
rect 7566 5403 7874 5412
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7668 4690 7696 5306
rect 7944 5234 7972 8366
rect 8036 6458 8064 9046
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8128 6390 8156 10202
rect 8220 8673 8248 11698
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8392 11280 8444 11286
rect 8392 11222 8444 11228
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8312 9586 8340 10678
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8206 8664 8262 8673
rect 8206 8599 8262 8608
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8312 7886 8340 8502
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 7410 8248 7686
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7944 4758 7972 5170
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7288 4548 7340 4554
rect 7668 4536 7696 4626
rect 7288 4490 7340 4496
rect 7392 4508 7696 4536
rect 7300 3126 7328 4490
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 6826 2952 6882 2961
rect 6826 2887 6882 2896
rect 6840 1970 6868 2887
rect 7392 2774 7420 4508
rect 7566 4380 7874 4389
rect 7566 4378 7572 4380
rect 7628 4378 7652 4380
rect 7708 4378 7732 4380
rect 7788 4378 7812 4380
rect 7868 4378 7874 4380
rect 7628 4326 7630 4378
rect 7810 4326 7812 4378
rect 7566 4324 7572 4326
rect 7628 4324 7652 4326
rect 7708 4324 7732 4326
rect 7788 4324 7812 4326
rect 7868 4324 7874 4326
rect 7566 4315 7874 4324
rect 7566 3292 7874 3301
rect 7566 3290 7572 3292
rect 7628 3290 7652 3292
rect 7708 3290 7732 3292
rect 7788 3290 7812 3292
rect 7868 3290 7874 3292
rect 7628 3238 7630 3290
rect 7810 3238 7812 3290
rect 7566 3236 7572 3238
rect 7628 3236 7652 3238
rect 7708 3236 7732 3238
rect 7788 3236 7812 3238
rect 7868 3236 7874 3238
rect 7566 3227 7874 3236
rect 7300 2746 7420 2774
rect 7300 2650 7328 2746
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7566 2204 7874 2213
rect 7566 2202 7572 2204
rect 7628 2202 7652 2204
rect 7708 2202 7732 2204
rect 7788 2202 7812 2204
rect 7868 2202 7874 2204
rect 7628 2150 7630 2202
rect 7810 2150 7812 2202
rect 7566 2148 7572 2150
rect 7628 2148 7652 2150
rect 7708 2148 7732 2150
rect 7788 2148 7812 2150
rect 7868 2148 7874 2150
rect 7566 2139 7874 2148
rect 6828 1964 6880 1970
rect 6828 1906 6880 1912
rect 8036 1902 8064 6054
rect 8220 5846 8248 6938
rect 8312 6934 8340 7822
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8128 5370 8156 5646
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8114 2544 8170 2553
rect 8312 2514 8340 5238
rect 8404 4622 8432 11222
rect 8496 10198 8524 11562
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8482 9616 8538 9625
rect 8482 9551 8538 9560
rect 8496 8430 8524 9551
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8484 8288 8536 8294
rect 8484 8230 8536 8236
rect 8496 7410 8524 8230
rect 8588 7546 8616 11086
rect 8668 10464 8720 10470
rect 8666 10432 8668 10441
rect 8720 10432 8722 10441
rect 8666 10367 8722 10376
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8680 8634 8708 10066
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8772 8514 8800 9862
rect 8864 9382 8892 11494
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8680 8486 8800 8514
rect 8864 8498 8892 8842
rect 8852 8492 8904 8498
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8576 7268 8628 7274
rect 8576 7210 8628 7216
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5098 8524 5510
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8588 4078 8616 7210
rect 8680 6322 8708 8486
rect 8852 8434 8904 8440
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8390 3632 8446 3641
rect 8390 3567 8446 3576
rect 8404 2514 8432 3567
rect 8680 2922 8708 6258
rect 8772 6118 8800 8366
rect 8864 6866 8892 8434
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 8956 6746 8984 11154
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9128 10600 9180 10606
rect 9588 10600 9640 10606
rect 9128 10542 9180 10548
rect 9586 10568 9588 10577
rect 9640 10568 9642 10577
rect 9140 9450 9168 10542
rect 9586 10503 9642 10512
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9140 7342 9168 9386
rect 9128 7336 9180 7342
rect 8864 6718 8984 6746
rect 9048 7296 9128 7324
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8772 5710 8800 6054
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8864 2582 8892 6718
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8852 2576 8904 2582
rect 8852 2518 8904 2524
rect 8114 2479 8170 2488
rect 8300 2508 8352 2514
rect 8128 2378 8156 2479
rect 8300 2450 8352 2456
rect 8392 2508 8444 2514
rect 8392 2450 8444 2456
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8116 2372 8168 2378
rect 8116 2314 8168 2320
rect 8772 2258 8800 2450
rect 8588 2230 8800 2258
rect 8116 2032 8168 2038
rect 8116 1974 8168 1980
rect 8024 1896 8076 1902
rect 8024 1838 8076 1844
rect 8128 1562 8156 1974
rect 8588 1834 8616 2230
rect 8576 1828 8628 1834
rect 8576 1770 8628 1776
rect 8116 1556 8168 1562
rect 8116 1498 8168 1504
rect 6184 1420 6236 1426
rect 6184 1362 6236 1368
rect 6092 1352 6144 1358
rect 6092 1294 6144 1300
rect 8588 1222 8616 1770
rect 8850 1728 8906 1737
rect 8850 1663 8906 1672
rect 8864 1426 8892 1663
rect 8956 1562 8984 6190
rect 9048 5681 9076 7296
rect 9128 7278 9180 7284
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9140 5778 9168 6666
rect 9232 6458 9260 9454
rect 9416 7954 9444 9998
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9402 7032 9458 7041
rect 9402 6967 9458 6976
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9034 5672 9090 5681
rect 9034 5607 9090 5616
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 9048 3670 9076 4966
rect 9036 3664 9088 3670
rect 9036 3606 9088 3612
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 8944 1556 8996 1562
rect 8944 1498 8996 1504
rect 8852 1420 8904 1426
rect 8852 1362 8904 1368
rect 8760 1284 8812 1290
rect 8760 1226 8812 1232
rect 8576 1216 8628 1222
rect 8576 1158 8628 1164
rect 7566 1116 7874 1125
rect 7566 1114 7572 1116
rect 7628 1114 7652 1116
rect 7708 1114 7732 1116
rect 7788 1114 7812 1116
rect 7868 1114 7874 1116
rect 7628 1062 7630 1114
rect 7810 1062 7812 1114
rect 7566 1060 7572 1062
rect 7628 1060 7652 1062
rect 7708 1060 7732 1062
rect 7788 1060 7812 1062
rect 7868 1060 7874 1062
rect 7566 1051 7874 1060
rect 8772 1018 8800 1226
rect 8760 1012 8812 1018
rect 8760 954 8812 960
rect 5908 876 5960 882
rect 5908 818 5960 824
rect 8864 746 8892 1362
rect 9048 1018 9076 2382
rect 9140 1562 9168 5510
rect 9232 3398 9260 6394
rect 9324 5846 9352 6802
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9312 5704 9364 5710
rect 9310 5672 9312 5681
rect 9364 5672 9366 5681
rect 9310 5607 9366 5616
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9324 5370 9352 5510
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9416 4146 9444 6967
rect 9508 6866 9536 9522
rect 9586 9480 9642 9489
rect 9586 9415 9642 9424
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9508 3738 9536 6666
rect 9600 4826 9628 9415
rect 9784 8838 9812 9998
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9692 8022 9720 8570
rect 9784 8430 9812 8774
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9692 6322 9720 7278
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9876 6254 9904 11018
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9588 4820 9640 4826
rect 9588 4762 9640 4768
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9494 3632 9550 3641
rect 9494 3567 9550 3576
rect 9588 3596 9640 3602
rect 9508 3398 9536 3567
rect 9588 3538 9640 3544
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9232 2446 9260 3062
rect 9600 2650 9628 3538
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9312 1828 9364 1834
rect 9312 1770 9364 1776
rect 9128 1556 9180 1562
rect 9128 1498 9180 1504
rect 9220 1488 9272 1494
rect 9220 1430 9272 1436
rect 9036 1012 9088 1018
rect 9036 954 9088 960
rect 3056 740 3108 746
rect 3056 682 3108 688
rect 5632 740 5684 746
rect 5632 682 5684 688
rect 8852 740 8904 746
rect 8852 682 8904 688
rect 9232 678 9260 1430
rect 9324 1358 9352 1770
rect 9600 1426 9628 2586
rect 9588 1420 9640 1426
rect 9588 1362 9640 1368
rect 9312 1352 9364 1358
rect 9312 1294 9364 1300
rect 9312 1216 9364 1222
rect 9312 1158 9364 1164
rect 9324 814 9352 1158
rect 9692 1018 9720 5646
rect 9784 5098 9812 6054
rect 9772 5092 9824 5098
rect 9772 5034 9824 5040
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9784 2446 9812 3538
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9680 1012 9732 1018
rect 9680 954 9732 960
rect 9784 882 9812 2246
rect 9876 1902 9904 6190
rect 9864 1896 9916 1902
rect 9864 1838 9916 1844
rect 9968 1018 9996 9522
rect 10060 5778 10088 12271
rect 13818 11928 13874 11937
rect 13818 11863 13820 11872
rect 13872 11863 13874 11872
rect 17960 11892 18012 11898
rect 13820 11834 13872 11840
rect 17960 11834 18012 11840
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10244 9382 10272 9998
rect 11058 9888 11114 9897
rect 11058 9823 11114 9832
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10244 8566 10272 9318
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10046 3768 10102 3777
rect 10046 3703 10102 3712
rect 10060 2650 10088 3703
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 10060 2106 10088 2450
rect 10152 2310 10180 5034
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10138 2136 10194 2145
rect 10048 2100 10100 2106
rect 10138 2071 10194 2080
rect 10048 2042 10100 2048
rect 10152 1986 10180 2071
rect 10060 1958 10180 1986
rect 10060 1766 10088 1958
rect 10048 1760 10100 1766
rect 10048 1702 10100 1708
rect 9956 1012 10008 1018
rect 9956 954 10008 960
rect 9772 876 9824 882
rect 9772 818 9824 824
rect 10060 814 10088 1702
rect 10244 1290 10272 8502
rect 11072 5914 11100 9823
rect 17972 7206 18000 11834
rect 22098 11112 22154 11121
rect 22098 11047 22154 11056
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 16578 6624 16634 6633
rect 16578 6559 16634 6568
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 16592 5574 16620 6559
rect 16854 6216 16910 6225
rect 16854 6151 16910 6160
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16578 5400 16634 5409
rect 16578 5335 16634 5344
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10336 1426 10364 5170
rect 16592 4010 16620 5335
rect 16670 4992 16726 5001
rect 16670 4927 16726 4936
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16684 3534 16712 4927
rect 16762 4584 16818 4593
rect 16762 4519 16818 4528
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 16578 2544 16634 2553
rect 16578 2479 16634 2488
rect 16592 2038 16620 2479
rect 16580 2032 16632 2038
rect 16580 1974 16632 1980
rect 16776 1834 16804 4519
rect 16868 2922 16896 6151
rect 16946 5808 17002 5817
rect 16946 5743 17002 5752
rect 16856 2916 16908 2922
rect 16856 2858 16908 2864
rect 16960 2514 16988 5743
rect 22112 3942 22140 11047
rect 22282 8256 22338 8265
rect 22282 8191 22338 8200
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 22296 1970 22324 8191
rect 22284 1964 22336 1970
rect 22284 1906 22336 1912
rect 16764 1828 16816 1834
rect 16764 1770 16816 1776
rect 10324 1420 10376 1426
rect 10324 1362 10376 1368
rect 10232 1284 10284 1290
rect 10232 1226 10284 1232
rect 13820 944 13872 950
rect 13818 912 13820 921
rect 13872 912 13874 921
rect 13818 847 13874 856
rect 9312 808 9364 814
rect 9312 750 9364 756
rect 10048 808 10100 814
rect 10048 750 10100 756
rect 2320 672 2372 678
rect 2320 614 2372 620
rect 5448 672 5500 678
rect 5448 614 5500 620
rect 9220 672 9272 678
rect 9220 614 9272 620
rect 5066 572 5374 581
rect 5066 570 5072 572
rect 5128 570 5152 572
rect 5208 570 5232 572
rect 5288 570 5312 572
rect 5368 570 5374 572
rect 5128 518 5130 570
rect 5310 518 5312 570
rect 5066 516 5072 518
rect 5128 516 5152 518
rect 5208 516 5232 518
rect 5288 516 5312 518
rect 5368 516 5374 518
rect 5066 507 5374 516
rect 5460 513 5488 614
rect 5446 504 5502 513
rect 5446 439 5502 448
<< via2 >>
rect 1398 11056 1454 11112
rect 1214 9288 1270 9344
rect 2572 11994 2628 11996
rect 2652 11994 2708 11996
rect 2732 11994 2788 11996
rect 2812 11994 2868 11996
rect 2572 11942 2618 11994
rect 2618 11942 2628 11994
rect 2652 11942 2682 11994
rect 2682 11942 2694 11994
rect 2694 11942 2708 11994
rect 2732 11942 2746 11994
rect 2746 11942 2758 11994
rect 2758 11942 2788 11994
rect 2812 11942 2822 11994
rect 2822 11942 2868 11994
rect 2572 11940 2628 11942
rect 2652 11940 2708 11942
rect 2732 11940 2788 11942
rect 2812 11940 2868 11942
rect 2502 11600 2558 11656
rect 2572 10906 2628 10908
rect 2652 10906 2708 10908
rect 2732 10906 2788 10908
rect 2812 10906 2868 10908
rect 2572 10854 2618 10906
rect 2618 10854 2628 10906
rect 2652 10854 2682 10906
rect 2682 10854 2694 10906
rect 2694 10854 2708 10906
rect 2732 10854 2746 10906
rect 2746 10854 2758 10906
rect 2758 10854 2788 10906
rect 2812 10854 2822 10906
rect 2822 10854 2868 10906
rect 2572 10852 2628 10854
rect 2652 10852 2708 10854
rect 2732 10852 2788 10854
rect 2812 10852 2868 10854
rect 2778 10648 2834 10704
rect 1306 8200 1362 8256
rect 2134 8472 2190 8528
rect 3054 10512 3110 10568
rect 2870 9968 2926 10024
rect 2962 9832 3018 9888
rect 2572 9818 2628 9820
rect 2652 9818 2708 9820
rect 2732 9818 2788 9820
rect 2812 9818 2868 9820
rect 2572 9766 2618 9818
rect 2618 9766 2628 9818
rect 2652 9766 2682 9818
rect 2682 9766 2694 9818
rect 2694 9766 2708 9818
rect 2732 9766 2746 9818
rect 2746 9766 2758 9818
rect 2758 9766 2788 9818
rect 2812 9766 2822 9818
rect 2822 9766 2868 9818
rect 2572 9764 2628 9766
rect 2652 9764 2708 9766
rect 2732 9764 2788 9766
rect 2812 9764 2868 9766
rect 2778 9424 2834 9480
rect 2572 8730 2628 8732
rect 2652 8730 2708 8732
rect 2732 8730 2788 8732
rect 2812 8730 2868 8732
rect 2572 8678 2618 8730
rect 2618 8678 2628 8730
rect 2652 8678 2682 8730
rect 2682 8678 2694 8730
rect 2694 8678 2708 8730
rect 2732 8678 2746 8730
rect 2746 8678 2758 8730
rect 2758 8678 2788 8730
rect 2812 8678 2822 8730
rect 2822 8678 2868 8730
rect 2572 8676 2628 8678
rect 2652 8676 2708 8678
rect 2732 8676 2788 8678
rect 2812 8676 2868 8678
rect 2502 7812 2558 7848
rect 2502 7792 2504 7812
rect 2504 7792 2556 7812
rect 2556 7792 2558 7812
rect 2572 7642 2628 7644
rect 2652 7642 2708 7644
rect 2732 7642 2788 7644
rect 2812 7642 2868 7644
rect 2572 7590 2618 7642
rect 2618 7590 2628 7642
rect 2652 7590 2682 7642
rect 2682 7590 2694 7642
rect 2694 7590 2708 7642
rect 2732 7590 2746 7642
rect 2746 7590 2758 7642
rect 2758 7590 2788 7642
rect 2812 7590 2822 7642
rect 2822 7590 2868 7642
rect 2572 7588 2628 7590
rect 2652 7588 2708 7590
rect 2732 7588 2788 7590
rect 2812 7588 2868 7590
rect 2572 6554 2628 6556
rect 2652 6554 2708 6556
rect 2732 6554 2788 6556
rect 2812 6554 2868 6556
rect 2572 6502 2618 6554
rect 2618 6502 2628 6554
rect 2652 6502 2682 6554
rect 2682 6502 2694 6554
rect 2694 6502 2708 6554
rect 2732 6502 2746 6554
rect 2746 6502 2758 6554
rect 2758 6502 2788 6554
rect 2812 6502 2822 6554
rect 2822 6502 2868 6554
rect 2572 6500 2628 6502
rect 2652 6500 2708 6502
rect 2732 6500 2788 6502
rect 2812 6500 2868 6502
rect 2778 6316 2834 6352
rect 2778 6296 2780 6316
rect 2780 6296 2832 6316
rect 2832 6296 2834 6316
rect 2572 5466 2628 5468
rect 2652 5466 2708 5468
rect 2732 5466 2788 5468
rect 2812 5466 2868 5468
rect 2572 5414 2618 5466
rect 2618 5414 2628 5466
rect 2652 5414 2682 5466
rect 2682 5414 2694 5466
rect 2694 5414 2708 5466
rect 2732 5414 2746 5466
rect 2746 5414 2758 5466
rect 2758 5414 2788 5466
rect 2812 5414 2822 5466
rect 2822 5414 2868 5466
rect 2572 5412 2628 5414
rect 2652 5412 2708 5414
rect 2732 5412 2788 5414
rect 2812 5412 2868 5414
rect 2686 3408 2688 3428
rect 2688 3408 2740 3428
rect 2740 3408 2742 3428
rect 2686 3372 2742 3408
rect 3606 11192 3662 11248
rect 3330 10784 3386 10840
rect 3330 8336 3386 8392
rect 2572 1114 2628 1116
rect 2652 1114 2708 1116
rect 2732 1114 2788 1116
rect 2812 1114 2868 1116
rect 2572 1062 2618 1114
rect 2618 1062 2628 1114
rect 2652 1062 2682 1114
rect 2682 1062 2694 1114
rect 2694 1062 2708 1114
rect 2732 1062 2746 1114
rect 2746 1062 2758 1114
rect 2758 1062 2788 1114
rect 2812 1062 2822 1114
rect 2822 1062 2868 1114
rect 2572 1060 2628 1062
rect 2652 1060 2708 1062
rect 2732 1060 2788 1062
rect 2812 1060 2868 1062
rect 3790 9016 3846 9072
rect 3882 8608 3938 8664
rect 3882 8336 3938 8392
rect 3882 6704 3938 6760
rect 4342 11056 4398 11112
rect 4250 8880 4306 8936
rect 4250 8608 4306 8664
rect 4066 7248 4122 7304
rect 4066 6704 4122 6760
rect 3790 2508 3846 2544
rect 3790 2488 3792 2508
rect 3792 2488 3844 2508
rect 3844 2488 3846 2508
rect 5072 11450 5128 11452
rect 5152 11450 5208 11452
rect 5232 11450 5288 11452
rect 5312 11450 5368 11452
rect 5072 11398 5118 11450
rect 5118 11398 5128 11450
rect 5152 11398 5182 11450
rect 5182 11398 5194 11450
rect 5194 11398 5208 11450
rect 5232 11398 5246 11450
rect 5246 11398 5258 11450
rect 5258 11398 5288 11450
rect 5312 11398 5322 11450
rect 5322 11398 5368 11450
rect 5072 11396 5128 11398
rect 5152 11396 5208 11398
rect 5232 11396 5288 11398
rect 5312 11396 5368 11398
rect 5354 10532 5410 10568
rect 5354 10512 5356 10532
rect 5356 10512 5408 10532
rect 5408 10512 5410 10532
rect 5072 10362 5128 10364
rect 5152 10362 5208 10364
rect 5232 10362 5288 10364
rect 5312 10362 5368 10364
rect 5072 10310 5118 10362
rect 5118 10310 5128 10362
rect 5152 10310 5182 10362
rect 5182 10310 5194 10362
rect 5194 10310 5208 10362
rect 5232 10310 5246 10362
rect 5246 10310 5258 10362
rect 5258 10310 5288 10362
rect 5312 10310 5322 10362
rect 5322 10310 5368 10362
rect 5072 10308 5128 10310
rect 5152 10308 5208 10310
rect 5232 10308 5288 10310
rect 5312 10308 5368 10310
rect 5538 10512 5594 10568
rect 5446 10240 5502 10296
rect 4894 9424 4950 9480
rect 4802 9288 4858 9344
rect 4434 8200 4490 8256
rect 4250 6840 4306 6896
rect 4158 6296 4214 6352
rect 5354 9560 5410 9616
rect 5072 9274 5128 9276
rect 5152 9274 5208 9276
rect 5232 9274 5288 9276
rect 5312 9274 5368 9276
rect 5072 9222 5118 9274
rect 5118 9222 5128 9274
rect 5152 9222 5182 9274
rect 5182 9222 5194 9274
rect 5194 9222 5208 9274
rect 5232 9222 5246 9274
rect 5246 9222 5258 9274
rect 5258 9222 5288 9274
rect 5312 9222 5322 9274
rect 5322 9222 5368 9274
rect 5072 9220 5128 9222
rect 5152 9220 5208 9222
rect 5232 9220 5288 9222
rect 5312 9220 5368 9222
rect 5072 8186 5128 8188
rect 5152 8186 5208 8188
rect 5232 8186 5288 8188
rect 5312 8186 5368 8188
rect 5072 8134 5118 8186
rect 5118 8134 5128 8186
rect 5152 8134 5182 8186
rect 5182 8134 5194 8186
rect 5194 8134 5208 8186
rect 5232 8134 5246 8186
rect 5246 8134 5258 8186
rect 5258 8134 5288 8186
rect 5312 8134 5322 8186
rect 5322 8134 5368 8186
rect 5072 8132 5128 8134
rect 5152 8132 5208 8134
rect 5232 8132 5288 8134
rect 5312 8132 5368 8134
rect 5446 7384 5502 7440
rect 5446 7112 5502 7168
rect 5072 7098 5128 7100
rect 5152 7098 5208 7100
rect 5232 7098 5288 7100
rect 5312 7098 5368 7100
rect 5072 7046 5118 7098
rect 5118 7046 5128 7098
rect 5152 7046 5182 7098
rect 5182 7046 5194 7098
rect 5194 7046 5208 7098
rect 5232 7046 5246 7098
rect 5246 7046 5258 7098
rect 5258 7046 5288 7098
rect 5312 7046 5322 7098
rect 5322 7046 5368 7098
rect 5072 7044 5128 7046
rect 5152 7044 5208 7046
rect 5232 7044 5288 7046
rect 5312 7044 5368 7046
rect 5072 6010 5128 6012
rect 5152 6010 5208 6012
rect 5232 6010 5288 6012
rect 5312 6010 5368 6012
rect 5072 5958 5118 6010
rect 5118 5958 5128 6010
rect 5152 5958 5182 6010
rect 5182 5958 5194 6010
rect 5194 5958 5208 6010
rect 5232 5958 5246 6010
rect 5246 5958 5258 6010
rect 5258 5958 5288 6010
rect 5312 5958 5322 6010
rect 5322 5958 5368 6010
rect 5072 5956 5128 5958
rect 5152 5956 5208 5958
rect 5232 5956 5288 5958
rect 5312 5956 5368 5958
rect 5072 4922 5128 4924
rect 5152 4922 5208 4924
rect 5232 4922 5288 4924
rect 5312 4922 5368 4924
rect 5072 4870 5118 4922
rect 5118 4870 5128 4922
rect 5152 4870 5182 4922
rect 5182 4870 5194 4922
rect 5194 4870 5208 4922
rect 5232 4870 5246 4922
rect 5246 4870 5258 4922
rect 5258 4870 5288 4922
rect 5312 4870 5322 4922
rect 5322 4870 5368 4922
rect 5072 4868 5128 4870
rect 5152 4868 5208 4870
rect 5232 4868 5288 4870
rect 5312 4868 5368 4870
rect 5354 4120 5410 4176
rect 5814 9560 5870 9616
rect 5722 8744 5778 8800
rect 5630 8472 5686 8528
rect 5814 7112 5870 7168
rect 5722 6568 5778 6624
rect 5538 3848 5594 3904
rect 5072 3834 5128 3836
rect 5152 3834 5208 3836
rect 5232 3834 5288 3836
rect 5312 3834 5368 3836
rect 5072 3782 5118 3834
rect 5118 3782 5128 3834
rect 5152 3782 5182 3834
rect 5182 3782 5194 3834
rect 5194 3782 5208 3834
rect 5232 3782 5246 3834
rect 5246 3782 5258 3834
rect 5258 3782 5288 3834
rect 5312 3782 5322 3834
rect 5322 3782 5368 3834
rect 5072 3780 5128 3782
rect 5152 3780 5208 3782
rect 5232 3780 5288 3782
rect 5312 3780 5368 3782
rect 5078 3476 5080 3496
rect 5080 3476 5132 3496
rect 5132 3476 5134 3496
rect 5078 3440 5134 3476
rect 5072 2746 5128 2748
rect 5152 2746 5208 2748
rect 5232 2746 5288 2748
rect 5312 2746 5368 2748
rect 5072 2694 5118 2746
rect 5118 2694 5128 2746
rect 5152 2694 5182 2746
rect 5182 2694 5194 2746
rect 5194 2694 5208 2746
rect 5232 2694 5246 2746
rect 5246 2694 5258 2746
rect 5258 2694 5288 2746
rect 5312 2694 5322 2746
rect 5322 2694 5368 2746
rect 5072 2692 5128 2694
rect 5152 2692 5208 2694
rect 5232 2692 5288 2694
rect 5312 2692 5368 2694
rect 5072 1658 5128 1660
rect 5152 1658 5208 1660
rect 5232 1658 5288 1660
rect 5312 1658 5368 1660
rect 5072 1606 5118 1658
rect 5118 1606 5128 1658
rect 5152 1606 5182 1658
rect 5182 1606 5194 1658
rect 5194 1606 5208 1658
rect 5232 1606 5246 1658
rect 5246 1606 5258 1658
rect 5258 1606 5288 1658
rect 5312 1606 5322 1658
rect 5322 1606 5368 1658
rect 5072 1604 5128 1606
rect 5152 1604 5208 1606
rect 5232 1604 5288 1606
rect 5312 1604 5368 1606
rect 5446 1300 5448 1320
rect 5448 1300 5500 1320
rect 5500 1300 5502 1320
rect 5446 1264 5502 1300
rect 10046 12280 10102 12336
rect 6090 10376 6146 10432
rect 7572 11994 7628 11996
rect 7652 11994 7708 11996
rect 7732 11994 7788 11996
rect 7812 11994 7868 11996
rect 7572 11942 7618 11994
rect 7618 11942 7628 11994
rect 7652 11942 7682 11994
rect 7682 11942 7694 11994
rect 7694 11942 7708 11994
rect 7732 11942 7746 11994
rect 7746 11942 7758 11994
rect 7758 11942 7788 11994
rect 7812 11942 7822 11994
rect 7822 11942 7868 11994
rect 7572 11940 7628 11942
rect 7652 11940 7708 11942
rect 7732 11940 7788 11942
rect 7812 11940 7868 11942
rect 5998 8608 6054 8664
rect 6550 9288 6606 9344
rect 6550 6740 6552 6760
rect 6552 6740 6604 6760
rect 6604 6740 6606 6760
rect 6550 6704 6606 6740
rect 6734 9288 6790 9344
rect 6918 10648 6974 10704
rect 7194 10804 7250 10840
rect 7194 10784 7196 10804
rect 7196 10784 7248 10804
rect 7248 10784 7250 10804
rect 7572 10906 7628 10908
rect 7652 10906 7708 10908
rect 7732 10906 7788 10908
rect 7812 10906 7868 10908
rect 7572 10854 7618 10906
rect 7618 10854 7628 10906
rect 7652 10854 7682 10906
rect 7682 10854 7694 10906
rect 7694 10854 7708 10906
rect 7732 10854 7746 10906
rect 7746 10854 7758 10906
rect 7758 10854 7788 10906
rect 7812 10854 7822 10906
rect 7822 10854 7868 10906
rect 7572 10852 7628 10854
rect 7652 10852 7708 10854
rect 7732 10852 7788 10854
rect 7812 10852 7868 10854
rect 7572 9818 7628 9820
rect 7652 9818 7708 9820
rect 7732 9818 7788 9820
rect 7812 9818 7868 9820
rect 7572 9766 7618 9818
rect 7618 9766 7628 9818
rect 7652 9766 7682 9818
rect 7682 9766 7694 9818
rect 7694 9766 7708 9818
rect 7732 9766 7746 9818
rect 7746 9766 7758 9818
rect 7758 9766 7788 9818
rect 7812 9766 7822 9818
rect 7822 9766 7868 9818
rect 7572 9764 7628 9766
rect 7652 9764 7708 9766
rect 7732 9764 7788 9766
rect 7812 9764 7868 9766
rect 7562 9424 7618 9480
rect 7102 8880 7158 8936
rect 7194 8744 7250 8800
rect 7102 6840 7158 6896
rect 6826 4120 6882 4176
rect 7102 3576 7158 3632
rect 7470 8880 7526 8936
rect 7572 8730 7628 8732
rect 7652 8730 7708 8732
rect 7732 8730 7788 8732
rect 7812 8730 7868 8732
rect 7572 8678 7618 8730
rect 7618 8678 7628 8730
rect 7652 8678 7682 8730
rect 7682 8678 7694 8730
rect 7694 8678 7708 8730
rect 7732 8678 7746 8730
rect 7746 8678 7758 8730
rect 7758 8678 7788 8730
rect 7812 8678 7822 8730
rect 7822 8678 7868 8730
rect 7572 8676 7628 8678
rect 7652 8676 7708 8678
rect 7732 8676 7788 8678
rect 7812 8676 7868 8678
rect 7572 7642 7628 7644
rect 7652 7642 7708 7644
rect 7732 7642 7788 7644
rect 7812 7642 7868 7644
rect 7572 7590 7618 7642
rect 7618 7590 7628 7642
rect 7652 7590 7682 7642
rect 7682 7590 7694 7642
rect 7694 7590 7708 7642
rect 7732 7590 7746 7642
rect 7746 7590 7758 7642
rect 7758 7590 7788 7642
rect 7812 7590 7822 7642
rect 7822 7590 7868 7642
rect 7572 7588 7628 7590
rect 7652 7588 7708 7590
rect 7732 7588 7788 7590
rect 7812 7588 7868 7590
rect 7572 6554 7628 6556
rect 7652 6554 7708 6556
rect 7732 6554 7788 6556
rect 7812 6554 7868 6556
rect 7572 6502 7618 6554
rect 7618 6502 7628 6554
rect 7652 6502 7682 6554
rect 7682 6502 7694 6554
rect 7694 6502 7708 6554
rect 7732 6502 7746 6554
rect 7746 6502 7758 6554
rect 7758 6502 7788 6554
rect 7812 6502 7822 6554
rect 7822 6502 7868 6554
rect 7572 6500 7628 6502
rect 7652 6500 7708 6502
rect 7732 6500 7788 6502
rect 7812 6500 7868 6502
rect 7572 5466 7628 5468
rect 7652 5466 7708 5468
rect 7732 5466 7788 5468
rect 7812 5466 7868 5468
rect 7572 5414 7618 5466
rect 7618 5414 7628 5466
rect 7652 5414 7682 5466
rect 7682 5414 7694 5466
rect 7694 5414 7708 5466
rect 7732 5414 7746 5466
rect 7746 5414 7758 5466
rect 7758 5414 7788 5466
rect 7812 5414 7822 5466
rect 7822 5414 7868 5466
rect 7572 5412 7628 5414
rect 7652 5412 7708 5414
rect 7732 5412 7788 5414
rect 7812 5412 7868 5414
rect 8206 8608 8262 8664
rect 6826 2896 6882 2952
rect 7572 4378 7628 4380
rect 7652 4378 7708 4380
rect 7732 4378 7788 4380
rect 7812 4378 7868 4380
rect 7572 4326 7618 4378
rect 7618 4326 7628 4378
rect 7652 4326 7682 4378
rect 7682 4326 7694 4378
rect 7694 4326 7708 4378
rect 7732 4326 7746 4378
rect 7746 4326 7758 4378
rect 7758 4326 7788 4378
rect 7812 4326 7822 4378
rect 7822 4326 7868 4378
rect 7572 4324 7628 4326
rect 7652 4324 7708 4326
rect 7732 4324 7788 4326
rect 7812 4324 7868 4326
rect 7572 3290 7628 3292
rect 7652 3290 7708 3292
rect 7732 3290 7788 3292
rect 7812 3290 7868 3292
rect 7572 3238 7618 3290
rect 7618 3238 7628 3290
rect 7652 3238 7682 3290
rect 7682 3238 7694 3290
rect 7694 3238 7708 3290
rect 7732 3238 7746 3290
rect 7746 3238 7758 3290
rect 7758 3238 7788 3290
rect 7812 3238 7822 3290
rect 7822 3238 7868 3290
rect 7572 3236 7628 3238
rect 7652 3236 7708 3238
rect 7732 3236 7788 3238
rect 7812 3236 7868 3238
rect 7572 2202 7628 2204
rect 7652 2202 7708 2204
rect 7732 2202 7788 2204
rect 7812 2202 7868 2204
rect 7572 2150 7618 2202
rect 7618 2150 7628 2202
rect 7652 2150 7682 2202
rect 7682 2150 7694 2202
rect 7694 2150 7708 2202
rect 7732 2150 7746 2202
rect 7746 2150 7758 2202
rect 7758 2150 7788 2202
rect 7812 2150 7822 2202
rect 7822 2150 7868 2202
rect 7572 2148 7628 2150
rect 7652 2148 7708 2150
rect 7732 2148 7788 2150
rect 7812 2148 7868 2150
rect 8114 2488 8170 2544
rect 8482 9560 8538 9616
rect 8666 10412 8668 10432
rect 8668 10412 8720 10432
rect 8720 10412 8722 10432
rect 8666 10376 8722 10412
rect 8390 3576 8446 3632
rect 9586 10548 9588 10568
rect 9588 10548 9640 10568
rect 9640 10548 9642 10568
rect 9586 10512 9642 10548
rect 8850 1672 8906 1728
rect 9402 6976 9458 7032
rect 9034 5616 9090 5672
rect 7572 1114 7628 1116
rect 7652 1114 7708 1116
rect 7732 1114 7788 1116
rect 7812 1114 7868 1116
rect 7572 1062 7618 1114
rect 7618 1062 7628 1114
rect 7652 1062 7682 1114
rect 7682 1062 7694 1114
rect 7694 1062 7708 1114
rect 7732 1062 7746 1114
rect 7746 1062 7758 1114
rect 7758 1062 7788 1114
rect 7812 1062 7822 1114
rect 7822 1062 7868 1114
rect 7572 1060 7628 1062
rect 7652 1060 7708 1062
rect 7732 1060 7788 1062
rect 7812 1060 7868 1062
rect 9310 5652 9312 5672
rect 9312 5652 9364 5672
rect 9364 5652 9366 5672
rect 9310 5616 9366 5652
rect 9586 9424 9642 9480
rect 9494 3576 9550 3632
rect 13818 11892 13874 11928
rect 13818 11872 13820 11892
rect 13820 11872 13872 11892
rect 13872 11872 13874 11892
rect 11058 9832 11114 9888
rect 10046 3712 10102 3768
rect 10138 2080 10194 2136
rect 22098 11056 22154 11112
rect 16578 6568 16634 6624
rect 16854 6160 16910 6216
rect 16578 5344 16634 5400
rect 16670 4936 16726 4992
rect 16762 4528 16818 4584
rect 16578 2488 16634 2544
rect 16946 5752 17002 5808
rect 22282 8200 22338 8256
rect 13818 892 13820 912
rect 13820 892 13872 912
rect 13872 892 13874 912
rect 13818 856 13874 892
rect 5072 570 5128 572
rect 5152 570 5208 572
rect 5232 570 5288 572
rect 5312 570 5368 572
rect 5072 518 5118 570
rect 5118 518 5128 570
rect 5152 518 5182 570
rect 5182 518 5194 570
rect 5194 518 5208 570
rect 5232 518 5246 570
rect 5246 518 5258 570
rect 5258 518 5288 570
rect 5312 518 5322 570
rect 5322 518 5368 570
rect 5072 516 5128 518
rect 5152 516 5208 518
rect 5232 516 5288 518
rect 5312 516 5368 518
rect 5446 448 5502 504
<< obsm2 >>
rect 24000 0 34000 13000
<< metal3 >>
rect 10041 12338 10107 12341
rect 14000 12338 34000 12368
rect 10041 12336 34000 12338
rect 10041 12280 10046 12336
rect 10102 12280 34000 12336
rect 10041 12278 34000 12280
rect 10041 12275 10107 12278
rect 14000 12248 34000 12278
rect 2562 12000 2878 12001
rect 2562 11936 2568 12000
rect 2632 11936 2648 12000
rect 2712 11936 2728 12000
rect 2792 11936 2808 12000
rect 2872 11936 2878 12000
rect 2562 11935 2878 11936
rect 7562 12000 7878 12001
rect 7562 11936 7568 12000
rect 7632 11936 7648 12000
rect 7712 11936 7728 12000
rect 7792 11936 7808 12000
rect 7872 11936 7878 12000
rect 7562 11935 7878 11936
rect 13813 11930 13879 11933
rect 14000 11930 34000 11960
rect 13813 11928 34000 11930
rect 13813 11872 13818 11928
rect 13874 11872 34000 11928
rect 13813 11870 34000 11872
rect 13813 11867 13879 11870
rect 14000 11840 34000 11870
rect 2497 11658 2563 11661
rect 2497 11656 12450 11658
rect 2497 11600 2502 11656
rect 2558 11600 12450 11656
rect 2497 11598 12450 11600
rect 2497 11595 2563 11598
rect 12390 11522 12450 11598
rect 14000 11522 34000 11552
rect 12390 11462 34000 11522
rect 5062 11456 5378 11457
rect 5062 11392 5068 11456
rect 5132 11392 5148 11456
rect 5212 11392 5228 11456
rect 5292 11392 5308 11456
rect 5372 11392 5378 11456
rect 14000 11432 34000 11462
rect 5062 11391 5378 11392
rect 3601 11250 3667 11253
rect 4470 11250 4476 11252
rect 3601 11248 4476 11250
rect 3601 11192 3606 11248
rect 3662 11192 4476 11248
rect 3601 11190 4476 11192
rect 3601 11187 3667 11190
rect 4470 11188 4476 11190
rect 4540 11188 4546 11252
rect 1393 11114 1459 11117
rect 4337 11114 4403 11117
rect 1393 11112 4403 11114
rect 1393 11056 1398 11112
rect 1454 11056 4342 11112
rect 4398 11056 4403 11112
rect 1393 11054 4403 11056
rect 1393 11051 1459 11054
rect 4337 11051 4403 11054
rect 14000 11112 34000 11144
rect 14000 11056 22098 11112
rect 22154 11056 34000 11112
rect 14000 11024 34000 11056
rect 2562 10912 2878 10913
rect 2562 10848 2568 10912
rect 2632 10848 2648 10912
rect 2712 10848 2728 10912
rect 2792 10848 2808 10912
rect 2872 10848 2878 10912
rect 2562 10847 2878 10848
rect 7562 10912 7878 10913
rect 7562 10848 7568 10912
rect 7632 10848 7648 10912
rect 7712 10848 7728 10912
rect 7792 10848 7808 10912
rect 7872 10848 7878 10912
rect 7562 10847 7878 10848
rect 3325 10842 3391 10845
rect 7189 10842 7255 10845
rect 3325 10840 7255 10842
rect 3325 10784 3330 10840
rect 3386 10784 7194 10840
rect 7250 10784 7255 10840
rect 3325 10782 7255 10784
rect 3325 10779 3391 10782
rect 7189 10779 7255 10782
rect 2773 10706 2839 10709
rect 6913 10706 6979 10709
rect 14000 10706 34000 10736
rect 2773 10704 5412 10706
rect 2773 10648 2778 10704
rect 2834 10648 5412 10704
rect 2773 10646 5412 10648
rect 2773 10643 2839 10646
rect 5352 10573 5412 10646
rect 6913 10704 34000 10706
rect 6913 10648 6918 10704
rect 6974 10648 34000 10704
rect 6913 10646 34000 10648
rect 6913 10643 6979 10646
rect 14000 10616 34000 10646
rect 3049 10572 3115 10573
rect 2998 10570 3004 10572
rect 2958 10510 3004 10570
rect 3068 10568 3115 10572
rect 3110 10512 3115 10568
rect 2998 10508 3004 10510
rect 3068 10508 3115 10512
rect 3049 10507 3115 10508
rect 5349 10570 5415 10573
rect 5533 10570 5599 10573
rect 9581 10570 9647 10573
rect 5349 10568 9647 10570
rect 5349 10512 5354 10568
rect 5410 10512 5538 10568
rect 5594 10512 9586 10568
rect 9642 10512 9647 10568
rect 5349 10510 9647 10512
rect 5349 10507 5415 10510
rect 5533 10507 5599 10510
rect 9581 10507 9647 10510
rect 6085 10434 6151 10437
rect 8661 10434 8727 10437
rect 6085 10432 8727 10434
rect 6085 10376 6090 10432
rect 6146 10376 8666 10432
rect 8722 10376 8727 10432
rect 6085 10374 8727 10376
rect 6085 10371 6151 10374
rect 8661 10371 8727 10374
rect 5062 10368 5378 10369
rect 5062 10304 5068 10368
rect 5132 10304 5148 10368
rect 5212 10304 5228 10368
rect 5292 10304 5308 10368
rect 5372 10304 5378 10368
rect 5062 10303 5378 10304
rect 5441 10298 5507 10301
rect 14000 10298 34000 10328
rect 5441 10296 34000 10298
rect 5441 10240 5446 10296
rect 5502 10240 34000 10296
rect 5441 10238 34000 10240
rect 5441 10235 5507 10238
rect 14000 10208 34000 10238
rect 2865 10026 2931 10029
rect 2865 10024 3066 10026
rect 2865 9968 2870 10024
rect 2926 9968 3066 10024
rect 2865 9966 3066 9968
rect 2865 9963 2931 9966
rect 3006 9893 3066 9966
rect 2957 9888 3066 9893
rect 2957 9832 2962 9888
rect 3018 9832 3066 9888
rect 2957 9830 3066 9832
rect 11053 9890 11119 9893
rect 14000 9890 34000 9920
rect 11053 9888 34000 9890
rect 11053 9832 11058 9888
rect 11114 9832 34000 9888
rect 11053 9830 34000 9832
rect 2957 9827 3023 9830
rect 11053 9827 11119 9830
rect 2562 9824 2878 9825
rect 2562 9760 2568 9824
rect 2632 9760 2648 9824
rect 2712 9760 2728 9824
rect 2792 9760 2808 9824
rect 2872 9760 2878 9824
rect 2562 9759 2878 9760
rect 7562 9824 7878 9825
rect 7562 9760 7568 9824
rect 7632 9760 7648 9824
rect 7712 9760 7728 9824
rect 7792 9760 7808 9824
rect 7872 9760 7878 9824
rect 14000 9800 34000 9830
rect 7562 9759 7878 9760
rect 4838 9556 4844 9620
rect 4908 9618 4914 9620
rect 5349 9618 5415 9621
rect 4908 9616 5415 9618
rect 4908 9560 5354 9616
rect 5410 9560 5415 9616
rect 4908 9558 5415 9560
rect 4908 9556 4914 9558
rect 5349 9555 5415 9558
rect 5809 9618 5875 9621
rect 8477 9618 8543 9621
rect 5809 9616 8543 9618
rect 5809 9560 5814 9616
rect 5870 9560 8482 9616
rect 8538 9560 8543 9616
rect 5809 9558 8543 9560
rect 5809 9555 5875 9558
rect 8477 9555 8543 9558
rect 2773 9482 2839 9485
rect 4889 9482 4955 9485
rect 7557 9482 7623 9485
rect 2773 9480 7623 9482
rect 2773 9424 2778 9480
rect 2834 9424 4894 9480
rect 4950 9424 7562 9480
rect 7618 9424 7623 9480
rect 2773 9422 7623 9424
rect 2773 9419 2839 9422
rect 4889 9419 4955 9422
rect 7557 9419 7623 9422
rect 9581 9482 9647 9485
rect 14000 9482 34000 9512
rect 9581 9480 34000 9482
rect 9581 9424 9586 9480
rect 9642 9424 34000 9480
rect 9581 9422 34000 9424
rect 9581 9419 9647 9422
rect 14000 9392 34000 9422
rect 1209 9346 1275 9349
rect 4797 9346 4863 9349
rect 1209 9344 4863 9346
rect 1209 9288 1214 9344
rect 1270 9288 4802 9344
rect 4858 9288 4863 9344
rect 1209 9286 4863 9288
rect 1209 9283 1275 9286
rect 4797 9283 4863 9286
rect 6545 9346 6611 9349
rect 6729 9346 6795 9349
rect 6545 9344 6795 9346
rect 6545 9288 6550 9344
rect 6606 9288 6734 9344
rect 6790 9288 6795 9344
rect 6545 9286 6795 9288
rect 6545 9283 6611 9286
rect 6729 9283 6795 9286
rect 5062 9280 5378 9281
rect 5062 9216 5068 9280
rect 5132 9216 5148 9280
rect 5212 9216 5228 9280
rect 5292 9216 5308 9280
rect 5372 9216 5378 9280
rect 5062 9215 5378 9216
rect 3785 9074 3851 9077
rect 14000 9074 34000 9104
rect 3785 9072 34000 9074
rect 3785 9016 3790 9072
rect 3846 9016 34000 9072
rect 3785 9014 34000 9016
rect 3785 9011 3851 9014
rect 14000 8984 34000 9014
rect 4245 8938 4311 8941
rect 7097 8938 7163 8941
rect 7465 8938 7531 8941
rect 4245 8936 7531 8938
rect 4245 8880 4250 8936
rect 4306 8880 7102 8936
rect 7158 8880 7470 8936
rect 7526 8880 7531 8936
rect 4245 8878 7531 8880
rect 4245 8875 4311 8878
rect 7097 8875 7163 8878
rect 7465 8875 7531 8878
rect 5717 8802 5783 8805
rect 7189 8802 7255 8805
rect 5717 8800 7255 8802
rect 5717 8744 5722 8800
rect 5778 8744 7194 8800
rect 7250 8744 7255 8800
rect 5717 8742 7255 8744
rect 5717 8739 5783 8742
rect 7189 8739 7255 8742
rect 2562 8736 2878 8737
rect 2562 8672 2568 8736
rect 2632 8672 2648 8736
rect 2712 8672 2728 8736
rect 2792 8672 2808 8736
rect 2872 8672 2878 8736
rect 2562 8671 2878 8672
rect 7562 8736 7878 8737
rect 7562 8672 7568 8736
rect 7632 8672 7648 8736
rect 7712 8672 7728 8736
rect 7792 8672 7808 8736
rect 7872 8672 7878 8736
rect 7562 8671 7878 8672
rect 3877 8666 3943 8669
rect 4245 8666 4311 8669
rect 3877 8664 4311 8666
rect 3877 8608 3882 8664
rect 3938 8608 4250 8664
rect 4306 8608 4311 8664
rect 3877 8606 4311 8608
rect 3877 8603 3943 8606
rect 4245 8603 4311 8606
rect 5758 8604 5764 8668
rect 5828 8666 5834 8668
rect 5993 8666 6059 8669
rect 5828 8664 6059 8666
rect 5828 8608 5998 8664
rect 6054 8608 6059 8664
rect 5828 8606 6059 8608
rect 5828 8604 5834 8606
rect 5993 8603 6059 8606
rect 8201 8666 8267 8669
rect 14000 8666 34000 8696
rect 8201 8664 34000 8666
rect 8201 8608 8206 8664
rect 8262 8608 34000 8664
rect 8201 8606 34000 8608
rect 8201 8603 8267 8606
rect 14000 8576 34000 8606
rect 2129 8530 2195 8533
rect 5625 8530 5691 8533
rect 2129 8528 5691 8530
rect 2129 8472 2134 8528
rect 2190 8472 5630 8528
rect 5686 8472 5691 8528
rect 2129 8470 5691 8472
rect 2129 8467 2195 8470
rect 5625 8467 5691 8470
rect 3325 8394 3391 8397
rect 3877 8394 3943 8397
rect 3325 8392 3943 8394
rect 3325 8336 3330 8392
rect 3386 8336 3882 8392
rect 3938 8336 3943 8392
rect 3325 8334 3943 8336
rect 3325 8331 3391 8334
rect 3877 8331 3943 8334
rect 1301 8258 1367 8261
rect 4429 8258 4495 8261
rect 1301 8256 4495 8258
rect 1301 8200 1306 8256
rect 1362 8200 4434 8256
rect 4490 8200 4495 8256
rect 1301 8198 4495 8200
rect 1301 8195 1367 8198
rect 4429 8195 4495 8198
rect 14000 8256 34000 8288
rect 14000 8200 22282 8256
rect 22338 8200 34000 8256
rect 5062 8192 5378 8193
rect 5062 8128 5068 8192
rect 5132 8128 5148 8192
rect 5212 8128 5228 8192
rect 5292 8128 5308 8192
rect 5372 8128 5378 8192
rect 14000 8168 34000 8200
rect 5062 8127 5378 8128
rect 2497 7850 2563 7853
rect 14000 7850 34000 7880
rect 2497 7848 34000 7850
rect 2497 7792 2502 7848
rect 2558 7792 34000 7848
rect 2497 7790 34000 7792
rect 2497 7787 2563 7790
rect 14000 7760 34000 7790
rect 2562 7648 2878 7649
rect 2562 7584 2568 7648
rect 2632 7584 2648 7648
rect 2712 7584 2728 7648
rect 2792 7584 2808 7648
rect 2872 7584 2878 7648
rect 2562 7583 2878 7584
rect 7562 7648 7878 7649
rect 7562 7584 7568 7648
rect 7632 7584 7648 7648
rect 7712 7584 7728 7648
rect 7792 7584 7808 7648
rect 7872 7584 7878 7648
rect 7562 7583 7878 7584
rect 5441 7442 5507 7445
rect 14000 7442 34000 7472
rect 5441 7440 34000 7442
rect 5441 7384 5446 7440
rect 5502 7384 34000 7440
rect 5441 7382 34000 7384
rect 5441 7379 5507 7382
rect 14000 7352 34000 7382
rect 4061 7306 4127 7309
rect 4061 7304 5504 7306
rect 4061 7248 4066 7304
rect 4122 7248 5504 7304
rect 4061 7246 5504 7248
rect 4061 7243 4127 7246
rect 5444 7173 5504 7246
rect 5441 7170 5507 7173
rect 5809 7170 5875 7173
rect 5441 7168 5875 7170
rect 5441 7112 5446 7168
rect 5502 7112 5814 7168
rect 5870 7112 5875 7168
rect 5441 7110 5875 7112
rect 5441 7107 5507 7110
rect 5809 7107 5875 7110
rect 5062 7104 5378 7105
rect 5062 7040 5068 7104
rect 5132 7040 5148 7104
rect 5212 7040 5228 7104
rect 5292 7040 5308 7104
rect 5372 7040 5378 7104
rect 5062 7039 5378 7040
rect 9397 7034 9463 7037
rect 14000 7034 34000 7064
rect 9397 7032 34000 7034
rect 9397 6976 9402 7032
rect 9458 6976 34000 7032
rect 9397 6974 34000 6976
rect 9397 6971 9463 6974
rect 14000 6944 34000 6974
rect 4245 6898 4311 6901
rect 7097 6898 7163 6901
rect 4245 6896 7163 6898
rect 4245 6840 4250 6896
rect 4306 6840 7102 6896
rect 7158 6840 7163 6896
rect 4245 6838 7163 6840
rect 4245 6835 4311 6838
rect 7097 6835 7163 6838
rect 3877 6762 3943 6765
rect 4061 6762 4127 6765
rect 3877 6760 4127 6762
rect 3877 6704 3882 6760
rect 3938 6704 4066 6760
rect 4122 6704 4127 6760
rect 3877 6702 4127 6704
rect 3877 6699 3943 6702
rect 4061 6699 4127 6702
rect 4470 6700 4476 6764
rect 4540 6762 4546 6764
rect 5574 6762 5580 6764
rect 4540 6702 5580 6762
rect 4540 6700 4546 6702
rect 5574 6700 5580 6702
rect 5644 6762 5650 6764
rect 6545 6762 6611 6765
rect 5644 6760 6611 6762
rect 5644 6704 6550 6760
rect 6606 6704 6611 6760
rect 5644 6702 6611 6704
rect 5644 6700 5650 6702
rect 6545 6699 6611 6702
rect 5717 6628 5783 6629
rect 5717 6624 5764 6628
rect 5828 6626 5834 6628
rect 5717 6568 5722 6624
rect 5717 6564 5764 6568
rect 5828 6566 5874 6626
rect 14000 6624 34000 6656
rect 14000 6568 16578 6624
rect 16634 6568 34000 6624
rect 5828 6564 5834 6566
rect 5717 6563 5783 6564
rect 2562 6560 2878 6561
rect 2562 6496 2568 6560
rect 2632 6496 2648 6560
rect 2712 6496 2728 6560
rect 2792 6496 2808 6560
rect 2872 6496 2878 6560
rect 2562 6495 2878 6496
rect 7562 6560 7878 6561
rect 7562 6496 7568 6560
rect 7632 6496 7648 6560
rect 7712 6496 7728 6560
rect 7792 6496 7808 6560
rect 7872 6496 7878 6560
rect 14000 6536 34000 6568
rect 7562 6495 7878 6496
rect 2773 6354 2839 6357
rect 2998 6354 3004 6356
rect 2773 6352 3004 6354
rect 2773 6296 2778 6352
rect 2834 6296 3004 6352
rect 2773 6294 3004 6296
rect 2773 6291 2839 6294
rect 2998 6292 3004 6294
rect 3068 6354 3074 6356
rect 4153 6354 4219 6357
rect 3068 6352 4219 6354
rect 3068 6296 4158 6352
rect 4214 6296 4219 6352
rect 3068 6294 4219 6296
rect 3068 6292 3074 6294
rect 4153 6291 4219 6294
rect 14000 6216 34000 6248
rect 14000 6160 16854 6216
rect 16910 6160 34000 6216
rect 14000 6128 34000 6160
rect 5062 6016 5378 6017
rect 5062 5952 5068 6016
rect 5132 5952 5148 6016
rect 5212 5952 5228 6016
rect 5292 5952 5308 6016
rect 5372 5952 5378 6016
rect 5062 5951 5378 5952
rect 14000 5808 34000 5840
rect 14000 5752 16946 5808
rect 17002 5752 34000 5808
rect 14000 5720 34000 5752
rect 9029 5674 9095 5677
rect 9305 5674 9371 5677
rect 9029 5672 9371 5674
rect 9029 5616 9034 5672
rect 9090 5616 9310 5672
rect 9366 5616 9371 5672
rect 9029 5614 9371 5616
rect 9029 5611 9095 5614
rect 9305 5611 9371 5614
rect 2562 5472 2878 5473
rect 2562 5408 2568 5472
rect 2632 5408 2648 5472
rect 2712 5408 2728 5472
rect 2792 5408 2808 5472
rect 2872 5408 2878 5472
rect 2562 5407 2878 5408
rect 7562 5472 7878 5473
rect 7562 5408 7568 5472
rect 7632 5408 7648 5472
rect 7712 5408 7728 5472
rect 7792 5408 7808 5472
rect 7872 5408 7878 5472
rect 7562 5407 7878 5408
rect 14000 5400 34000 5432
rect 14000 5344 16578 5400
rect 16634 5344 34000 5400
rect 14000 5312 34000 5344
rect 14000 4992 34000 5024
rect 14000 4936 16670 4992
rect 16726 4936 34000 4992
rect 5062 4928 5378 4929
rect 5062 4864 5068 4928
rect 5132 4864 5148 4928
rect 5212 4864 5228 4928
rect 5292 4864 5308 4928
rect 5372 4864 5378 4928
rect 14000 4904 34000 4936
rect 5062 4863 5378 4864
rect 14000 4584 34000 4616
rect 14000 4528 16762 4584
rect 16818 4528 34000 4584
rect 14000 4496 34000 4528
rect 7562 4384 7878 4385
rect 7562 4320 7568 4384
rect 7632 4320 7648 4384
rect 7712 4320 7728 4384
rect 7792 4320 7808 4384
rect 7872 4320 7878 4384
rect 7562 4319 7878 4320
rect 4838 4116 4844 4180
rect 4908 4178 4914 4180
rect 5349 4178 5415 4181
rect 4908 4176 5415 4178
rect 4908 4120 5354 4176
rect 5410 4120 5415 4176
rect 4908 4118 5415 4120
rect 4908 4116 4914 4118
rect 5349 4115 5415 4118
rect 6821 4178 6887 4181
rect 14000 4178 34000 4208
rect 6821 4176 34000 4178
rect 6821 4120 6826 4176
rect 6882 4120 34000 4176
rect 6821 4118 34000 4120
rect 6821 4115 6887 4118
rect 14000 4088 34000 4118
rect 5533 3908 5599 3909
rect 5533 3904 5580 3908
rect 5644 3906 5650 3908
rect 5533 3848 5538 3904
rect 5533 3844 5580 3848
rect 5644 3846 5690 3906
rect 5644 3844 5650 3846
rect 5533 3843 5599 3844
rect 5062 3840 5378 3841
rect 5062 3776 5068 3840
rect 5132 3776 5148 3840
rect 5212 3776 5228 3840
rect 5292 3776 5308 3840
rect 5372 3776 5378 3840
rect 5062 3775 5378 3776
rect 10041 3770 10107 3773
rect 14000 3770 34000 3800
rect 10041 3768 34000 3770
rect 10041 3712 10046 3768
rect 10102 3712 34000 3768
rect 10041 3710 34000 3712
rect 10041 3707 10107 3710
rect 14000 3680 34000 3710
rect 7097 3634 7163 3637
rect 8385 3634 8451 3637
rect 9489 3634 9555 3637
rect 7097 3632 9555 3634
rect 7097 3576 7102 3632
rect 7158 3576 8390 3632
rect 8446 3576 9494 3632
rect 9550 3576 9555 3632
rect 7097 3574 9555 3576
rect 7097 3571 7163 3574
rect 8385 3571 8451 3574
rect 9489 3571 9555 3574
rect 5073 3498 5139 3501
rect 5073 3496 12450 3498
rect 5073 3440 5078 3496
rect 5134 3440 12450 3496
rect 5073 3438 12450 3440
rect 5073 3435 5139 3438
rect 2681 3430 2747 3433
rect 2484 3428 2747 3430
rect 2484 3372 2686 3428
rect 2742 3372 2747 3428
rect 2484 3370 2747 3372
rect 2681 3367 2747 3370
rect 12390 3362 12450 3438
rect 14000 3362 34000 3392
rect 12390 3302 34000 3362
rect 7562 3296 7878 3297
rect 7562 3232 7568 3296
rect 7632 3232 7648 3296
rect 7712 3232 7728 3296
rect 7792 3232 7808 3296
rect 7872 3232 7878 3296
rect 14000 3272 34000 3302
rect 7562 3231 7878 3232
rect 6821 2954 6887 2957
rect 14000 2954 34000 2984
rect 6821 2952 34000 2954
rect 6821 2896 6826 2952
rect 6882 2896 34000 2952
rect 6821 2894 34000 2896
rect 6821 2891 6887 2894
rect 14000 2864 34000 2894
rect 5062 2752 5378 2753
rect 5062 2688 5068 2752
rect 5132 2688 5148 2752
rect 5212 2688 5228 2752
rect 5292 2688 5308 2752
rect 5372 2688 5378 2752
rect 5062 2687 5378 2688
rect 3785 2546 3851 2549
rect 4838 2546 4844 2548
rect 3785 2544 4844 2546
rect 3785 2488 3790 2544
rect 3846 2488 4844 2544
rect 3785 2486 4844 2488
rect 3785 2483 3851 2486
rect 4838 2484 4844 2486
rect 4908 2546 4914 2548
rect 8109 2546 8175 2549
rect 4908 2544 8175 2546
rect 4908 2488 8114 2544
rect 8170 2488 8175 2544
rect 4908 2486 8175 2488
rect 4908 2484 4914 2486
rect 8109 2483 8175 2486
rect 14000 2544 34000 2576
rect 14000 2488 16578 2544
rect 16634 2488 34000 2544
rect 14000 2456 34000 2488
rect 7562 2208 7878 2209
rect 7562 2144 7568 2208
rect 7632 2144 7648 2208
rect 7712 2144 7728 2208
rect 7792 2144 7808 2208
rect 7872 2144 7878 2208
rect 7562 2143 7878 2144
rect 10133 2138 10199 2141
rect 14000 2138 34000 2168
rect 10133 2136 34000 2138
rect 10133 2080 10138 2136
rect 10194 2080 34000 2136
rect 10133 2078 34000 2080
rect 10133 2075 10199 2078
rect 14000 2048 34000 2078
rect 8845 1730 8911 1733
rect 14000 1730 34000 1760
rect 8845 1728 34000 1730
rect 8845 1672 8850 1728
rect 8906 1672 34000 1728
rect 8845 1670 34000 1672
rect 8845 1667 8911 1670
rect 5062 1664 5378 1665
rect 5062 1600 5068 1664
rect 5132 1600 5148 1664
rect 5212 1600 5228 1664
rect 5292 1600 5308 1664
rect 5372 1600 5378 1664
rect 14000 1640 34000 1670
rect 5062 1599 5378 1600
rect 5441 1322 5507 1325
rect 14000 1322 34000 1352
rect 5441 1320 34000 1322
rect 5441 1264 5446 1320
rect 5502 1264 34000 1320
rect 5441 1262 34000 1264
rect 5441 1259 5507 1262
rect 14000 1232 34000 1262
rect 2562 1120 2878 1121
rect 2562 1056 2568 1120
rect 2632 1056 2648 1120
rect 2712 1056 2728 1120
rect 2792 1056 2808 1120
rect 2872 1056 2878 1120
rect 2562 1055 2878 1056
rect 7562 1120 7878 1121
rect 7562 1056 7568 1120
rect 7632 1056 7648 1120
rect 7712 1056 7728 1120
rect 7792 1056 7808 1120
rect 7872 1056 7878 1120
rect 7562 1055 7878 1056
rect 13813 914 13879 917
rect 14000 914 34000 944
rect 13813 912 34000 914
rect 13813 856 13818 912
rect 13874 856 34000 912
rect 13813 854 34000 856
rect 13813 851 13879 854
rect 14000 824 34000 854
rect 5062 576 5378 577
rect 5062 512 5068 576
rect 5132 512 5148 576
rect 5212 512 5228 576
rect 5292 512 5308 576
rect 5372 512 5378 576
rect 5062 511 5378 512
rect 5441 506 5507 509
rect 14000 506 34000 536
rect 5441 504 34000 506
rect 5441 448 5446 504
rect 5502 448 34000 504
rect 5441 446 34000 448
rect 5441 443 5507 446
rect 14000 416 34000 446
<< via3 >>
rect 2568 11996 2632 12000
rect 2568 11940 2572 11996
rect 2572 11940 2628 11996
rect 2628 11940 2632 11996
rect 2568 11936 2632 11940
rect 2648 11996 2712 12000
rect 2648 11940 2652 11996
rect 2652 11940 2708 11996
rect 2708 11940 2712 11996
rect 2648 11936 2712 11940
rect 2728 11996 2792 12000
rect 2728 11940 2732 11996
rect 2732 11940 2788 11996
rect 2788 11940 2792 11996
rect 2728 11936 2792 11940
rect 2808 11996 2872 12000
rect 2808 11940 2812 11996
rect 2812 11940 2868 11996
rect 2868 11940 2872 11996
rect 2808 11936 2872 11940
rect 7568 11996 7632 12000
rect 7568 11940 7572 11996
rect 7572 11940 7628 11996
rect 7628 11940 7632 11996
rect 7568 11936 7632 11940
rect 7648 11996 7712 12000
rect 7648 11940 7652 11996
rect 7652 11940 7708 11996
rect 7708 11940 7712 11996
rect 7648 11936 7712 11940
rect 7728 11996 7792 12000
rect 7728 11940 7732 11996
rect 7732 11940 7788 11996
rect 7788 11940 7792 11996
rect 7728 11936 7792 11940
rect 7808 11996 7872 12000
rect 7808 11940 7812 11996
rect 7812 11940 7868 11996
rect 7868 11940 7872 11996
rect 7808 11936 7872 11940
rect 5068 11452 5132 11456
rect 5068 11396 5072 11452
rect 5072 11396 5128 11452
rect 5128 11396 5132 11452
rect 5068 11392 5132 11396
rect 5148 11452 5212 11456
rect 5148 11396 5152 11452
rect 5152 11396 5208 11452
rect 5208 11396 5212 11452
rect 5148 11392 5212 11396
rect 5228 11452 5292 11456
rect 5228 11396 5232 11452
rect 5232 11396 5288 11452
rect 5288 11396 5292 11452
rect 5228 11392 5292 11396
rect 5308 11452 5372 11456
rect 5308 11396 5312 11452
rect 5312 11396 5368 11452
rect 5368 11396 5372 11452
rect 5308 11392 5372 11396
rect 4476 11188 4540 11252
rect 2568 10908 2632 10912
rect 2568 10852 2572 10908
rect 2572 10852 2628 10908
rect 2628 10852 2632 10908
rect 2568 10848 2632 10852
rect 2648 10908 2712 10912
rect 2648 10852 2652 10908
rect 2652 10852 2708 10908
rect 2708 10852 2712 10908
rect 2648 10848 2712 10852
rect 2728 10908 2792 10912
rect 2728 10852 2732 10908
rect 2732 10852 2788 10908
rect 2788 10852 2792 10908
rect 2728 10848 2792 10852
rect 2808 10908 2872 10912
rect 2808 10852 2812 10908
rect 2812 10852 2868 10908
rect 2868 10852 2872 10908
rect 2808 10848 2872 10852
rect 7568 10908 7632 10912
rect 7568 10852 7572 10908
rect 7572 10852 7628 10908
rect 7628 10852 7632 10908
rect 7568 10848 7632 10852
rect 7648 10908 7712 10912
rect 7648 10852 7652 10908
rect 7652 10852 7708 10908
rect 7708 10852 7712 10908
rect 7648 10848 7712 10852
rect 7728 10908 7792 10912
rect 7728 10852 7732 10908
rect 7732 10852 7788 10908
rect 7788 10852 7792 10908
rect 7728 10848 7792 10852
rect 7808 10908 7872 10912
rect 7808 10852 7812 10908
rect 7812 10852 7868 10908
rect 7868 10852 7872 10908
rect 7808 10848 7872 10852
rect 3004 10568 3068 10572
rect 3004 10512 3054 10568
rect 3054 10512 3068 10568
rect 3004 10508 3068 10512
rect 5068 10364 5132 10368
rect 5068 10308 5072 10364
rect 5072 10308 5128 10364
rect 5128 10308 5132 10364
rect 5068 10304 5132 10308
rect 5148 10364 5212 10368
rect 5148 10308 5152 10364
rect 5152 10308 5208 10364
rect 5208 10308 5212 10364
rect 5148 10304 5212 10308
rect 5228 10364 5292 10368
rect 5228 10308 5232 10364
rect 5232 10308 5288 10364
rect 5288 10308 5292 10364
rect 5228 10304 5292 10308
rect 5308 10364 5372 10368
rect 5308 10308 5312 10364
rect 5312 10308 5368 10364
rect 5368 10308 5372 10364
rect 5308 10304 5372 10308
rect 2568 9820 2632 9824
rect 2568 9764 2572 9820
rect 2572 9764 2628 9820
rect 2628 9764 2632 9820
rect 2568 9760 2632 9764
rect 2648 9820 2712 9824
rect 2648 9764 2652 9820
rect 2652 9764 2708 9820
rect 2708 9764 2712 9820
rect 2648 9760 2712 9764
rect 2728 9820 2792 9824
rect 2728 9764 2732 9820
rect 2732 9764 2788 9820
rect 2788 9764 2792 9820
rect 2728 9760 2792 9764
rect 2808 9820 2872 9824
rect 2808 9764 2812 9820
rect 2812 9764 2868 9820
rect 2868 9764 2872 9820
rect 2808 9760 2872 9764
rect 7568 9820 7632 9824
rect 7568 9764 7572 9820
rect 7572 9764 7628 9820
rect 7628 9764 7632 9820
rect 7568 9760 7632 9764
rect 7648 9820 7712 9824
rect 7648 9764 7652 9820
rect 7652 9764 7708 9820
rect 7708 9764 7712 9820
rect 7648 9760 7712 9764
rect 7728 9820 7792 9824
rect 7728 9764 7732 9820
rect 7732 9764 7788 9820
rect 7788 9764 7792 9820
rect 7728 9760 7792 9764
rect 7808 9820 7872 9824
rect 7808 9764 7812 9820
rect 7812 9764 7868 9820
rect 7868 9764 7872 9820
rect 7808 9760 7872 9764
rect 4844 9556 4908 9620
rect 5068 9276 5132 9280
rect 5068 9220 5072 9276
rect 5072 9220 5128 9276
rect 5128 9220 5132 9276
rect 5068 9216 5132 9220
rect 5148 9276 5212 9280
rect 5148 9220 5152 9276
rect 5152 9220 5208 9276
rect 5208 9220 5212 9276
rect 5148 9216 5212 9220
rect 5228 9276 5292 9280
rect 5228 9220 5232 9276
rect 5232 9220 5288 9276
rect 5288 9220 5292 9276
rect 5228 9216 5292 9220
rect 5308 9276 5372 9280
rect 5308 9220 5312 9276
rect 5312 9220 5368 9276
rect 5368 9220 5372 9276
rect 5308 9216 5372 9220
rect 2568 8732 2632 8736
rect 2568 8676 2572 8732
rect 2572 8676 2628 8732
rect 2628 8676 2632 8732
rect 2568 8672 2632 8676
rect 2648 8732 2712 8736
rect 2648 8676 2652 8732
rect 2652 8676 2708 8732
rect 2708 8676 2712 8732
rect 2648 8672 2712 8676
rect 2728 8732 2792 8736
rect 2728 8676 2732 8732
rect 2732 8676 2788 8732
rect 2788 8676 2792 8732
rect 2728 8672 2792 8676
rect 2808 8732 2872 8736
rect 2808 8676 2812 8732
rect 2812 8676 2868 8732
rect 2868 8676 2872 8732
rect 2808 8672 2872 8676
rect 7568 8732 7632 8736
rect 7568 8676 7572 8732
rect 7572 8676 7628 8732
rect 7628 8676 7632 8732
rect 7568 8672 7632 8676
rect 7648 8732 7712 8736
rect 7648 8676 7652 8732
rect 7652 8676 7708 8732
rect 7708 8676 7712 8732
rect 7648 8672 7712 8676
rect 7728 8732 7792 8736
rect 7728 8676 7732 8732
rect 7732 8676 7788 8732
rect 7788 8676 7792 8732
rect 7728 8672 7792 8676
rect 7808 8732 7872 8736
rect 7808 8676 7812 8732
rect 7812 8676 7868 8732
rect 7868 8676 7872 8732
rect 7808 8672 7872 8676
rect 5764 8604 5828 8668
rect 5068 8188 5132 8192
rect 5068 8132 5072 8188
rect 5072 8132 5128 8188
rect 5128 8132 5132 8188
rect 5068 8128 5132 8132
rect 5148 8188 5212 8192
rect 5148 8132 5152 8188
rect 5152 8132 5208 8188
rect 5208 8132 5212 8188
rect 5148 8128 5212 8132
rect 5228 8188 5292 8192
rect 5228 8132 5232 8188
rect 5232 8132 5288 8188
rect 5288 8132 5292 8188
rect 5228 8128 5292 8132
rect 5308 8188 5372 8192
rect 5308 8132 5312 8188
rect 5312 8132 5368 8188
rect 5368 8132 5372 8188
rect 5308 8128 5372 8132
rect 2568 7644 2632 7648
rect 2568 7588 2572 7644
rect 2572 7588 2628 7644
rect 2628 7588 2632 7644
rect 2568 7584 2632 7588
rect 2648 7644 2712 7648
rect 2648 7588 2652 7644
rect 2652 7588 2708 7644
rect 2708 7588 2712 7644
rect 2648 7584 2712 7588
rect 2728 7644 2792 7648
rect 2728 7588 2732 7644
rect 2732 7588 2788 7644
rect 2788 7588 2792 7644
rect 2728 7584 2792 7588
rect 2808 7644 2872 7648
rect 2808 7588 2812 7644
rect 2812 7588 2868 7644
rect 2868 7588 2872 7644
rect 2808 7584 2872 7588
rect 7568 7644 7632 7648
rect 7568 7588 7572 7644
rect 7572 7588 7628 7644
rect 7628 7588 7632 7644
rect 7568 7584 7632 7588
rect 7648 7644 7712 7648
rect 7648 7588 7652 7644
rect 7652 7588 7708 7644
rect 7708 7588 7712 7644
rect 7648 7584 7712 7588
rect 7728 7644 7792 7648
rect 7728 7588 7732 7644
rect 7732 7588 7788 7644
rect 7788 7588 7792 7644
rect 7728 7584 7792 7588
rect 7808 7644 7872 7648
rect 7808 7588 7812 7644
rect 7812 7588 7868 7644
rect 7868 7588 7872 7644
rect 7808 7584 7872 7588
rect 5068 7100 5132 7104
rect 5068 7044 5072 7100
rect 5072 7044 5128 7100
rect 5128 7044 5132 7100
rect 5068 7040 5132 7044
rect 5148 7100 5212 7104
rect 5148 7044 5152 7100
rect 5152 7044 5208 7100
rect 5208 7044 5212 7100
rect 5148 7040 5212 7044
rect 5228 7100 5292 7104
rect 5228 7044 5232 7100
rect 5232 7044 5288 7100
rect 5288 7044 5292 7100
rect 5228 7040 5292 7044
rect 5308 7100 5372 7104
rect 5308 7044 5312 7100
rect 5312 7044 5368 7100
rect 5368 7044 5372 7100
rect 5308 7040 5372 7044
rect 4476 6700 4540 6764
rect 5580 6700 5644 6764
rect 5764 6624 5828 6628
rect 5764 6568 5778 6624
rect 5778 6568 5828 6624
rect 5764 6564 5828 6568
rect 2568 6556 2632 6560
rect 2568 6500 2572 6556
rect 2572 6500 2628 6556
rect 2628 6500 2632 6556
rect 2568 6496 2632 6500
rect 2648 6556 2712 6560
rect 2648 6500 2652 6556
rect 2652 6500 2708 6556
rect 2708 6500 2712 6556
rect 2648 6496 2712 6500
rect 2728 6556 2792 6560
rect 2728 6500 2732 6556
rect 2732 6500 2788 6556
rect 2788 6500 2792 6556
rect 2728 6496 2792 6500
rect 2808 6556 2872 6560
rect 2808 6500 2812 6556
rect 2812 6500 2868 6556
rect 2868 6500 2872 6556
rect 2808 6496 2872 6500
rect 7568 6556 7632 6560
rect 7568 6500 7572 6556
rect 7572 6500 7628 6556
rect 7628 6500 7632 6556
rect 7568 6496 7632 6500
rect 7648 6556 7712 6560
rect 7648 6500 7652 6556
rect 7652 6500 7708 6556
rect 7708 6500 7712 6556
rect 7648 6496 7712 6500
rect 7728 6556 7792 6560
rect 7728 6500 7732 6556
rect 7732 6500 7788 6556
rect 7788 6500 7792 6556
rect 7728 6496 7792 6500
rect 7808 6556 7872 6560
rect 7808 6500 7812 6556
rect 7812 6500 7868 6556
rect 7868 6500 7872 6556
rect 7808 6496 7872 6500
rect 3004 6292 3068 6356
rect 5068 6012 5132 6016
rect 5068 5956 5072 6012
rect 5072 5956 5128 6012
rect 5128 5956 5132 6012
rect 5068 5952 5132 5956
rect 5148 6012 5212 6016
rect 5148 5956 5152 6012
rect 5152 5956 5208 6012
rect 5208 5956 5212 6012
rect 5148 5952 5212 5956
rect 5228 6012 5292 6016
rect 5228 5956 5232 6012
rect 5232 5956 5288 6012
rect 5288 5956 5292 6012
rect 5228 5952 5292 5956
rect 5308 6012 5372 6016
rect 5308 5956 5312 6012
rect 5312 5956 5368 6012
rect 5368 5956 5372 6012
rect 5308 5952 5372 5956
rect 2568 5468 2632 5472
rect 2568 5412 2572 5468
rect 2572 5412 2628 5468
rect 2628 5412 2632 5468
rect 2568 5408 2632 5412
rect 2648 5468 2712 5472
rect 2648 5412 2652 5468
rect 2652 5412 2708 5468
rect 2708 5412 2712 5468
rect 2648 5408 2712 5412
rect 2728 5468 2792 5472
rect 2728 5412 2732 5468
rect 2732 5412 2788 5468
rect 2788 5412 2792 5468
rect 2728 5408 2792 5412
rect 2808 5468 2872 5472
rect 2808 5412 2812 5468
rect 2812 5412 2868 5468
rect 2868 5412 2872 5468
rect 2808 5408 2872 5412
rect 7568 5468 7632 5472
rect 7568 5412 7572 5468
rect 7572 5412 7628 5468
rect 7628 5412 7632 5468
rect 7568 5408 7632 5412
rect 7648 5468 7712 5472
rect 7648 5412 7652 5468
rect 7652 5412 7708 5468
rect 7708 5412 7712 5468
rect 7648 5408 7712 5412
rect 7728 5468 7792 5472
rect 7728 5412 7732 5468
rect 7732 5412 7788 5468
rect 7788 5412 7792 5468
rect 7728 5408 7792 5412
rect 7808 5468 7872 5472
rect 7808 5412 7812 5468
rect 7812 5412 7868 5468
rect 7868 5412 7872 5468
rect 7808 5408 7872 5412
rect 5068 4924 5132 4928
rect 5068 4868 5072 4924
rect 5072 4868 5128 4924
rect 5128 4868 5132 4924
rect 5068 4864 5132 4868
rect 5148 4924 5212 4928
rect 5148 4868 5152 4924
rect 5152 4868 5208 4924
rect 5208 4868 5212 4924
rect 5148 4864 5212 4868
rect 5228 4924 5292 4928
rect 5228 4868 5232 4924
rect 5232 4868 5288 4924
rect 5288 4868 5292 4924
rect 5228 4864 5292 4868
rect 5308 4924 5372 4928
rect 5308 4868 5312 4924
rect 5312 4868 5368 4924
rect 5368 4868 5372 4924
rect 5308 4864 5372 4868
rect 7568 4380 7632 4384
rect 7568 4324 7572 4380
rect 7572 4324 7628 4380
rect 7628 4324 7632 4380
rect 7568 4320 7632 4324
rect 7648 4380 7712 4384
rect 7648 4324 7652 4380
rect 7652 4324 7708 4380
rect 7708 4324 7712 4380
rect 7648 4320 7712 4324
rect 7728 4380 7792 4384
rect 7728 4324 7732 4380
rect 7732 4324 7788 4380
rect 7788 4324 7792 4380
rect 7728 4320 7792 4324
rect 7808 4380 7872 4384
rect 7808 4324 7812 4380
rect 7812 4324 7868 4380
rect 7868 4324 7872 4380
rect 7808 4320 7872 4324
rect 4844 4116 4908 4180
rect 5580 3904 5644 3908
rect 5580 3848 5594 3904
rect 5594 3848 5644 3904
rect 5580 3844 5644 3848
rect 5068 3836 5132 3840
rect 5068 3780 5072 3836
rect 5072 3780 5128 3836
rect 5128 3780 5132 3836
rect 5068 3776 5132 3780
rect 5148 3836 5212 3840
rect 5148 3780 5152 3836
rect 5152 3780 5208 3836
rect 5208 3780 5212 3836
rect 5148 3776 5212 3780
rect 5228 3836 5292 3840
rect 5228 3780 5232 3836
rect 5232 3780 5288 3836
rect 5288 3780 5292 3836
rect 5228 3776 5292 3780
rect 5308 3836 5372 3840
rect 5308 3780 5312 3836
rect 5312 3780 5368 3836
rect 5368 3780 5372 3836
rect 5308 3776 5372 3780
rect 7568 3292 7632 3296
rect 7568 3236 7572 3292
rect 7572 3236 7628 3292
rect 7628 3236 7632 3292
rect 7568 3232 7632 3236
rect 7648 3292 7712 3296
rect 7648 3236 7652 3292
rect 7652 3236 7708 3292
rect 7708 3236 7712 3292
rect 7648 3232 7712 3236
rect 7728 3292 7792 3296
rect 7728 3236 7732 3292
rect 7732 3236 7788 3292
rect 7788 3236 7792 3292
rect 7728 3232 7792 3236
rect 7808 3292 7872 3296
rect 7808 3236 7812 3292
rect 7812 3236 7868 3292
rect 7868 3236 7872 3292
rect 7808 3232 7872 3236
rect 5068 2748 5132 2752
rect 5068 2692 5072 2748
rect 5072 2692 5128 2748
rect 5128 2692 5132 2748
rect 5068 2688 5132 2692
rect 5148 2748 5212 2752
rect 5148 2692 5152 2748
rect 5152 2692 5208 2748
rect 5208 2692 5212 2748
rect 5148 2688 5212 2692
rect 5228 2748 5292 2752
rect 5228 2692 5232 2748
rect 5232 2692 5288 2748
rect 5288 2692 5292 2748
rect 5228 2688 5292 2692
rect 5308 2748 5372 2752
rect 5308 2692 5312 2748
rect 5312 2692 5368 2748
rect 5368 2692 5372 2748
rect 5308 2688 5372 2692
rect 4844 2484 4908 2548
rect 7568 2204 7632 2208
rect 7568 2148 7572 2204
rect 7572 2148 7628 2204
rect 7628 2148 7632 2204
rect 7568 2144 7632 2148
rect 7648 2204 7712 2208
rect 7648 2148 7652 2204
rect 7652 2148 7708 2204
rect 7708 2148 7712 2204
rect 7648 2144 7712 2148
rect 7728 2204 7792 2208
rect 7728 2148 7732 2204
rect 7732 2148 7788 2204
rect 7788 2148 7792 2204
rect 7728 2144 7792 2148
rect 7808 2204 7872 2208
rect 7808 2148 7812 2204
rect 7812 2148 7868 2204
rect 7868 2148 7872 2204
rect 7808 2144 7872 2148
rect 5068 1660 5132 1664
rect 5068 1604 5072 1660
rect 5072 1604 5128 1660
rect 5128 1604 5132 1660
rect 5068 1600 5132 1604
rect 5148 1660 5212 1664
rect 5148 1604 5152 1660
rect 5152 1604 5208 1660
rect 5208 1604 5212 1660
rect 5148 1600 5212 1604
rect 5228 1660 5292 1664
rect 5228 1604 5232 1660
rect 5232 1604 5288 1660
rect 5288 1604 5292 1660
rect 5228 1600 5292 1604
rect 5308 1660 5372 1664
rect 5308 1604 5312 1660
rect 5312 1604 5368 1660
rect 5368 1604 5372 1660
rect 5308 1600 5372 1604
rect 2568 1116 2632 1120
rect 2568 1060 2572 1116
rect 2572 1060 2628 1116
rect 2628 1060 2632 1116
rect 2568 1056 2632 1060
rect 2648 1116 2712 1120
rect 2648 1060 2652 1116
rect 2652 1060 2708 1116
rect 2708 1060 2712 1116
rect 2648 1056 2712 1060
rect 2728 1116 2792 1120
rect 2728 1060 2732 1116
rect 2732 1060 2788 1116
rect 2788 1060 2792 1116
rect 2728 1056 2792 1060
rect 2808 1116 2872 1120
rect 2808 1060 2812 1116
rect 2812 1060 2868 1116
rect 2868 1060 2872 1116
rect 2808 1056 2872 1060
rect 7568 1116 7632 1120
rect 7568 1060 7572 1116
rect 7572 1060 7628 1116
rect 7628 1060 7632 1116
rect 7568 1056 7632 1060
rect 7648 1116 7712 1120
rect 7648 1060 7652 1116
rect 7652 1060 7708 1116
rect 7708 1060 7712 1116
rect 7648 1056 7712 1060
rect 7728 1116 7792 1120
rect 7728 1060 7732 1116
rect 7732 1060 7788 1116
rect 7788 1060 7792 1116
rect 7728 1056 7792 1060
rect 7808 1116 7872 1120
rect 7808 1060 7812 1116
rect 7812 1060 7868 1116
rect 7868 1060 7872 1116
rect 7808 1056 7872 1060
rect 5068 572 5132 576
rect 5068 516 5072 572
rect 5072 516 5128 572
rect 5128 516 5132 572
rect 5068 512 5132 516
rect 5148 572 5212 576
rect 5148 516 5152 572
rect 5152 516 5208 572
rect 5208 516 5212 572
rect 5148 512 5212 516
rect 5228 572 5292 576
rect 5228 516 5232 572
rect 5232 516 5288 572
rect 5288 516 5292 572
rect 5228 512 5292 516
rect 5308 572 5372 576
rect 5308 516 5312 572
rect 5312 516 5368 572
rect 5368 516 5372 572
rect 5308 512 5372 516
<< metal4 >>
rect 2560 12000 2880 12016
rect 2560 11936 2568 12000
rect 2632 11936 2648 12000
rect 2712 11936 2728 12000
rect 2792 11936 2808 12000
rect 2872 11936 2880 12000
rect 2560 11598 2880 11936
rect 2560 11362 2602 11598
rect 2838 11362 2880 11598
rect 2560 10912 2880 11362
rect 2560 10848 2568 10912
rect 2632 10848 2648 10912
rect 2712 10848 2728 10912
rect 2792 10848 2808 10912
rect 2872 10848 2880 10912
rect 2560 9824 2880 10848
rect 3003 10572 3069 10573
rect 3003 10508 3004 10572
rect 3068 10508 3069 10572
rect 3003 10507 3069 10508
rect 2560 9760 2568 9824
rect 2632 9760 2648 9824
rect 2712 9760 2728 9824
rect 2792 9760 2808 9824
rect 2872 9760 2880 9824
rect 2560 8736 2880 9760
rect 2560 8672 2568 8736
rect 2632 8672 2648 8736
rect 2712 8672 2728 8736
rect 2792 8672 2808 8736
rect 2872 8672 2880 8736
rect 2560 8218 2880 8672
rect 2560 7982 2602 8218
rect 2838 7982 2880 8218
rect 2560 7648 2880 7982
rect 2560 7584 2568 7648
rect 2632 7584 2648 7648
rect 2712 7584 2728 7648
rect 2792 7584 2808 7648
rect 2872 7584 2880 7648
rect 2560 6560 2880 7584
rect 2560 6496 2568 6560
rect 2632 6496 2648 6560
rect 2712 6496 2728 6560
rect 2792 6496 2808 6560
rect 2872 6496 2880 6560
rect 2560 5472 2880 6496
rect 3006 6357 3066 10507
rect 3560 9266 3880 12016
rect 5060 11456 5380 12016
rect 5060 11392 5068 11456
rect 5132 11392 5148 11456
rect 5212 11392 5228 11456
rect 5292 11392 5308 11456
rect 5372 11392 5380 11456
rect 4475 11252 4541 11253
rect 4475 11188 4476 11252
rect 4540 11188 4541 11252
rect 4475 11187 4541 11188
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3003 6356 3069 6357
rect 3003 6292 3004 6356
rect 3068 6292 3069 6356
rect 3003 6291 3069 6292
rect 2560 5408 2568 5472
rect 2632 5408 2648 5472
rect 2712 5408 2728 5472
rect 2792 5408 2808 5472
rect 2872 5408 2880 5472
rect 2560 4838 2880 5408
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1120 2880 1222
rect 2560 1056 2568 1120
rect 2632 1056 2648 1120
rect 2712 1056 2728 1120
rect 2792 1056 2808 1120
rect 2872 1056 2880 1120
rect 2560 496 2880 1056
rect 3560 5886 3880 9030
rect 4478 6765 4538 11187
rect 5060 10368 5380 11392
rect 5060 10304 5068 10368
rect 5132 10304 5148 10368
rect 5212 10304 5228 10368
rect 5292 10304 5308 10368
rect 5372 10304 5380 10368
rect 5060 9908 5380 10304
rect 5060 9672 5102 9908
rect 5338 9672 5380 9908
rect 4843 9620 4909 9621
rect 4843 9556 4844 9620
rect 4908 9556 4909 9620
rect 4843 9555 4909 9556
rect 4475 6764 4541 6765
rect 4475 6700 4476 6764
rect 4540 6700 4541 6764
rect 4475 6699 4541 6700
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 3560 2506 3880 5650
rect 4846 4181 4906 9555
rect 5060 9280 5380 9672
rect 5060 9216 5068 9280
rect 5132 9216 5148 9280
rect 5212 9216 5228 9280
rect 5292 9216 5308 9280
rect 5372 9216 5380 9280
rect 5060 8192 5380 9216
rect 6060 10956 6380 12016
rect 6060 10720 6102 10956
rect 6338 10720 6380 10956
rect 5763 8668 5829 8669
rect 5763 8604 5764 8668
rect 5828 8604 5829 8668
rect 5763 8603 5829 8604
rect 5060 8128 5068 8192
rect 5132 8128 5148 8192
rect 5212 8128 5228 8192
rect 5292 8128 5308 8192
rect 5372 8128 5380 8192
rect 5060 7104 5380 8128
rect 5060 7040 5068 7104
rect 5132 7040 5148 7104
rect 5212 7040 5228 7104
rect 5292 7040 5308 7104
rect 5372 7040 5380 7104
rect 5060 6528 5380 7040
rect 5579 6764 5645 6765
rect 5579 6700 5580 6764
rect 5644 6700 5645 6764
rect 5579 6699 5645 6700
rect 5060 6292 5102 6528
rect 5338 6292 5380 6528
rect 5060 6016 5380 6292
rect 5060 5952 5068 6016
rect 5132 5952 5148 6016
rect 5212 5952 5228 6016
rect 5292 5952 5308 6016
rect 5372 5952 5380 6016
rect 5060 4928 5380 5952
rect 5060 4864 5068 4928
rect 5132 4864 5148 4928
rect 5212 4864 5228 4928
rect 5292 4864 5308 4928
rect 5372 4864 5380 4928
rect 4843 4180 4909 4181
rect 4843 4116 4844 4180
rect 4908 4116 4909 4180
rect 4843 4115 4909 4116
rect 4846 2549 4906 4115
rect 5060 3840 5380 4864
rect 5582 3909 5642 6699
rect 5766 6629 5826 8603
rect 6060 7576 6380 10720
rect 6060 7340 6102 7576
rect 6338 7340 6380 7576
rect 5763 6628 5829 6629
rect 5763 6564 5764 6628
rect 5828 6564 5829 6628
rect 5763 6563 5829 6564
rect 6060 4196 6380 7340
rect 6060 3960 6102 4196
rect 6338 3960 6380 4196
rect 5579 3908 5645 3909
rect 5579 3844 5580 3908
rect 5644 3844 5645 3908
rect 5579 3843 5645 3844
rect 5060 3776 5068 3840
rect 5132 3776 5148 3840
rect 5212 3776 5228 3840
rect 5292 3776 5308 3840
rect 5372 3776 5380 3840
rect 5060 3148 5380 3776
rect 5060 2912 5102 3148
rect 5338 2912 5380 3148
rect 5060 2752 5380 2912
rect 5060 2688 5068 2752
rect 5132 2688 5148 2752
rect 5212 2688 5228 2752
rect 5292 2688 5308 2752
rect 5372 2688 5380 2752
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 4843 2548 4909 2549
rect 4843 2484 4844 2548
rect 4908 2484 4909 2548
rect 4843 2483 4909 2484
rect 3560 496 3880 2270
rect 5060 1664 5380 2688
rect 5060 1600 5068 1664
rect 5132 1600 5148 1664
rect 5212 1600 5228 1664
rect 5292 1600 5308 1664
rect 5372 1600 5380 1664
rect 5060 576 5380 1600
rect 5060 512 5068 576
rect 5132 512 5148 576
rect 5212 512 5228 576
rect 5292 512 5308 576
rect 5372 512 5380 576
rect 5060 496 5380 512
rect 6060 496 6380 3960
rect 7560 12000 7880 12016
rect 7560 11936 7568 12000
rect 7632 11936 7648 12000
rect 7712 11936 7728 12000
rect 7792 11936 7808 12000
rect 7872 11936 7880 12000
rect 7560 11598 7880 11936
rect 7560 11362 7602 11598
rect 7838 11362 7880 11598
rect 7560 10912 7880 11362
rect 7560 10848 7568 10912
rect 7632 10848 7648 10912
rect 7712 10848 7728 10912
rect 7792 10848 7808 10912
rect 7872 10848 7880 10912
rect 7560 9824 7880 10848
rect 7560 9760 7568 9824
rect 7632 9760 7648 9824
rect 7712 9760 7728 9824
rect 7792 9760 7808 9824
rect 7872 9760 7880 9824
rect 7560 8736 7880 9760
rect 7560 8672 7568 8736
rect 7632 8672 7648 8736
rect 7712 8672 7728 8736
rect 7792 8672 7808 8736
rect 7872 8672 7880 8736
rect 7560 8218 7880 8672
rect 7560 7982 7602 8218
rect 7838 7982 7880 8218
rect 7560 7648 7880 7982
rect 7560 7584 7568 7648
rect 7632 7584 7648 7648
rect 7712 7584 7728 7648
rect 7792 7584 7808 7648
rect 7872 7584 7880 7648
rect 7560 6560 7880 7584
rect 7560 6496 7568 6560
rect 7632 6496 7648 6560
rect 7712 6496 7728 6560
rect 7792 6496 7808 6560
rect 7872 6496 7880 6560
rect 7560 5472 7880 6496
rect 7560 5408 7568 5472
rect 7632 5408 7648 5472
rect 7712 5408 7728 5472
rect 7792 5408 7808 5472
rect 7872 5408 7880 5472
rect 7560 4838 7880 5408
rect 7560 4602 7602 4838
rect 7838 4602 7880 4838
rect 7560 4384 7880 4602
rect 7560 4320 7568 4384
rect 7632 4320 7648 4384
rect 7712 4320 7728 4384
rect 7792 4320 7808 4384
rect 7872 4320 7880 4384
rect 7560 3296 7880 4320
rect 7560 3232 7568 3296
rect 7632 3232 7648 3296
rect 7712 3232 7728 3296
rect 7792 3232 7808 3296
rect 7872 3232 7880 3296
rect 7560 2208 7880 3232
rect 7560 2144 7568 2208
rect 7632 2144 7648 2208
rect 7712 2144 7728 2208
rect 7792 2144 7808 2208
rect 7872 2144 7880 2208
rect 7560 1458 7880 2144
rect 7560 1222 7602 1458
rect 7838 1222 7880 1458
rect 7560 1120 7880 1222
rect 7560 1056 7568 1120
rect 7632 1056 7648 1120
rect 7712 1056 7728 1120
rect 7792 1056 7808 1120
rect 7872 1056 7880 1120
rect 7560 496 7880 1056
rect 8560 9266 8880 12016
rect 8560 9030 8602 9266
rect 8838 9030 8880 9266
rect 8560 5886 8880 9030
rect 8560 5650 8602 5886
rect 8838 5650 8880 5886
rect 8560 2506 8880 5650
rect 8560 2270 8602 2506
rect 8838 2270 8880 2506
rect 8560 496 8880 2270
<< obsm4 >>
rect 9800 0 34000 13000
<< via4 >>
rect 2602 11362 2838 11598
rect 2602 7982 2838 8218
rect 3602 9030 3838 9266
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 2602 1222 2838 1458
rect 5102 9672 5338 9908
rect 3602 5650 3838 5886
rect 6102 10720 6338 10956
rect 5102 6292 5338 6528
rect 6102 7340 6338 7576
rect 6102 3960 6338 4196
rect 5102 2912 5338 3148
rect 3602 2270 3838 2506
rect 7602 11362 7838 11598
rect 7602 7982 7838 8218
rect 7602 4602 7838 4838
rect 7602 1222 7838 1458
rect 8602 9030 8838 9266
rect 8602 5650 8838 5886
rect 8602 2270 8838 2506
<< metal5 >>
rect 872 11598 10000 11640
rect 872 11362 2602 11598
rect 2838 11362 7602 11598
rect 7838 11362 10000 11598
rect 872 11320 10000 11362
rect 872 10956 10000 10998
rect 872 10720 6102 10956
rect 6338 10720 10000 10956
rect 872 10678 10000 10720
rect 872 9908 10000 9950
rect 872 9672 5102 9908
rect 5338 9672 10000 9908
rect 872 9630 10000 9672
rect 872 9266 10000 9308
rect 872 9030 3602 9266
rect 3838 9030 8602 9266
rect 8838 9030 10000 9266
rect 872 8988 10000 9030
rect 872 8218 10000 8260
rect 872 7982 2602 8218
rect 2838 7982 7602 8218
rect 7838 7982 10000 8218
rect 872 7940 10000 7982
rect 872 7576 10000 7618
rect 872 7340 6102 7576
rect 6338 7340 10000 7576
rect 872 7298 10000 7340
rect 872 6528 10000 6570
rect 872 6292 5102 6528
rect 5338 6292 10000 6528
rect 872 6250 10000 6292
rect 872 5886 10000 5928
rect 872 5650 3602 5886
rect 3838 5650 8602 5886
rect 8838 5650 10000 5886
rect 872 5608 10000 5650
rect 872 4838 10000 4880
rect 872 4602 2602 4838
rect 2838 4602 7602 4838
rect 7838 4602 10000 4838
rect 872 4560 10000 4602
rect 872 4196 10000 4238
rect 872 3960 2018 4196
rect 2254 3960 6102 4196
rect 6338 3960 10000 4196
rect 872 3918 10000 3960
rect 872 3148 10000 3190
rect 872 2912 5102 3148
rect 5338 2912 10000 3148
rect 872 2870 10000 2912
rect 872 2506 10000 2548
rect 872 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 8602 2506
rect 8838 2270 10000 2506
rect 872 2228 10000 2270
rect 872 1458 10000 1500
rect 872 1222 2602 1458
rect 2838 1222 7602 1458
rect 7838 1222 10000 1458
rect 872 1180 10000 1222
<< obsm5 >>
rect 10000 0 34000 13000
use sky130_fd_sc_hd__diode_2  ANTENNA__058__1_A deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3036 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A0
timestamp 1662439860
transform -1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__B
timestamp 1662439860
transform -1 0 9752 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__B
timestamp 1662439860
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__B
timestamp 1662439860
transform -1 0 8648 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__B
timestamp 1662439860
transform -1 0 2484 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__B
timestamp 1662439860
transform 1 0 3680 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__B
timestamp 1662439860
transform -1 0 3772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__B
timestamp 1662439860
transform -1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__B
timestamp 1662439860
transform -1 0 8832 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__B
timestamp 1662439860
transform -1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__B
timestamp 1662439860
transform -1 0 3680 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__B
timestamp 1662439860
transform -1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__B
timestamp 1662439860
transform 1 0 3312 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__B
timestamp 1662439860
transform -1 0 3496 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__B
timestamp 1662439860
transform -1 0 5152 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__B
timestamp 1662439860
transform -1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1662439860
transform -1 0 10120 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__B
timestamp 1662439860
transform -1 0 9568 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__B
timestamp 1662439860
transform -1 0 9752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__B
timestamp 1662439860
transform -1 0 2668 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__B
timestamp 1662439860
transform -1 0 8924 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__B
timestamp 1662439860
transform -1 0 9108 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__B
timestamp 1662439860
transform -1 0 5612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__B
timestamp 1662439860
transform -1 0 4508 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__B
timestamp 1662439860
transform 1 0 1196 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__B
timestamp 1662439860
transform 1 0 5704 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__B
timestamp 1662439860
transform -1 0 4324 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__B
timestamp 1662439860
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__B
timestamp 1662439860
transform -1 0 6164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__2_A
timestamp 1662439860
transform 1 0 5336 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__5_A
timestamp 1662439860
transform 1 0 3220 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__6_A
timestamp 1662439860
transform 1 0 3772 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__7_A
timestamp 1662439860
transform 1 0 3588 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__9_A
timestamp 1662439860
transform 1 0 2852 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__10_A
timestamp 1662439860
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__RESET_B
timestamp 1662439860
transform -1 0 2852 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1662439860
transform 1 0 5520 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A
timestamp 1662439860
transform -1 0 1380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_load_A
timestamp 1662439860
transform -1 0 3680 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout27_A
timestamp 1662439860
transform -1 0 6440 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout28_A
timestamp 1662439860
transform 1 0 8280 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1662439860
transform -1 0 6624 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1662439860
transform -1 0 5888 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1662439860
transform -1 0 6072 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1662439860
transform -1 0 4692 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1662439860
transform -1 0 4140 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_serial_load_out_buffer_A
timestamp 1662439860
transform 1 0 5152 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3404 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33
timestamp 1662439860
transform 1 0 3956 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 1662439860
transform 1 0 6164 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30 deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3680 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_34
timestamp 1662439860
transform 1 0 4048 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp 1662439860
transform 1 0 3864 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_41 deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 4692 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49 deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 5428 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_43
timestamp 1662439860
transform 1 0 4876 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_52
timestamp 1662439860
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_84
timestamp 1662439860
transform 1 0 8648 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_26
timestamp 1662439860
transform 1 0 3312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_34
timestamp 1662439860
transform 1 0 4048 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_80
timestamp 1662439860
transform 1 0 8280 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_26
timestamp 1662439860
transform 1 0 3312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_65
timestamp 1662439860
transform 1 0 6900 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1662439860
transform 1 0 10028 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_99
timestamp 1662439860
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1662439860
transform 1 0 8556 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_50
timestamp 1662439860
transform 1 0 5520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1662439860
transform 1 0 6164 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_99
timestamp 1662439860
transform 1 0 10028 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0 deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 920 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1662439860
transform -1 0 10396 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1662439860
transform 1 0 3036 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1662439860
transform -1 0 10396 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1662439860
transform 1 0 3036 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1662439860
transform -1 0 10396 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1662439860
transform 1 0 3036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1662439860
transform -1 0 10396 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1662439860
transform 1 0 3036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1662439860
transform -1 0 10396 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1662439860
transform 1 0 3036 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1662439860
transform -1 0 10396 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1662439860
transform 1 0 3036 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1662439860
transform -1 0 10396 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1662439860
transform 1 0 3036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1662439860
transform -1 0 10396 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1662439860
transform 1 0 3036 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1662439860
transform -1 0 10396 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1662439860
transform 1 0 920 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1662439860
transform -1 0 10396 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1662439860
transform 1 0 920 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1662439860
transform -1 0 10396 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1662439860
transform 1 0 920 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1662439860
transform -1 0 10396 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1662439860
transform 1 0 920 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1662439860
transform -1 0 10396 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1662439860
transform 1 0 920 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1662439860
transform -1 0 10396 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1662439860
transform 1 0 920 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1662439860
transform -1 0 10396 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1662439860
transform 1 0 920 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1662439860
transform -1 0 10396 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1662439860
transform 1 0 920 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1662439860
transform -1 0 10396 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1662439860
transform 1 0 920 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1662439860
transform -1 0 10396 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1662439860
transform 1 0 920 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1662439860
transform -1 0 10396 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1662439860
transform 1 0 920 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1662439860
transform -1 0 10396 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1662439860
transform 1 0 920 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1662439860
transform -1 0 10396 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42 deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3496 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1662439860
transform 1 0 6072 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1662439860
transform 1 0 8648 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1662439860
transform 1 0 8188 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1662439860
transform 1 0 5612 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1662439860
transform 1 0 8188 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1662439860
transform 1 0 5612 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1662439860
transform 1 0 8188 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1662439860
transform 1 0 5612 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1662439860
transform 1 0 8188 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1662439860
transform 1 0 5612 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1662439860
transform 1 0 3496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1662439860
transform 1 0 6072 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1662439860
transform 1 0 8648 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1662439860
transform 1 0 3496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1662439860
transform 1 0 8648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1662439860
transform 1 0 6072 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1662439860
transform 1 0 3496 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1662439860
transform 1 0 8648 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1662439860
transform 1 0 6072 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1662439860
transform 1 0 3496 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1662439860
transform 1 0 8648 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1662439860
transform 1 0 6072 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1662439860
transform 1 0 3496 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1662439860
transform 1 0 8648 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1662439860
transform 1 0 6072 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1662439860
transform 1 0 3496 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1662439860
transform 1 0 8648 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1662439860
transform 1 0 6072 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1662439860
transform 1 0 3496 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1662439860
transform 1 0 6072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1662439860
transform 1 0 8648 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _058__1 deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 2024 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059__14
timestamp 1662439860
transform -1 0 4876 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and2_0  _060_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 8740 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _061_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2b_2  _062_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 9384 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _063_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9936 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _064_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 9108 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _065_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 10120 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _066_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 10120 0 -1 7072
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _067_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 8556 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__or2_0  _068_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 6164 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _069_
timestamp 1662439860
transform 1 0 9476 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _070_
timestamp 1662439860
transform -1 0 1656 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _071_
timestamp 1662439860
transform -1 0 4232 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _072_
timestamp 1662439860
transform 1 0 5612 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _073_
timestamp 1662439860
transform 1 0 6900 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _074_
timestamp 1662439860
transform -1 0 10028 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _075_
timestamp 1662439860
transform -1 0 10120 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _076_
timestamp 1662439860
transform 1 0 3588 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _077_
timestamp 1662439860
transform -1 0 6808 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _078_
timestamp 1662439860
transform 1 0 3312 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _079_
timestamp 1662439860
transform -1 0 4048 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _080_
timestamp 1662439860
transform 1 0 5152 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _081_
timestamp 1662439860
transform 1 0 6900 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _082_
timestamp 1662439860
transform -1 0 10028 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _083_
timestamp 1662439860
transform -1 0 9384 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _084_
timestamp 1662439860
transform -1 0 1656 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _085_
timestamp 1662439860
transform 1 0 9476 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _086_
timestamp 1662439860
transform 1 0 9108 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _087_
timestamp 1662439860
transform 1 0 7544 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _088_
timestamp 1662439860
transform 1 0 1196 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _089_
timestamp 1662439860
transform -1 0 5244 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _090_
timestamp 1662439860
transform 1 0 6440 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _091_
timestamp 1662439860
transform 1 0 3404 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__or2_0  _092_
timestamp 1662439860
transform 1 0 6164 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _093_
timestamp 1662439860
transform 1 0 6624 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _094__2
timestamp 1662439860
transform -1 0 5428 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095__3
timestamp 1662439860
transform 1 0 8372 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096__4
timestamp 1662439860
transform -1 0 1472 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097__5
timestamp 1662439860
transform 1 0 1748 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098__6
timestamp 1662439860
transform 1 0 1196 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099__7
timestamp 1662439860
transform 1 0 1472 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100__8
timestamp 1662439860
transform -1 0 7544 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101__9
timestamp 1662439860
transform 1 0 1196 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102__10
timestamp 1662439860
transform 1 0 8740 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103__11
timestamp 1662439860
transform -1 0 3864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _104__12
timestamp 1662439860
transform -1 0 4600 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105__13
timestamp 1662439860
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_2  _106_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 5888 0 1 10336
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _107_
timestamp 1662439860
transform 1 0 3496 0 -1 11424
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _108_
timestamp 1662439860
transform -1 0 8648 0 1 7072
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _109_
timestamp 1662439860
transform 1 0 7544 0 -1 8160
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _110_
timestamp 1662439860
transform 1 0 3588 0 1 9248
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _111_
timestamp 1662439860
transform 1 0 3496 0 -1 8160
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _112_
timestamp 1662439860
transform 1 0 3496 0 -1 10336
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _113_
timestamp 1662439860
transform 1 0 6992 0 1 4896
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _114_
timestamp 1662439860
transform 1 0 6992 0 -1 10336
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _115_
timestamp 1662439860
transform 1 0 7544 0 -1 11424
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _116_
timestamp 1662439860
transform 1 0 3496 0 -1 7072
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _117_
timestamp 1662439860
transform 1 0 4048 0 -1 4896
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _118_
timestamp 1662439860
transform 1 0 5244 0 1 5984
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_4  _119_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 3772 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _120_
timestamp 1662439860
transform 1 0 1380 0 -1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _121_
timestamp 1662439860
transform 1 0 1380 0 1 10336
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _122_
timestamp 1662439860
transform -1 0 3496 0 1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _123_
timestamp 1662439860
transform 1 0 2668 0 -1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _124_
timestamp 1662439860
transform -1 0 3496 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _125_
timestamp 1662439860
transform 1 0 1380 0 -1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _126_
timestamp 1662439860
transform 1 0 3956 0 -1 5984
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _127_
timestamp 1662439860
transform -1 0 6072 0 1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _128_
timestamp 1662439860
transform 1 0 6256 0 1 8160
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _129_
timestamp 1662439860
transform -1 0 8924 0 -1 7072
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _130_
timestamp 1662439860
transform -1 0 8280 0 -1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _131_
timestamp 1662439860
transform 1 0 6532 0 1 9248
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _132_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 3496 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _133_ deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9568 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1662439860
transform 1 0 5704 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 3496 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_load
timestamp 1662439860
transform -1 0 3496 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_clock
timestamp 1662439860
transform -1 0 3496 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_serial_load
timestamp 1662439860
transform 1 0 3772 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_clock
timestamp 1662439860
transform 1 0 8280 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_serial_load
timestamp 1662439860
transform 1 0 3312 0 1 2720
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  const_source deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 9384 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1662439860
transform -1 0 6532 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1662439860
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1662439860
transform -1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 1662439860
transform -1 0 8648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1662439860
transform -1 0 9936 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1662439860
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1662439860
transform -1 0 1564 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout30
timestamp 1662439860
transform 1 0 9752 0 -1 3808
box -38 -48 406 592
use gpio_logic_high  gpio_logic_high
timestamp 0
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform 1 0 6256 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1662439860
transform -1 0 9476 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1662439860
transform -1 0 9476 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1662439860
transform -1 0 9476 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1662439860
transform -1 0 6900 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1662439860
transform 1 0 1196 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1662439860
transform 1 0 6164 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1662439860
transform -1 0 9476 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1662439860
transform 1 0 7820 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1662439860
transform -1 0 5520 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1662439860
transform -1 0 6440 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1662439860
transform 1 0 3864 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1662439860
transform 1 0 1932 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1662439860
transform 1 0 8832 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1662439860
transform -1 0 10120 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1662439860
transform -1 0 10120 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1662439860
transform -1 0 3680 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1662439860
transform -1 0 3956 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_16  one_buffer deps/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1662439860
transform -1 0 6164 0 -1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output6
timestamp 1662439860
transform -1 0 8648 0 1 544
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output7
timestamp 1662439860
transform 1 0 6164 0 -1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output8
timestamp 1662439860
transform -1 0 8096 0 1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output9
timestamp 1662439860
transform -1 0 6164 0 -1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output10
timestamp 1662439860
transform -1 0 8188 0 -1 2720
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output11
timestamp 1662439860
transform -1 0 8096 0 1 2720
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output12
timestamp 1662439860
transform -1 0 10120 0 1 1632
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output13
timestamp 1662439860
transform 1 0 6164 0 -1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output14
timestamp 1662439860
transform 1 0 6072 0 1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output15
timestamp 1662439860
transform 1 0 8096 0 1 2720
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output16
timestamp 1662439860
transform -1 0 8648 0 -1 5984
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output17
timestamp 1662439860
transform 1 0 8096 0 1 3808
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output18
timestamp 1662439860
transform -1 0 6256 0 1 8160
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output19
timestamp 1662439860
transform -1 0 3496 0 -1 8160
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output20
timestamp 1662439860
transform 1 0 6624 0 1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output21
timestamp 1662439860
transform 1 0 4048 0 1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_16  output22
timestamp 1662439860
transform -1 0 3496 0 1 11424
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_16  serial_clock_out_buffer
timestamp 1662439860
transform 1 0 8280 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  serial_load_out_buffer
timestamp 1662439860
transform 1 0 3312 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_16  zero_buffer
timestamp 1662439860
transform -1 0 6072 0 1 544
box -38 -48 2062 592
<< labels >>
flabel metal2 s 938 12200 994 13000 0 FreeSans 224 90 0 0 gpio_defaults[0]
port 0 nsew signal input
flabel metal2 s 5538 12200 5594 13000 0 FreeSans 224 90 0 0 gpio_defaults[10]
port 1 nsew signal input
flabel metal2 s 5998 12200 6054 13000 0 FreeSans 224 90 0 0 gpio_defaults[11]
port 2 nsew signal input
flabel metal2 s 6458 12200 6514 13000 0 FreeSans 224 90 0 0 gpio_defaults[12]
port 3 nsew signal input
flabel metal2 s 1398 12200 1454 13000 0 FreeSans 224 90 0 0 gpio_defaults[1]
port 4 nsew signal input
flabel metal2 s 1858 12200 1914 13000 0 FreeSans 224 90 0 0 gpio_defaults[2]
port 5 nsew signal input
flabel metal2 s 2318 12200 2374 13000 0 FreeSans 224 90 0 0 gpio_defaults[3]
port 6 nsew signal input
flabel metal2 s 2778 12200 2834 13000 0 FreeSans 224 90 0 0 gpio_defaults[4]
port 7 nsew signal input
flabel metal2 s 3238 12200 3294 13000 0 FreeSans 224 90 0 0 gpio_defaults[5]
port 8 nsew signal input
flabel metal2 s 3698 12200 3754 13000 0 FreeSans 224 90 0 0 gpio_defaults[6]
port 9 nsew signal input
flabel metal2 s 4158 12200 4214 13000 0 FreeSans 224 90 0 0 gpio_defaults[7]
port 10 nsew signal input
flabel metal2 s 4618 12200 4674 13000 0 FreeSans 224 90 0 0 gpio_defaults[8]
port 11 nsew signal input
flabel metal2 s 5078 12200 5134 13000 0 FreeSans 224 90 0 0 gpio_defaults[9]
port 12 nsew signal input
flabel metal3 s 14000 824 34000 944 0 FreeSans 480 0 0 0 mgmt_gpio_in
port 13 nsew signal tristate
flabel metal3 s 14000 1640 34000 1760 0 FreeSans 480 0 0 0 mgmt_gpio_oeb
port 14 nsew signal input
flabel metal3 s 14000 2048 34000 2168 0 FreeSans 480 0 0 0 mgmt_gpio_out
port 15 nsew signal input
flabel metal3 s 14000 1232 34000 1352 0 FreeSans 480 0 0 0 one
port 16 nsew signal tristate
flabel metal3 s 14000 2456 34000 2576 0 FreeSans 480 0 0 0 pad_gpio_ana_en
port 17 nsew signal tristate
flabel metal3 s 14000 2864 34000 2984 0 FreeSans 480 0 0 0 pad_gpio_ana_pol
port 18 nsew signal tristate
flabel metal3 s 14000 3272 34000 3392 0 FreeSans 480 0 0 0 pad_gpio_ana_sel
port 19 nsew signal tristate
flabel metal3 s 14000 3680 34000 3800 0 FreeSans 480 0 0 0 pad_gpio_dm[0]
port 20 nsew signal tristate
flabel metal3 s 14000 4088 34000 4208 0 FreeSans 480 0 0 0 pad_gpio_dm[1]
port 21 nsew signal tristate
flabel metal3 s 14000 4496 34000 4616 0 FreeSans 480 0 0 0 pad_gpio_dm[2]
port 22 nsew signal tristate
flabel metal3 s 14000 4904 34000 5024 0 FreeSans 480 0 0 0 pad_gpio_holdover
port 23 nsew signal tristate
flabel metal3 s 14000 5312 34000 5432 0 FreeSans 480 0 0 0 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
flabel metal3 s 14000 5720 34000 5840 0 FreeSans 480 0 0 0 pad_gpio_in
port 25 nsew signal input
flabel metal3 s 14000 6128 34000 6248 0 FreeSans 480 0 0 0 pad_gpio_inenb
port 26 nsew signal tristate
flabel metal3 s 14000 6536 34000 6656 0 FreeSans 480 0 0 0 pad_gpio_out
port 27 nsew signal tristate
flabel metal3 s 14000 6944 34000 7064 0 FreeSans 480 0 0 0 pad_gpio_outenb
port 28 nsew signal tristate
flabel metal3 s 14000 7352 34000 7472 0 FreeSans 480 0 0 0 pad_gpio_slow_sel
port 29 nsew signal tristate
flabel metal3 s 14000 7760 34000 7880 0 FreeSans 480 0 0 0 pad_gpio_vtrip_sel
port 30 nsew signal tristate
flabel metal3 s 14000 8168 34000 8288 0 FreeSans 480 0 0 0 resetn
port 31 nsew signal input
flabel metal3 s 14000 8576 34000 8696 0 FreeSans 480 0 0 0 resetn_out
port 32 nsew signal tristate
flabel metal3 s 14000 8984 34000 9104 0 FreeSans 480 0 0 0 serial_clock
port 33 nsew signal input
flabel metal3 s 14000 9392 34000 9512 0 FreeSans 480 0 0 0 serial_clock_out
port 34 nsew signal tristate
flabel metal3 s 14000 9800 34000 9920 0 FreeSans 480 0 0 0 serial_data_in
port 35 nsew signal input
flabel metal3 s 14000 10208 34000 10328 0 FreeSans 480 0 0 0 serial_data_out
port 36 nsew signal tristate
flabel metal3 s 14000 10616 34000 10736 0 FreeSans 480 0 0 0 serial_load
port 37 nsew signal input
flabel metal3 s 14000 11024 34000 11144 0 FreeSans 480 0 0 0 serial_load_out
port 38 nsew signal tristate
flabel metal3 s 14000 11432 34000 11552 0 FreeSans 480 0 0 0 user_gpio_in
port 39 nsew signal tristate
flabel metal3 s 14000 11840 34000 11960 0 FreeSans 480 0 0 0 user_gpio_oeb
port 40 nsew signal input
flabel metal3 s 14000 12248 34000 12368 0 FreeSans 480 0 0 0 user_gpio_out
port 41 nsew signal input
flabel metal4 s 2560 496 2880 12016 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 7560 496 7880 12016 0 FreeSans 1920 90 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 1180 10000 1500 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 4560 10000 4880 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 7940 10000 8260 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal5 s 872 11320 10000 11640 0 FreeSans 2560 0 0 0 vccd
port 42 nsew power bidirectional
flabel metal4 s 3560 496 3880 12016 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 8560 496 8880 12016 0 FreeSans 1920 90 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 2228 10000 2548 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 5608 10000 5928 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal5 s 872 8988 10000 9308 0 FreeSans 2560 0 0 0 vccd1
port 43 nsew power bidirectional
flabel metal4 s 5060 496 5380 12016 0 FreeSans 1920 90 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 2870 10000 3190 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 6250 10000 6570 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal5 s 872 9630 10000 9950 0 FreeSans 2560 0 0 0 vssd
port 44 nsew ground bidirectional
flabel metal4 s 6060 496 6380 12016 0 FreeSans 1920 90 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 3918 10000 4238 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 7298 10000 7618 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal5 s 872 10678 10000 10998 0 FreeSans 2560 0 0 0 vssd1
port 45 nsew ground bidirectional
flabel metal3 s 14000 416 34000 536 0 FreeSans 480 0 0 0 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
