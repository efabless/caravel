magic
tech sky130A
magscale 1 2
timestamp 1503891474
<< checkpaint >>
rect -1260 -1260 1261 1261
<< properties >>
string FIXED_BBOX 0 0 600000 5000
<< end >>
