magic
tech sky130A
magscale 1 2
timestamp 1608132867
<< obsli1 >>
rect 960 797 29952 3273
<< obsm1 >>
rect 784 763 29952 3307
<< metal2 >>
rect 2930 763 2990 3307
rect 3330 814 3390 3256
rect 3730 814 3790 3256
rect 10930 763 10990 3307
rect 11330 814 11390 3256
rect 11730 814 11790 3256
rect 18930 763 18990 3307
rect 19330 814 19390 3256
rect 19730 814 19790 3256
rect 26930 763 26990 3307
rect 27330 814 27390 3256
rect 27730 814 27790 3256
<< obsm2 >>
rect 788 925 2874 2923
rect 3046 925 3274 2923
rect 3446 925 3674 2923
rect 3846 925 10874 2923
rect 11046 925 11274 2923
rect 11446 925 11674 2923
rect 11846 925 18218 2923
<< metal3 >>
rect 960 3093 29952 3153
rect 0 2826 800 2946
rect 960 2864 29952 2924
rect 960 2464 29952 2524
rect 960 2013 29952 2073
rect 960 1784 29952 1844
rect 960 1384 29952 1444
rect 0 902 800 1022
rect 960 933 29952 993
<< obsm3 >>
rect 800 3026 880 3156
rect 880 3004 27793 3013
rect 880 2746 27793 2784
rect 800 2604 27793 2746
rect 800 2384 880 2604
rect 800 2153 27793 2384
rect 800 1933 880 2153
rect 800 1924 27793 1933
rect 800 1704 880 1924
rect 800 1524 27793 1704
rect 800 1304 880 1524
rect 800 1102 27793 1304
rect 880 1073 27793 1102
<< labels >>
rlabel metal3 s 0 902 800 1022 6 mprj2_vdd_logic1
port 1 nsew signal output
rlabel metal3 s 0 2826 800 2946 6 mprj_vdd_logic1
port 2 nsew signal output
rlabel metal2 s 18930 763 18990 3307 6 vccd
port 3 nsew power bidirectional
rlabel metal2 s 2930 763 2990 3307 6 vccd
port 4 nsew power bidirectional
rlabel metal3 s 960 3093 29952 3153 6 vccd
port 5 nsew power bidirectional
rlabel metal3 s 960 933 29952 993 6 vccd
port 6 nsew power bidirectional
rlabel metal2 s 26930 763 26990 3307 6 vssd
port 7 nsew ground bidirectional
rlabel metal2 s 10930 763 10990 3307 6 vssd
port 8 nsew ground bidirectional
rlabel metal3 s 960 2013 29952 2073 6 vssd
port 9 nsew ground bidirectional
rlabel metal2 s 19330 814 19390 3256 6 vdda1
port 10 nsew power bidirectional
rlabel metal2 s 3330 814 3390 3256 6 vdda1
port 11 nsew power bidirectional
rlabel metal3 s 960 1384 29952 1444 6 vdda1
port 12 nsew power bidirectional
rlabel metal2 s 27330 814 27390 3256 6 vssa1
port 13 nsew ground bidirectional
rlabel metal2 s 11330 814 11390 3256 6 vssa1
port 14 nsew ground bidirectional
rlabel metal3 s 960 2464 29952 2524 6 vssa1
port 15 nsew ground bidirectional
rlabel metal2 s 19730 814 19790 3256 6 vdda2
port 16 nsew power bidirectional
rlabel metal2 s 3730 814 3790 3256 6 vdda2
port 17 nsew power bidirectional
rlabel metal3 s 960 1784 29952 1844 6 vdda2
port 18 nsew power bidirectional
rlabel metal2 s 27730 814 27790 3256 6 vssa2
port 19 nsew ground bidirectional
rlabel metal2 s 11730 814 11790 3256 6 vssa2
port 20 nsew ground bidirectional
rlabel metal3 s 960 2864 29952 2924 6 vssa2
port 21 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 30000 4000
string LEFview TRUE
string GDS_FILE ../gds/mgmt_protect_hv.gds
string GDS_END 64368
string GDS_START 42692
<< end >>
