* NGSPICE file created from caravan.ext - technology: sky130A

* Black-box entry subcircuit for gpio_control_block abstract view
.subckt gpio_control_block gpio_defaults[0] gpio_defaults[10] gpio_defaults[11] gpio_defaults[12]
+ gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4] gpio_defaults[5]
+ gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in
+ mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en pad_gpio_ana_pol pad_gpio_ana_sel
+ pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover pad_gpio_ib_mode_sel
+ pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel pad_gpio_vtrip_sel
+ resetn resetn_out serial_clock serial_clock_out serial_data_in serial_data_out serial_load
+ serial_load_out user_gpio_in user_gpio_oeb user_gpio_out vccd vccd1 vssd vssd1 zero
.ends

* Black-box entry subcircuit for gpio_defaults_block abstract view
.subckt gpio_defaults_block VGND VPWR gpio_defaults[0] gpio_defaults[10] gpio_defaults[11]
+ gpio_defaults[12] gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4]
+ gpio_defaults[5] gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9]
.ends

* Black-box entry subcircuit for digital_pll abstract view
.subckt digital_pll VGND VPWR clockp[0] clockp[1] dco div[0] div[1] div[2] div[3]
+ div[4] enable ext_trim[0] ext_trim[10] ext_trim[11] ext_trim[12] ext_trim[13] ext_trim[14]
+ ext_trim[15] ext_trim[16] ext_trim[17] ext_trim[18] ext_trim[19] ext_trim[1] ext_trim[20]
+ ext_trim[21] ext_trim[22] ext_trim[23] ext_trim[24] ext_trim[25] ext_trim[2] ext_trim[3]
+ ext_trim[4] ext_trim[5] ext_trim[6] ext_trim[7] ext_trim[8] ext_trim[9] osc resetb
.ends

* Black-box entry subcircuit for chip_io_alt abstract view
.subckt chip_io_alt clock clock_core por flash_clk flash_csb flash_io0 flash_io0_di_core
+ flash_io0_do_core flash_io0_ieb_core flash_io0_oeb_core flash_io1 flash_io1_di_core
+ flash_io1_do_core flash_io1_ieb_core flash_io1_oeb_core gpio gpio_in_core gpio_inenb_core
+ gpio_mode0_core gpio_out_core gpio_outenb_core vccd_pad vdda_pad vddio_pad vddio_pad2
+ vssa_pad vssd_pad vssio_pad vssio_pad2 mprj_io[0] mprj_io_analog_en[0] mprj_io_analog_pol[0]
+ mprj_io_analog_sel[0] mprj_io_dm[0] mprj_io_dm[1] mprj_io_dm[2] mprj_io_holdover[0]
+ mprj_io_ib_mode_sel[0] mprj_io_inp_dis[0] mprj_io_oeb[0] mprj_io_out[0] mprj_io_slow_sel[0]
+ mprj_io_vtrip_sel[0] mprj_io_in[0] mprj_io_in_3v3[0] mprj_gpio_analog[3] mprj_gpio_noesd[3]
+ mprj_io[10] mprj_io_analog_en[10] mprj_io_analog_pol[10] mprj_io_analog_sel[10]
+ mprj_io_dm[30] mprj_io_dm[31] mprj_io_dm[32] mprj_io_holdover[10] mprj_io_ib_mode_sel[10]
+ mprj_io_inp_dis[10] mprj_io_oeb[10] mprj_io_out[10] mprj_io_slow_sel[10] mprj_io_vtrip_sel[10]
+ mprj_io_in[10] mprj_io_in_3v3[10] mprj_gpio_analog[4] mprj_gpio_noesd[4] mprj_io[11]
+ mprj_io_analog_en[11] mprj_io_analog_pol[11] mprj_io_analog_sel[11] mprj_io_dm[33]
+ mprj_io_dm[34] mprj_io_dm[35] mprj_io_holdover[11] mprj_io_ib_mode_sel[11] mprj_io_inp_dis[11]
+ mprj_io_oeb[11] mprj_io_out[11] mprj_io_slow_sel[11] mprj_io_vtrip_sel[11] mprj_io_in[11]
+ mprj_io_in_3v3[11] mprj_gpio_analog[5] mprj_gpio_noesd[5] mprj_io[12] mprj_io_analog_en[12]
+ mprj_io_analog_pol[12] mprj_io_analog_sel[12] mprj_io_dm[36] mprj_io_dm[37] mprj_io_dm[38]
+ mprj_io_holdover[12] mprj_io_ib_mode_sel[12] mprj_io_inp_dis[12] mprj_io_oeb[12]
+ mprj_io_out[12] mprj_io_slow_sel[12] mprj_io_vtrip_sel[12] mprj_io_in[12] mprj_io_in_3v3[12]
+ mprj_gpio_analog[6] mprj_gpio_noesd[6] mprj_io[13] mprj_io_analog_en[13] mprj_io_analog_pol[13]
+ mprj_io_analog_sel[13] mprj_io_dm[39] mprj_io_dm[40] mprj_io_dm[41] mprj_io_holdover[13]
+ mprj_io_ib_mode_sel[13] mprj_io_inp_dis[13] mprj_io_oeb[13] mprj_io_out[13] mprj_io_slow_sel[13]
+ mprj_io_vtrip_sel[13] mprj_io_in[13] mprj_io_in_3v3[13] mprj_io[1] mprj_io_analog_en[1]
+ mprj_io_analog_pol[1] mprj_io_analog_sel[1] mprj_io_dm[3] mprj_io_dm[4] mprj_io_dm[5]
+ mprj_io_holdover[1] mprj_io_ib_mode_sel[1] mprj_io_inp_dis[1] mprj_io_oeb[1] mprj_io_out[1]
+ mprj_io_slow_sel[1] mprj_io_vtrip_sel[1] mprj_io_in[1] mprj_io_in_3v3[1] mprj_io[2]
+ mprj_io_analog_en[2] mprj_io_analog_pol[2] mprj_io_analog_sel[2] mprj_io_dm[6] mprj_io_dm[7]
+ mprj_io_dm[8] mprj_io_holdover[2] mprj_io_ib_mode_sel[2] mprj_io_inp_dis[2] mprj_io_oeb[2]
+ mprj_io_out[2] mprj_io_slow_sel[2] mprj_io_vtrip_sel[2] mprj_io_in[2] mprj_io_in_3v3[2]
+ mprj_io[3] mprj_io_analog_en[3] mprj_io_analog_pol[3] mprj_io_analog_sel[3] mprj_io_dm[10]
+ mprj_io_dm[11] mprj_io_dm[9] mprj_io_holdover[3] mprj_io_ib_mode_sel[3] mprj_io_inp_dis[3]
+ mprj_io_oeb[3] mprj_io_out[3] mprj_io_slow_sel[3] mprj_io_vtrip_sel[3] mprj_io_in[3]
+ mprj_io_in_3v3[3] mprj_io[4] mprj_io_analog_en[4] mprj_io_analog_pol[4] mprj_io_analog_sel[4]
+ mprj_io_dm[12] mprj_io_dm[13] mprj_io_dm[14] mprj_io_holdover[4] mprj_io_ib_mode_sel[4]
+ mprj_io_inp_dis[4] mprj_io_oeb[4] mprj_io_out[4] mprj_io_slow_sel[4] mprj_io_vtrip_sel[4]
+ mprj_io_in[4] mprj_io_in_3v3[4] mprj_io[5] mprj_io_analog_en[5] mprj_io_analog_pol[5]
+ mprj_io_analog_sel[5] mprj_io_dm[15] mprj_io_dm[16] mprj_io_dm[17] mprj_io_holdover[5]
+ mprj_io_ib_mode_sel[5] mprj_io_inp_dis[5] mprj_io_oeb[5] mprj_io_out[5] mprj_io_slow_sel[5]
+ mprj_io_vtrip_sel[5] mprj_io_in[5] mprj_io_in_3v3[5] mprj_io[6] mprj_io_analog_en[6]
+ mprj_io_analog_pol[6] mprj_io_analog_sel[6] mprj_io_dm[18] mprj_io_dm[19] mprj_io_dm[20]
+ mprj_io_holdover[6] mprj_io_ib_mode_sel[6] mprj_io_inp_dis[6] mprj_io_oeb[6] mprj_io_out[6]
+ mprj_io_slow_sel[6] mprj_io_vtrip_sel[6] mprj_io_in[6] mprj_io_in_3v3[6] mprj_gpio_analog[0]
+ mprj_gpio_noesd[0] mprj_io[7] mprj_io_analog_en[7] mprj_io_analog_pol[7] mprj_io_analog_sel[7]
+ mprj_io_dm[21] mprj_io_dm[22] mprj_io_dm[23] mprj_io_holdover[7] mprj_io_ib_mode_sel[7]
+ mprj_io_inp_dis[7] mprj_io_oeb[7] mprj_io_out[7] mprj_io_slow_sel[7] mprj_io_vtrip_sel[7]
+ mprj_io_in[7] mprj_io_in_3v3[7] mprj_gpio_analog[1] mprj_gpio_noesd[1] mprj_io[8]
+ mprj_io_analog_en[8] mprj_io_analog_pol[8] mprj_io_analog_sel[8] mprj_io_dm[24]
+ mprj_io_dm[25] mprj_io_dm[26] mprj_io_holdover[8] mprj_io_ib_mode_sel[8] mprj_io_inp_dis[8]
+ mprj_io_oeb[8] mprj_io_out[8] mprj_io_slow_sel[8] mprj_io_vtrip_sel[8] mprj_io_in[8]
+ mprj_io_in_3v3[8] mprj_gpio_analog[2] mprj_gpio_noesd[2] mprj_io[9] mprj_io_analog_en[9]
+ mprj_io_analog_pol[9] mprj_io_analog_sel[9] mprj_io_dm[27] mprj_io_dm[28] mprj_io_dm[29]
+ mprj_io_holdover[9] mprj_io_ib_mode_sel[9] mprj_io_inp_dis[9] mprj_io_oeb[9] mprj_io_out[9]
+ mprj_io_slow_sel[9] mprj_io_vtrip_sel[9] mprj_io_in[9] mprj_io_in_3v3[9] mprj_gpio_analog[7]
+ mprj_gpio_noesd[7] mprj_io[25] mprj_io_analog_en[14] mprj_io_analog_pol[14] mprj_io_analog_sel[14]
+ mprj_io_dm[42] mprj_io_dm[43] mprj_io_dm[44] mprj_io_holdover[14] mprj_io_ib_mode_sel[14]
+ mprj_io_inp_dis[14] mprj_io_oeb[14] mprj_io_out[14] mprj_io_slow_sel[14] mprj_io_vtrip_sel[14]
+ mprj_io_in[14] mprj_io_in_3v3[14] mprj_gpio_analog[17] mprj_gpio_noesd[17] mprj_io[35]
+ mprj_io_analog_en[24] mprj_io_analog_pol[24] mprj_io_analog_sel[24] mprj_io_dm[72]
+ mprj_io_dm[73] mprj_io_dm[74] mprj_io_holdover[24] mprj_io_ib_mode_sel[24] mprj_io_inp_dis[24]
+ mprj_io_oeb[24] mprj_io_out[24] mprj_io_slow_sel[24] mprj_io_vtrip_sel[24] mprj_io_in[24]
+ mprj_io_in_3v3[24] mprj_io[36] mprj_io_analog_en[25] mprj_io_analog_pol[25] mprj_io_analog_sel[25]
+ mprj_io_dm[75] mprj_io_dm[76] mprj_io_dm[77] mprj_io_holdover[25] mprj_io_ib_mode_sel[25]
+ mprj_io_inp_dis[25] mprj_io_oeb[25] mprj_io_out[25] mprj_io_slow_sel[25] mprj_io_vtrip_sel[25]
+ mprj_io_in[25] mprj_io_in_3v3[25] mprj_io[37] mprj_io_analog_en[26] mprj_io_analog_pol[26]
+ mprj_io_analog_sel[26] mprj_io_dm[78] mprj_io_dm[79] mprj_io_dm[80] mprj_io_holdover[26]
+ mprj_io_ib_mode_sel[26] mprj_io_inp_dis[26] mprj_io_oeb[26] mprj_io_out[26] mprj_io_slow_sel[26]
+ mprj_io_vtrip_sel[26] mprj_io_in[26] mprj_io_in_3v3[26] mprj_gpio_analog[8] mprj_gpio_noesd[8]
+ mprj_io[26] mprj_io_analog_en[15] mprj_io_analog_pol[15] mprj_io_analog_sel[15]
+ mprj_io_dm[45] mprj_io_dm[46] mprj_io_dm[47] mprj_io_holdover[15] mprj_io_ib_mode_sel[15]
+ mprj_io_inp_dis[15] mprj_io_oeb[15] mprj_io_out[15] mprj_io_slow_sel[15] mprj_io_vtrip_sel[15]
+ mprj_io_in[15] mprj_io_in_3v3[15] mprj_gpio_analog[9] mprj_gpio_noesd[9] mprj_io[27]
+ mprj_io_analog_en[16] mprj_io_analog_pol[16] mprj_io_analog_sel[16] mprj_io_dm[48]
+ mprj_io_dm[49] mprj_io_dm[50] mprj_io_holdover[16] mprj_io_ib_mode_sel[16] mprj_io_inp_dis[16]
+ mprj_io_oeb[16] mprj_io_out[16] mprj_io_slow_sel[16] mprj_io_vtrip_sel[16] mprj_io_in[16]
+ mprj_io_in_3v3[16] mprj_gpio_analog[10] mprj_gpio_noesd[10] mprj_io[28] mprj_io_analog_en[17]
+ mprj_io_analog_pol[17] mprj_io_analog_sel[17] mprj_io_dm[51] mprj_io_dm[52] mprj_io_dm[53]
+ mprj_io_holdover[17] mprj_io_ib_mode_sel[17] mprj_io_inp_dis[17] mprj_io_oeb[17]
+ mprj_io_out[17] mprj_io_slow_sel[17] mprj_io_vtrip_sel[17] mprj_io_in[17] mprj_io_in_3v3[17]
+ mprj_gpio_analog[11] mprj_gpio_noesd[11] mprj_io[29] mprj_io_analog_en[18] mprj_io_analog_pol[18]
+ mprj_io_analog_sel[18] mprj_io_dm[54] mprj_io_dm[55] mprj_io_dm[56] mprj_io_holdover[18]
+ mprj_io_ib_mode_sel[18] mprj_io_inp_dis[18] mprj_io_oeb[18] mprj_io_out[18] mprj_io_slow_sel[18]
+ mprj_io_vtrip_sel[18] mprj_io_in[18] mprj_io_in_3v3[18] mprj_gpio_analog[12] mprj_gpio_noesd[12]
+ mprj_io[30] mprj_io_analog_en[19] mprj_io_analog_pol[19] mprj_io_analog_sel[19]
+ mprj_io_dm[57] mprj_io_dm[58] mprj_io_dm[59] mprj_io_holdover[19] mprj_io_ib_mode_sel[19]
+ mprj_io_inp_dis[19] mprj_io_oeb[19] mprj_io_out[19] mprj_io_slow_sel[19] mprj_io_vtrip_sel[19]
+ mprj_io_in[19] mprj_io_in_3v3[19] mprj_gpio_analog[13] mprj_gpio_noesd[13] mprj_io[31]
+ mprj_io_analog_en[20] mprj_io_analog_pol[20] mprj_io_analog_sel[20] mprj_io_dm[60]
+ mprj_io_dm[61] mprj_io_dm[62] mprj_io_holdover[20] mprj_io_ib_mode_sel[20] mprj_io_inp_dis[20]
+ mprj_io_oeb[20] mprj_io_out[20] mprj_io_slow_sel[20] mprj_io_vtrip_sel[20] mprj_io_in[20]
+ mprj_io_in_3v3[20] mprj_gpio_analog[14] mprj_gpio_noesd[14] mprj_io[32] mprj_io_analog_en[21]
+ mprj_io_analog_pol[21] mprj_io_analog_sel[21] mprj_io_dm[63] mprj_io_dm[64] mprj_io_dm[65]
+ mprj_io_holdover[21] mprj_io_ib_mode_sel[21] mprj_io_inp_dis[21] mprj_io_oeb[21]
+ mprj_io_out[21] mprj_io_slow_sel[21] mprj_io_vtrip_sel[21] mprj_io_in[21] mprj_io_in_3v3[21]
+ mprj_gpio_analog[15] mprj_gpio_noesd[15] mprj_io[33] mprj_io_analog_en[22] mprj_io_analog_pol[22]
+ mprj_io_analog_sel[22] mprj_io_dm[66] mprj_io_dm[67] mprj_io_dm[68] mprj_io_holdover[22]
+ mprj_io_ib_mode_sel[22] mprj_io_inp_dis[22] mprj_io_oeb[22] mprj_io_out[22] mprj_io_slow_sel[22]
+ mprj_io_vtrip_sel[22] mprj_io_in[22] mprj_io_in_3v3[22] mprj_gpio_analog[16] mprj_gpio_noesd[16]
+ mprj_io[34] mprj_io_analog_en[23] mprj_io_analog_pol[23] mprj_io_analog_sel[23]
+ mprj_io_dm[69] mprj_io_dm[70] mprj_io_dm[71] mprj_io_holdover[23] mprj_io_ib_mode_sel[23]
+ mprj_io_inp_dis[23] mprj_io_oeb[23] mprj_io_out[23] mprj_io_slow_sel[23] mprj_io_vtrip_sel[23]
+ mprj_io_in[23] mprj_io_in_3v3[23] resetb resetb_core_h vdda mprj_analog[1] mprj_io[15]
+ mprj_analog[2] mprj_io[16] mprj_analog[3] mprj_io[17] mprj_analog[0] mprj_io[14]
+ mprj_analog[4] mprj_clamp_high[0] mprj_clamp_low[0] mprj_io[18] vccd1_pad vdda1_pad
+ vdda1_pad2 vssa1_pad vssa1_pad2 vccd1 vdda1 vssa1 vssd1 vssd1_pad mprj_analog[7]
+ mprj_io[21] mprj_analog[8] mprj_io[22] mprj_analog[9] mprj_io[23] mprj_analog[10]
+ mprj_io[24] mprj_analog[5] mprj_clamp_high[1] mprj_clamp_low[1] mprj_io[19] mprj_analog[6]
+ mprj_clamp_high[2] mprj_clamp_low[2] mprj_io[20] vccd2_pad vdda2_pad vssa2_pad vccd2
+ vdda2 vssa2 vssd2 vssd2_pad flash_csb_core flash_clk_oeb_core flash_clk_core flash_csb_oeb_core
+ mprj_io_one[0] mprj_io_one[1] mprj_io_one[2] mprj_io_one[3] mprj_io_one[4] mprj_io_one[5]
+ mprj_io_one[6] mprj_io_one[7] mprj_io_one[8] mprj_io_one[9] mprj_io_one[10] mprj_io_one[11]
+ mprj_io_one[12] mprj_io_one[13] mprj_io_one[14] mprj_io_one[15] mprj_io_one[16]
+ mprj_io_one[17] mprj_io_one[18] mprj_io_one[19] mprj_io_one[20] mprj_io_one[21]
+ mprj_io_one[22] mprj_io_one[23] mprj_io_one[24] mprj_io_one[25] mprj_io_one[26]
+ porb_h gpio_mode1_core vccd vddio vssa vssd vssio
.ends

* Black-box entry subcircuit for mgmt_core_wrapper abstract view
.subckt mgmt_core_wrapper VGND VPWR clk_in clk_out core_clk core_rstn debug_in debug_mode
+ debug_oeb debug_out flash_clk flash_csb flash_io0_di flash_io0_do flash_io0_oeb
+ flash_io1_di flash_io1_do flash_io1_oeb flash_io2_di flash_io2_do flash_io2_oeb
+ flash_io3_di flash_io3_do flash_io3_oeb gpio_in_pad gpio_inenb_pad gpio_mode0_pad
+ gpio_mode1_pad gpio_out_pad gpio_outenb_pad hk_ack_i hk_cyc_o hk_dat_i[0] hk_dat_i[10]
+ hk_dat_i[11] hk_dat_i[12] hk_dat_i[13] hk_dat_i[14] hk_dat_i[15] hk_dat_i[16] hk_dat_i[17]
+ hk_dat_i[18] hk_dat_i[19] hk_dat_i[1] hk_dat_i[20] hk_dat_i[21] hk_dat_i[22] hk_dat_i[23]
+ hk_dat_i[24] hk_dat_i[25] hk_dat_i[26] hk_dat_i[27] hk_dat_i[28] hk_dat_i[29] hk_dat_i[2]
+ hk_dat_i[30] hk_dat_i[31] hk_dat_i[3] hk_dat_i[4] hk_dat_i[5] hk_dat_i[6] hk_dat_i[7]
+ hk_dat_i[8] hk_dat_i[9] hk_stb_o irq[0] irq[1] irq[2] irq[3] irq[4] irq[5] la_iena[0]
+ la_iena[100] la_iena[101] la_iena[102] la_iena[103] la_iena[104] la_iena[105] la_iena[106]
+ la_iena[107] la_iena[108] la_iena[109] la_iena[10] la_iena[110] la_iena[111] la_iena[112]
+ la_iena[113] la_iena[114] la_iena[115] la_iena[116] la_iena[117] la_iena[118] la_iena[119]
+ la_iena[11] la_iena[120] la_iena[121] la_iena[122] la_iena[123] la_iena[124] la_iena[125]
+ la_iena[126] la_iena[127] la_iena[12] la_iena[13] la_iena[14] la_iena[15] la_iena[16]
+ la_iena[17] la_iena[18] la_iena[19] la_iena[1] la_iena[20] la_iena[21] la_iena[22]
+ la_iena[23] la_iena[24] la_iena[25] la_iena[26] la_iena[27] la_iena[28] la_iena[29]
+ la_iena[2] la_iena[30] la_iena[31] la_iena[32] la_iena[33] la_iena[34] la_iena[35]
+ la_iena[36] la_iena[37] la_iena[38] la_iena[39] la_iena[3] la_iena[40] la_iena[41]
+ la_iena[42] la_iena[43] la_iena[44] la_iena[45] la_iena[46] la_iena[47] la_iena[48]
+ la_iena[49] la_iena[4] la_iena[50] la_iena[51] la_iena[52] la_iena[53] la_iena[54]
+ la_iena[55] la_iena[56] la_iena[57] la_iena[58] la_iena[59] la_iena[5] la_iena[60]
+ la_iena[61] la_iena[62] la_iena[63] la_iena[64] la_iena[65] la_iena[66] la_iena[67]
+ la_iena[68] la_iena[69] la_iena[6] la_iena[70] la_iena[71] la_iena[72] la_iena[73]
+ la_iena[74] la_iena[75] la_iena[76] la_iena[77] la_iena[78] la_iena[79] la_iena[7]
+ la_iena[80] la_iena[81] la_iena[82] la_iena[83] la_iena[84] la_iena[85] la_iena[86]
+ la_iena[87] la_iena[88] la_iena[89] la_iena[8] la_iena[90] la_iena[91] la_iena[92]
+ la_iena[93] la_iena[94] la_iena[95] la_iena[96] la_iena[97] la_iena[98] la_iena[99]
+ la_iena[9] la_input[0] la_input[100] la_input[101] la_input[102] la_input[103] la_input[104]
+ la_input[105] la_input[106] la_input[107] la_input[108] la_input[109] la_input[10]
+ la_input[110] la_input[111] la_input[112] la_input[113] la_input[114] la_input[115]
+ la_input[116] la_input[117] la_input[118] la_input[119] la_input[11] la_input[120]
+ la_input[121] la_input[122] la_input[123] la_input[124] la_input[125] la_input[126]
+ la_input[127] la_input[12] la_input[13] la_input[14] la_input[15] la_input[16] la_input[17]
+ la_input[18] la_input[19] la_input[1] la_input[20] la_input[21] la_input[22] la_input[23]
+ la_input[24] la_input[25] la_input[26] la_input[27] la_input[28] la_input[29] la_input[2]
+ la_input[30] la_input[31] la_input[32] la_input[33] la_input[34] la_input[35] la_input[36]
+ la_input[37] la_input[38] la_input[39] la_input[3] la_input[40] la_input[41] la_input[42]
+ la_input[43] la_input[44] la_input[45] la_input[46] la_input[47] la_input[48] la_input[49]
+ la_input[4] la_input[50] la_input[51] la_input[52] la_input[53] la_input[54] la_input[55]
+ la_input[56] la_input[57] la_input[58] la_input[59] la_input[5] la_input[60] la_input[61]
+ la_input[62] la_input[63] la_input[64] la_input[65] la_input[66] la_input[67] la_input[68]
+ la_input[69] la_input[6] la_input[70] la_input[71] la_input[72] la_input[73] la_input[74]
+ la_input[75] la_input[76] la_input[77] la_input[78] la_input[79] la_input[7] la_input[80]
+ la_input[81] la_input[82] la_input[83] la_input[84] la_input[85] la_input[86] la_input[87]
+ la_input[88] la_input[89] la_input[8] la_input[90] la_input[91] la_input[92] la_input[93]
+ la_input[94] la_input[95] la_input[96] la_input[97] la_input[98] la_input[99] la_input[9]
+ la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105]
+ la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111]
+ la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118]
+ la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124]
+ la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15]
+ la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21]
+ la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28]
+ la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34]
+ la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40]
+ la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47]
+ la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53]
+ la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5]
+ la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66]
+ la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72]
+ la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79]
+ la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85]
+ la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91]
+ la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98]
+ la_oenb[99] la_oenb[9] la_output[0] la_output[100] la_output[101] la_output[102]
+ la_output[103] la_output[104] la_output[105] la_output[106] la_output[107] la_output[108]
+ la_output[109] la_output[10] la_output[110] la_output[111] la_output[112] la_output[113]
+ la_output[114] la_output[115] la_output[116] la_output[117] la_output[118] la_output[119]
+ la_output[11] la_output[120] la_output[121] la_output[122] la_output[123] la_output[124]
+ la_output[125] la_output[126] la_output[127] la_output[12] la_output[13] la_output[14]
+ la_output[15] la_output[16] la_output[17] la_output[18] la_output[19] la_output[1]
+ la_output[20] la_output[21] la_output[22] la_output[23] la_output[24] la_output[25]
+ la_output[26] la_output[27] la_output[28] la_output[29] la_output[2] la_output[30]
+ la_output[31] la_output[32] la_output[33] la_output[34] la_output[35] la_output[36]
+ la_output[37] la_output[38] la_output[39] la_output[3] la_output[40] la_output[41]
+ la_output[42] la_output[43] la_output[44] la_output[45] la_output[46] la_output[47]
+ la_output[48] la_output[49] la_output[4] la_output[50] la_output[51] la_output[52]
+ la_output[53] la_output[54] la_output[55] la_output[56] la_output[57] la_output[58]
+ la_output[59] la_output[5] la_output[60] la_output[61] la_output[62] la_output[63]
+ la_output[64] la_output[65] la_output[66] la_output[67] la_output[68] la_output[69]
+ la_output[6] la_output[70] la_output[71] la_output[72] la_output[73] la_output[74]
+ la_output[75] la_output[76] la_output[77] la_output[78] la_output[79] la_output[7]
+ la_output[80] la_output[81] la_output[82] la_output[83] la_output[84] la_output[85]
+ la_output[86] la_output[87] la_output[88] la_output[89] la_output[8] la_output[90]
+ la_output[91] la_output[92] la_output[93] la_output[94] la_output[95] la_output[96]
+ la_output[97] la_output[98] la_output[99] la_output[9] mprj_ack_i mprj_adr_o[0]
+ mprj_adr_o[10] mprj_adr_o[11] mprj_adr_o[12] mprj_adr_o[13] mprj_adr_o[14] mprj_adr_o[15]
+ mprj_adr_o[16] mprj_adr_o[17] mprj_adr_o[18] mprj_adr_o[19] mprj_adr_o[1] mprj_adr_o[20]
+ mprj_adr_o[21] mprj_adr_o[22] mprj_adr_o[23] mprj_adr_o[24] mprj_adr_o[25] mprj_adr_o[26]
+ mprj_adr_o[27] mprj_adr_o[28] mprj_adr_o[29] mprj_adr_o[2] mprj_adr_o[30] mprj_adr_o[31]
+ mprj_adr_o[3] mprj_adr_o[4] mprj_adr_o[5] mprj_adr_o[6] mprj_adr_o[7] mprj_adr_o[8]
+ mprj_adr_o[9] mprj_cyc_o mprj_dat_i[0] mprj_dat_i[10] mprj_dat_i[11] mprj_dat_i[12]
+ mprj_dat_i[13] mprj_dat_i[14] mprj_dat_i[15] mprj_dat_i[16] mprj_dat_i[17] mprj_dat_i[18]
+ mprj_dat_i[19] mprj_dat_i[1] mprj_dat_i[20] mprj_dat_i[21] mprj_dat_i[22] mprj_dat_i[23]
+ mprj_dat_i[24] mprj_dat_i[25] mprj_dat_i[26] mprj_dat_i[27] mprj_dat_i[28] mprj_dat_i[29]
+ mprj_dat_i[2] mprj_dat_i[30] mprj_dat_i[31] mprj_dat_i[3] mprj_dat_i[4] mprj_dat_i[5]
+ mprj_dat_i[6] mprj_dat_i[7] mprj_dat_i[8] mprj_dat_i[9] mprj_dat_o[0] mprj_dat_o[10]
+ mprj_dat_o[11] mprj_dat_o[12] mprj_dat_o[13] mprj_dat_o[14] mprj_dat_o[15] mprj_dat_o[16]
+ mprj_dat_o[17] mprj_dat_o[18] mprj_dat_o[19] mprj_dat_o[1] mprj_dat_o[20] mprj_dat_o[21]
+ mprj_dat_o[22] mprj_dat_o[23] mprj_dat_o[24] mprj_dat_o[25] mprj_dat_o[26] mprj_dat_o[27]
+ mprj_dat_o[28] mprj_dat_o[29] mprj_dat_o[2] mprj_dat_o[30] mprj_dat_o[31] mprj_dat_o[3]
+ mprj_dat_o[4] mprj_dat_o[5] mprj_dat_o[6] mprj_dat_o[7] mprj_dat_o[8] mprj_dat_o[9]
+ mprj_sel_o[0] mprj_sel_o[1] mprj_sel_o[2] mprj_sel_o[3] mprj_stb_o mprj_wb_iena
+ mprj_we_o por_l_in por_l_out porb_h_in porb_h_out qspi_enabled resetn_in resetn_out
+ rstb_l_in rstb_l_out ser_rx ser_tx serial_clock_in serial_clock_out serial_data_2_in
+ serial_data_2_out serial_load_in serial_load_out serial_resetn_in serial_resetn_out
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb trap uart_enabled user_irq_ena[0]
+ user_irq_ena[1] user_irq_ena[2]
.ends

* Black-box entry subcircuit for simple_por abstract view
.subckt simple_por vdd1v8 vdd3v3 vss3v3 porb_h por_l porb_l vss1v8
.ends

* Black-box entry subcircuit for caravel_clocking abstract view
.subckt caravel_clocking VGND VPWR core_clk ext_clk ext_clk_sel ext_reset pll_clk
+ pll_clk90 resetb resetb_sync sel2[0] sel2[1] sel2[2] sel[0] sel[1] sel[2] user_clk
.ends

* Black-box entry subcircuit for spare_logic_block abstract view
.subckt spare_logic_block spare_xfq[0] spare_xfq[1] spare_xfqn[0] spare_xfqn[1] spare_xi[0]
+ spare_xi[1] spare_xi[2] spare_xi[3] spare_xib spare_xmx[0] spare_xmx[1] spare_xna[0]
+ spare_xna[1] spare_xno[0] spare_xno[1] spare_xz[0] spare_xz[10] spare_xz[11] spare_xz[12]
+ spare_xz[13] spare_xz[14] spare_xz[15] spare_xz[16] spare_xz[17] spare_xz[18] spare_xz[19]
+ spare_xz[1] spare_xz[20] spare_xz[21] spare_xz[22] spare_xz[23] spare_xz[24] spare_xz[25]
+ spare_xz[26] spare_xz[2] spare_xz[3] spare_xz[4] spare_xz[5] spare_xz[6] spare_xz[7]
+ spare_xz[8] spare_xz[9] vccd vssd
.ends

* Black-box entry subcircuit for user_id_programming abstract view
.subckt user_id_programming mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13]
+ mask_rev[14] mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1]
+ mask_rev[20] mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26]
+ mask_rev[27] mask_rev[28] mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3]
+ mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] VPWR VGND
.ends

.subckt sky130_fd_sc_hd__buf_8 A VGND VPWR X VNB VPB
X0 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X2 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X16 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=4.73e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=4.73e+06u
.ends

.subckt gpio_signal_buffering_alt mgmt_io_in_unbuf[6] mgmt_io_out_buf[6] mgmt_io_in_unbuf[5]
+ mgmt_io_in_unbuf[4] mgmt_io_in_unbuf[3] mgmt_io_in_unbuf[2] mgmt_io_in_unbuf[1]
+ mgmt_io_in_unbuf[0] mgmt_io_out_buf[0] mgmt_io_out_buf[1] mgmt_io_out_buf[2] mgmt_io_out_buf[3]
+ mgmt_io_out_buf[4] mgmt_io_out_buf[5] mgmt_io_out_unbuf[0] mgmt_io_out_unbuf[1]
+ mgmt_io_out_unbuf[2] mgmt_io_out_unbuf[3] mgmt_io_out_unbuf[4] mgmt_io_out_unbuf[5]
+ mgmt_io_out_unbuf[6] mgmt_io_in_buf[6] mgmt_io_in_buf[5] mgmt_io_in_buf[4] mgmt_io_in_buf[3]
+ mgmt_io_in_buf[2] mgmt_io_in_buf[1] mgmt_io_in_buf[0] mgmt_io_out_buf[10] mgmt_io_out_buf[11]
+ mgmt_io_in_unbuf[11] mgmt_io_in_unbuf[10] mgmt_io_out_buf[12] mgmt_io_out_buf[13]
+ mgmt_io_out_buf[14] mgmt_io_out_buf[15] mgmt_io_in_unbuf[15] mgmt_io_in_unbuf[14]
+ mgmt_io_in_unbuf[13] mgmt_io_in_unbuf[12] mgmt_io_out_buf[16] mgmt_io_out_buf[17]
+ mgmt_io_out_buf[18] mgmt_io_out_buf[19] mgmt_io_in_unbuf[19] mgmt_io_in_unbuf[18]
+ mgmt_io_in_unbuf[17] mgmt_io_in_unbuf[16] mgmt_io_oeb_buf[0] mgmt_io_oeb_buf[1]
+ mgmt_io_oeb_buf[2] mgmt_io_oeb_unbuf[2] mgmt_io_oeb_unbuf[1] mgmt_io_oeb_unbuf[0]
+ mgmt_io_in_buf[19] mgmt_io_in_buf[18] mgmt_io_in_buf[17] mgmt_io_in_buf[16] mgmt_io_out_unbuf[16]
+ mgmt_io_out_unbuf[17] mgmt_io_out_unbuf[18] mgmt_io_out_unbuf[19] mgmt_io_out_unbuf[15]
+ mgmt_io_out_unbuf[14] mgmt_io_out_unbuf[13] mgmt_io_out_unbuf[12] mgmt_io_out_unbuf[11]
+ mgmt_io_out_unbuf[10] mgmt_io_out_unbuf[9] mgmt_io_out_unbuf[8] mgmt_io_out_unbuf[7]
+ mgmt_io_in_buf[7] mgmt_io_in_buf[8] mgmt_io_in_buf[9] mgmt_io_in_buf[10] mgmt_io_in_buf[11]
+ mgmt_io_in_buf[12] mgmt_io_in_buf[13] mgmt_io_in_buf[14] mgmt_io_in_buf[15] vccd
+ mgmt_io_out_buf[9] mgmt_io_in_unbuf[9] mgmt_io_out_buf[8] mgmt_io_in_unbuf[8] mgmt_io_out_buf[7]
+ mgmt_io_in_unbuf[7] vssd
Xsky130_fd_sc_hd__buf_8_1 sky130_fd_sc_hd__buf_8_1/A vssd vccd sky130_fd_sc_hd__buf_8_1/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_2 mgmt_io_in_unbuf[16] vssd vccd sky130_fd_sc_hd__buf_8_2/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_3 sky130_fd_sc_hd__buf_8_3/A vssd vccd mgmt_io_out_buf[17]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_4 mgmt_io_in_unbuf[18] vssd vccd sky130_fd_sc_hd__buf_8_4/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_5 sky130_fd_sc_hd__buf_8_5/A vssd vccd mgmt_io_out_buf[19]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_6 mgmt_io_in_unbuf[19] vssd vccd sky130_fd_sc_hd__buf_8_6/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_7 sky130_fd_sc_hd__buf_8_7/A vssd vccd mgmt_io_oeb_buf[0]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_8 sky130_fd_sc_hd__buf_8_8/A vssd vccd mgmt_io_oeb_buf[1]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_0 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_9 sky130_fd_sc_hd__buf_8_9/A vssd vccd mgmt_io_oeb_buf[2]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_1 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_2 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_3 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_50 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_4 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_51 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_40 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_90 sky130_fd_sc_hd__buf_8_90/A vssd vccd mgmt_io_in_buf[14]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_5 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_170 sky130_fd_sc_hd__buf_8_170/A vssd vccd mgmt_io_out_buf[7]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_52 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_41 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_30 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_6 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_91 mgmt_io_out_unbuf[13] vssd vccd sky130_fd_sc_hd__buf_8_91/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_80 sky130_fd_sc_hd__buf_8_80/A vssd vccd sky130_fd_sc_hd__buf_8_90/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_53 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_42 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_31 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_20 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_171 mgmt_io_in_unbuf[7] vssd vccd sky130_fd_sc_hd__buf_8_171/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_7 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_92 mgmt_io_out_unbuf[12] vssd vccd sky130_fd_sc_hd__buf_8_92/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_81 sky130_fd_sc_hd__buf_8_91/X vssd vccd sky130_fd_sc_hd__buf_8_81/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_70 sky130_fd_sc_hd__buf_8_70/A vssd vccd sky130_fd_sc_hd__buf_8_70/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_172 mgmt_io_in_unbuf[8] vssd vccd sky130_fd_sc_hd__buf_8_172/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_54 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_43 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_32 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_21 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_10 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_8 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_93 sky130_fd_sc_hd__buf_8_93/A vssd vccd mgmt_io_in_buf[13]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_82 sky130_fd_sc_hd__buf_8_82/A vssd vccd sky130_fd_sc_hd__buf_8_89/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_71 sky130_fd_sc_hd__buf_8_71/A vssd vccd sky130_fd_sc_hd__buf_8_71/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_55 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_44 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_33 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_22 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_11 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_173 sky130_fd_sc_hd__buf_8_173/A vssd vccd mgmt_io_out_buf[8]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_140 sky130_fd_sc_hd__buf_8_71/X vssd vccd sky130_fd_sc_hd__buf_8_173/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_9 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_94 mgmt_io_out_unbuf[11] vssd vccd sky130_fd_sc_hd__buf_8_94/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_83 sky130_fd_sc_hd__buf_8_88/X vssd vccd sky130_fd_sc_hd__buf_8_83/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_72 sky130_fd_sc_hd__buf_8_72/A vssd vccd sky130_fd_sc_hd__buf_8_97/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_50 mgmt_io_out_unbuf[3] vssd vccd mgmt_io_out_buf[3] vssd
+ vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_141 sky130_fd_sc_hd__buf_8_172/X vssd vccd sky130_fd_sc_hd__buf_8_68/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_130 mgmt_io_in_unbuf[14] vssd vccd sky130_fd_sc_hd__buf_8_80/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_56 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_45 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_34 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_23 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_12 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_174 sky130_fd_sc_hd__buf_8_174/A vssd vccd mgmt_io_out_buf[9]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_95 sky130_fd_sc_hd__buf_8_95/A vssd vccd mgmt_io_in_buf[12]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_84 sky130_fd_sc_hd__buf_8_84/A vssd vccd mgmt_io_out_buf[18]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_73 sky130_fd_sc_hd__buf_8_99/X vssd vccd sky130_fd_sc_hd__buf_8_73/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_51 mgmt_io_in_unbuf[3] vssd vccd mgmt_io_in_buf[3] vssd vccd
+ sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_57 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_46 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_35 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_24 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_13 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_175 mgmt_io_in_unbuf[9] vssd vccd sky130_fd_sc_hd__buf_8_175/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_142 sky130_fd_sc_hd__buf_8_73/X vssd vccd sky130_fd_sc_hd__buf_8_174/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_131 sky130_fd_sc_hd__buf_8_83/X vssd vccd mgmt_io_out_buf[14]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_120 mgmt_io_out_unbuf[18] vssd vccd sky130_fd_sc_hd__buf_8_84/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_96 sky130_fd_sc_hd__buf_8_96/A vssd vccd mgmt_io_in_buf[11]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_85 mgmt_io_in_unbuf[17] vssd vccd sky130_fd_sc_hd__buf_8_85/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_74 sky130_fd_sc_hd__buf_8_74/A vssd vccd sky130_fd_sc_hd__buf_8_96/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_52 mgmt_io_out_unbuf[4] vssd vccd mgmt_io_out_buf[4] vssd
+ vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_58 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_47 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_36 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_25 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_14 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_176 sky130_fd_sc_hd__buf_8_176/A vssd vccd mgmt_io_out_buf[10]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_143 sky130_fd_sc_hd__buf_8_175/X vssd vccd sky130_fd_sc_hd__buf_8_70/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_132 mgmt_io_in_unbuf[13] vssd vccd sky130_fd_sc_hd__buf_8_79/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_121 sky130_fd_sc_hd__buf_8_85/X vssd vccd mgmt_io_in_buf[17]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_97 sky130_fd_sc_hd__buf_8_97/A vssd vccd mgmt_io_in_buf[10]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_86 mgmt_io_out_unbuf[15] vssd vccd sky130_fd_sc_hd__buf_8_1/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_75 sky130_fd_sc_hd__buf_8_98/X vssd vccd sky130_fd_sc_hd__buf_8_75/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_53 mgmt_io_in_unbuf[4] vssd vccd mgmt_io_in_buf[4] vssd vccd
+ sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_59 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_48 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_37 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_26 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_15 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_177 mgmt_io_in_unbuf[10] vssd vccd sky130_fd_sc_hd__buf_8_177/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_133 sky130_fd_sc_hd__buf_8_81/X vssd vccd mgmt_io_out_buf[13]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_122 sky130_fd_sc_hd__buf_8_4/X vssd vccd mgmt_io_in_buf[18]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_100 sky130_fd_sc_hd__buf_8_70/X vssd vccd mgmt_io_in_buf[9]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_98 mgmt_io_out_unbuf[10] vssd vccd sky130_fd_sc_hd__buf_8_98/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_76 sky130_fd_sc_hd__buf_8_76/A vssd vccd sky130_fd_sc_hd__buf_8_95/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_49 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_38 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_27 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_16 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_178 sky130_fd_sc_hd__buf_8_178/A vssd vccd mgmt_io_out_buf[11]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_134 sky130_fd_sc_hd__buf_8_177/X vssd vccd sky130_fd_sc_hd__buf_8_72/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_123 mgmt_io_out_unbuf[19] vssd vccd sky130_fd_sc_hd__buf_8_5/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_101 sky130_fd_sc_hd__buf_8_68/X vssd vccd mgmt_io_in_buf[8]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_99 mgmt_io_out_unbuf[9] vssd vccd sky130_fd_sc_hd__buf_8_99/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_88 mgmt_io_out_unbuf[14] vssd vccd sky130_fd_sc_hd__buf_8_88/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_77 sky130_fd_sc_hd__buf_8_94/X vssd vccd sky130_fd_sc_hd__buf_8_77/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_55 sky130_fd_sc_hd__buf_8_55/A vssd vccd mgmt_io_out_buf[16]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_39 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_28 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_17 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_179 mgmt_io_in_unbuf[11] vssd vccd sky130_fd_sc_hd__buf_8_179/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_135 sky130_fd_sc_hd__buf_8_75/X vssd vccd sky130_fd_sc_hd__buf_8_176/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_124 sky130_fd_sc_hd__buf_8_6/X vssd vccd mgmt_io_in_buf[19]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_102 sky130_fd_sc_hd__buf_8_67/X vssd vccd mgmt_io_in_buf[7]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_89 sky130_fd_sc_hd__buf_8_89/A vssd vccd mgmt_io_in_buf[15]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_78 sky130_fd_sc_hd__buf_8_92/X vssd vccd sky130_fd_sc_hd__buf_8_78/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_67 sky130_fd_sc_hd__buf_8_67/A vssd vccd sky130_fd_sc_hd__buf_8_67/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_34 mgmt_io_in_unbuf[5] vssd vccd mgmt_io_in_buf[5] vssd vccd
+ sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_12 mgmt_io_out_unbuf[0] vssd vccd mgmt_io_out_buf[0] vssd
+ vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_29 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_18 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_136 sky130_fd_sc_hd__buf_8_179/X vssd vccd sky130_fd_sc_hd__buf_8_74/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_125 mgmt_io_oeb_unbuf[1] vssd vccd sky130_fd_sc_hd__buf_8_8/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_103 mgmt_io_out_unbuf[8] vssd vccd sky130_fd_sc_hd__buf_8_71/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_24 sky130_fd_sc_hd__buf_8_37/X vssd vccd mgmt_io_out_buf[6]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_13 mgmt_io_in_unbuf[0] vssd vccd mgmt_io_in_buf[0] vssd vccd
+ sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_79 sky130_fd_sc_hd__buf_8_79/A vssd vccd sky130_fd_sc_hd__buf_8_93/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_68 sky130_fd_sc_hd__buf_8_68/A vssd vccd sky130_fd_sc_hd__buf_8_68/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_46 mgmt_io_in_unbuf[1] vssd vccd mgmt_io_in_buf[1] vssd vccd
+ sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_35 mgmt_io_out_unbuf[5] vssd vccd mgmt_io_out_buf[5] vssd
+ vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_148 sky130_fd_sc_hd__buf_8_69/X vssd vccd sky130_fd_sc_hd__buf_8_170/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_137 sky130_fd_sc_hd__buf_8_77/X vssd vccd sky130_fd_sc_hd__buf_8_178/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_126 mgmt_io_oeb_unbuf[0] vssd vccd sky130_fd_sc_hd__buf_8_7/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_104 mgmt_io_out_unbuf[7] vssd vccd sky130_fd_sc_hd__buf_8_69/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_ef_sc_hd__decap_12_19 vssd vccd vssd vccd sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_8_69 sky130_fd_sc_hd__buf_8_69/A vssd vccd sky130_fd_sc_hd__buf_8_69/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_47 mgmt_io_out_unbuf[1] vssd vccd mgmt_io_out_buf[1] vssd
+ vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_36 sky130_fd_sc_hd__buf_8_36/A vssd vccd mgmt_io_in_buf[6]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_25 mgmt_io_in_unbuf[6] vssd vccd sky130_fd_sc_hd__buf_8_36/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_149 sky130_fd_sc_hd__buf_8_171/X vssd vccd sky130_fd_sc_hd__buf_8_67/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_138 sky130_fd_sc_hd__buf_8_78/X vssd vccd mgmt_io_out_buf[12]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_127 mgmt_io_oeb_unbuf[2] vssd vccd sky130_fd_sc_hd__buf_8_9/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_48 mgmt_io_out_unbuf[2] vssd vccd mgmt_io_out_buf[2] vssd
+ vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_37 mgmt_io_out_unbuf[6] vssd vccd sky130_fd_sc_hd__buf_8_37/X
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_139 mgmt_io_in_unbuf[12] vssd vccd sky130_fd_sc_hd__buf_8_76/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_128 mgmt_io_in_unbuf[15] vssd vccd sky130_fd_sc_hd__buf_8_82/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_117 mgmt_io_out_unbuf[16] vssd vccd sky130_fd_sc_hd__buf_8_55/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_49 mgmt_io_in_unbuf[2] vssd vccd mgmt_io_in_buf[2] vssd vccd
+ sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_129 sky130_fd_sc_hd__buf_8_1/X vssd vccd mgmt_io_out_buf[15]
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_118 mgmt_io_out_unbuf[17] vssd vccd sky130_fd_sc_hd__buf_8_3/A
+ vssd vccd sky130_fd_sc_hd__buf_8
Xsky130_fd_sc_hd__buf_8_119 sky130_fd_sc_hd__buf_8_2/X vssd vccd mgmt_io_in_buf[16]
+ vssd vccd sky130_fd_sc_hd__buf_8
.ends

* Black-box entry subcircuit for mgmt_protect abstract view
.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_ack_i_core mprj_ack_i_user mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11]
+ mprj_adr_o_core[12] mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15]
+ mprj_adr_o_core[16] mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19]
+ mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23]
+ mprj_adr_o_core[24] mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27]
+ mprj_adr_o_core[28] mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31]
+ mprj_adr_o_core[3] mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7]
+ mprj_adr_o_core[8] mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11]
+ mprj_adr_o_user[12] mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15]
+ mprj_adr_o_user[16] mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19]
+ mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23]
+ mprj_adr_o_user[24] mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27]
+ mprj_adr_o_user[28] mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31]
+ mprj_adr_o_user[3] mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7]
+ mprj_adr_o_user[8] mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_i_core[0]
+ mprj_dat_i_core[10] mprj_dat_i_core[11] mprj_dat_i_core[12] mprj_dat_i_core[13]
+ mprj_dat_i_core[14] mprj_dat_i_core[15] mprj_dat_i_core[16] mprj_dat_i_core[17]
+ mprj_dat_i_core[18] mprj_dat_i_core[19] mprj_dat_i_core[1] mprj_dat_i_core[20] mprj_dat_i_core[21]
+ mprj_dat_i_core[22] mprj_dat_i_core[23] mprj_dat_i_core[24] mprj_dat_i_core[25]
+ mprj_dat_i_core[26] mprj_dat_i_core[27] mprj_dat_i_core[28] mprj_dat_i_core[29]
+ mprj_dat_i_core[2] mprj_dat_i_core[30] mprj_dat_i_core[31] mprj_dat_i_core[3] mprj_dat_i_core[4]
+ mprj_dat_i_core[5] mprj_dat_i_core[6] mprj_dat_i_core[7] mprj_dat_i_core[8] mprj_dat_i_core[9]
+ mprj_dat_i_user[0] mprj_dat_i_user[10] mprj_dat_i_user[11] mprj_dat_i_user[12] mprj_dat_i_user[13]
+ mprj_dat_i_user[14] mprj_dat_i_user[15] mprj_dat_i_user[16] mprj_dat_i_user[17]
+ mprj_dat_i_user[18] mprj_dat_i_user[19] mprj_dat_i_user[1] mprj_dat_i_user[20] mprj_dat_i_user[21]
+ mprj_dat_i_user[22] mprj_dat_i_user[23] mprj_dat_i_user[24] mprj_dat_i_user[25]
+ mprj_dat_i_user[26] mprj_dat_i_user[27] mprj_dat_i_user[28] mprj_dat_i_user[29]
+ mprj_dat_i_user[2] mprj_dat_i_user[30] mprj_dat_i_user[31] mprj_dat_i_user[3] mprj_dat_i_user[4]
+ mprj_dat_i_user[5] mprj_dat_i_user[6] mprj_dat_i_user[7] mprj_dat_i_user[8] mprj_dat_i_user[9]
+ mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13]
+ mprj_dat_o_core[14] mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17]
+ mprj_dat_o_core[18] mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21]
+ mprj_dat_o_core[22] mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25]
+ mprj_dat_o_core[26] mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29]
+ mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4]
+ mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9]
+ mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13]
+ mprj_dat_o_user[14] mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17]
+ mprj_dat_o_user[18] mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21]
+ mprj_dat_o_user[22] mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25]
+ mprj_dat_o_user[26] mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29]
+ mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4]
+ mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9]
+ mprj_iena_wb mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2] mprj_sel_o_core[3]
+ mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3] mprj_stb_o_core
+ mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood user1_vdd_powergood
+ user2_vcc_powergood user2_vdd_powergood user_clock user_clock2 user_irq[0] user_irq[1]
+ user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2] user_irq_ena[0] user_irq_ena[1]
+ user_irq_ena[2] user_reset vccd vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd vssd1 vssd2
.ends

* Black-box entry subcircuit for xres_buf abstract view
.subckt xres_buf A X VPWR VGND LVPWR LVGND
.ends

* Black-box entry subcircuit for user_analog_project_wrapper abstract view
.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[10]
+ io_analog[1] io_analog[2] io_analog[3] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_analog[6] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for housekeeping abstract view
.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
.ends

* Black-box entry subcircuit for buff_flash_clkrst abstract view
.subckt buff_flash_clkrst VGND VPWR in_n[0] in_n[10] in_n[11] in_n[1] in_n[2] in_n[3]
+ in_n[4] in_n[5] in_n[6] in_n[7] in_n[8] in_n[9] in_s[0] in_s[1] in_s[2] out_n[0]
+ out_n[1] out_n[2] out_s[0] out_s[10] out_s[11] out_s[1] out_s[2] out_s[3] out_s[4]
+ out_s[5] out_s[6] out_s[7] out_s[8] out_s[9]
.ends

.subckt caravan clock flash_clk flash_csb flash_io0 flash_io1 gpio mprj_io[0] mprj_io[10]
+ mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] mprj_io[15] mprj_io[16] mprj_io[17]
+ mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20] mprj_io[21] mprj_io[22] mprj_io[23]
+ mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27] mprj_io[28] mprj_io[29] mprj_io[2]
+ mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33] mprj_io[34] mprj_io[35] mprj_io[36]
+ mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] mprj_io[7] mprj_io[8] mprj_io[9]
+ resetb vccd vccd1 vccd2 vdda vdda1 vdda1_2 vdda2 vddio vddio_2 vssa vssa1 vssa1_2
+ vssa2 vssd vssd1 vssd2 vssio vssio_2
Xgpio_control_in_2\[0\] gpio_defaults_block_25/gpio_defaults[0] gpio_defaults_block_25/gpio_defaults[10]
+ gpio_defaults_block_25/gpio_defaults[11] gpio_defaults_block_25/gpio_defaults[12]
+ gpio_defaults_block_25/gpio_defaults[1] gpio_defaults_block_25/gpio_defaults[2]
+ gpio_defaults_block_25/gpio_defaults[3] gpio_defaults_block_25/gpio_defaults[4]
+ gpio_defaults_block_25/gpio_defaults[5] gpio_defaults_block_25/gpio_defaults[6]
+ gpio_defaults_block_25/gpio_defaults[7] gpio_defaults_block_25/gpio_defaults[8]
+ gpio_defaults_block_25/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[7] padframe/mprj_io_one[14]
+ sigbuf/mgmt_io_out_buf[7] padframe/mprj_io_one[14] padframe/mprj_io_analog_en[14]
+ padframe/mprj_io_analog_pol[14] padframe/mprj_io_analog_sel[14] padframe/mprj_io_dm[42]
+ padframe/mprj_io_dm[43] padframe/mprj_io_dm[44] padframe/mprj_io_holdover[14] padframe/mprj_io_ib_mode_sel[14]
+ padframe/mprj_io_in[14] padframe/mprj_io_inp_dis[14] padframe/mprj_io_out[14] padframe/mprj_io_oeb[14]
+ padframe/mprj_io_slow_sel[14] padframe/mprj_io_vtrip_sel[14] gpio_control_in_2\[0\]/resetn
+ gpio_control_in_2\[0\]/resetn_out gpio_control_in_2\[0\]/serial_clock gpio_control_in_2\[0\]/serial_clock_out
+ gpio_control_in_2\[0\]/serial_data_in gpio_control_in_2\[0\]/serial_data_out gpio_control_in_2\[0\]/serial_load
+ gpio_control_in_2\[0\]/serial_load_out mprj/io_in[14] mprj/io_oeb[14] mprj/io_out[14]
+ gpio_defaults_block_25/VPWR vccd1_core gpio_defaults_block_25/VGND vssd1_core gpio_control_in_2\[0\]/zero
+ gpio_control_block
Xgpio_defaults_block_11 gpio_defaults_block_11/VGND gpio_defaults_block_11/VPWR gpio_defaults_block_11/gpio_defaults[0]
+ gpio_defaults_block_11/gpio_defaults[10] gpio_defaults_block_11/gpio_defaults[11]
+ gpio_defaults_block_11/gpio_defaults[12] gpio_defaults_block_11/gpio_defaults[1]
+ gpio_defaults_block_11/gpio_defaults[2] gpio_defaults_block_11/gpio_defaults[3]
+ gpio_defaults_block_11/gpio_defaults[4] gpio_defaults_block_11/gpio_defaults[5]
+ gpio_defaults_block_11/gpio_defaults[6] gpio_defaults_block_11/gpio_defaults[7]
+ gpio_defaults_block_11/gpio_defaults[8] gpio_defaults_block_11/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_defaults_block_33 gpio_defaults_block_33/VGND gpio_defaults_block_33/VPWR gpio_defaults_block_33/gpio_defaults[0]
+ gpio_defaults_block_33/gpio_defaults[10] gpio_defaults_block_33/gpio_defaults[11]
+ gpio_defaults_block_33/gpio_defaults[12] gpio_defaults_block_33/gpio_defaults[1]
+ gpio_defaults_block_33/gpio_defaults[2] gpio_defaults_block_33/gpio_defaults[3]
+ gpio_defaults_block_33/gpio_defaults[4] gpio_defaults_block_33/gpio_defaults[5]
+ gpio_defaults_block_33/gpio_defaults[6] gpio_defaults_block_33/gpio_defaults[7]
+ gpio_defaults_block_33/gpio_defaults[8] gpio_defaults_block_33/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_defaults_block_12 gpio_defaults_block_12/VGND gpio_defaults_block_12/VPWR gpio_defaults_block_12/gpio_defaults[0]
+ gpio_defaults_block_12/gpio_defaults[10] gpio_defaults_block_12/gpio_defaults[11]
+ gpio_defaults_block_12/gpio_defaults[12] gpio_defaults_block_12/gpio_defaults[1]
+ gpio_defaults_block_12/gpio_defaults[2] gpio_defaults_block_12/gpio_defaults[3]
+ gpio_defaults_block_12/gpio_defaults[4] gpio_defaults_block_12/gpio_defaults[5]
+ gpio_defaults_block_12/gpio_defaults[6] gpio_defaults_block_12/gpio_defaults[7]
+ gpio_defaults_block_12/gpio_defaults[8] gpio_defaults_block_12/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_defaults_block_34 VSUBS sigbuf/vccd gpio_defaults_block_34/gpio_defaults[0]
+ gpio_defaults_block_34/gpio_defaults[10] gpio_defaults_block_34/gpio_defaults[11]
+ gpio_defaults_block_34/gpio_defaults[12] gpio_defaults_block_34/gpio_defaults[1]
+ gpio_defaults_block_34/gpio_defaults[2] gpio_defaults_block_34/gpio_defaults[3]
+ gpio_defaults_block_34/gpio_defaults[4] gpio_defaults_block_34/gpio_defaults[5]
+ gpio_defaults_block_34/gpio_defaults[6] gpio_defaults_block_34/gpio_defaults[7]
+ gpio_defaults_block_34/gpio_defaults[8] gpio_defaults_block_34/gpio_defaults[9]
+ gpio_defaults_block
Xpll soc/VGND soc/VPWR pll/clockp[0] pll/clockp[1] pll/dco pll/div[0] pll/div[1] pll/div[2]
+ pll/div[3] pll/div[4] pll/enable pll/ext_trim[0] pll/ext_trim[10] pll/ext_trim[11]
+ pll/ext_trim[12] pll/ext_trim[13] pll/ext_trim[14] pll/ext_trim[15] pll/ext_trim[16]
+ pll/ext_trim[17] pll/ext_trim[18] pll/ext_trim[19] pll/ext_trim[1] pll/ext_trim[20]
+ pll/ext_trim[21] pll/ext_trim[22] pll/ext_trim[23] pll/ext_trim[24] pll/ext_trim[25]
+ pll/ext_trim[2] pll/ext_trim[3] pll/ext_trim[4] pll/ext_trim[5] pll/ext_trim[6]
+ pll/ext_trim[7] pll/ext_trim[8] pll/ext_trim[9] pll/osc pll/resetb digital_pll
Xpadframe clock padframe/clock_core padframe/por flash_clk flash_csb flash_io0 padframe/flash_io0_di_core
+ padframe/flash_io0_do_core padframe/flash_io0_ieb_core padframe/flash_io0_oeb_core
+ flash_io1 padframe/flash_io1_di_core padframe/flash_io1_do_core padframe/flash_io1_ieb_core
+ padframe/flash_io1_oeb_core gpio soc/gpio_in_pad soc/gpio_inenb_pad soc/gpio_mode0_pad
+ soc/gpio_out_pad soc/gpio_outenb_pad vccd vdda vddio vddio_2 vssa vssd vssio vssio_2
+ mprj_io[0] padframe/mprj_io_analog_en[0] padframe/mprj_io_analog_pol[0] padframe/mprj_io_analog_sel[0]
+ padframe/mprj_io_dm[0] padframe/mprj_io_dm[1] padframe/mprj_io_dm[2] padframe/mprj_io_holdover[0]
+ padframe/mprj_io_ib_mode_sel[0] padframe/mprj_io_inp_dis[0] padframe/mprj_io_oeb[0]
+ padframe/mprj_io_out[0] padframe/mprj_io_slow_sel[0] padframe/mprj_io_vtrip_sel[0]
+ padframe/mprj_io_in[0] mprj/io_in_3v3[0] mprj/gpio_analog[3] mprj/gpio_noesd[3]
+ mprj_io[10] padframe/mprj_io_analog_en[10] padframe/mprj_io_analog_pol[10] padframe/mprj_io_analog_sel[10]
+ padframe/mprj_io_dm[30] padframe/mprj_io_dm[31] padframe/mprj_io_dm[32] padframe/mprj_io_holdover[10]
+ padframe/mprj_io_ib_mode_sel[10] padframe/mprj_io_inp_dis[10] padframe/mprj_io_oeb[10]
+ padframe/mprj_io_out[10] padframe/mprj_io_slow_sel[10] padframe/mprj_io_vtrip_sel[10]
+ padframe/mprj_io_in[10] mprj/io_in_3v3[10] mprj/gpio_analog[4] mprj/gpio_noesd[4]
+ mprj_io[11] padframe/mprj_io_analog_en[11] padframe/mprj_io_analog_pol[11] padframe/mprj_io_analog_sel[11]
+ padframe/mprj_io_dm[33] padframe/mprj_io_dm[34] padframe/mprj_io_dm[35] padframe/mprj_io_holdover[11]
+ padframe/mprj_io_ib_mode_sel[11] padframe/mprj_io_inp_dis[11] padframe/mprj_io_oeb[11]
+ padframe/mprj_io_out[11] padframe/mprj_io_slow_sel[11] padframe/mprj_io_vtrip_sel[11]
+ padframe/mprj_io_in[11] mprj/io_in_3v3[11] mprj/gpio_analog[5] mprj/gpio_noesd[5]
+ mprj_io[12] padframe/mprj_io_analog_en[12] padframe/mprj_io_analog_pol[12] padframe/mprj_io_analog_sel[12]
+ padframe/mprj_io_dm[36] padframe/mprj_io_dm[37] padframe/mprj_io_dm[38] padframe/mprj_io_holdover[12]
+ padframe/mprj_io_ib_mode_sel[12] padframe/mprj_io_inp_dis[12] padframe/mprj_io_oeb[12]
+ padframe/mprj_io_out[12] padframe/mprj_io_slow_sel[12] padframe/mprj_io_vtrip_sel[12]
+ padframe/mprj_io_in[12] mprj/io_in_3v3[12] mprj/gpio_analog[6] mprj/gpio_noesd[6]
+ mprj_io[13] padframe/mprj_io_analog_en[13] padframe/mprj_io_analog_pol[13] padframe/mprj_io_analog_sel[13]
+ padframe/mprj_io_dm[39] padframe/mprj_io_dm[40] padframe/mprj_io_dm[41] padframe/mprj_io_holdover[13]
+ padframe/mprj_io_ib_mode_sel[13] padframe/mprj_io_inp_dis[13] padframe/mprj_io_oeb[13]
+ padframe/mprj_io_out[13] padframe/mprj_io_slow_sel[13] padframe/mprj_io_vtrip_sel[13]
+ padframe/mprj_io_in[13] mprj/io_in_3v3[13] mprj_io[1] padframe/mprj_io_analog_en[1]
+ padframe/mprj_io_analog_pol[1] padframe/mprj_io_analog_sel[1] padframe/mprj_io_dm[3]
+ padframe/mprj_io_dm[4] padframe/mprj_io_dm[5] padframe/mprj_io_holdover[1] padframe/mprj_io_ib_mode_sel[1]
+ padframe/mprj_io_inp_dis[1] padframe/mprj_io_oeb[1] padframe/mprj_io_out[1] padframe/mprj_io_slow_sel[1]
+ padframe/mprj_io_vtrip_sel[1] padframe/mprj_io_in[1] mprj/io_in_3v3[1] mprj_io[2]
+ padframe/mprj_io_analog_en[2] padframe/mprj_io_analog_pol[2] padframe/mprj_io_analog_sel[2]
+ padframe/mprj_io_dm[6] padframe/mprj_io_dm[7] padframe/mprj_io_dm[8] padframe/mprj_io_holdover[2]
+ padframe/mprj_io_ib_mode_sel[2] padframe/mprj_io_inp_dis[2] padframe/mprj_io_oeb[2]
+ padframe/mprj_io_out[2] padframe/mprj_io_slow_sel[2] padframe/mprj_io_vtrip_sel[2]
+ padframe/mprj_io_in[2] mprj/io_in_3v3[2] mprj_io[3] padframe/mprj_io_analog_en[3]
+ padframe/mprj_io_analog_pol[3] padframe/mprj_io_analog_sel[3] padframe/mprj_io_dm[10]
+ padframe/mprj_io_dm[11] padframe/mprj_io_dm[9] padframe/mprj_io_holdover[3] padframe/mprj_io_ib_mode_sel[3]
+ padframe/mprj_io_inp_dis[3] padframe/mprj_io_oeb[3] padframe/mprj_io_out[3] padframe/mprj_io_slow_sel[3]
+ padframe/mprj_io_vtrip_sel[3] padframe/mprj_io_in[3] mprj/io_in_3v3[3] mprj_io[4]
+ padframe/mprj_io_analog_en[4] padframe/mprj_io_analog_pol[4] padframe/mprj_io_analog_sel[4]
+ padframe/mprj_io_dm[12] padframe/mprj_io_dm[13] padframe/mprj_io_dm[14] padframe/mprj_io_holdover[4]
+ padframe/mprj_io_ib_mode_sel[4] padframe/mprj_io_inp_dis[4] padframe/mprj_io_oeb[4]
+ padframe/mprj_io_out[4] padframe/mprj_io_slow_sel[4] padframe/mprj_io_vtrip_sel[4]
+ padframe/mprj_io_in[4] mprj/io_in_3v3[4] mprj_io[5] padframe/mprj_io_analog_en[5]
+ padframe/mprj_io_analog_pol[5] padframe/mprj_io_analog_sel[5] padframe/mprj_io_dm[15]
+ padframe/mprj_io_dm[16] padframe/mprj_io_dm[17] padframe/mprj_io_holdover[5] padframe/mprj_io_ib_mode_sel[5]
+ padframe/mprj_io_inp_dis[5] padframe/mprj_io_oeb[5] padframe/mprj_io_out[5] padframe/mprj_io_slow_sel[5]
+ padframe/mprj_io_vtrip_sel[5] padframe/mprj_io_in[5] mprj/io_in_3v3[5] mprj_io[6]
+ padframe/mprj_io_analog_en[6] padframe/mprj_io_analog_pol[6] padframe/mprj_io_analog_sel[6]
+ padframe/mprj_io_dm[18] padframe/mprj_io_dm[19] padframe/mprj_io_dm[20] padframe/mprj_io_holdover[6]
+ padframe/mprj_io_ib_mode_sel[6] padframe/mprj_io_inp_dis[6] padframe/mprj_io_oeb[6]
+ padframe/mprj_io_out[6] padframe/mprj_io_slow_sel[6] padframe/mprj_io_vtrip_sel[6]
+ padframe/mprj_io_in[6] mprj/io_in_3v3[6] mprj/gpio_analog[0] mprj/gpio_noesd[0]
+ mprj_io[7] padframe/mprj_io_analog_en[7] padframe/mprj_io_analog_pol[7] padframe/mprj_io_analog_sel[7]
+ padframe/mprj_io_dm[21] padframe/mprj_io_dm[22] padframe/mprj_io_dm[23] padframe/mprj_io_holdover[7]
+ padframe/mprj_io_ib_mode_sel[7] padframe/mprj_io_inp_dis[7] padframe/mprj_io_oeb[7]
+ padframe/mprj_io_out[7] padframe/mprj_io_slow_sel[7] padframe/mprj_io_vtrip_sel[7]
+ padframe/mprj_io_in[7] mprj/io_in_3v3[7] mprj/gpio_analog[1] mprj/gpio_noesd[1]
+ mprj_io[8] padframe/mprj_io_analog_en[8] padframe/mprj_io_analog_pol[8] padframe/mprj_io_analog_sel[8]
+ padframe/mprj_io_dm[24] padframe/mprj_io_dm[25] padframe/mprj_io_dm[26] padframe/mprj_io_holdover[8]
+ padframe/mprj_io_ib_mode_sel[8] padframe/mprj_io_inp_dis[8] padframe/mprj_io_oeb[8]
+ padframe/mprj_io_out[8] padframe/mprj_io_slow_sel[8] padframe/mprj_io_vtrip_sel[8]
+ padframe/mprj_io_in[8] mprj/io_in_3v3[8] mprj/gpio_analog[2] mprj/gpio_noesd[2]
+ mprj_io[9] padframe/mprj_io_analog_en[9] padframe/mprj_io_analog_pol[9] padframe/mprj_io_analog_sel[9]
+ padframe/mprj_io_dm[27] padframe/mprj_io_dm[28] padframe/mprj_io_dm[29] padframe/mprj_io_holdover[9]
+ padframe/mprj_io_ib_mode_sel[9] padframe/mprj_io_inp_dis[9] padframe/mprj_io_oeb[9]
+ padframe/mprj_io_out[9] padframe/mprj_io_slow_sel[9] padframe/mprj_io_vtrip_sel[9]
+ padframe/mprj_io_in[9] mprj/io_in_3v3[9] mprj/gpio_analog[7] mprj/gpio_noesd[7]
+ mprj_io[25] padframe/mprj_io_analog_en[14] padframe/mprj_io_analog_pol[14] padframe/mprj_io_analog_sel[14]
+ padframe/mprj_io_dm[42] padframe/mprj_io_dm[43] padframe/mprj_io_dm[44] padframe/mprj_io_holdover[14]
+ padframe/mprj_io_ib_mode_sel[14] padframe/mprj_io_inp_dis[14] padframe/mprj_io_oeb[14]
+ padframe/mprj_io_out[14] padframe/mprj_io_slow_sel[14] padframe/mprj_io_vtrip_sel[14]
+ padframe/mprj_io_in[14] mprj/io_in_3v3[14] mprj/gpio_analog[17] mprj/gpio_noesd[17]
+ mprj_io[35] padframe/mprj_io_analog_en[24] padframe/mprj_io_analog_pol[24] padframe/mprj_io_analog_sel[24]
+ padframe/mprj_io_dm[72] padframe/mprj_io_dm[73] padframe/mprj_io_dm[74] padframe/mprj_io_holdover[24]
+ padframe/mprj_io_ib_mode_sel[24] padframe/mprj_io_inp_dis[24] padframe/mprj_io_oeb[24]
+ padframe/mprj_io_out[24] padframe/mprj_io_slow_sel[24] padframe/mprj_io_vtrip_sel[24]
+ padframe/mprj_io_in[24] mprj/io_in_3v3[24] mprj_io[36] padframe/mprj_io_analog_en[25]
+ padframe/mprj_io_analog_pol[25] padframe/mprj_io_analog_sel[25] padframe/mprj_io_dm[75]
+ padframe/mprj_io_dm[76] padframe/mprj_io_dm[77] padframe/mprj_io_holdover[25] padframe/mprj_io_ib_mode_sel[25]
+ padframe/mprj_io_inp_dis[25] padframe/mprj_io_oeb[25] padframe/mprj_io_out[25] padframe/mprj_io_slow_sel[25]
+ padframe/mprj_io_vtrip_sel[25] padframe/mprj_io_in[25] mprj/io_in_3v3[25] mprj_io[37]
+ padframe/mprj_io_analog_en[26] padframe/mprj_io_analog_pol[26] padframe/mprj_io_analog_sel[26]
+ padframe/mprj_io_dm[78] padframe/mprj_io_dm[79] padframe/mprj_io_dm[80] padframe/mprj_io_holdover[26]
+ padframe/mprj_io_ib_mode_sel[26] padframe/mprj_io_inp_dis[26] padframe/mprj_io_oeb[26]
+ padframe/mprj_io_out[26] padframe/mprj_io_slow_sel[26] padframe/mprj_io_vtrip_sel[26]
+ padframe/mprj_io_in[26] mprj/io_in_3v3[26] mprj/gpio_analog[8] mprj/gpio_noesd[8]
+ mprj_io[26] padframe/mprj_io_analog_en[15] padframe/mprj_io_analog_pol[15] padframe/mprj_io_analog_sel[15]
+ padframe/mprj_io_dm[45] padframe/mprj_io_dm[46] padframe/mprj_io_dm[47] padframe/mprj_io_holdover[15]
+ padframe/mprj_io_ib_mode_sel[15] padframe/mprj_io_inp_dis[15] padframe/mprj_io_oeb[15]
+ padframe/mprj_io_out[15] padframe/mprj_io_slow_sel[15] padframe/mprj_io_vtrip_sel[15]
+ padframe/mprj_io_in[15] mprj/io_in_3v3[15] mprj/gpio_analog[9] mprj/gpio_noesd[9]
+ mprj_io[27] padframe/mprj_io_analog_en[16] padframe/mprj_io_analog_pol[16] padframe/mprj_io_analog_sel[16]
+ padframe/mprj_io_dm[48] padframe/mprj_io_dm[49] padframe/mprj_io_dm[50] padframe/mprj_io_holdover[16]
+ padframe/mprj_io_ib_mode_sel[16] padframe/mprj_io_inp_dis[16] padframe/mprj_io_oeb[16]
+ padframe/mprj_io_out[16] padframe/mprj_io_slow_sel[16] padframe/mprj_io_vtrip_sel[16]
+ padframe/mprj_io_in[16] mprj/io_in_3v3[16] mprj/gpio_analog[10] mprj/gpio_noesd[10]
+ mprj_io[28] padframe/mprj_io_analog_en[17] padframe/mprj_io_analog_pol[17] padframe/mprj_io_analog_sel[17]
+ padframe/mprj_io_dm[51] padframe/mprj_io_dm[52] padframe/mprj_io_dm[53] padframe/mprj_io_holdover[17]
+ padframe/mprj_io_ib_mode_sel[17] padframe/mprj_io_inp_dis[17] padframe/mprj_io_oeb[17]
+ padframe/mprj_io_out[17] padframe/mprj_io_slow_sel[17] padframe/mprj_io_vtrip_sel[17]
+ padframe/mprj_io_in[17] mprj/io_in_3v3[17] mprj/gpio_analog[11] mprj/gpio_noesd[11]
+ mprj_io[29] padframe/mprj_io_analog_en[18] padframe/mprj_io_analog_pol[18] padframe/mprj_io_analog_sel[18]
+ padframe/mprj_io_dm[54] padframe/mprj_io_dm[55] padframe/mprj_io_dm[56] padframe/mprj_io_holdover[18]
+ padframe/mprj_io_ib_mode_sel[18] padframe/mprj_io_inp_dis[18] padframe/mprj_io_oeb[18]
+ padframe/mprj_io_out[18] padframe/mprj_io_slow_sel[18] padframe/mprj_io_vtrip_sel[18]
+ padframe/mprj_io_in[18] mprj/io_in_3v3[18] mprj/gpio_analog[12] mprj/gpio_noesd[12]
+ mprj_io[30] padframe/mprj_io_analog_en[19] padframe/mprj_io_analog_pol[19] padframe/mprj_io_analog_sel[19]
+ padframe/mprj_io_dm[57] padframe/mprj_io_dm[58] padframe/mprj_io_dm[59] padframe/mprj_io_holdover[19]
+ padframe/mprj_io_ib_mode_sel[19] padframe/mprj_io_inp_dis[19] padframe/mprj_io_oeb[19]
+ padframe/mprj_io_out[19] padframe/mprj_io_slow_sel[19] padframe/mprj_io_vtrip_sel[19]
+ padframe/mprj_io_in[19] mprj/io_in_3v3[19] mprj/gpio_analog[13] mprj/gpio_noesd[13]
+ mprj_io[31] padframe/mprj_io_analog_en[20] padframe/mprj_io_analog_pol[20] padframe/mprj_io_analog_sel[20]
+ padframe/mprj_io_dm[60] padframe/mprj_io_dm[61] padframe/mprj_io_dm[62] padframe/mprj_io_holdover[20]
+ padframe/mprj_io_ib_mode_sel[20] padframe/mprj_io_inp_dis[20] padframe/mprj_io_oeb[20]
+ padframe/mprj_io_out[20] padframe/mprj_io_slow_sel[20] padframe/mprj_io_vtrip_sel[20]
+ padframe/mprj_io_in[20] mprj/io_in_3v3[20] mprj/gpio_analog[14] mprj/gpio_noesd[14]
+ mprj_io[32] padframe/mprj_io_analog_en[21] padframe/mprj_io_analog_pol[21] padframe/mprj_io_analog_sel[21]
+ padframe/mprj_io_dm[63] padframe/mprj_io_dm[64] padframe/mprj_io_dm[65] padframe/mprj_io_holdover[21]
+ padframe/mprj_io_ib_mode_sel[21] padframe/mprj_io_inp_dis[21] padframe/mprj_io_oeb[21]
+ padframe/mprj_io_out[21] padframe/mprj_io_slow_sel[21] padframe/mprj_io_vtrip_sel[21]
+ padframe/mprj_io_in[21] mprj/io_in_3v3[21] mprj/gpio_analog[15] mprj/gpio_noesd[15]
+ mprj_io[33] padframe/mprj_io_analog_en[22] padframe/mprj_io_analog_pol[22] padframe/mprj_io_analog_sel[22]
+ padframe/mprj_io_dm[66] padframe/mprj_io_dm[67] padframe/mprj_io_dm[68] padframe/mprj_io_holdover[22]
+ padframe/mprj_io_ib_mode_sel[22] padframe/mprj_io_inp_dis[22] padframe/mprj_io_oeb[22]
+ padframe/mprj_io_out[22] padframe/mprj_io_slow_sel[22] padframe/mprj_io_vtrip_sel[22]
+ padframe/mprj_io_in[22] mprj/io_in_3v3[22] mprj/gpio_analog[16] mprj/gpio_noesd[16]
+ mprj_io[34] padframe/mprj_io_analog_en[23] padframe/mprj_io_analog_pol[23] padframe/mprj_io_analog_sel[23]
+ padframe/mprj_io_dm[69] padframe/mprj_io_dm[70] padframe/mprj_io_dm[71] padframe/mprj_io_holdover[23]
+ padframe/mprj_io_ib_mode_sel[23] padframe/mprj_io_inp_dis[23] padframe/mprj_io_oeb[23]
+ padframe/mprj_io_out[23] padframe/mprj_io_slow_sel[23] padframe/mprj_io_vtrip_sel[23]
+ padframe/mprj_io_in[23] mprj/io_in_3v3[23] resetb rstb_level/A padframe/vdda mprj/io_analog[1]
+ mprj_io[15] mprj/io_analog[2] mprj_io[16] mprj/io_analog[3] mprj_io[17] mprj/io_analog[0]
+ mprj_io[14] mprj/io_analog[4] padframe/mprj_clamp_high[0] padframe/mprj_clamp_low[0]
+ mprj_io[18] vccd1 vdda1 vdda1_2 vssa1 vssa1_2 vccd1_core padframe/vdda1 padframe/vssa1
+ vssd1_core vssd1 mprj/io_analog[7] mprj_io[21] mprj/io_analog[8] mprj_io[22] mprj/io_analog[9]
+ mprj_io[23] mprj/io_analog[10] mprj_io[24] mprj/io_analog[5] padframe/mprj_clamp_high[1]
+ padframe/mprj_clamp_low[1] mprj_io[19] mprj/io_analog[6] padframe/mprj_clamp_high[2]
+ padframe/mprj_clamp_low[2] mprj_io[20] vccd2 vdda2 vssa2 vccd2_core padframe/vdda2
+ padframe/vssa2 vssd2_core vssd2 padframe/flash_csb_core padframe/flash_clk_oeb_core
+ padframe/flash_clk_core padframe/flash_csb_oeb_core padframe/mprj_io_one[0] padframe/mprj_io_one[1]
+ padframe/mprj_io_one[2] padframe/mprj_io_one[3] padframe/mprj_io_one[4] padframe/mprj_io_one[5]
+ padframe/mprj_io_one[6] padframe/mprj_io_one[7] padframe/mprj_io_one[8] padframe/mprj_io_one[9]
+ padframe/mprj_io_one[10] padframe/mprj_io_one[11] padframe/mprj_io_one[12] padframe/mprj_io_one[13]
+ padframe/mprj_io_one[14] padframe/mprj_io_one[15] padframe/mprj_io_one[16] padframe/mprj_io_one[17]
+ padframe/mprj_io_one[18] padframe/mprj_io_one[19] padframe/mprj_io_one[20] padframe/mprj_io_one[21]
+ padframe/mprj_io_one[22] padframe/mprj_io_one[23] padframe/mprj_io_one[24] padframe/mprj_io_one[25]
+ padframe/mprj_io_one[26] por/porb_h soc/gpio_mode1_pad padframe/vccd padframe/vddio
+ padframe/vssa padframe/vssd padframe/vssio chip_io_alt
Xgpio_defaults_block_13 gpio_defaults_block_13/VGND gpio_defaults_block_13/VPWR gpio_defaults_block_13/gpio_defaults[0]
+ gpio_defaults_block_13/gpio_defaults[10] gpio_defaults_block_13/gpio_defaults[11]
+ gpio_defaults_block_13/gpio_defaults[12] gpio_defaults_block_13/gpio_defaults[1]
+ gpio_defaults_block_13/gpio_defaults[2] gpio_defaults_block_13/gpio_defaults[3]
+ gpio_defaults_block_13/gpio_defaults[4] gpio_defaults_block_13/gpio_defaults[5]
+ gpio_defaults_block_13/gpio_defaults[6] gpio_defaults_block_13/gpio_defaults[7]
+ gpio_defaults_block_13/gpio_defaults[8] gpio_defaults_block_13/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_control_in_1a\[3\] gpio_defaults_block_5/gpio_defaults[0] gpio_defaults_block_5/gpio_defaults[10]
+ gpio_defaults_block_5/gpio_defaults[11] gpio_defaults_block_5/gpio_defaults[12]
+ gpio_defaults_block_5/gpio_defaults[1] gpio_defaults_block_5/gpio_defaults[2] gpio_defaults_block_5/gpio_defaults[3]
+ gpio_defaults_block_5/gpio_defaults[4] gpio_defaults_block_5/gpio_defaults[5] gpio_defaults_block_5/gpio_defaults[6]
+ gpio_defaults_block_5/gpio_defaults[7] gpio_defaults_block_5/gpio_defaults[8] gpio_defaults_block_5/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[5] padframe/mprj_io_one[5] housekeeping/mgmt_gpio_out[5]
+ padframe/mprj_io_one[5] padframe/mprj_io_analog_en[5] padframe/mprj_io_analog_pol[5]
+ padframe/mprj_io_analog_sel[5] padframe/mprj_io_dm[15] padframe/mprj_io_dm[16] padframe/mprj_io_dm[17]
+ padframe/mprj_io_holdover[5] padframe/mprj_io_ib_mode_sel[5] padframe/mprj_io_in[5]
+ padframe/mprj_io_inp_dis[5] padframe/mprj_io_out[5] padframe/mprj_io_oeb[5] padframe/mprj_io_slow_sel[5]
+ padframe/mprj_io_vtrip_sel[5] gpio_control_in_1a\[3\]/resetn gpio_control_in_1a\[4\]/resetn
+ gpio_control_in_1a\[3\]/serial_clock gpio_control_in_1a\[4\]/serial_clock gpio_control_in_1a\[3\]/serial_data_in
+ gpio_control_in_1a\[4\]/serial_data_in gpio_control_in_1a\[3\]/serial_load gpio_control_in_1a\[4\]/serial_load
+ mprj/io_in[5] mprj/io_oeb[5] mprj/io_out[5] gpio_defaults_block_5/VPWR vccd1_core
+ gpio_defaults_block_5/VGND vssd1_core gpio_control_in_1a\[3\]/zero gpio_control_block
Xgpio_defaults_block_35 gpio_defaults_block_35/VGND gpio_defaults_block_35/VPWR gpio_defaults_block_35/gpio_defaults[0]
+ gpio_defaults_block_35/gpio_defaults[10] gpio_defaults_block_35/gpio_defaults[11]
+ gpio_defaults_block_35/gpio_defaults[12] gpio_defaults_block_35/gpio_defaults[1]
+ gpio_defaults_block_35/gpio_defaults[2] gpio_defaults_block_35/gpio_defaults[3]
+ gpio_defaults_block_35/gpio_defaults[4] gpio_defaults_block_35/gpio_defaults[5]
+ gpio_defaults_block_35/gpio_defaults[6] gpio_defaults_block_35/gpio_defaults[7]
+ gpio_defaults_block_35/gpio_defaults[8] gpio_defaults_block_35/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_control_bidir_2\[0\] gpio_defaults_block_35/gpio_defaults[0] gpio_defaults_block_35/gpio_defaults[10]
+ gpio_defaults_block_35/gpio_defaults[11] gpio_defaults_block_35/gpio_defaults[12]
+ gpio_defaults_block_35/gpio_defaults[1] gpio_defaults_block_35/gpio_defaults[2]
+ gpio_defaults_block_35/gpio_defaults[3] gpio_defaults_block_35/gpio_defaults[4]
+ gpio_defaults_block_35/gpio_defaults[5] gpio_defaults_block_35/gpio_defaults[6]
+ gpio_defaults_block_35/gpio_defaults[7] gpio_defaults_block_35/gpio_defaults[8]
+ gpio_defaults_block_35/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[17] sigbuf/mgmt_io_oeb_buf[0]
+ sigbuf/mgmt_io_out_buf[17] padframe/mprj_io_one[24] padframe/mprj_io_analog_en[24]
+ padframe/mprj_io_analog_pol[24] padframe/mprj_io_analog_sel[24] padframe/mprj_io_dm[72]
+ padframe/mprj_io_dm[73] padframe/mprj_io_dm[74] padframe/mprj_io_holdover[24] padframe/mprj_io_ib_mode_sel[24]
+ padframe/mprj_io_in[24] padframe/mprj_io_inp_dis[24] padframe/mprj_io_out[24] padframe/mprj_io_oeb[24]
+ padframe/mprj_io_slow_sel[24] padframe/mprj_io_vtrip_sel[24] gpio_control_bidir_2\[0\]/resetn
+ gpio_control_in_2\[9\]/resetn gpio_control_bidir_2\[0\]/serial_clock gpio_control_in_2\[9\]/serial_clock
+ gpio_control_bidir_2\[0\]/serial_data_in gpio_control_in_2\[9\]/serial_data_in gpio_control_bidir_2\[0\]/serial_load
+ gpio_control_in_2\[9\]/serial_load mprj/io_in[24] mprj/io_oeb[24] mprj/io_out[24]
+ gpio_defaults_block_35/VPWR vccd1_core gpio_defaults_block_35/VGND vssd1_core gpio_control_bidir_2\[0\]/zero
+ gpio_control_block
Xsoc soc/VGND soc/VPWR soc/clk_in soc/clk_out soc/clk_in soc/resetn_in soc/debug_in
+ soc/debug_mode soc/debug_oeb soc/debug_out soc/flash_clk soc/flash_csb soc/flash_io0_di
+ soc/flash_io0_do soc/flash_io0_oeb soc/flash_io1_di soc/flash_io1_do soc/flash_io1_oeb
+ soc/flash_io2_di soc/flash_io2_do soc/flash_io2_oeb soc/flash_io3_di soc/flash_io3_do
+ soc/flash_io3_oeb soc/gpio_in_pad soc/gpio_inenb_pad soc/gpio_mode0_pad soc/gpio_mode1_pad
+ soc/gpio_out_pad soc/gpio_outenb_pad soc/hk_ack_i soc/hk_cyc_o soc/hk_dat_i[0] soc/hk_dat_i[10]
+ soc/hk_dat_i[11] soc/hk_dat_i[12] soc/hk_dat_i[13] soc/hk_dat_i[14] soc/hk_dat_i[15]
+ soc/hk_dat_i[16] soc/hk_dat_i[17] soc/hk_dat_i[18] soc/hk_dat_i[19] soc/hk_dat_i[1]
+ soc/hk_dat_i[20] soc/hk_dat_i[21] soc/hk_dat_i[22] soc/hk_dat_i[23] soc/hk_dat_i[24]
+ soc/hk_dat_i[25] soc/hk_dat_i[26] soc/hk_dat_i[27] soc/hk_dat_i[28] soc/hk_dat_i[29]
+ soc/hk_dat_i[2] soc/hk_dat_i[30] soc/hk_dat_i[31] soc/hk_dat_i[3] soc/hk_dat_i[4]
+ soc/hk_dat_i[5] soc/hk_dat_i[6] soc/hk_dat_i[7] soc/hk_dat_i[8] soc/hk_dat_i[9]
+ soc/hk_stb_o soc/irq[0] soc/irq[1] soc/irq[2] soc/irq[3] soc/irq[4] soc/irq[5] soc/la_iena[0]
+ soc/la_iena[100] soc/la_iena[101] soc/la_iena[102] soc/la_iena[103] soc/la_iena[104]
+ soc/la_iena[105] soc/la_iena[106] soc/la_iena[107] soc/la_iena[108] soc/la_iena[109]
+ soc/la_iena[10] soc/la_iena[110] soc/la_iena[111] soc/la_iena[112] soc/la_iena[113]
+ soc/la_iena[114] soc/la_iena[115] soc/la_iena[116] soc/la_iena[117] soc/la_iena[118]
+ soc/la_iena[119] soc/la_iena[11] soc/la_iena[120] soc/la_iena[121] soc/la_iena[122]
+ soc/la_iena[123] soc/la_iena[124] soc/la_iena[125] soc/la_iena[126] soc/la_iena[127]
+ soc/la_iena[12] soc/la_iena[13] soc/la_iena[14] soc/la_iena[15] soc/la_iena[16]
+ soc/la_iena[17] soc/la_iena[18] soc/la_iena[19] soc/la_iena[1] soc/la_iena[20] soc/la_iena[21]
+ soc/la_iena[22] soc/la_iena[23] soc/la_iena[24] soc/la_iena[25] soc/la_iena[26]
+ soc/la_iena[27] soc/la_iena[28] soc/la_iena[29] soc/la_iena[2] soc/la_iena[30] soc/la_iena[31]
+ soc/la_iena[32] soc/la_iena[33] soc/la_iena[34] soc/la_iena[35] soc/la_iena[36]
+ soc/la_iena[37] soc/la_iena[38] soc/la_iena[39] soc/la_iena[3] soc/la_iena[40] soc/la_iena[41]
+ soc/la_iena[42] soc/la_iena[43] soc/la_iena[44] soc/la_iena[45] soc/la_iena[46]
+ soc/la_iena[47] soc/la_iena[48] soc/la_iena[49] soc/la_iena[4] soc/la_iena[50] soc/la_iena[51]
+ soc/la_iena[52] soc/la_iena[53] soc/la_iena[54] soc/la_iena[55] soc/la_iena[56]
+ soc/la_iena[57] soc/la_iena[58] soc/la_iena[59] soc/la_iena[5] soc/la_iena[60] soc/la_iena[61]
+ soc/la_iena[62] soc/la_iena[63] soc/la_iena[64] soc/la_iena[65] soc/la_iena[66]
+ soc/la_iena[67] soc/la_iena[68] soc/la_iena[69] soc/la_iena[6] soc/la_iena[70] soc/la_iena[71]
+ soc/la_iena[72] soc/la_iena[73] soc/la_iena[74] soc/la_iena[75] soc/la_iena[76]
+ soc/la_iena[77] soc/la_iena[78] soc/la_iena[79] soc/la_iena[7] soc/la_iena[80] soc/la_iena[81]
+ soc/la_iena[82] soc/la_iena[83] soc/la_iena[84] soc/la_iena[85] soc/la_iena[86]
+ soc/la_iena[87] soc/la_iena[88] soc/la_iena[89] soc/la_iena[8] soc/la_iena[90] soc/la_iena[91]
+ soc/la_iena[92] soc/la_iena[93] soc/la_iena[94] soc/la_iena[95] soc/la_iena[96]
+ soc/la_iena[97] soc/la_iena[98] soc/la_iena[99] soc/la_iena[9] soc/la_input[0] soc/la_input[100]
+ soc/la_input[101] soc/la_input[102] soc/la_input[103] soc/la_input[104] soc/la_input[105]
+ soc/la_input[106] soc/la_input[107] soc/la_input[108] soc/la_input[109] soc/la_input[10]
+ soc/la_input[110] soc/la_input[111] soc/la_input[112] soc/la_input[113] soc/la_input[114]
+ soc/la_input[115] soc/la_input[116] soc/la_input[117] soc/la_input[118] soc/la_input[119]
+ soc/la_input[11] soc/la_input[120] soc/la_input[121] soc/la_input[122] soc/la_input[123]
+ soc/la_input[124] soc/la_input[125] soc/la_input[126] soc/la_input[127] soc/la_input[12]
+ soc/la_input[13] soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17]
+ soc/la_input[18] soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21]
+ soc/la_input[22] soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26]
+ soc/la_input[27] soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30]
+ soc/la_input[31] soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35]
+ soc/la_input[36] soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3]
+ soc/la_input[40] soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44]
+ soc/la_input[45] soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49]
+ soc/la_input[4] soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53]
+ soc/la_input[54] soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58]
+ soc/la_input[59] soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62]
+ soc/la_input[63] soc/la_input[64] soc/la_input[65] soc/la_input[66] soc/la_input[67]
+ soc/la_input[68] soc/la_input[69] soc/la_input[6] soc/la_input[70] soc/la_input[71]
+ soc/la_input[72] soc/la_input[73] soc/la_input[74] soc/la_input[75] soc/la_input[76]
+ soc/la_input[77] soc/la_input[78] soc/la_input[79] soc/la_input[7] soc/la_input[80]
+ soc/la_input[81] soc/la_input[82] soc/la_input[83] soc/la_input[84] soc/la_input[85]
+ soc/la_input[86] soc/la_input[87] soc/la_input[88] soc/la_input[89] soc/la_input[8]
+ soc/la_input[90] soc/la_input[91] soc/la_input[92] soc/la_input[93] soc/la_input[94]
+ soc/la_input[95] soc/la_input[96] soc/la_input[97] soc/la_input[98] soc/la_input[99]
+ soc/la_input[9] soc/la_oenb[0] soc/la_oenb[100] soc/la_oenb[101] soc/la_oenb[102]
+ soc/la_oenb[103] soc/la_oenb[104] soc/la_oenb[105] soc/la_oenb[106] soc/la_oenb[107]
+ soc/la_oenb[108] soc/la_oenb[109] soc/la_oenb[10] soc/la_oenb[110] soc/la_oenb[111]
+ soc/la_oenb[112] soc/la_oenb[113] soc/la_oenb[114] soc/la_oenb[115] soc/la_oenb[116]
+ soc/la_oenb[117] soc/la_oenb[118] soc/la_oenb[119] soc/la_oenb[11] soc/la_oenb[120]
+ soc/la_oenb[121] soc/la_oenb[122] soc/la_oenb[123] soc/la_oenb[124] soc/la_oenb[125]
+ soc/la_oenb[126] soc/la_oenb[127] soc/la_oenb[12] soc/la_oenb[13] soc/la_oenb[14]
+ soc/la_oenb[15] soc/la_oenb[16] soc/la_oenb[17] soc/la_oenb[18] soc/la_oenb[19]
+ soc/la_oenb[1] soc/la_oenb[20] soc/la_oenb[21] soc/la_oenb[22] soc/la_oenb[23] soc/la_oenb[24]
+ soc/la_oenb[25] soc/la_oenb[26] soc/la_oenb[27] soc/la_oenb[28] soc/la_oenb[29]
+ soc/la_oenb[2] soc/la_oenb[30] soc/la_oenb[31] soc/la_oenb[32] soc/la_oenb[33] soc/la_oenb[34]
+ soc/la_oenb[35] soc/la_oenb[36] soc/la_oenb[37] soc/la_oenb[38] soc/la_oenb[39]
+ soc/la_oenb[3] soc/la_oenb[40] soc/la_oenb[41] soc/la_oenb[42] soc/la_oenb[43] soc/la_oenb[44]
+ soc/la_oenb[45] soc/la_oenb[46] soc/la_oenb[47] soc/la_oenb[48] soc/la_oenb[49]
+ soc/la_oenb[4] soc/la_oenb[50] soc/la_oenb[51] soc/la_oenb[52] soc/la_oenb[53] soc/la_oenb[54]
+ soc/la_oenb[55] soc/la_oenb[56] soc/la_oenb[57] soc/la_oenb[58] soc/la_oenb[59]
+ soc/la_oenb[5] soc/la_oenb[60] soc/la_oenb[61] soc/la_oenb[62] soc/la_oenb[63] soc/la_oenb[64]
+ soc/la_oenb[65] soc/la_oenb[66] soc/la_oenb[67] soc/la_oenb[68] soc/la_oenb[69]
+ soc/la_oenb[6] soc/la_oenb[70] soc/la_oenb[71] soc/la_oenb[72] soc/la_oenb[73] soc/la_oenb[74]
+ soc/la_oenb[75] soc/la_oenb[76] soc/la_oenb[77] soc/la_oenb[78] soc/la_oenb[79]
+ soc/la_oenb[7] soc/la_oenb[80] soc/la_oenb[81] soc/la_oenb[82] soc/la_oenb[83] soc/la_oenb[84]
+ soc/la_oenb[85] soc/la_oenb[86] soc/la_oenb[87] soc/la_oenb[88] soc/la_oenb[89]
+ soc/la_oenb[8] soc/la_oenb[90] soc/la_oenb[91] soc/la_oenb[92] soc/la_oenb[93] soc/la_oenb[94]
+ soc/la_oenb[95] soc/la_oenb[96] soc/la_oenb[97] soc/la_oenb[98] soc/la_oenb[99]
+ soc/la_oenb[9] soc/la_output[0] soc/la_output[100] soc/la_output[101] soc/la_output[102]
+ soc/la_output[103] soc/la_output[104] soc/la_output[105] soc/la_output[106] soc/la_output[107]
+ soc/la_output[108] soc/la_output[109] soc/la_output[10] soc/la_output[110] soc/la_output[111]
+ soc/la_output[112] soc/la_output[113] soc/la_output[114] soc/la_output[115] soc/la_output[116]
+ soc/la_output[117] soc/la_output[118] soc/la_output[119] soc/la_output[11] soc/la_output[120]
+ soc/la_output[121] soc/la_output[122] soc/la_output[123] soc/la_output[124] soc/la_output[125]
+ soc/la_output[126] soc/la_output[127] soc/la_output[12] soc/la_output[13] soc/la_output[14]
+ soc/la_output[15] soc/la_output[16] soc/la_output[17] soc/la_output[18] soc/la_output[19]
+ soc/la_output[1] soc/la_output[20] soc/la_output[21] soc/la_output[22] soc/la_output[23]
+ soc/la_output[24] soc/la_output[25] soc/la_output[26] soc/la_output[27] soc/la_output[28]
+ soc/la_output[29] soc/la_output[2] soc/la_output[30] soc/la_output[31] soc/la_output[32]
+ soc/la_output[33] soc/la_output[34] soc/la_output[35] soc/la_output[36] soc/la_output[37]
+ soc/la_output[38] soc/la_output[39] soc/la_output[3] soc/la_output[40] soc/la_output[41]
+ soc/la_output[42] soc/la_output[43] soc/la_output[44] soc/la_output[45] soc/la_output[46]
+ soc/la_output[47] soc/la_output[48] soc/la_output[49] soc/la_output[4] soc/la_output[50]
+ soc/la_output[51] soc/la_output[52] soc/la_output[53] soc/la_output[54] soc/la_output[55]
+ soc/la_output[56] soc/la_output[57] soc/la_output[58] soc/la_output[59] soc/la_output[5]
+ soc/la_output[60] soc/la_output[61] soc/la_output[62] soc/la_output[63] soc/la_output[64]
+ soc/la_output[65] soc/la_output[66] soc/la_output[67] soc/la_output[68] soc/la_output[69]
+ soc/la_output[6] soc/la_output[70] soc/la_output[71] soc/la_output[72] soc/la_output[73]
+ soc/la_output[74] soc/la_output[75] soc/la_output[76] soc/la_output[77] soc/la_output[78]
+ soc/la_output[79] soc/la_output[7] soc/la_output[80] soc/la_output[81] soc/la_output[82]
+ soc/la_output[83] soc/la_output[84] soc/la_output[85] soc/la_output[86] soc/la_output[87]
+ soc/la_output[88] soc/la_output[89] soc/la_output[8] soc/la_output[90] soc/la_output[91]
+ soc/la_output[92] soc/la_output[93] soc/la_output[94] soc/la_output[95] soc/la_output[96]
+ soc/la_output[97] soc/la_output[98] soc/la_output[99] soc/la_output[9] soc/mprj_ack_i
+ soc/mprj_adr_o[0] soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13]
+ soc/mprj_adr_o[14] soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18]
+ soc/mprj_adr_o[19] soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22]
+ soc/mprj_adr_o[23] soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27]
+ soc/mprj_adr_o[28] soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31]
+ soc/mprj_adr_o[3] soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7]
+ soc/mprj_adr_o[8] soc/mprj_adr_o[9] soc/mprj_cyc_o soc/mprj_dat_i[0] soc/mprj_dat_i[10]
+ soc/mprj_dat_i[11] soc/mprj_dat_i[12] soc/mprj_dat_i[13] soc/mprj_dat_i[14] soc/mprj_dat_i[15]
+ soc/mprj_dat_i[16] soc/mprj_dat_i[17] soc/mprj_dat_i[18] soc/mprj_dat_i[19] soc/mprj_dat_i[1]
+ soc/mprj_dat_i[20] soc/mprj_dat_i[21] soc/mprj_dat_i[22] soc/mprj_dat_i[23] soc/mprj_dat_i[24]
+ soc/mprj_dat_i[25] soc/mprj_dat_i[26] soc/mprj_dat_i[27] soc/mprj_dat_i[28] soc/mprj_dat_i[29]
+ soc/mprj_dat_i[2] soc/mprj_dat_i[30] soc/mprj_dat_i[31] soc/mprj_dat_i[3] soc/mprj_dat_i[4]
+ soc/mprj_dat_i[5] soc/mprj_dat_i[6] soc/mprj_dat_i[7] soc/mprj_dat_i[8] soc/mprj_dat_i[9]
+ soc/mprj_dat_o[0] soc/mprj_dat_o[10] soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13]
+ soc/mprj_dat_o[14] soc/mprj_dat_o[15] soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18]
+ soc/mprj_dat_o[19] soc/mprj_dat_o[1] soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22]
+ soc/mprj_dat_o[23] soc/mprj_dat_o[24] soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27]
+ soc/mprj_dat_o[28] soc/mprj_dat_o[29] soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31]
+ soc/mprj_dat_o[3] soc/mprj_dat_o[4] soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7]
+ soc/mprj_dat_o[8] soc/mprj_dat_o[9] soc/mprj_sel_o[0] soc/mprj_sel_o[1] soc/mprj_sel_o[2]
+ soc/mprj_sel_o[3] soc/mprj_stb_o soc/mprj_wb_iena soc/mprj_we_o por/por_l padframe/por
+ por/por_l soc/porb_h_out soc/qspi_enabled soc/resetn_in soc/resetn_out rstb_level/X
+ pll/resetb soc/ser_rx soc/ser_tx soc/serial_clock_in soc/serial_clock_out soc/serial_data_2_in
+ soc/serial_data_2_out soc/serial_load_in soc/serial_load_out soc/serial_resetn_in
+ soc/serial_resetn_out soc/spi_csb soc/spi_enabled soc/spi_sck soc/spi_sdi soc/spi_sdo
+ soc/spi_sdoenb soc/trap soc/uart_enabled soc/user_irq_ena[0] soc/user_irq_ena[1]
+ soc/user_irq_ena[2] mgmt_core_wrapper
Xgpio_defaults_block_25 gpio_defaults_block_25/VGND gpio_defaults_block_25/VPWR gpio_defaults_block_25/gpio_defaults[0]
+ gpio_defaults_block_25/gpio_defaults[10] gpio_defaults_block_25/gpio_defaults[11]
+ gpio_defaults_block_25/gpio_defaults[12] gpio_defaults_block_25/gpio_defaults[1]
+ gpio_defaults_block_25/gpio_defaults[2] gpio_defaults_block_25/gpio_defaults[3]
+ gpio_defaults_block_25/gpio_defaults[4] gpio_defaults_block_25/gpio_defaults[5]
+ gpio_defaults_block_25/gpio_defaults[6] gpio_defaults_block_25/gpio_defaults[7]
+ gpio_defaults_block_25/gpio_defaults[8] gpio_defaults_block_25/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_control_in_2\[9\] gpio_defaults_block_34/gpio_defaults[0] gpio_defaults_block_34/gpio_defaults[10]
+ gpio_defaults_block_34/gpio_defaults[11] gpio_defaults_block_34/gpio_defaults[12]
+ gpio_defaults_block_34/gpio_defaults[1] gpio_defaults_block_34/gpio_defaults[2]
+ gpio_defaults_block_34/gpio_defaults[3] gpio_defaults_block_34/gpio_defaults[4]
+ gpio_defaults_block_34/gpio_defaults[5] gpio_defaults_block_34/gpio_defaults[6]
+ gpio_defaults_block_34/gpio_defaults[7] gpio_defaults_block_34/gpio_defaults[8]
+ gpio_defaults_block_34/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[16] padframe/mprj_io_one[23]
+ sigbuf/mgmt_io_out_buf[16] padframe/mprj_io_one[23] padframe/mprj_io_analog_en[23]
+ padframe/mprj_io_analog_pol[23] padframe/mprj_io_analog_sel[23] padframe/mprj_io_dm[69]
+ padframe/mprj_io_dm[70] padframe/mprj_io_dm[71] padframe/mprj_io_holdover[23] padframe/mprj_io_ib_mode_sel[23]
+ padframe/mprj_io_in[23] padframe/mprj_io_inp_dis[23] padframe/mprj_io_out[23] padframe/mprj_io_oeb[23]
+ padframe/mprj_io_slow_sel[23] padframe/mprj_io_vtrip_sel[23] gpio_control_in_2\[9\]/resetn
+ gpio_control_in_2\[8\]/resetn gpio_control_in_2\[9\]/serial_clock gpio_control_in_2\[8\]/serial_clock
+ gpio_control_in_2\[9\]/serial_data_in gpio_control_in_2\[8\]/serial_data_in gpio_control_in_2\[9\]/serial_load
+ gpio_control_in_2\[8\]/serial_load mprj/io_in[23] mprj/io_oeb[23] mprj/io_out[23]
+ sigbuf/vccd vccd1_core VSUBS vssd1_core gpio_control_in_2\[9\]/zero gpio_control_block
Xgpio_defaults_block_36 gpio_defaults_block_36/VGND gpio_defaults_block_36/VPWR gpio_defaults_block_36/gpio_defaults[0]
+ gpio_defaults_block_36/gpio_defaults[10] gpio_defaults_block_36/gpio_defaults[11]
+ gpio_defaults_block_36/gpio_defaults[12] gpio_defaults_block_36/gpio_defaults[1]
+ gpio_defaults_block_36/gpio_defaults[2] gpio_defaults_block_36/gpio_defaults[3]
+ gpio_defaults_block_36/gpio_defaults[4] gpio_defaults_block_36/gpio_defaults[5]
+ gpio_defaults_block_36/gpio_defaults[6] gpio_defaults_block_36/gpio_defaults[7]
+ gpio_defaults_block_36/gpio_defaults[8] gpio_defaults_block_36/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_defaults_block_26 gpio_defaults_block_26/VGND gpio_defaults_block_26/VPWR gpio_defaults_block_26/gpio_defaults[0]
+ gpio_defaults_block_26/gpio_defaults[10] gpio_defaults_block_26/gpio_defaults[11]
+ gpio_defaults_block_26/gpio_defaults[12] gpio_defaults_block_26/gpio_defaults[1]
+ gpio_defaults_block_26/gpio_defaults[2] gpio_defaults_block_26/gpio_defaults[3]
+ gpio_defaults_block_26/gpio_defaults[4] gpio_defaults_block_26/gpio_defaults[5]
+ gpio_defaults_block_26/gpio_defaults[6] gpio_defaults_block_26/gpio_defaults[7]
+ gpio_defaults_block_26/gpio_defaults[8] gpio_defaults_block_26/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_control_in_1\[4\] gpio_defaults_block_12/gpio_defaults[0] gpio_defaults_block_12/gpio_defaults[10]
+ gpio_defaults_block_12/gpio_defaults[11] gpio_defaults_block_12/gpio_defaults[12]
+ gpio_defaults_block_12/gpio_defaults[1] gpio_defaults_block_12/gpio_defaults[2]
+ gpio_defaults_block_12/gpio_defaults[3] gpio_defaults_block_12/gpio_defaults[4]
+ gpio_defaults_block_12/gpio_defaults[5] gpio_defaults_block_12/gpio_defaults[6]
+ gpio_defaults_block_12/gpio_defaults[7] gpio_defaults_block_12/gpio_defaults[8]
+ gpio_defaults_block_12/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[5] padframe/mprj_io_one[12]
+ sigbuf/mgmt_io_out_buf[5] padframe/mprj_io_one[12] padframe/mprj_io_analog_en[12]
+ padframe/mprj_io_analog_pol[12] padframe/mprj_io_analog_sel[12] padframe/mprj_io_dm[36]
+ padframe/mprj_io_dm[37] padframe/mprj_io_dm[38] padframe/mprj_io_holdover[12] padframe/mprj_io_ib_mode_sel[12]
+ padframe/mprj_io_in[12] padframe/mprj_io_inp_dis[12] padframe/mprj_io_out[12] padframe/mprj_io_oeb[12]
+ padframe/mprj_io_slow_sel[12] padframe/mprj_io_vtrip_sel[12] gpio_control_in_1\[4\]/resetn
+ gpio_control_in_1\[5\]/resetn gpio_control_in_1\[4\]/serial_clock gpio_control_in_1\[5\]/serial_clock
+ gpio_control_in_1\[4\]/serial_data_in gpio_control_in_1\[5\]/serial_data_in gpio_control_in_1\[4\]/serial_load
+ gpio_control_in_1\[5\]/serial_load mprj/io_in[12] mprj/io_oeb[12] mprj/io_out[12]
+ gpio_defaults_block_12/VPWR vccd1_core gpio_defaults_block_12/VGND vssd1_core gpio_control_in_1\[4\]/zero
+ gpio_control_block
Xgpio_defaults_block_37 gpio_defaults_block_37/VGND gpio_defaults_block_37/VPWR gpio_defaults_block_37/gpio_defaults[0]
+ gpio_defaults_block_37/gpio_defaults[10] gpio_defaults_block_37/gpio_defaults[11]
+ gpio_defaults_block_37/gpio_defaults[12] gpio_defaults_block_37/gpio_defaults[1]
+ gpio_defaults_block_37/gpio_defaults[2] gpio_defaults_block_37/gpio_defaults[3]
+ gpio_defaults_block_37/gpio_defaults[4] gpio_defaults_block_37/gpio_defaults[5]
+ gpio_defaults_block_37/gpio_defaults[6] gpio_defaults_block_37/gpio_defaults[7]
+ gpio_defaults_block_37/gpio_defaults[8] gpio_defaults_block_37/gpio_defaults[9]
+ gpio_defaults_block
Xpor soc/VPWR por/vdd3v3 por/vss3v3 por/porb_h por/por_l por/porb_l soc/VGND simple_por
Xgpio_defaults_block_27 gpio_defaults_block_27/VGND gpio_defaults_block_27/VPWR gpio_defaults_block_27/gpio_defaults[0]
+ gpio_defaults_block_27/gpio_defaults[10] gpio_defaults_block_27/gpio_defaults[11]
+ gpio_defaults_block_27/gpio_defaults[12] gpio_defaults_block_27/gpio_defaults[1]
+ gpio_defaults_block_27/gpio_defaults[2] gpio_defaults_block_27/gpio_defaults[3]
+ gpio_defaults_block_27/gpio_defaults[4] gpio_defaults_block_27/gpio_defaults[5]
+ gpio_defaults_block_27/gpio_defaults[6] gpio_defaults_block_27/gpio_defaults[7]
+ gpio_defaults_block_27/gpio_defaults[8] gpio_defaults_block_27/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_control_in_1a\[1\] gpio_defaults_block_3/gpio_defaults[0] gpio_defaults_block_3/gpio_defaults[10]
+ gpio_defaults_block_3/gpio_defaults[11] gpio_defaults_block_3/gpio_defaults[12]
+ gpio_defaults_block_3/gpio_defaults[1] gpio_defaults_block_3/gpio_defaults[2] gpio_defaults_block_3/gpio_defaults[3]
+ gpio_defaults_block_3/gpio_defaults[4] gpio_defaults_block_3/gpio_defaults[5] gpio_defaults_block_3/gpio_defaults[6]
+ gpio_defaults_block_3/gpio_defaults[7] gpio_defaults_block_3/gpio_defaults[8] gpio_defaults_block_3/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[3] padframe/mprj_io_one[3] housekeeping/mgmt_gpio_out[3]
+ padframe/mprj_io_one[3] padframe/mprj_io_analog_en[3] padframe/mprj_io_analog_pol[3]
+ padframe/mprj_io_analog_sel[3] padframe/mprj_io_dm[9] padframe/mprj_io_dm[10] padframe/mprj_io_dm[11]
+ padframe/mprj_io_holdover[3] padframe/mprj_io_ib_mode_sel[3] padframe/mprj_io_in[3]
+ padframe/mprj_io_inp_dis[3] padframe/mprj_io_out[3] padframe/mprj_io_oeb[3] padframe/mprj_io_slow_sel[3]
+ padframe/mprj_io_vtrip_sel[3] gpio_control_in_1a\[1\]/resetn gpio_control_in_1a\[2\]/resetn
+ gpio_control_in_1a\[1\]/serial_clock gpio_control_in_1a\[2\]/serial_clock gpio_control_in_1a\[1\]/serial_data_in
+ gpio_control_in_1a\[2\]/serial_data_in gpio_control_in_1a\[1\]/serial_load gpio_control_in_1a\[2\]/serial_load
+ mprj/io_in[3] mprj/io_oeb[3] mprj/io_out[3] gpio_defaults_block_3/VPWR vccd1_core
+ gpio_defaults_block_3/VGND vssd1_core gpio_control_in_1a\[1\]/zero gpio_control_block
Xclock_ctrl soc/VGND soc/VPWR clock_ctrl/core_clk pll/osc clock_ctrl/ext_clk_sel housekeeping/reset
+ pll/clockp[1] pll/clockp[0] pll/resetb housekeeping/wb_rstn_i clock_ctrl/sel2[0]
+ clock_ctrl/sel2[1] clock_ctrl/sel2[2] clock_ctrl/sel[0] clock_ctrl/sel[1] clock_ctrl/sel[2]
+ clock_ctrl/user_clk caravel_clocking
Xgpio_defaults_block_28 gpio_defaults_block_28/VGND gpio_defaults_block_28/VPWR gpio_defaults_block_28/gpio_defaults[0]
+ gpio_defaults_block_28/gpio_defaults[10] gpio_defaults_block_28/gpio_defaults[11]
+ gpio_defaults_block_28/gpio_defaults[12] gpio_defaults_block_28/gpio_defaults[1]
+ gpio_defaults_block_28/gpio_defaults[2] gpio_defaults_block_28/gpio_defaults[3]
+ gpio_defaults_block_28/gpio_defaults[4] gpio_defaults_block_28/gpio_defaults[5]
+ gpio_defaults_block_28/gpio_defaults[6] gpio_defaults_block_28/gpio_defaults[7]
+ gpio_defaults_block_28/gpio_defaults[8] gpio_defaults_block_28/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_control_in_2\[7\] gpio_defaults_block_32/gpio_defaults[0] gpio_defaults_block_32/gpio_defaults[10]
+ gpio_defaults_block_32/gpio_defaults[11] gpio_defaults_block_32/gpio_defaults[12]
+ gpio_defaults_block_32/gpio_defaults[1] gpio_defaults_block_32/gpio_defaults[2]
+ gpio_defaults_block_32/gpio_defaults[3] gpio_defaults_block_32/gpio_defaults[4]
+ gpio_defaults_block_32/gpio_defaults[5] gpio_defaults_block_32/gpio_defaults[6]
+ gpio_defaults_block_32/gpio_defaults[7] gpio_defaults_block_32/gpio_defaults[8]
+ gpio_defaults_block_32/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[14] padframe/mprj_io_one[21]
+ sigbuf/mgmt_io_out_buf[14] padframe/mprj_io_one[21] padframe/mprj_io_analog_en[21]
+ padframe/mprj_io_analog_pol[21] padframe/mprj_io_analog_sel[21] padframe/mprj_io_dm[63]
+ padframe/mprj_io_dm[64] padframe/mprj_io_dm[65] padframe/mprj_io_holdover[21] padframe/mprj_io_ib_mode_sel[21]
+ padframe/mprj_io_in[21] padframe/mprj_io_inp_dis[21] padframe/mprj_io_out[21] padframe/mprj_io_oeb[21]
+ padframe/mprj_io_slow_sel[21] padframe/mprj_io_vtrip_sel[21] gpio_control_in_2\[7\]/resetn
+ gpio_control_in_2\[6\]/resetn gpio_control_in_2\[7\]/serial_clock gpio_control_in_2\[6\]/serial_clock
+ gpio_control_in_2\[7\]/serial_data_in gpio_control_in_2\[6\]/serial_data_in gpio_control_in_2\[7\]/serial_load
+ gpio_control_in_2\[6\]/serial_load mprj/io_in[21] mprj/io_oeb[21] mprj/io_out[21]
+ gpio_defaults_block_32/VPWR vccd1_core gpio_defaults_block_32/VGND vssd1_core gpio_control_in_2\[7\]/zero
+ gpio_control_block
Xgpio_defaults_block_29 gpio_defaults_block_29/VGND gpio_defaults_block_29/VPWR gpio_defaults_block_29/gpio_defaults[0]
+ gpio_defaults_block_29/gpio_defaults[10] gpio_defaults_block_29/gpio_defaults[11]
+ gpio_defaults_block_29/gpio_defaults[12] gpio_defaults_block_29/gpio_defaults[1]
+ gpio_defaults_block_29/gpio_defaults[2] gpio_defaults_block_29/gpio_defaults[3]
+ gpio_defaults_block_29/gpio_defaults[4] gpio_defaults_block_29/gpio_defaults[5]
+ gpio_defaults_block_29/gpio_defaults[6] gpio_defaults_block_29/gpio_defaults[7]
+ gpio_defaults_block_29/gpio_defaults[8] gpio_defaults_block_29/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_control_in_1\[2\] gpio_defaults_block_10/gpio_defaults[0] gpio_defaults_block_10/gpio_defaults[10]
+ gpio_defaults_block_10/gpio_defaults[11] gpio_defaults_block_10/gpio_defaults[12]
+ gpio_defaults_block_10/gpio_defaults[1] gpio_defaults_block_10/gpio_defaults[2]
+ gpio_defaults_block_10/gpio_defaults[3] gpio_defaults_block_10/gpio_defaults[4]
+ gpio_defaults_block_10/gpio_defaults[5] gpio_defaults_block_10/gpio_defaults[6]
+ gpio_defaults_block_10/gpio_defaults[7] gpio_defaults_block_10/gpio_defaults[8]
+ gpio_defaults_block_10/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[3] padframe/mprj_io_one[10]
+ sigbuf/mgmt_io_out_buf[3] padframe/mprj_io_one[10] padframe/mprj_io_analog_en[10]
+ padframe/mprj_io_analog_pol[10] padframe/mprj_io_analog_sel[10] padframe/mprj_io_dm[30]
+ padframe/mprj_io_dm[31] padframe/mprj_io_dm[32] padframe/mprj_io_holdover[10] padframe/mprj_io_ib_mode_sel[10]
+ padframe/mprj_io_in[10] padframe/mprj_io_inp_dis[10] padframe/mprj_io_out[10] padframe/mprj_io_oeb[10]
+ padframe/mprj_io_slow_sel[10] padframe/mprj_io_vtrip_sel[10] gpio_control_in_1\[2\]/resetn
+ gpio_control_in_1\[3\]/resetn gpio_control_in_1\[2\]/serial_clock gpio_control_in_1\[3\]/serial_clock
+ gpio_control_in_1\[2\]/serial_data_in gpio_control_in_1\[3\]/serial_data_in gpio_control_in_1\[2\]/serial_load
+ gpio_control_in_1\[3\]/serial_load mprj/io_in[10] mprj/io_oeb[10] mprj/io_out[10]
+ gpio_defaults_block_10/VPWR vccd1_core gpio_defaults_block_10/VGND vssd1_core gpio_control_in_1\[2\]/zero
+ gpio_control_block
Xgpio_control_in_1\[0\] gpio_defaults_block_8/gpio_defaults[0] gpio_defaults_block_8/gpio_defaults[10]
+ gpio_defaults_block_8/gpio_defaults[11] gpio_defaults_block_8/gpio_defaults[12]
+ gpio_defaults_block_8/gpio_defaults[1] gpio_defaults_block_8/gpio_defaults[2] gpio_defaults_block_8/gpio_defaults[3]
+ gpio_defaults_block_8/gpio_defaults[4] gpio_defaults_block_8/gpio_defaults[5] gpio_defaults_block_8/gpio_defaults[6]
+ gpio_defaults_block_8/gpio_defaults[7] gpio_defaults_block_8/gpio_defaults[8] gpio_defaults_block_8/gpio_defaults[9]
+ sigbuf/mgmt_io_in_unbuf[1] padframe/mprj_io_one[8] sigbuf/mgmt_io_out_buf[1] padframe/mprj_io_one[8]
+ padframe/mprj_io_analog_en[8] padframe/mprj_io_analog_pol[8] padframe/mprj_io_analog_sel[8]
+ padframe/mprj_io_dm[24] padframe/mprj_io_dm[25] padframe/mprj_io_dm[26] padframe/mprj_io_holdover[8]
+ padframe/mprj_io_ib_mode_sel[8] padframe/mprj_io_in[8] padframe/mprj_io_inp_dis[8]
+ padframe/mprj_io_out[8] padframe/mprj_io_oeb[8] padframe/mprj_io_slow_sel[8] padframe/mprj_io_vtrip_sel[8]
+ gpio_control_in_1\[0\]/resetn gpio_control_in_1\[1\]/resetn gpio_control_in_1\[0\]/serial_clock
+ gpio_control_in_1\[1\]/serial_clock gpio_control_in_1\[0\]/serial_data_in gpio_control_in_1\[1\]/serial_data_in
+ gpio_control_in_1\[0\]/serial_load gpio_control_in_1\[1\]/serial_load mprj/io_in[8]
+ mprj/io_oeb[8] mprj/io_out[8] gpio_defaults_block_8/VPWR vccd1_core gpio_defaults_block_8/VGND
+ vssd1_core gpio_control_in_1\[0\]/zero gpio_control_block
Xgpio_control_in_2\[5\] gpio_defaults_block_30/gpio_defaults[0] gpio_defaults_block_30/gpio_defaults[10]
+ gpio_defaults_block_30/gpio_defaults[11] gpio_defaults_block_30/gpio_defaults[12]
+ gpio_defaults_block_30/gpio_defaults[1] gpio_defaults_block_30/gpio_defaults[2]
+ gpio_defaults_block_30/gpio_defaults[3] gpio_defaults_block_30/gpio_defaults[4]
+ gpio_defaults_block_30/gpio_defaults[5] gpio_defaults_block_30/gpio_defaults[6]
+ gpio_defaults_block_30/gpio_defaults[7] gpio_defaults_block_30/gpio_defaults[8]
+ gpio_defaults_block_30/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[12] padframe/mprj_io_one[19]
+ sigbuf/mgmt_io_out_buf[12] padframe/mprj_io_one[19] padframe/mprj_io_analog_en[19]
+ padframe/mprj_io_analog_pol[19] padframe/mprj_io_analog_sel[19] padframe/mprj_io_dm[57]
+ padframe/mprj_io_dm[58] padframe/mprj_io_dm[59] padframe/mprj_io_holdover[19] padframe/mprj_io_ib_mode_sel[19]
+ padframe/mprj_io_in[19] padframe/mprj_io_inp_dis[19] padframe/mprj_io_out[19] padframe/mprj_io_oeb[19]
+ padframe/mprj_io_slow_sel[19] padframe/mprj_io_vtrip_sel[19] gpio_control_in_2\[5\]/resetn
+ gpio_control_in_2\[4\]/resetn gpio_control_in_2\[5\]/serial_clock gpio_control_in_2\[4\]/serial_clock
+ gpio_control_in_2\[5\]/serial_data_in gpio_control_in_2\[4\]/serial_data_in gpio_control_in_2\[5\]/serial_load
+ gpio_control_in_2\[4\]/serial_load mprj/io_in[19] mprj/io_oeb[19] mprj/io_out[19]
+ sigbuf/vccd vccd1_core VSUBS vssd1_core gpio_control_in_2\[5\]/zero gpio_control_block
Xgpio_defaults_block_0 gpio_defaults_block_0/VGND gpio_defaults_block_0/VPWR gpio_defaults_block_0/gpio_defaults[0]
+ gpio_defaults_block_0/gpio_defaults[10] gpio_defaults_block_0/gpio_defaults[11]
+ gpio_defaults_block_0/gpio_defaults[12] gpio_defaults_block_0/gpio_defaults[1] gpio_defaults_block_0/gpio_defaults[2]
+ gpio_defaults_block_0/gpio_defaults[3] gpio_defaults_block_0/gpio_defaults[4] gpio_defaults_block_0/gpio_defaults[5]
+ gpio_defaults_block_0/gpio_defaults[6] gpio_defaults_block_0/gpio_defaults[7] gpio_defaults_block_0/gpio_defaults[8]
+ gpio_defaults_block_0/gpio_defaults[9] gpio_defaults_block
Xspare_logic\[3\] spare_logic\[3\]/spare_xfq[0] spare_logic\[3\]/spare_xfq[1] spare_logic\[3\]/spare_xfqn[0]
+ spare_logic\[3\]/spare_xfqn[1] spare_logic\[3\]/spare_xi[0] spare_logic\[3\]/spare_xi[1]
+ spare_logic\[3\]/spare_xi[2] spare_logic\[3\]/spare_xi[3] spare_logic\[3\]/spare_xib
+ spare_logic\[3\]/spare_xmx[0] spare_logic\[3\]/spare_xmx[1] spare_logic\[3\]/spare_xna[0]
+ spare_logic\[3\]/spare_xna[1] spare_logic\[3\]/spare_xno[0] spare_logic\[3\]/spare_xno[1]
+ spare_logic\[3\]/spare_xz[0] spare_logic\[3\]/spare_xz[10] spare_logic\[3\]/spare_xz[11]
+ spare_logic\[3\]/spare_xz[12] spare_logic\[3\]/spare_xz[13] spare_logic\[3\]/spare_xz[14]
+ spare_logic\[3\]/spare_xz[15] spare_logic\[3\]/spare_xz[16] spare_logic\[3\]/spare_xz[17]
+ spare_logic\[3\]/spare_xz[18] spare_logic\[3\]/spare_xz[19] spare_logic\[3\]/spare_xz[1]
+ spare_logic\[3\]/spare_xz[20] spare_logic\[3\]/spare_xz[21] spare_logic\[3\]/spare_xz[22]
+ spare_logic\[3\]/spare_xz[23] spare_logic\[3\]/spare_xz[24] spare_logic\[3\]/spare_xz[25]
+ spare_logic\[3\]/spare_xz[26] spare_logic\[3\]/spare_xz[2] spare_logic\[3\]/spare_xz[3]
+ spare_logic\[3\]/spare_xz[4] spare_logic\[3\]/spare_xz[5] spare_logic\[3\]/spare_xz[6]
+ spare_logic\[3\]/spare_xz[7] spare_logic\[3\]/spare_xz[8] spare_logic\[3\]/spare_xz[9]
+ soc/VPWR soc/VGND spare_logic_block
Xgpio_defaults_block_1 gpio_defaults_block_1/VGND gpio_defaults_block_1/VPWR gpio_defaults_block_1/gpio_defaults[0]
+ gpio_defaults_block_1/gpio_defaults[10] gpio_defaults_block_1/gpio_defaults[11]
+ gpio_defaults_block_1/gpio_defaults[12] gpio_defaults_block_1/gpio_defaults[1] gpio_defaults_block_1/gpio_defaults[2]
+ gpio_defaults_block_1/gpio_defaults[3] gpio_defaults_block_1/gpio_defaults[4] gpio_defaults_block_1/gpio_defaults[5]
+ gpio_defaults_block_1/gpio_defaults[6] gpio_defaults_block_1/gpio_defaults[7] gpio_defaults_block_1/gpio_defaults[8]
+ gpio_defaults_block_1/gpio_defaults[9] gpio_defaults_block
Xuser_id_value user_id_value/mask_rev[0] user_id_value/mask_rev[10] user_id_value/mask_rev[11]
+ user_id_value/mask_rev[12] user_id_value/mask_rev[13] user_id_value/mask_rev[14]
+ user_id_value/mask_rev[15] user_id_value/mask_rev[16] user_id_value/mask_rev[17]
+ user_id_value/mask_rev[18] user_id_value/mask_rev[19] user_id_value/mask_rev[1]
+ user_id_value/mask_rev[20] user_id_value/mask_rev[21] user_id_value/mask_rev[22]
+ user_id_value/mask_rev[23] user_id_value/mask_rev[24] user_id_value/mask_rev[25]
+ user_id_value/mask_rev[26] user_id_value/mask_rev[27] user_id_value/mask_rev[28]
+ user_id_value/mask_rev[29] user_id_value/mask_rev[2] user_id_value/mask_rev[30]
+ user_id_value/mask_rev[31] user_id_value/mask_rev[3] user_id_value/mask_rev[4] user_id_value/mask_rev[5]
+ user_id_value/mask_rev[6] user_id_value/mask_rev[7] user_id_value/mask_rev[8] user_id_value/mask_rev[9]
+ soc/VPWR soc/VGND user_id_programming
Xgpio_control_in_2\[3\] gpio_defaults_block_28/gpio_defaults[0] gpio_defaults_block_28/gpio_defaults[10]
+ gpio_defaults_block_28/gpio_defaults[11] gpio_defaults_block_28/gpio_defaults[12]
+ gpio_defaults_block_28/gpio_defaults[1] gpio_defaults_block_28/gpio_defaults[2]
+ gpio_defaults_block_28/gpio_defaults[3] gpio_defaults_block_28/gpio_defaults[4]
+ gpio_defaults_block_28/gpio_defaults[5] gpio_defaults_block_28/gpio_defaults[6]
+ gpio_defaults_block_28/gpio_defaults[7] gpio_defaults_block_28/gpio_defaults[8]
+ gpio_defaults_block_28/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[10] padframe/mprj_io_one[17]
+ sigbuf/mgmt_io_out_buf[10] padframe/mprj_io_one[17] padframe/mprj_io_analog_en[17]
+ padframe/mprj_io_analog_pol[17] padframe/mprj_io_analog_sel[17] padframe/mprj_io_dm[51]
+ padframe/mprj_io_dm[52] padframe/mprj_io_dm[53] padframe/mprj_io_holdover[17] padframe/mprj_io_ib_mode_sel[17]
+ padframe/mprj_io_in[17] padframe/mprj_io_inp_dis[17] padframe/mprj_io_out[17] padframe/mprj_io_oeb[17]
+ padframe/mprj_io_slow_sel[17] padframe/mprj_io_vtrip_sel[17] gpio_control_in_2\[3\]/resetn
+ gpio_control_in_2\[2\]/resetn gpio_control_in_2\[3\]/serial_clock gpio_control_in_2\[2\]/serial_clock
+ gpio_control_in_2\[3\]/serial_data_in gpio_control_in_2\[2\]/serial_data_in gpio_control_in_2\[3\]/serial_load
+ gpio_control_in_2\[2\]/serial_load mprj/io_in[17] mprj/io_oeb[17] mprj/io_out[17]
+ gpio_defaults_block_28/VPWR vccd1_core gpio_defaults_block_28/VGND vssd1_core gpio_control_in_2\[3\]/zero
+ gpio_control_block
Xgpio_defaults_block_2 gpio_defaults_block_2/VGND gpio_defaults_block_2/VPWR gpio_defaults_block_2/gpio_defaults[0]
+ gpio_defaults_block_2/gpio_defaults[10] gpio_defaults_block_2/gpio_defaults[11]
+ gpio_defaults_block_2/gpio_defaults[12] gpio_defaults_block_2/gpio_defaults[1] gpio_defaults_block_2/gpio_defaults[2]
+ gpio_defaults_block_2/gpio_defaults[3] gpio_defaults_block_2/gpio_defaults[4] gpio_defaults_block_2/gpio_defaults[5]
+ gpio_defaults_block_2/gpio_defaults[6] gpio_defaults_block_2/gpio_defaults[7] gpio_defaults_block_2/gpio_defaults[8]
+ gpio_defaults_block_2/gpio_defaults[9] gpio_defaults_block
Xgpio_defaults_block_3 gpio_defaults_block_3/VGND gpio_defaults_block_3/VPWR gpio_defaults_block_3/gpio_defaults[0]
+ gpio_defaults_block_3/gpio_defaults[10] gpio_defaults_block_3/gpio_defaults[11]
+ gpio_defaults_block_3/gpio_defaults[12] gpio_defaults_block_3/gpio_defaults[1] gpio_defaults_block_3/gpio_defaults[2]
+ gpio_defaults_block_3/gpio_defaults[3] gpio_defaults_block_3/gpio_defaults[4] gpio_defaults_block_3/gpio_defaults[5]
+ gpio_defaults_block_3/gpio_defaults[6] gpio_defaults_block_3/gpio_defaults[7] gpio_defaults_block_3/gpio_defaults[8]
+ gpio_defaults_block_3/gpio_defaults[9] gpio_defaults_block
Xgpio_control_bidir_1\[0\] gpio_defaults_block_0/gpio_defaults[0] gpio_defaults_block_0/gpio_defaults[10]
+ gpio_defaults_block_0/gpio_defaults[11] gpio_defaults_block_0/gpio_defaults[12]
+ gpio_defaults_block_0/gpio_defaults[1] gpio_defaults_block_0/gpio_defaults[2] gpio_defaults_block_0/gpio_defaults[3]
+ gpio_defaults_block_0/gpio_defaults[4] gpio_defaults_block_0/gpio_defaults[5] gpio_defaults_block_0/gpio_defaults[6]
+ gpio_defaults_block_0/gpio_defaults[7] gpio_defaults_block_0/gpio_defaults[8] gpio_defaults_block_0/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[0] housekeeping/mgmt_gpio_oeb[0] housekeeping/mgmt_gpio_out[0]
+ padframe/mprj_io_one[0] padframe/mprj_io_analog_en[0] padframe/mprj_io_analog_pol[0]
+ padframe/mprj_io_analog_sel[0] padframe/mprj_io_dm[0] padframe/mprj_io_dm[1] padframe/mprj_io_dm[2]
+ padframe/mprj_io_holdover[0] padframe/mprj_io_ib_mode_sel[0] padframe/mprj_io_in[0]
+ padframe/mprj_io_inp_dis[0] padframe/mprj_io_out[0] padframe/mprj_io_oeb[0] padframe/mprj_io_slow_sel[0]
+ padframe/mprj_io_vtrip_sel[0] soc/serial_resetn_in gpio_control_bidir_1\[1\]/resetn
+ soc/serial_clock_in gpio_control_bidir_1\[1\]/serial_clock housekeeping/serial_data_1
+ gpio_control_bidir_1\[1\]/serial_data_in soc/serial_load_in gpio_control_bidir_1\[1\]/serial_load
+ mprj/io_in[0] mprj/io_oeb[0] mprj/io_out[0] gpio_defaults_block_0/VPWR vccd1_core
+ gpio_defaults_block_0/VGND vssd1_core housekeeping/mgmt_gpio_in[15] gpio_control_block
Xgpio_defaults_block_5 gpio_defaults_block_5/VGND gpio_defaults_block_5/VPWR gpio_defaults_block_5/gpio_defaults[0]
+ gpio_defaults_block_5/gpio_defaults[10] gpio_defaults_block_5/gpio_defaults[11]
+ gpio_defaults_block_5/gpio_defaults[12] gpio_defaults_block_5/gpio_defaults[1] gpio_defaults_block_5/gpio_defaults[2]
+ gpio_defaults_block_5/gpio_defaults[3] gpio_defaults_block_5/gpio_defaults[4] gpio_defaults_block_5/gpio_defaults[5]
+ gpio_defaults_block_5/gpio_defaults[6] gpio_defaults_block_5/gpio_defaults[7] gpio_defaults_block_5/gpio_defaults[8]
+ gpio_defaults_block_5/gpio_defaults[9] gpio_defaults_block
Xgpio_defaults_block_4 gpio_defaults_block_4/VGND gpio_defaults_block_4/VPWR gpio_defaults_block_4/gpio_defaults[0]
+ gpio_defaults_block_4/gpio_defaults[10] gpio_defaults_block_4/gpio_defaults[11]
+ gpio_defaults_block_4/gpio_defaults[12] gpio_defaults_block_4/gpio_defaults[1] gpio_defaults_block_4/gpio_defaults[2]
+ gpio_defaults_block_4/gpio_defaults[3] gpio_defaults_block_4/gpio_defaults[4] gpio_defaults_block_4/gpio_defaults[5]
+ gpio_defaults_block_4/gpio_defaults[6] gpio_defaults_block_4/gpio_defaults[7] gpio_defaults_block_4/gpio_defaults[8]
+ gpio_defaults_block_4/gpio_defaults[9] gpio_defaults_block
Xspare_logic\[1\] spare_logic\[1\]/spare_xfq[0] spare_logic\[1\]/spare_xfq[1] spare_logic\[1\]/spare_xfqn[0]
+ spare_logic\[1\]/spare_xfqn[1] spare_logic\[1\]/spare_xi[0] spare_logic\[1\]/spare_xi[1]
+ spare_logic\[1\]/spare_xi[2] spare_logic\[1\]/spare_xi[3] spare_logic\[1\]/spare_xib
+ spare_logic\[1\]/spare_xmx[0] spare_logic\[1\]/spare_xmx[1] spare_logic\[1\]/spare_xna[0]
+ spare_logic\[1\]/spare_xna[1] spare_logic\[1\]/spare_xno[0] spare_logic\[1\]/spare_xno[1]
+ spare_logic\[1\]/spare_xz[0] spare_logic\[1\]/spare_xz[10] spare_logic\[1\]/spare_xz[11]
+ spare_logic\[1\]/spare_xz[12] spare_logic\[1\]/spare_xz[13] spare_logic\[1\]/spare_xz[14]
+ spare_logic\[1\]/spare_xz[15] spare_logic\[1\]/spare_xz[16] spare_logic\[1\]/spare_xz[17]
+ spare_logic\[1\]/spare_xz[18] spare_logic\[1\]/spare_xz[19] spare_logic\[1\]/spare_xz[1]
+ spare_logic\[1\]/spare_xz[20] spare_logic\[1\]/spare_xz[21] spare_logic\[1\]/spare_xz[22]
+ spare_logic\[1\]/spare_xz[23] spare_logic\[1\]/spare_xz[24] spare_logic\[1\]/spare_xz[25]
+ spare_logic\[1\]/spare_xz[26] spare_logic\[1\]/spare_xz[2] spare_logic\[1\]/spare_xz[3]
+ spare_logic\[1\]/spare_xz[4] spare_logic\[1\]/spare_xz[5] spare_logic\[1\]/spare_xz[6]
+ spare_logic\[1\]/spare_xz[7] spare_logic\[1\]/spare_xz[8] spare_logic\[1\]/spare_xz[9]
+ soc/VPWR soc/VGND spare_logic_block
Xgpio_control_in_2\[1\] gpio_defaults_block_26/gpio_defaults[0] gpio_defaults_block_26/gpio_defaults[10]
+ gpio_defaults_block_26/gpio_defaults[11] gpio_defaults_block_26/gpio_defaults[12]
+ gpio_defaults_block_26/gpio_defaults[1] gpio_defaults_block_26/gpio_defaults[2]
+ gpio_defaults_block_26/gpio_defaults[3] gpio_defaults_block_26/gpio_defaults[4]
+ gpio_defaults_block_26/gpio_defaults[5] gpio_defaults_block_26/gpio_defaults[6]
+ gpio_defaults_block_26/gpio_defaults[7] gpio_defaults_block_26/gpio_defaults[8]
+ gpio_defaults_block_26/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[8] padframe/mprj_io_one[15]
+ sigbuf/mgmt_io_out_buf[8] padframe/mprj_io_one[15] padframe/mprj_io_analog_en[15]
+ padframe/mprj_io_analog_pol[15] padframe/mprj_io_analog_sel[15] padframe/mprj_io_dm[45]
+ padframe/mprj_io_dm[46] padframe/mprj_io_dm[47] padframe/mprj_io_holdover[15] padframe/mprj_io_ib_mode_sel[15]
+ padframe/mprj_io_in[15] padframe/mprj_io_inp_dis[15] padframe/mprj_io_out[15] padframe/mprj_io_oeb[15]
+ padframe/mprj_io_slow_sel[15] padframe/mprj_io_vtrip_sel[15] gpio_control_in_2\[1\]/resetn
+ gpio_control_in_2\[0\]/resetn gpio_control_in_2\[1\]/serial_clock gpio_control_in_2\[0\]/serial_clock
+ gpio_control_in_2\[1\]/serial_data_in gpio_control_in_2\[0\]/serial_data_in gpio_control_in_2\[1\]/serial_load
+ gpio_control_in_2\[0\]/serial_load mprj/io_in[15] mprj/io_oeb[15] mprj/io_out[15]
+ gpio_defaults_block_26/VPWR vccd1_core gpio_defaults_block_26/VGND vssd1_core gpio_control_in_2\[1\]/zero
+ gpio_control_block
Xgpio_defaults_block_6 gpio_defaults_block_6/VGND gpio_defaults_block_6/VPWR gpio_defaults_block_6/gpio_defaults[0]
+ gpio_defaults_block_6/gpio_defaults[10] gpio_defaults_block_6/gpio_defaults[11]
+ gpio_defaults_block_6/gpio_defaults[12] gpio_defaults_block_6/gpio_defaults[1] gpio_defaults_block_6/gpio_defaults[2]
+ gpio_defaults_block_6/gpio_defaults[3] gpio_defaults_block_6/gpio_defaults[4] gpio_defaults_block_6/gpio_defaults[5]
+ gpio_defaults_block_6/gpio_defaults[6] gpio_defaults_block_6/gpio_defaults[7] gpio_defaults_block_6/gpio_defaults[8]
+ gpio_defaults_block_6/gpio_defaults[9] gpio_defaults_block
Xgpio_defaults_block_7 gpio_defaults_block_7/VGND gpio_defaults_block_7/VPWR gpio_defaults_block_7/gpio_defaults[0]
+ gpio_defaults_block_7/gpio_defaults[10] gpio_defaults_block_7/gpio_defaults[11]
+ gpio_defaults_block_7/gpio_defaults[12] gpio_defaults_block_7/gpio_defaults[1] gpio_defaults_block_7/gpio_defaults[2]
+ gpio_defaults_block_7/gpio_defaults[3] gpio_defaults_block_7/gpio_defaults[4] gpio_defaults_block_7/gpio_defaults[5]
+ gpio_defaults_block_7/gpio_defaults[6] gpio_defaults_block_7/gpio_defaults[7] gpio_defaults_block_7/gpio_defaults[8]
+ gpio_defaults_block_7/gpio_defaults[9] gpio_defaults_block
Xsigbuf sigbuf/mgmt_io_in_unbuf[6] sigbuf/mgmt_io_out_buf[6] sigbuf/mgmt_io_in_unbuf[5]
+ sigbuf/mgmt_io_in_unbuf[4] sigbuf/mgmt_io_in_unbuf[3] sigbuf/mgmt_io_in_unbuf[2]
+ sigbuf/mgmt_io_in_unbuf[1] sigbuf/mgmt_io_in_unbuf[0] sigbuf/mgmt_io_out_buf[0]
+ sigbuf/mgmt_io_out_buf[1] sigbuf/mgmt_io_out_buf[2] sigbuf/mgmt_io_out_buf[3] sigbuf/mgmt_io_out_buf[4]
+ sigbuf/mgmt_io_out_buf[5] sigbuf/mgmt_io_out_unbuf[0] sigbuf/mgmt_io_out_unbuf[1]
+ sigbuf/mgmt_io_out_unbuf[2] sigbuf/mgmt_io_out_unbuf[3] sigbuf/mgmt_io_out_unbuf[4]
+ sigbuf/mgmt_io_out_unbuf[5] sigbuf/mgmt_io_out_unbuf[6] sigbuf/mgmt_io_in_buf[6]
+ sigbuf/mgmt_io_in_buf[5] sigbuf/mgmt_io_in_buf[4] sigbuf/mgmt_io_in_buf[3] sigbuf/mgmt_io_in_buf[2]
+ sigbuf/mgmt_io_in_buf[1] sigbuf/mgmt_io_in_buf[0] sigbuf/mgmt_io_out_buf[10] sigbuf/mgmt_io_out_buf[11]
+ sigbuf/mgmt_io_in_unbuf[11] sigbuf/mgmt_io_in_unbuf[10] sigbuf/mgmt_io_out_buf[12]
+ sigbuf/mgmt_io_out_buf[13] sigbuf/mgmt_io_out_buf[14] sigbuf/mgmt_io_out_buf[15]
+ sigbuf/mgmt_io_in_unbuf[15] sigbuf/mgmt_io_in_unbuf[14] sigbuf/mgmt_io_in_unbuf[13]
+ sigbuf/mgmt_io_in_unbuf[12] sigbuf/mgmt_io_out_buf[16] sigbuf/mgmt_io_out_buf[17]
+ sigbuf/mgmt_io_out_buf[18] sigbuf/mgmt_io_out_buf[19] sigbuf/mgmt_io_in_unbuf[19]
+ sigbuf/mgmt_io_in_unbuf[18] sigbuf/mgmt_io_in_unbuf[17] sigbuf/mgmt_io_in_unbuf[16]
+ sigbuf/mgmt_io_oeb_buf[0] sigbuf/mgmt_io_oeb_buf[1] sigbuf/mgmt_io_oeb_buf[2] sigbuf/mgmt_io_oeb_unbuf[2]
+ sigbuf/mgmt_io_oeb_unbuf[1] sigbuf/mgmt_io_oeb_unbuf[0] sigbuf/mgmt_io_in_buf[19]
+ sigbuf/mgmt_io_in_buf[18] sigbuf/mgmt_io_in_buf[17] sigbuf/mgmt_io_in_buf[16] sigbuf/mgmt_io_out_unbuf[16]
+ sigbuf/mgmt_io_out_unbuf[17] sigbuf/mgmt_io_out_unbuf[18] sigbuf/mgmt_io_out_unbuf[19]
+ sigbuf/mgmt_io_out_unbuf[15] sigbuf/mgmt_io_out_unbuf[14] sigbuf/mgmt_io_out_unbuf[13]
+ sigbuf/mgmt_io_out_unbuf[12] sigbuf/mgmt_io_out_unbuf[11] sigbuf/mgmt_io_out_unbuf[10]
+ sigbuf/mgmt_io_out_unbuf[9] sigbuf/mgmt_io_out_unbuf[8] sigbuf/mgmt_io_out_unbuf[7]
+ sigbuf/mgmt_io_in_buf[7] sigbuf/mgmt_io_in_buf[8] sigbuf/mgmt_io_in_buf[9] sigbuf/mgmt_io_in_buf[10]
+ sigbuf/mgmt_io_in_buf[11] sigbuf/mgmt_io_in_buf[12] sigbuf/mgmt_io_in_buf[13] sigbuf/mgmt_io_in_buf[14]
+ sigbuf/mgmt_io_in_buf[15] sigbuf/vccd sigbuf/mgmt_io_out_buf[9] sigbuf/mgmt_io_in_unbuf[9]
+ sigbuf/mgmt_io_out_buf[8] sigbuf/mgmt_io_in_unbuf[8] sigbuf/mgmt_io_out_buf[7] sigbuf/mgmt_io_in_unbuf[7]
+ VSUBS gpio_signal_buffering_alt
Xgpio_defaults_block_8 gpio_defaults_block_8/VGND gpio_defaults_block_8/VPWR gpio_defaults_block_8/gpio_defaults[0]
+ gpio_defaults_block_8/gpio_defaults[10] gpio_defaults_block_8/gpio_defaults[11]
+ gpio_defaults_block_8/gpio_defaults[12] gpio_defaults_block_8/gpio_defaults[1] gpio_defaults_block_8/gpio_defaults[2]
+ gpio_defaults_block_8/gpio_defaults[3] gpio_defaults_block_8/gpio_defaults[4] gpio_defaults_block_8/gpio_defaults[5]
+ gpio_defaults_block_8/gpio_defaults[6] gpio_defaults_block_8/gpio_defaults[7] gpio_defaults_block_8/gpio_defaults[8]
+ gpio_defaults_block_8/gpio_defaults[9] gpio_defaults_block
Xgpio_control_in_1a\[4\] gpio_defaults_block_6/gpio_defaults[0] gpio_defaults_block_6/gpio_defaults[10]
+ gpio_defaults_block_6/gpio_defaults[11] gpio_defaults_block_6/gpio_defaults[12]
+ gpio_defaults_block_6/gpio_defaults[1] gpio_defaults_block_6/gpio_defaults[2] gpio_defaults_block_6/gpio_defaults[3]
+ gpio_defaults_block_6/gpio_defaults[4] gpio_defaults_block_6/gpio_defaults[5] gpio_defaults_block_6/gpio_defaults[6]
+ gpio_defaults_block_6/gpio_defaults[7] gpio_defaults_block_6/gpio_defaults[8] gpio_defaults_block_6/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[6] padframe/mprj_io_one[6] housekeeping/mgmt_gpio_out[6]
+ padframe/mprj_io_one[6] padframe/mprj_io_analog_en[6] padframe/mprj_io_analog_pol[6]
+ padframe/mprj_io_analog_sel[6] padframe/mprj_io_dm[18] padframe/mprj_io_dm[19] padframe/mprj_io_dm[20]
+ padframe/mprj_io_holdover[6] padframe/mprj_io_ib_mode_sel[6] padframe/mprj_io_in[6]
+ padframe/mprj_io_inp_dis[6] padframe/mprj_io_out[6] padframe/mprj_io_oeb[6] padframe/mprj_io_slow_sel[6]
+ padframe/mprj_io_vtrip_sel[6] gpio_control_in_1a\[4\]/resetn gpio_control_in_1a\[5\]/resetn
+ gpio_control_in_1a\[4\]/serial_clock gpio_control_in_1a\[5\]/serial_clock gpio_control_in_1a\[4\]/serial_data_in
+ gpio_control_in_1a\[5\]/serial_data_in gpio_control_in_1a\[4\]/serial_load gpio_control_in_1a\[5\]/serial_load
+ mprj/io_in[6] mprj/io_oeb[6] mprj/io_out[6] gpio_defaults_block_6/VPWR vccd1_core
+ gpio_defaults_block_6/VGND vssd1_core gpio_control_in_1a\[4\]/zero gpio_control_block
Xmgmt_buffers soc/clk_out clock_ctrl/user_clk soc/resetn_out mprj/la_data_in[0] mprj/la_data_in[100]
+ mprj/la_data_in[101] mprj/la_data_in[102] mprj/la_data_in[103] mprj/la_data_in[104]
+ mprj/la_data_in[105] mprj/la_data_in[106] mprj/la_data_in[107] mprj/la_data_in[108]
+ mprj/la_data_in[109] mprj/la_data_in[10] mprj/la_data_in[110] mprj/la_data_in[111]
+ mprj/la_data_in[112] mprj/la_data_in[113] mprj/la_data_in[114] mprj/la_data_in[115]
+ mprj/la_data_in[116] mprj/la_data_in[117] mprj/la_data_in[118] mprj/la_data_in[119]
+ mprj/la_data_in[11] mprj/la_data_in[120] mprj/la_data_in[121] mprj/la_data_in[122]
+ mprj/la_data_in[123] mprj/la_data_in[124] mprj/la_data_in[125] mprj/la_data_in[126]
+ mprj/la_data_in[127] mprj/la_data_in[12] mprj/la_data_in[13] mprj/la_data_in[14]
+ mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17] mprj/la_data_in[18]
+ mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21] mprj/la_data_in[22]
+ mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25] mprj/la_data_in[26]
+ mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29] mprj/la_data_in[2] mprj/la_data_in[30]
+ mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33] mprj/la_data_in[34]
+ mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37] mprj/la_data_in[38]
+ mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41] mprj/la_data_in[42]
+ mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45] mprj/la_data_in[46]
+ mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49] mprj/la_data_in[4] mprj/la_data_in[50]
+ mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53] mprj/la_data_in[54]
+ mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57] mprj/la_data_in[58]
+ mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61] mprj/la_data_in[62]
+ mprj/la_data_in[63] mprj/la_data_in[64] mprj/la_data_in[65] mprj/la_data_in[66]
+ mprj/la_data_in[67] mprj/la_data_in[68] mprj/la_data_in[69] mprj/la_data_in[6] mprj/la_data_in[70]
+ mprj/la_data_in[71] mprj/la_data_in[72] mprj/la_data_in[73] mprj/la_data_in[74]
+ mprj/la_data_in[75] mprj/la_data_in[76] mprj/la_data_in[77] mprj/la_data_in[78]
+ mprj/la_data_in[79] mprj/la_data_in[7] mprj/la_data_in[80] mprj/la_data_in[81] mprj/la_data_in[82]
+ mprj/la_data_in[83] mprj/la_data_in[84] mprj/la_data_in[85] mprj/la_data_in[86]
+ mprj/la_data_in[87] mprj/la_data_in[88] mprj/la_data_in[89] mprj/la_data_in[8] mprj/la_data_in[90]
+ mprj/la_data_in[91] mprj/la_data_in[92] mprj/la_data_in[93] mprj/la_data_in[94]
+ mprj/la_data_in[95] mprj/la_data_in[96] mprj/la_data_in[97] mprj/la_data_in[98]
+ mprj/la_data_in[99] mprj/la_data_in[9] soc/la_input[0] soc/la_input[100] soc/la_input[101]
+ soc/la_input[102] soc/la_input[103] soc/la_input[104] soc/la_input[105] soc/la_input[106]
+ soc/la_input[107] soc/la_input[108] soc/la_input[109] soc/la_input[10] soc/la_input[110]
+ soc/la_input[111] soc/la_input[112] soc/la_input[113] soc/la_input[114] soc/la_input[115]
+ soc/la_input[116] soc/la_input[117] soc/la_input[118] soc/la_input[119] soc/la_input[11]
+ soc/la_input[120] soc/la_input[121] soc/la_input[122] soc/la_input[123] soc/la_input[124]
+ soc/la_input[125] soc/la_input[126] soc/la_input[127] soc/la_input[12] soc/la_input[13]
+ soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17] soc/la_input[18]
+ soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21] soc/la_input[22]
+ soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26] soc/la_input[27]
+ soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30] soc/la_input[31]
+ soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35] soc/la_input[36]
+ soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3] soc/la_input[40]
+ soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44] soc/la_input[45]
+ soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49] soc/la_input[4]
+ soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53] soc/la_input[54]
+ soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58] soc/la_input[59]
+ soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62] soc/la_input[63]
+ soc/la_input[64] soc/la_input[65] soc/la_input[66] soc/la_input[67] soc/la_input[68]
+ soc/la_input[69] soc/la_input[6] soc/la_input[70] soc/la_input[71] soc/la_input[72]
+ soc/la_input[73] soc/la_input[74] soc/la_input[75] soc/la_input[76] soc/la_input[77]
+ soc/la_input[78] soc/la_input[79] soc/la_input[7] soc/la_input[80] soc/la_input[81]
+ soc/la_input[82] soc/la_input[83] soc/la_input[84] soc/la_input[85] soc/la_input[86]
+ soc/la_input[87] soc/la_input[88] soc/la_input[89] soc/la_input[8] soc/la_input[90]
+ soc/la_input[91] soc/la_input[92] soc/la_input[93] soc/la_input[94] soc/la_input[95]
+ soc/la_input[96] soc/la_input[97] soc/la_input[98] soc/la_input[99] soc/la_input[9]
+ mprj/la_data_out[0] mprj/la_data_out[100] mprj/la_data_out[101] mprj/la_data_out[102]
+ mprj/la_data_out[103] mprj/la_data_out[104] mprj/la_data_out[105] mprj/la_data_out[106]
+ mprj/la_data_out[107] mprj/la_data_out[108] mprj/la_data_out[109] mprj/la_data_out[10]
+ mprj/la_data_out[110] mprj/la_data_out[111] mprj/la_data_out[112] mprj/la_data_out[113]
+ mprj/la_data_out[114] mprj/la_data_out[115] mprj/la_data_out[116] mprj/la_data_out[117]
+ mprj/la_data_out[118] mprj/la_data_out[119] mprj/la_data_out[11] mprj/la_data_out[120]
+ mprj/la_data_out[121] mprj/la_data_out[122] mprj/la_data_out[123] mprj/la_data_out[124]
+ mprj/la_data_out[125] mprj/la_data_out[126] mprj/la_data_out[127] mprj/la_data_out[12]
+ mprj/la_data_out[13] mprj/la_data_out[14] mprj/la_data_out[15] mprj/la_data_out[16]
+ mprj/la_data_out[17] mprj/la_data_out[18] mprj/la_data_out[19] mprj/la_data_out[1]
+ mprj/la_data_out[20] mprj/la_data_out[21] mprj/la_data_out[22] mprj/la_data_out[23]
+ mprj/la_data_out[24] mprj/la_data_out[25] mprj/la_data_out[26] mprj/la_data_out[27]
+ mprj/la_data_out[28] mprj/la_data_out[29] mprj/la_data_out[2] mprj/la_data_out[30]
+ mprj/la_data_out[31] mprj/la_data_out[32] mprj/la_data_out[33] mprj/la_data_out[34]
+ mprj/la_data_out[35] mprj/la_data_out[36] mprj/la_data_out[37] mprj/la_data_out[38]
+ mprj/la_data_out[39] mprj/la_data_out[3] mprj/la_data_out[40] mprj/la_data_out[41]
+ mprj/la_data_out[42] mprj/la_data_out[43] mprj/la_data_out[44] mprj/la_data_out[45]
+ mprj/la_data_out[46] mprj/la_data_out[47] mprj/la_data_out[48] mprj/la_data_out[49]
+ mprj/la_data_out[4] mprj/la_data_out[50] mprj/la_data_out[51] mprj/la_data_out[52]
+ mprj/la_data_out[53] mprj/la_data_out[54] mprj/la_data_out[55] mprj/la_data_out[56]
+ mprj/la_data_out[57] mprj/la_data_out[58] mprj/la_data_out[59] mprj/la_data_out[5]
+ mprj/la_data_out[60] mprj/la_data_out[61] mprj/la_data_out[62] mprj/la_data_out[63]
+ mprj/la_data_out[64] mprj/la_data_out[65] mprj/la_data_out[66] mprj/la_data_out[67]
+ mprj/la_data_out[68] mprj/la_data_out[69] mprj/la_data_out[6] mprj/la_data_out[70]
+ mprj/la_data_out[71] mprj/la_data_out[72] mprj/la_data_out[73] mprj/la_data_out[74]
+ mprj/la_data_out[75] mprj/la_data_out[76] mprj/la_data_out[77] mprj/la_data_out[78]
+ mprj/la_data_out[79] mprj/la_data_out[7] mprj/la_data_out[80] mprj/la_data_out[81]
+ mprj/la_data_out[82] mprj/la_data_out[83] mprj/la_data_out[84] mprj/la_data_out[85]
+ mprj/la_data_out[86] mprj/la_data_out[87] mprj/la_data_out[88] mprj/la_data_out[89]
+ mprj/la_data_out[8] mprj/la_data_out[90] mprj/la_data_out[91] mprj/la_data_out[92]
+ mprj/la_data_out[93] mprj/la_data_out[94] mprj/la_data_out[95] mprj/la_data_out[96]
+ mprj/la_data_out[97] mprj/la_data_out[98] mprj/la_data_out[99] mprj/la_data_out[9]
+ soc/la_output[0] soc/la_output[100] soc/la_output[101] soc/la_output[102] soc/la_output[103]
+ soc/la_output[104] soc/la_output[105] soc/la_output[106] soc/la_output[107] soc/la_output[108]
+ soc/la_output[109] soc/la_output[10] soc/la_output[110] soc/la_output[111] soc/la_output[112]
+ soc/la_output[113] soc/la_output[114] soc/la_output[115] soc/la_output[116] soc/la_output[117]
+ soc/la_output[118] soc/la_output[119] soc/la_output[11] soc/la_output[120] soc/la_output[121]
+ soc/la_output[122] soc/la_output[123] soc/la_output[124] soc/la_output[125] soc/la_output[126]
+ soc/la_output[127] soc/la_output[12] soc/la_output[13] soc/la_output[14] soc/la_output[15]
+ soc/la_output[16] soc/la_output[17] soc/la_output[18] soc/la_output[19] soc/la_output[1]
+ soc/la_output[20] soc/la_output[21] soc/la_output[22] soc/la_output[23] soc/la_output[24]
+ soc/la_output[25] soc/la_output[26] soc/la_output[27] soc/la_output[28] soc/la_output[29]
+ soc/la_output[2] soc/la_output[30] soc/la_output[31] soc/la_output[32] soc/la_output[33]
+ soc/la_output[34] soc/la_output[35] soc/la_output[36] soc/la_output[37] soc/la_output[38]
+ soc/la_output[39] soc/la_output[3] soc/la_output[40] soc/la_output[41] soc/la_output[42]
+ soc/la_output[43] soc/la_output[44] soc/la_output[45] soc/la_output[46] soc/la_output[47]
+ soc/la_output[48] soc/la_output[49] soc/la_output[4] soc/la_output[50] soc/la_output[51]
+ soc/la_output[52] soc/la_output[53] soc/la_output[54] soc/la_output[55] soc/la_output[56]
+ soc/la_output[57] soc/la_output[58] soc/la_output[59] soc/la_output[5] soc/la_output[60]
+ soc/la_output[61] soc/la_output[62] soc/la_output[63] soc/la_output[64] soc/la_output[65]
+ soc/la_output[66] soc/la_output[67] soc/la_output[68] soc/la_output[69] soc/la_output[6]
+ soc/la_output[70] soc/la_output[71] soc/la_output[72] soc/la_output[73] soc/la_output[74]
+ soc/la_output[75] soc/la_output[76] soc/la_output[77] soc/la_output[78] soc/la_output[79]
+ soc/la_output[7] soc/la_output[80] soc/la_output[81] soc/la_output[82] soc/la_output[83]
+ soc/la_output[84] soc/la_output[85] soc/la_output[86] soc/la_output[87] soc/la_output[88]
+ soc/la_output[89] soc/la_output[8] soc/la_output[90] soc/la_output[91] soc/la_output[92]
+ soc/la_output[93] soc/la_output[94] soc/la_output[95] soc/la_output[96] soc/la_output[97]
+ soc/la_output[98] soc/la_output[99] soc/la_output[9] soc/la_iena[0] soc/la_iena[100]
+ soc/la_iena[101] soc/la_iena[102] soc/la_iena[103] soc/la_iena[104] soc/la_iena[105]
+ soc/la_iena[106] soc/la_iena[107] soc/la_iena[108] soc/la_iena[109] soc/la_iena[10]
+ soc/la_iena[110] soc/la_iena[111] soc/la_iena[112] soc/la_iena[113] soc/la_iena[114]
+ soc/la_iena[115] soc/la_iena[116] soc/la_iena[117] soc/la_iena[118] soc/la_iena[119]
+ soc/la_iena[11] soc/la_iena[120] soc/la_iena[121] soc/la_iena[122] soc/la_iena[123]
+ soc/la_iena[124] soc/la_iena[125] soc/la_iena[126] soc/la_iena[127] soc/la_iena[12]
+ soc/la_iena[13] soc/la_iena[14] soc/la_iena[15] soc/la_iena[16] soc/la_iena[17]
+ soc/la_iena[18] soc/la_iena[19] soc/la_iena[1] soc/la_iena[20] soc/la_iena[21] soc/la_iena[22]
+ soc/la_iena[23] soc/la_iena[24] soc/la_iena[25] soc/la_iena[26] soc/la_iena[27]
+ soc/la_iena[28] soc/la_iena[29] soc/la_iena[2] soc/la_iena[30] soc/la_iena[31] soc/la_iena[32]
+ soc/la_iena[33] soc/la_iena[34] soc/la_iena[35] soc/la_iena[36] soc/la_iena[37]
+ soc/la_iena[38] soc/la_iena[39] soc/la_iena[3] soc/la_iena[40] soc/la_iena[41] soc/la_iena[42]
+ soc/la_iena[43] soc/la_iena[44] soc/la_iena[45] soc/la_iena[46] soc/la_iena[47]
+ soc/la_iena[48] soc/la_iena[49] soc/la_iena[4] soc/la_iena[50] soc/la_iena[51] soc/la_iena[52]
+ soc/la_iena[53] soc/la_iena[54] soc/la_iena[55] soc/la_iena[56] soc/la_iena[57]
+ soc/la_iena[58] soc/la_iena[59] soc/la_iena[5] soc/la_iena[60] soc/la_iena[61] soc/la_iena[62]
+ soc/la_iena[63] soc/la_iena[64] soc/la_iena[65] soc/la_iena[66] soc/la_iena[67]
+ soc/la_iena[68] soc/la_iena[69] soc/la_iena[6] soc/la_iena[70] soc/la_iena[71] soc/la_iena[72]
+ soc/la_iena[73] soc/la_iena[74] soc/la_iena[75] soc/la_iena[76] soc/la_iena[77]
+ soc/la_iena[78] soc/la_iena[79] soc/la_iena[7] soc/la_iena[80] soc/la_iena[81] soc/la_iena[82]
+ soc/la_iena[83] soc/la_iena[84] soc/la_iena[85] soc/la_iena[86] soc/la_iena[87]
+ soc/la_iena[88] soc/la_iena[89] soc/la_iena[8] soc/la_iena[90] soc/la_iena[91] soc/la_iena[92]
+ soc/la_iena[93] soc/la_iena[94] soc/la_iena[95] soc/la_iena[96] soc/la_iena[97]
+ soc/la_iena[98] soc/la_iena[99] soc/la_iena[9] mprj/la_oenb[0] mprj/la_oenb[100]
+ mprj/la_oenb[101] mprj/la_oenb[102] mprj/la_oenb[103] mprj/la_oenb[104] mprj/la_oenb[105]
+ mprj/la_oenb[106] mprj/la_oenb[107] mprj/la_oenb[108] mprj/la_oenb[109] mprj/la_oenb[10]
+ mprj/la_oenb[110] mprj/la_oenb[111] mprj/la_oenb[112] mprj/la_oenb[113] mprj/la_oenb[114]
+ mprj/la_oenb[115] mprj/la_oenb[116] mprj/la_oenb[117] mprj/la_oenb[118] mprj/la_oenb[119]
+ mprj/la_oenb[11] mprj/la_oenb[120] mprj/la_oenb[121] mprj/la_oenb[122] mprj/la_oenb[123]
+ mprj/la_oenb[124] mprj/la_oenb[125] mprj/la_oenb[126] mprj/la_oenb[127] mprj/la_oenb[12]
+ mprj/la_oenb[13] mprj/la_oenb[14] mprj/la_oenb[15] mprj/la_oenb[16] mprj/la_oenb[17]
+ mprj/la_oenb[18] mprj/la_oenb[19] mprj/la_oenb[1] mprj/la_oenb[20] mprj/la_oenb[21]
+ mprj/la_oenb[22] mprj/la_oenb[23] mprj/la_oenb[24] mprj/la_oenb[25] mprj/la_oenb[26]
+ mprj/la_oenb[27] mprj/la_oenb[28] mprj/la_oenb[29] mprj/la_oenb[2] mprj/la_oenb[30]
+ mprj/la_oenb[31] mprj/la_oenb[32] mprj/la_oenb[33] mprj/la_oenb[34] mprj/la_oenb[35]
+ mprj/la_oenb[36] mprj/la_oenb[37] mprj/la_oenb[38] mprj/la_oenb[39] mprj/la_oenb[3]
+ mprj/la_oenb[40] mprj/la_oenb[41] mprj/la_oenb[42] mprj/la_oenb[43] mprj/la_oenb[44]
+ mprj/la_oenb[45] mprj/la_oenb[46] mprj/la_oenb[47] mprj/la_oenb[48] mprj/la_oenb[49]
+ mprj/la_oenb[4] mprj/la_oenb[50] mprj/la_oenb[51] mprj/la_oenb[52] mprj/la_oenb[53]
+ mprj/la_oenb[54] mprj/la_oenb[55] mprj/la_oenb[56] mprj/la_oenb[57] mprj/la_oenb[58]
+ mprj/la_oenb[59] mprj/la_oenb[5] mprj/la_oenb[60] mprj/la_oenb[61] mprj/la_oenb[62]
+ mprj/la_oenb[63] mprj/la_oenb[64] mprj/la_oenb[65] mprj/la_oenb[66] mprj/la_oenb[67]
+ mprj/la_oenb[68] mprj/la_oenb[69] mprj/la_oenb[6] mprj/la_oenb[70] mprj/la_oenb[71]
+ mprj/la_oenb[72] mprj/la_oenb[73] mprj/la_oenb[74] mprj/la_oenb[75] mprj/la_oenb[76]
+ mprj/la_oenb[77] mprj/la_oenb[78] mprj/la_oenb[79] mprj/la_oenb[7] mprj/la_oenb[80]
+ mprj/la_oenb[81] mprj/la_oenb[82] mprj/la_oenb[83] mprj/la_oenb[84] mprj/la_oenb[85]
+ mprj/la_oenb[86] mprj/la_oenb[87] mprj/la_oenb[88] mprj/la_oenb[89] mprj/la_oenb[8]
+ mprj/la_oenb[90] mprj/la_oenb[91] mprj/la_oenb[92] mprj/la_oenb[93] mprj/la_oenb[94]
+ mprj/la_oenb[95] mprj/la_oenb[96] mprj/la_oenb[97] mprj/la_oenb[98] mprj/la_oenb[99]
+ mprj/la_oenb[9] soc/la_oenb[0] soc/la_oenb[100] soc/la_oenb[101] soc/la_oenb[102]
+ soc/la_oenb[103] soc/la_oenb[104] soc/la_oenb[105] soc/la_oenb[106] soc/la_oenb[107]
+ soc/la_oenb[108] soc/la_oenb[109] soc/la_oenb[10] soc/la_oenb[110] soc/la_oenb[111]
+ soc/la_oenb[112] soc/la_oenb[113] soc/la_oenb[114] soc/la_oenb[115] soc/la_oenb[116]
+ soc/la_oenb[117] soc/la_oenb[118] soc/la_oenb[119] soc/la_oenb[11] soc/la_oenb[120]
+ soc/la_oenb[121] soc/la_oenb[122] soc/la_oenb[123] soc/la_oenb[124] soc/la_oenb[125]
+ soc/la_oenb[126] soc/la_oenb[127] soc/la_oenb[12] soc/la_oenb[13] soc/la_oenb[14]
+ soc/la_oenb[15] soc/la_oenb[16] soc/la_oenb[17] soc/la_oenb[18] soc/la_oenb[19]
+ soc/la_oenb[1] soc/la_oenb[20] soc/la_oenb[21] soc/la_oenb[22] soc/la_oenb[23] soc/la_oenb[24]
+ soc/la_oenb[25] soc/la_oenb[26] soc/la_oenb[27] soc/la_oenb[28] soc/la_oenb[29]
+ soc/la_oenb[2] soc/la_oenb[30] soc/la_oenb[31] soc/la_oenb[32] soc/la_oenb[33] soc/la_oenb[34]
+ soc/la_oenb[35] soc/la_oenb[36] soc/la_oenb[37] soc/la_oenb[38] soc/la_oenb[39]
+ soc/la_oenb[3] soc/la_oenb[40] soc/la_oenb[41] soc/la_oenb[42] soc/la_oenb[43] soc/la_oenb[44]
+ soc/la_oenb[45] soc/la_oenb[46] soc/la_oenb[47] soc/la_oenb[48] soc/la_oenb[49]
+ soc/la_oenb[4] soc/la_oenb[50] soc/la_oenb[51] soc/la_oenb[52] soc/la_oenb[53] soc/la_oenb[54]
+ soc/la_oenb[55] soc/la_oenb[56] soc/la_oenb[57] soc/la_oenb[58] soc/la_oenb[59]
+ soc/la_oenb[5] soc/la_oenb[60] soc/la_oenb[61] soc/la_oenb[62] soc/la_oenb[63] soc/la_oenb[64]
+ soc/la_oenb[65] soc/la_oenb[66] soc/la_oenb[67] soc/la_oenb[68] soc/la_oenb[69]
+ soc/la_oenb[6] soc/la_oenb[70] soc/la_oenb[71] soc/la_oenb[72] soc/la_oenb[73] soc/la_oenb[74]
+ soc/la_oenb[75] soc/la_oenb[76] soc/la_oenb[77] soc/la_oenb[78] soc/la_oenb[79]
+ soc/la_oenb[7] soc/la_oenb[80] soc/la_oenb[81] soc/la_oenb[82] soc/la_oenb[83] soc/la_oenb[84]
+ soc/la_oenb[85] soc/la_oenb[86] soc/la_oenb[87] soc/la_oenb[88] soc/la_oenb[89]
+ soc/la_oenb[8] soc/la_oenb[90] soc/la_oenb[91] soc/la_oenb[92] soc/la_oenb[93] soc/la_oenb[94]
+ soc/la_oenb[95] soc/la_oenb[96] soc/la_oenb[97] soc/la_oenb[98] soc/la_oenb[99]
+ soc/la_oenb[9] soc/mprj_ack_i mprj/wbs_ack_o soc/mprj_adr_o[0] soc/mprj_adr_o[10]
+ soc/mprj_adr_o[11] soc/mprj_adr_o[12] soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15]
+ soc/mprj_adr_o[16] soc/mprj_adr_o[17] soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1]
+ soc/mprj_adr_o[20] soc/mprj_adr_o[21] soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24]
+ soc/mprj_adr_o[25] soc/mprj_adr_o[26] soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29]
+ soc/mprj_adr_o[2] soc/mprj_adr_o[30] soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4]
+ soc/mprj_adr_o[5] soc/mprj_adr_o[6] soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9]
+ mprj/wbs_adr_i[0] mprj/wbs_adr_i[10] mprj/wbs_adr_i[11] mprj/wbs_adr_i[12] mprj/wbs_adr_i[13]
+ mprj/wbs_adr_i[14] mprj/wbs_adr_i[15] mprj/wbs_adr_i[16] mprj/wbs_adr_i[17] mprj/wbs_adr_i[18]
+ mprj/wbs_adr_i[19] mprj/wbs_adr_i[1] mprj/wbs_adr_i[20] mprj/wbs_adr_i[21] mprj/wbs_adr_i[22]
+ mprj/wbs_adr_i[23] mprj/wbs_adr_i[24] mprj/wbs_adr_i[25] mprj/wbs_adr_i[26] mprj/wbs_adr_i[27]
+ mprj/wbs_adr_i[28] mprj/wbs_adr_i[29] mprj/wbs_adr_i[2] mprj/wbs_adr_i[30] mprj/wbs_adr_i[31]
+ mprj/wbs_adr_i[3] mprj/wbs_adr_i[4] mprj/wbs_adr_i[5] mprj/wbs_adr_i[6] mprj/wbs_adr_i[7]
+ mprj/wbs_adr_i[8] mprj/wbs_adr_i[9] soc/mprj_cyc_o mprj/wbs_cyc_i soc/mprj_dat_i[0]
+ soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12] soc/mprj_dat_i[13] soc/mprj_dat_i[14]
+ soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17] soc/mprj_dat_i[18] soc/mprj_dat_i[19]
+ soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21] soc/mprj_dat_i[22] soc/mprj_dat_i[23]
+ soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26] soc/mprj_dat_i[27] soc/mprj_dat_i[28]
+ soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30] soc/mprj_dat_i[31] soc/mprj_dat_i[3]
+ soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6] soc/mprj_dat_i[7] soc/mprj_dat_i[8]
+ soc/mprj_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10] mprj/wbs_dat_o[11] mprj/wbs_dat_o[12]
+ mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15] mprj/wbs_dat_o[16] mprj/wbs_dat_o[17]
+ mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1] mprj/wbs_dat_o[20] mprj/wbs_dat_o[21]
+ mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24] mprj/wbs_dat_o[25] mprj/wbs_dat_o[26]
+ mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29] mprj/wbs_dat_o[2] mprj/wbs_dat_o[30]
+ mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4] mprj/wbs_dat_o[5] mprj/wbs_dat_o[6]
+ mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9] soc/mprj_dat_o[0] soc/mprj_dat_o[10]
+ soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15]
+ soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1]
+ soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24]
+ soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29]
+ soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4]
+ soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9]
+ mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12] mprj/wbs_dat_i[13]
+ mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17] mprj/wbs_dat_i[18]
+ mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21] mprj/wbs_dat_i[22]
+ mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26] mprj/wbs_dat_i[27]
+ mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30] mprj/wbs_dat_i[31]
+ mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6] mprj/wbs_dat_i[7]
+ mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] soc/mprj_wb_iena soc/mprj_sel_o[0] soc/mprj_sel_o[1]
+ soc/mprj_sel_o[2] soc/mprj_sel_o[3] mprj/wbs_sel_i[0] mprj/wbs_sel_i[1] mprj/wbs_sel_i[2]
+ mprj/wbs_sel_i[3] soc/mprj_stb_o mprj/wbs_stb_i soc/mprj_we_o mprj/wbs_we_i housekeeping/usr1_vcc_pwrgood
+ housekeeping/usr1_vdd_pwrgood housekeeping/usr2_vcc_pwrgood housekeeping/usr2_vdd_pwrgood
+ mprj/wb_clk_i mprj/user_clock2 soc/irq[0] soc/irq[1] soc/irq[2] mprj/user_irq[0]
+ mprj/user_irq[1] mprj/user_irq[2] soc/user_irq_ena[0] soc/user_irq_ena[1] soc/user_irq_ena[2]
+ mprj/wb_rst_i soc/VPWR vccd1_core vccd2_core vdda1_core vdda2_core vssa1_core vssa2_core
+ soc/VGND vssd1_core vssd2_core mgmt_protect
Xrstb_level rstb_level/A rstb_level/X rstb_level/VPWR rstb_level/VGND soc/VPWR soc/VGND
+ xres_buf
Xgpio_defaults_block_9 gpio_defaults_block_9/VGND gpio_defaults_block_9/VPWR gpio_defaults_block_9/gpio_defaults[0]
+ gpio_defaults_block_9/gpio_defaults[10] gpio_defaults_block_9/gpio_defaults[11]
+ gpio_defaults_block_9/gpio_defaults[12] gpio_defaults_block_9/gpio_defaults[1] gpio_defaults_block_9/gpio_defaults[2]
+ gpio_defaults_block_9/gpio_defaults[3] gpio_defaults_block_9/gpio_defaults[4] gpio_defaults_block_9/gpio_defaults[5]
+ gpio_defaults_block_9/gpio_defaults[6] gpio_defaults_block_9/gpio_defaults[7] gpio_defaults_block_9/gpio_defaults[8]
+ gpio_defaults_block_9/gpio_defaults[9] gpio_defaults_block
Xgpio_control_bidir_2\[1\] gpio_defaults_block_36/gpio_defaults[0] gpio_defaults_block_36/gpio_defaults[10]
+ gpio_defaults_block_36/gpio_defaults[11] gpio_defaults_block_36/gpio_defaults[12]
+ gpio_defaults_block_36/gpio_defaults[1] gpio_defaults_block_36/gpio_defaults[2]
+ gpio_defaults_block_36/gpio_defaults[3] gpio_defaults_block_36/gpio_defaults[4]
+ gpio_defaults_block_36/gpio_defaults[5] gpio_defaults_block_36/gpio_defaults[6]
+ gpio_defaults_block_36/gpio_defaults[7] gpio_defaults_block_36/gpio_defaults[8]
+ gpio_defaults_block_36/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[18] sigbuf/mgmt_io_oeb_buf[1]
+ sigbuf/mgmt_io_out_buf[18] padframe/mprj_io_one[25] padframe/mprj_io_analog_en[25]
+ padframe/mprj_io_analog_pol[25] padframe/mprj_io_analog_sel[25] padframe/mprj_io_dm[75]
+ padframe/mprj_io_dm[76] padframe/mprj_io_dm[77] padframe/mprj_io_holdover[25] padframe/mprj_io_ib_mode_sel[25]
+ padframe/mprj_io_in[25] padframe/mprj_io_inp_dis[25] padframe/mprj_io_out[25] padframe/mprj_io_oeb[25]
+ padframe/mprj_io_slow_sel[25] padframe/mprj_io_vtrip_sel[25] gpio_control_bidir_2\[1\]/resetn
+ gpio_control_bidir_2\[0\]/resetn gpio_control_bidir_2\[1\]/serial_clock gpio_control_bidir_2\[0\]/serial_clock
+ gpio_control_bidir_2\[1\]/serial_data_in gpio_control_bidir_2\[0\]/serial_data_in
+ gpio_control_bidir_2\[1\]/serial_load gpio_control_bidir_2\[0\]/serial_load mprj/io_in[25]
+ mprj/io_oeb[25] mprj/io_out[25] gpio_defaults_block_36/VPWR vccd1_core gpio_defaults_block_36/VGND
+ vssd1_core gpio_control_bidir_2\[1\]/zero gpio_control_block
Xgpio_control_in_1\[5\] gpio_defaults_block_13/gpio_defaults[0] gpio_defaults_block_13/gpio_defaults[10]
+ gpio_defaults_block_13/gpio_defaults[11] gpio_defaults_block_13/gpio_defaults[12]
+ gpio_defaults_block_13/gpio_defaults[1] gpio_defaults_block_13/gpio_defaults[2]
+ gpio_defaults_block_13/gpio_defaults[3] gpio_defaults_block_13/gpio_defaults[4]
+ gpio_defaults_block_13/gpio_defaults[5] gpio_defaults_block_13/gpio_defaults[6]
+ gpio_defaults_block_13/gpio_defaults[7] gpio_defaults_block_13/gpio_defaults[8]
+ gpio_defaults_block_13/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[6] padframe/mprj_io_one[13]
+ sigbuf/mgmt_io_out_buf[6] padframe/mprj_io_one[13] padframe/mprj_io_analog_en[13]
+ padframe/mprj_io_analog_pol[13] padframe/mprj_io_analog_sel[13] padframe/mprj_io_dm[39]
+ padframe/mprj_io_dm[40] padframe/mprj_io_dm[41] padframe/mprj_io_holdover[13] padframe/mprj_io_ib_mode_sel[13]
+ padframe/mprj_io_in[13] padframe/mprj_io_inp_dis[13] padframe/mprj_io_out[13] padframe/mprj_io_oeb[13]
+ padframe/mprj_io_slow_sel[13] padframe/mprj_io_vtrip_sel[13] gpio_control_in_1\[5\]/resetn
+ gpio_control_in_1\[5\]/resetn_out gpio_control_in_1\[5\]/serial_clock gpio_control_in_1\[5\]/serial_clock_out
+ gpio_control_in_1\[5\]/serial_data_in gpio_control_in_1\[5\]/serial_data_out gpio_control_in_1\[5\]/serial_load
+ gpio_control_in_1\[5\]/serial_load_out mprj/io_in[13] mprj/io_oeb[13] mprj/io_out[13]
+ gpio_defaults_block_13/VPWR vccd1_core gpio_defaults_block_13/VGND vssd1_core gpio_control_in_1\[5\]/zero
+ gpio_control_block
Xgpio_control_in_1a\[2\] gpio_defaults_block_4/gpio_defaults[0] gpio_defaults_block_4/gpio_defaults[10]
+ gpio_defaults_block_4/gpio_defaults[11] gpio_defaults_block_4/gpio_defaults[12]
+ gpio_defaults_block_4/gpio_defaults[1] gpio_defaults_block_4/gpio_defaults[2] gpio_defaults_block_4/gpio_defaults[3]
+ gpio_defaults_block_4/gpio_defaults[4] gpio_defaults_block_4/gpio_defaults[5] gpio_defaults_block_4/gpio_defaults[6]
+ gpio_defaults_block_4/gpio_defaults[7] gpio_defaults_block_4/gpio_defaults[8] gpio_defaults_block_4/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[4] padframe/mprj_io_one[4] housekeeping/mgmt_gpio_out[4]
+ padframe/mprj_io_one[4] padframe/mprj_io_analog_en[4] padframe/mprj_io_analog_pol[4]
+ padframe/mprj_io_analog_sel[4] padframe/mprj_io_dm[12] padframe/mprj_io_dm[13] padframe/mprj_io_dm[14]
+ padframe/mprj_io_holdover[4] padframe/mprj_io_ib_mode_sel[4] padframe/mprj_io_in[4]
+ padframe/mprj_io_inp_dis[4] padframe/mprj_io_out[4] padframe/mprj_io_oeb[4] padframe/mprj_io_slow_sel[4]
+ padframe/mprj_io_vtrip_sel[4] gpio_control_in_1a\[2\]/resetn gpio_control_in_1a\[3\]/resetn
+ gpio_control_in_1a\[2\]/serial_clock gpio_control_in_1a\[3\]/serial_clock gpio_control_in_1a\[2\]/serial_data_in
+ gpio_control_in_1a\[3\]/serial_data_in gpio_control_in_1a\[2\]/serial_load gpio_control_in_1a\[3\]/serial_load
+ mprj/io_in[4] mprj/io_oeb[4] mprj/io_out[4] gpio_defaults_block_4/VPWR vccd1_core
+ gpio_defaults_block_4/VGND vssd1_core gpio_control_in_1a\[2\]/zero gpio_control_block
Xgpio_control_in_2\[8\] gpio_defaults_block_33/gpio_defaults[0] gpio_defaults_block_33/gpio_defaults[10]
+ gpio_defaults_block_33/gpio_defaults[11] gpio_defaults_block_33/gpio_defaults[12]
+ gpio_defaults_block_33/gpio_defaults[1] gpio_defaults_block_33/gpio_defaults[2]
+ gpio_defaults_block_33/gpio_defaults[3] gpio_defaults_block_33/gpio_defaults[4]
+ gpio_defaults_block_33/gpio_defaults[5] gpio_defaults_block_33/gpio_defaults[6]
+ gpio_defaults_block_33/gpio_defaults[7] gpio_defaults_block_33/gpio_defaults[8]
+ gpio_defaults_block_33/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[15] padframe/mprj_io_one[22]
+ sigbuf/mgmt_io_out_buf[15] padframe/mprj_io_one[22] padframe/mprj_io_analog_en[22]
+ padframe/mprj_io_analog_pol[22] padframe/mprj_io_analog_sel[22] padframe/mprj_io_dm[66]
+ padframe/mprj_io_dm[67] padframe/mprj_io_dm[68] padframe/mprj_io_holdover[22] padframe/mprj_io_ib_mode_sel[22]
+ padframe/mprj_io_in[22] padframe/mprj_io_inp_dis[22] padframe/mprj_io_out[22] padframe/mprj_io_oeb[22]
+ padframe/mprj_io_slow_sel[22] padframe/mprj_io_vtrip_sel[22] gpio_control_in_2\[8\]/resetn
+ gpio_control_in_2\[7\]/resetn gpio_control_in_2\[8\]/serial_clock gpio_control_in_2\[7\]/serial_clock
+ gpio_control_in_2\[8\]/serial_data_in gpio_control_in_2\[7\]/serial_data_in gpio_control_in_2\[8\]/serial_load
+ gpio_control_in_2\[7\]/serial_load mprj/io_in[22] mprj/io_oeb[22] mprj/io_out[22]
+ gpio_defaults_block_33/VPWR vccd1_core gpio_defaults_block_33/VGND vssd1_core gpio_control_in_2\[8\]/zero
+ gpio_control_block
Xgpio_control_in_1\[3\] gpio_defaults_block_11/gpio_defaults[0] gpio_defaults_block_11/gpio_defaults[10]
+ gpio_defaults_block_11/gpio_defaults[11] gpio_defaults_block_11/gpio_defaults[12]
+ gpio_defaults_block_11/gpio_defaults[1] gpio_defaults_block_11/gpio_defaults[2]
+ gpio_defaults_block_11/gpio_defaults[3] gpio_defaults_block_11/gpio_defaults[4]
+ gpio_defaults_block_11/gpio_defaults[5] gpio_defaults_block_11/gpio_defaults[6]
+ gpio_defaults_block_11/gpio_defaults[7] gpio_defaults_block_11/gpio_defaults[8]
+ gpio_defaults_block_11/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[4] padframe/mprj_io_one[11]
+ sigbuf/mgmt_io_out_buf[4] padframe/mprj_io_one[11] padframe/mprj_io_analog_en[11]
+ padframe/mprj_io_analog_pol[11] padframe/mprj_io_analog_sel[11] padframe/mprj_io_dm[33]
+ padframe/mprj_io_dm[34] padframe/mprj_io_dm[35] padframe/mprj_io_holdover[11] padframe/mprj_io_ib_mode_sel[11]
+ padframe/mprj_io_in[11] padframe/mprj_io_inp_dis[11] padframe/mprj_io_out[11] padframe/mprj_io_oeb[11]
+ padframe/mprj_io_slow_sel[11] padframe/mprj_io_vtrip_sel[11] gpio_control_in_1\[3\]/resetn
+ gpio_control_in_1\[4\]/resetn gpio_control_in_1\[3\]/serial_clock gpio_control_in_1\[4\]/serial_clock
+ gpio_control_in_1\[3\]/serial_data_in gpio_control_in_1\[4\]/serial_data_in gpio_control_in_1\[3\]/serial_load
+ gpio_control_in_1\[4\]/serial_load mprj/io_in[11] mprj/io_oeb[11] mprj/io_out[11]
+ gpio_defaults_block_11/VPWR vccd1_core gpio_defaults_block_11/VGND vssd1_core gpio_control_in_1\[3\]/zero
+ gpio_control_block
Xgpio_control_in_1a\[0\] gpio_defaults_block_2/gpio_defaults[0] gpio_defaults_block_2/gpio_defaults[10]
+ gpio_defaults_block_2/gpio_defaults[11] gpio_defaults_block_2/gpio_defaults[12]
+ gpio_defaults_block_2/gpio_defaults[1] gpio_defaults_block_2/gpio_defaults[2] gpio_defaults_block_2/gpio_defaults[3]
+ gpio_defaults_block_2/gpio_defaults[4] gpio_defaults_block_2/gpio_defaults[5] gpio_defaults_block_2/gpio_defaults[6]
+ gpio_defaults_block_2/gpio_defaults[7] gpio_defaults_block_2/gpio_defaults[8] gpio_defaults_block_2/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[2] padframe/mprj_io_one[2] housekeeping/mgmt_gpio_out[2]
+ padframe/mprj_io_one[2] padframe/mprj_io_analog_en[2] padframe/mprj_io_analog_pol[2]
+ padframe/mprj_io_analog_sel[2] padframe/mprj_io_dm[6] padframe/mprj_io_dm[7] padframe/mprj_io_dm[8]
+ padframe/mprj_io_holdover[2] padframe/mprj_io_ib_mode_sel[2] padframe/mprj_io_in[2]
+ padframe/mprj_io_inp_dis[2] padframe/mprj_io_out[2] padframe/mprj_io_oeb[2] padframe/mprj_io_slow_sel[2]
+ padframe/mprj_io_vtrip_sel[2] gpio_control_in_1a\[0\]/resetn gpio_control_in_1a\[1\]/resetn
+ gpio_control_in_1a\[0\]/serial_clock gpio_control_in_1a\[1\]/serial_clock gpio_control_in_1a\[0\]/serial_data_in
+ gpio_control_in_1a\[1\]/serial_data_in gpio_control_in_1a\[0\]/serial_load gpio_control_in_1a\[1\]/serial_load
+ mprj/io_in[2] mprj/io_oeb[2] mprj/io_out[2] gpio_defaults_block_2/VPWR vccd1_core
+ gpio_defaults_block_2/VGND vssd1_core gpio_control_in_1a\[0\]/zero gpio_control_block
Xgpio_control_in_2\[6\] gpio_defaults_block_31/gpio_defaults[0] gpio_defaults_block_31/gpio_defaults[10]
+ gpio_defaults_block_31/gpio_defaults[11] gpio_defaults_block_31/gpio_defaults[12]
+ gpio_defaults_block_31/gpio_defaults[1] gpio_defaults_block_31/gpio_defaults[2]
+ gpio_defaults_block_31/gpio_defaults[3] gpio_defaults_block_31/gpio_defaults[4]
+ gpio_defaults_block_31/gpio_defaults[5] gpio_defaults_block_31/gpio_defaults[6]
+ gpio_defaults_block_31/gpio_defaults[7] gpio_defaults_block_31/gpio_defaults[8]
+ gpio_defaults_block_31/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[13] padframe/mprj_io_one[20]
+ sigbuf/mgmt_io_out_buf[13] padframe/mprj_io_one[20] padframe/mprj_io_analog_en[20]
+ padframe/mprj_io_analog_pol[20] padframe/mprj_io_analog_sel[20] padframe/mprj_io_dm[60]
+ padframe/mprj_io_dm[61] padframe/mprj_io_dm[62] padframe/mprj_io_holdover[20] padframe/mprj_io_ib_mode_sel[20]
+ padframe/mprj_io_in[20] padframe/mprj_io_inp_dis[20] padframe/mprj_io_out[20] padframe/mprj_io_oeb[20]
+ padframe/mprj_io_slow_sel[20] padframe/mprj_io_vtrip_sel[20] gpio_control_in_2\[6\]/resetn
+ gpio_control_in_2\[5\]/resetn gpio_control_in_2\[6\]/serial_clock gpio_control_in_2\[5\]/serial_clock
+ gpio_control_in_2\[6\]/serial_data_in gpio_control_in_2\[5\]/serial_data_in gpio_control_in_2\[6\]/serial_load
+ gpio_control_in_2\[5\]/serial_load mprj/io_in[20] mprj/io_oeb[20] mprj/io_out[20]
+ gpio_defaults_block_31/VPWR vccd1_core gpio_defaults_block_31/VGND vssd1_core gpio_control_in_2\[6\]/zero
+ gpio_control_block
Xgpio_control_in_1\[1\] gpio_defaults_block_9/gpio_defaults[0] gpio_defaults_block_9/gpio_defaults[10]
+ gpio_defaults_block_9/gpio_defaults[11] gpio_defaults_block_9/gpio_defaults[12]
+ gpio_defaults_block_9/gpio_defaults[1] gpio_defaults_block_9/gpio_defaults[2] gpio_defaults_block_9/gpio_defaults[3]
+ gpio_defaults_block_9/gpio_defaults[4] gpio_defaults_block_9/gpio_defaults[5] gpio_defaults_block_9/gpio_defaults[6]
+ gpio_defaults_block_9/gpio_defaults[7] gpio_defaults_block_9/gpio_defaults[8] gpio_defaults_block_9/gpio_defaults[9]
+ sigbuf/mgmt_io_in_unbuf[2] padframe/mprj_io_one[9] sigbuf/mgmt_io_out_buf[2] padframe/mprj_io_one[9]
+ padframe/mprj_io_analog_en[9] padframe/mprj_io_analog_pol[9] padframe/mprj_io_analog_sel[9]
+ padframe/mprj_io_dm[27] padframe/mprj_io_dm[28] padframe/mprj_io_dm[29] padframe/mprj_io_holdover[9]
+ padframe/mprj_io_ib_mode_sel[9] padframe/mprj_io_in[9] padframe/mprj_io_inp_dis[9]
+ padframe/mprj_io_out[9] padframe/mprj_io_oeb[9] padframe/mprj_io_slow_sel[9] padframe/mprj_io_vtrip_sel[9]
+ gpio_control_in_1\[1\]/resetn gpio_control_in_1\[2\]/resetn gpio_control_in_1\[1\]/serial_clock
+ gpio_control_in_1\[2\]/serial_clock gpio_control_in_1\[1\]/serial_data_in gpio_control_in_1\[2\]/serial_data_in
+ gpio_control_in_1\[1\]/serial_load gpio_control_in_1\[2\]/serial_load mprj/io_in[9]
+ mprj/io_oeb[9] mprj/io_out[9] gpio_defaults_block_9/VPWR vccd1_core gpio_defaults_block_9/VGND
+ vssd1_core gpio_control_in_1\[1\]/zero gpio_control_block
Xmprj mprj/gpio_analog[0] mprj/gpio_analog[10] mprj/gpio_analog[11] mprj/gpio_analog[12]
+ mprj/gpio_analog[13] mprj/gpio_analog[14] mprj/gpio_analog[15] mprj/gpio_analog[16]
+ mprj/gpio_analog[17] mprj/gpio_analog[1] mprj/gpio_analog[2] mprj/gpio_analog[3]
+ mprj/gpio_analog[4] mprj/gpio_analog[5] mprj/gpio_analog[6] mprj/gpio_analog[7]
+ mprj/gpio_analog[8] mprj/gpio_analog[9] mprj/gpio_noesd[0] mprj/gpio_noesd[10] mprj/gpio_noesd[11]
+ mprj/gpio_noesd[12] mprj/gpio_noesd[13] mprj/gpio_noesd[14] mprj/gpio_noesd[15]
+ mprj/gpio_noesd[16] mprj/gpio_noesd[17] mprj/gpio_noesd[1] mprj/gpio_noesd[2] mprj/gpio_noesd[3]
+ mprj/gpio_noesd[4] mprj/gpio_noesd[5] mprj/gpio_noesd[6] mprj/gpio_noesd[7] mprj/gpio_noesd[8]
+ mprj/gpio_noesd[9] mprj/io_analog[0] mprj/io_analog[10] mprj/io_analog[1] mprj/io_analog[2]
+ mprj/io_analog[3] mprj/io_analog[7] mprj/io_analog[8] mprj/io_analog[9] mprj/io_analog[4]
+ mprj/io_analog[5] mprj/io_analog[6] mprj/io_clamp_high[0] mprj/io_clamp_high[1]
+ mprj/io_clamp_high[2] mprj/io_clamp_low[0] mprj/io_clamp_low[1] mprj/io_clamp_low[2]
+ mprj/io_in[0] mprj/io_in[10] mprj/io_in[11] mprj/io_in[12] mprj/io_in[13] mprj/io_in[14]
+ mprj/io_in[15] mprj/io_in[16] mprj/io_in[17] mprj/io_in[18] mprj/io_in[19] mprj/io_in[1]
+ mprj/io_in[20] mprj/io_in[21] mprj/io_in[22] mprj/io_in[23] mprj/io_in[24] mprj/io_in[25]
+ mprj/io_in[26] mprj/io_in[2] mprj/io_in[3] mprj/io_in[4] mprj/io_in[5] mprj/io_in[6]
+ mprj/io_in[7] mprj/io_in[8] mprj/io_in[9] mprj/io_in_3v3[0] mprj/io_in_3v3[10] mprj/io_in_3v3[11]
+ mprj/io_in_3v3[12] mprj/io_in_3v3[13] mprj/io_in_3v3[14] mprj/io_in_3v3[15] mprj/io_in_3v3[16]
+ mprj/io_in_3v3[17] mprj/io_in_3v3[18] mprj/io_in_3v3[19] mprj/io_in_3v3[1] mprj/io_in_3v3[20]
+ mprj/io_in_3v3[21] mprj/io_in_3v3[22] mprj/io_in_3v3[23] mprj/io_in_3v3[24] mprj/io_in_3v3[25]
+ mprj/io_in_3v3[26] mprj/io_in_3v3[2] mprj/io_in_3v3[3] mprj/io_in_3v3[4] mprj/io_in_3v3[5]
+ mprj/io_in_3v3[6] mprj/io_in_3v3[7] mprj/io_in_3v3[8] mprj/io_in_3v3[9] mprj/io_oeb[0]
+ mprj/io_oeb[10] mprj/io_oeb[11] mprj/io_oeb[12] mprj/io_oeb[13] mprj/io_oeb[14]
+ mprj/io_oeb[15] mprj/io_oeb[16] mprj/io_oeb[17] mprj/io_oeb[18] mprj/io_oeb[19]
+ mprj/io_oeb[1] mprj/io_oeb[20] mprj/io_oeb[21] mprj/io_oeb[22] mprj/io_oeb[23] mprj/io_oeb[24]
+ mprj/io_oeb[25] mprj/io_oeb[26] mprj/io_oeb[2] mprj/io_oeb[3] mprj/io_oeb[4] mprj/io_oeb[5]
+ mprj/io_oeb[6] mprj/io_oeb[7] mprj/io_oeb[8] mprj/io_oeb[9] mprj/io_out[0] mprj/io_out[10]
+ mprj/io_out[11] mprj/io_out[12] mprj/io_out[13] mprj/io_out[14] mprj/io_out[15]
+ mprj/io_out[16] mprj/io_out[17] mprj/io_out[18] mprj/io_out[19] mprj/io_out[1] mprj/io_out[20]
+ mprj/io_out[21] mprj/io_out[22] mprj/io_out[23] mprj/io_out[24] mprj/io_out[25]
+ mprj/io_out[26] mprj/io_out[2] mprj/io_out[3] mprj/io_out[4] mprj/io_out[5] mprj/io_out[6]
+ mprj/io_out[7] mprj/io_out[8] mprj/io_out[9] mprj/la_data_in[0] mprj/la_data_in[100]
+ mprj/la_data_in[101] mprj/la_data_in[102] mprj/la_data_in[103] mprj/la_data_in[104]
+ mprj/la_data_in[105] mprj/la_data_in[106] mprj/la_data_in[107] mprj/la_data_in[108]
+ mprj/la_data_in[109] mprj/la_data_in[10] mprj/la_data_in[110] mprj/la_data_in[111]
+ mprj/la_data_in[112] mprj/la_data_in[113] mprj/la_data_in[114] mprj/la_data_in[115]
+ mprj/la_data_in[116] mprj/la_data_in[117] mprj/la_data_in[118] mprj/la_data_in[119]
+ mprj/la_data_in[11] mprj/la_data_in[120] mprj/la_data_in[121] mprj/la_data_in[122]
+ mprj/la_data_in[123] mprj/la_data_in[124] mprj/la_data_in[125] mprj/la_data_in[126]
+ mprj/la_data_in[127] mprj/la_data_in[12] mprj/la_data_in[13] mprj/la_data_in[14]
+ mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17] mprj/la_data_in[18]
+ mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21] mprj/la_data_in[22]
+ mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25] mprj/la_data_in[26]
+ mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29] mprj/la_data_in[2] mprj/la_data_in[30]
+ mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33] mprj/la_data_in[34]
+ mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37] mprj/la_data_in[38]
+ mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41] mprj/la_data_in[42]
+ mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45] mprj/la_data_in[46]
+ mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49] mprj/la_data_in[4] mprj/la_data_in[50]
+ mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53] mprj/la_data_in[54]
+ mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57] mprj/la_data_in[58]
+ mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61] mprj/la_data_in[62]
+ mprj/la_data_in[63] mprj/la_data_in[64] mprj/la_data_in[65] mprj/la_data_in[66]
+ mprj/la_data_in[67] mprj/la_data_in[68] mprj/la_data_in[69] mprj/la_data_in[6] mprj/la_data_in[70]
+ mprj/la_data_in[71] mprj/la_data_in[72] mprj/la_data_in[73] mprj/la_data_in[74]
+ mprj/la_data_in[75] mprj/la_data_in[76] mprj/la_data_in[77] mprj/la_data_in[78]
+ mprj/la_data_in[79] mprj/la_data_in[7] mprj/la_data_in[80] mprj/la_data_in[81] mprj/la_data_in[82]
+ mprj/la_data_in[83] mprj/la_data_in[84] mprj/la_data_in[85] mprj/la_data_in[86]
+ mprj/la_data_in[87] mprj/la_data_in[88] mprj/la_data_in[89] mprj/la_data_in[8] mprj/la_data_in[90]
+ mprj/la_data_in[91] mprj/la_data_in[92] mprj/la_data_in[93] mprj/la_data_in[94]
+ mprj/la_data_in[95] mprj/la_data_in[96] mprj/la_data_in[97] mprj/la_data_in[98]
+ mprj/la_data_in[99] mprj/la_data_in[9] mprj/la_data_out[0] mprj/la_data_out[100]
+ mprj/la_data_out[101] mprj/la_data_out[102] mprj/la_data_out[103] mprj/la_data_out[104]
+ mprj/la_data_out[105] mprj/la_data_out[106] mprj/la_data_out[107] mprj/la_data_out[108]
+ mprj/la_data_out[109] mprj/la_data_out[10] mprj/la_data_out[110] mprj/la_data_out[111]
+ mprj/la_data_out[112] mprj/la_data_out[113] mprj/la_data_out[114] mprj/la_data_out[115]
+ mprj/la_data_out[116] mprj/la_data_out[117] mprj/la_data_out[118] mprj/la_data_out[119]
+ mprj/la_data_out[11] mprj/la_data_out[120] mprj/la_data_out[121] mprj/la_data_out[122]
+ mprj/la_data_out[123] mprj/la_data_out[124] mprj/la_data_out[125] mprj/la_data_out[126]
+ mprj/la_data_out[127] mprj/la_data_out[12] mprj/la_data_out[13] mprj/la_data_out[14]
+ mprj/la_data_out[15] mprj/la_data_out[16] mprj/la_data_out[17] mprj/la_data_out[18]
+ mprj/la_data_out[19] mprj/la_data_out[1] mprj/la_data_out[20] mprj/la_data_out[21]
+ mprj/la_data_out[22] mprj/la_data_out[23] mprj/la_data_out[24] mprj/la_data_out[25]
+ mprj/la_data_out[26] mprj/la_data_out[27] mprj/la_data_out[28] mprj/la_data_out[29]
+ mprj/la_data_out[2] mprj/la_data_out[30] mprj/la_data_out[31] mprj/la_data_out[32]
+ mprj/la_data_out[33] mprj/la_data_out[34] mprj/la_data_out[35] mprj/la_data_out[36]
+ mprj/la_data_out[37] mprj/la_data_out[38] mprj/la_data_out[39] mprj/la_data_out[3]
+ mprj/la_data_out[40] mprj/la_data_out[41] mprj/la_data_out[42] mprj/la_data_out[43]
+ mprj/la_data_out[44] mprj/la_data_out[45] mprj/la_data_out[46] mprj/la_data_out[47]
+ mprj/la_data_out[48] mprj/la_data_out[49] mprj/la_data_out[4] mprj/la_data_out[50]
+ mprj/la_data_out[51] mprj/la_data_out[52] mprj/la_data_out[53] mprj/la_data_out[54]
+ mprj/la_data_out[55] mprj/la_data_out[56] mprj/la_data_out[57] mprj/la_data_out[58]
+ mprj/la_data_out[59] mprj/la_data_out[5] mprj/la_data_out[60] mprj/la_data_out[61]
+ mprj/la_data_out[62] mprj/la_data_out[63] mprj/la_data_out[64] mprj/la_data_out[65]
+ mprj/la_data_out[66] mprj/la_data_out[67] mprj/la_data_out[68] mprj/la_data_out[69]
+ mprj/la_data_out[6] mprj/la_data_out[70] mprj/la_data_out[71] mprj/la_data_out[72]
+ mprj/la_data_out[73] mprj/la_data_out[74] mprj/la_data_out[75] mprj/la_data_out[76]
+ mprj/la_data_out[77] mprj/la_data_out[78] mprj/la_data_out[79] mprj/la_data_out[7]
+ mprj/la_data_out[80] mprj/la_data_out[81] mprj/la_data_out[82] mprj/la_data_out[83]
+ mprj/la_data_out[84] mprj/la_data_out[85] mprj/la_data_out[86] mprj/la_data_out[87]
+ mprj/la_data_out[88] mprj/la_data_out[89] mprj/la_data_out[8] mprj/la_data_out[90]
+ mprj/la_data_out[91] mprj/la_data_out[92] mprj/la_data_out[93] mprj/la_data_out[94]
+ mprj/la_data_out[95] mprj/la_data_out[96] mprj/la_data_out[97] mprj/la_data_out[98]
+ mprj/la_data_out[99] mprj/la_data_out[9] mprj/la_oenb[0] mprj/la_oenb[100] mprj/la_oenb[101]
+ mprj/la_oenb[102] mprj/la_oenb[103] mprj/la_oenb[104] mprj/la_oenb[105] mprj/la_oenb[106]
+ mprj/la_oenb[107] mprj/la_oenb[108] mprj/la_oenb[109] mprj/la_oenb[10] mprj/la_oenb[110]
+ mprj/la_oenb[111] mprj/la_oenb[112] mprj/la_oenb[113] mprj/la_oenb[114] mprj/la_oenb[115]
+ mprj/la_oenb[116] mprj/la_oenb[117] mprj/la_oenb[118] mprj/la_oenb[119] mprj/la_oenb[11]
+ mprj/la_oenb[120] mprj/la_oenb[121] mprj/la_oenb[122] mprj/la_oenb[123] mprj/la_oenb[124]
+ mprj/la_oenb[125] mprj/la_oenb[126] mprj/la_oenb[127] mprj/la_oenb[12] mprj/la_oenb[13]
+ mprj/la_oenb[14] mprj/la_oenb[15] mprj/la_oenb[16] mprj/la_oenb[17] mprj/la_oenb[18]
+ mprj/la_oenb[19] mprj/la_oenb[1] mprj/la_oenb[20] mprj/la_oenb[21] mprj/la_oenb[22]
+ mprj/la_oenb[23] mprj/la_oenb[24] mprj/la_oenb[25] mprj/la_oenb[26] mprj/la_oenb[27]
+ mprj/la_oenb[28] mprj/la_oenb[29] mprj/la_oenb[2] mprj/la_oenb[30] mprj/la_oenb[31]
+ mprj/la_oenb[32] mprj/la_oenb[33] mprj/la_oenb[34] mprj/la_oenb[35] mprj/la_oenb[36]
+ mprj/la_oenb[37] mprj/la_oenb[38] mprj/la_oenb[39] mprj/la_oenb[3] mprj/la_oenb[40]
+ mprj/la_oenb[41] mprj/la_oenb[42] mprj/la_oenb[43] mprj/la_oenb[44] mprj/la_oenb[45]
+ mprj/la_oenb[46] mprj/la_oenb[47] mprj/la_oenb[48] mprj/la_oenb[49] mprj/la_oenb[4]
+ mprj/la_oenb[50] mprj/la_oenb[51] mprj/la_oenb[52] mprj/la_oenb[53] mprj/la_oenb[54]
+ mprj/la_oenb[55] mprj/la_oenb[56] mprj/la_oenb[57] mprj/la_oenb[58] mprj/la_oenb[59]
+ mprj/la_oenb[5] mprj/la_oenb[60] mprj/la_oenb[61] mprj/la_oenb[62] mprj/la_oenb[63]
+ mprj/la_oenb[64] mprj/la_oenb[65] mprj/la_oenb[66] mprj/la_oenb[67] mprj/la_oenb[68]
+ mprj/la_oenb[69] mprj/la_oenb[6] mprj/la_oenb[70] mprj/la_oenb[71] mprj/la_oenb[72]
+ mprj/la_oenb[73] mprj/la_oenb[74] mprj/la_oenb[75] mprj/la_oenb[76] mprj/la_oenb[77]
+ mprj/la_oenb[78] mprj/la_oenb[79] mprj/la_oenb[7] mprj/la_oenb[80] mprj/la_oenb[81]
+ mprj/la_oenb[82] mprj/la_oenb[83] mprj/la_oenb[84] mprj/la_oenb[85] mprj/la_oenb[86]
+ mprj/la_oenb[87] mprj/la_oenb[88] mprj/la_oenb[89] mprj/la_oenb[8] mprj/la_oenb[90]
+ mprj/la_oenb[91] mprj/la_oenb[92] mprj/la_oenb[93] mprj/la_oenb[94] mprj/la_oenb[95]
+ mprj/la_oenb[96] mprj/la_oenb[97] mprj/la_oenb[98] mprj/la_oenb[99] mprj/la_oenb[9]
+ mprj/user_clock2 mprj/user_irq[0] mprj/user_irq[1] mprj/user_irq[2] vccd1_core vccd2_core
+ vdda1_core vdda2_core vssa1_core vssa2_core vssd1_core vssd2_core mprj/wb_clk_i
+ mprj/wb_rst_i mprj/wbs_ack_o mprj/wbs_adr_i[0] mprj/wbs_adr_i[10] mprj/wbs_adr_i[11]
+ mprj/wbs_adr_i[12] mprj/wbs_adr_i[13] mprj/wbs_adr_i[14] mprj/wbs_adr_i[15] mprj/wbs_adr_i[16]
+ mprj/wbs_adr_i[17] mprj/wbs_adr_i[18] mprj/wbs_adr_i[19] mprj/wbs_adr_i[1] mprj/wbs_adr_i[20]
+ mprj/wbs_adr_i[21] mprj/wbs_adr_i[22] mprj/wbs_adr_i[23] mprj/wbs_adr_i[24] mprj/wbs_adr_i[25]
+ mprj/wbs_adr_i[26] mprj/wbs_adr_i[27] mprj/wbs_adr_i[28] mprj/wbs_adr_i[29] mprj/wbs_adr_i[2]
+ mprj/wbs_adr_i[30] mprj/wbs_adr_i[31] mprj/wbs_adr_i[3] mprj/wbs_adr_i[4] mprj/wbs_adr_i[5]
+ mprj/wbs_adr_i[6] mprj/wbs_adr_i[7] mprj/wbs_adr_i[8] mprj/wbs_adr_i[9] mprj/wbs_cyc_i
+ mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12] mprj/wbs_dat_i[13]
+ mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17] mprj/wbs_dat_i[18]
+ mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21] mprj/wbs_dat_i[22]
+ mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26] mprj/wbs_dat_i[27]
+ mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30] mprj/wbs_dat_i[31]
+ mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6] mprj/wbs_dat_i[7]
+ mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] mprj/wbs_dat_o[0] mprj/wbs_dat_o[10] mprj/wbs_dat_o[11]
+ mprj/wbs_dat_o[12] mprj/wbs_dat_o[13] mprj/wbs_dat_o[14] mprj/wbs_dat_o[15] mprj/wbs_dat_o[16]
+ mprj/wbs_dat_o[17] mprj/wbs_dat_o[18] mprj/wbs_dat_o[19] mprj/wbs_dat_o[1] mprj/wbs_dat_o[20]
+ mprj/wbs_dat_o[21] mprj/wbs_dat_o[22] mprj/wbs_dat_o[23] mprj/wbs_dat_o[24] mprj/wbs_dat_o[25]
+ mprj/wbs_dat_o[26] mprj/wbs_dat_o[27] mprj/wbs_dat_o[28] mprj/wbs_dat_o[29] mprj/wbs_dat_o[2]
+ mprj/wbs_dat_o[30] mprj/wbs_dat_o[31] mprj/wbs_dat_o[3] mprj/wbs_dat_o[4] mprj/wbs_dat_o[5]
+ mprj/wbs_dat_o[6] mprj/wbs_dat_o[7] mprj/wbs_dat_o[8] mprj/wbs_dat_o[9] mprj/wbs_sel_i[0]
+ mprj/wbs_sel_i[1] mprj/wbs_sel_i[2] mprj/wbs_sel_i[3] mprj/wbs_stb_i mprj/wbs_we_i
+ user_analog_project_wrapper
Xgpio_control_in_2\[4\] gpio_defaults_block_29/gpio_defaults[0] gpio_defaults_block_29/gpio_defaults[10]
+ gpio_defaults_block_29/gpio_defaults[11] gpio_defaults_block_29/gpio_defaults[12]
+ gpio_defaults_block_29/gpio_defaults[1] gpio_defaults_block_29/gpio_defaults[2]
+ gpio_defaults_block_29/gpio_defaults[3] gpio_defaults_block_29/gpio_defaults[4]
+ gpio_defaults_block_29/gpio_defaults[5] gpio_defaults_block_29/gpio_defaults[6]
+ gpio_defaults_block_29/gpio_defaults[7] gpio_defaults_block_29/gpio_defaults[8]
+ gpio_defaults_block_29/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[11] padframe/mprj_io_one[18]
+ sigbuf/mgmt_io_out_buf[11] padframe/mprj_io_one[18] padframe/mprj_io_analog_en[18]
+ padframe/mprj_io_analog_pol[18] padframe/mprj_io_analog_sel[18] padframe/mprj_io_dm[54]
+ padframe/mprj_io_dm[55] padframe/mprj_io_dm[56] padframe/mprj_io_holdover[18] padframe/mprj_io_ib_mode_sel[18]
+ padframe/mprj_io_in[18] padframe/mprj_io_inp_dis[18] padframe/mprj_io_out[18] padframe/mprj_io_oeb[18]
+ padframe/mprj_io_slow_sel[18] padframe/mprj_io_vtrip_sel[18] gpio_control_in_2\[4\]/resetn
+ gpio_control_in_2\[3\]/resetn gpio_control_in_2\[4\]/serial_clock gpio_control_in_2\[3\]/serial_clock
+ gpio_control_in_2\[4\]/serial_data_in gpio_control_in_2\[3\]/serial_data_in gpio_control_in_2\[4\]/serial_load
+ gpio_control_in_2\[3\]/serial_load mprj/io_in[18] mprj/io_oeb[18] mprj/io_out[18]
+ gpio_defaults_block_29/VPWR vccd1_core gpio_defaults_block_29/VGND vssd1_core gpio_control_in_2\[4\]/zero
+ gpio_control_block
Xgpio_control_bidir_1\[1\] gpio_defaults_block_1/gpio_defaults[0] gpio_defaults_block_1/gpio_defaults[10]
+ gpio_defaults_block_1/gpio_defaults[11] gpio_defaults_block_1/gpio_defaults[12]
+ gpio_defaults_block_1/gpio_defaults[1] gpio_defaults_block_1/gpio_defaults[2] gpio_defaults_block_1/gpio_defaults[3]
+ gpio_defaults_block_1/gpio_defaults[4] gpio_defaults_block_1/gpio_defaults[5] gpio_defaults_block_1/gpio_defaults[6]
+ gpio_defaults_block_1/gpio_defaults[7] gpio_defaults_block_1/gpio_defaults[8] gpio_defaults_block_1/gpio_defaults[9]
+ housekeeping/mgmt_gpio_in[1] housekeeping/mgmt_gpio_oeb[1] housekeeping/mgmt_gpio_out[1]
+ padframe/mprj_io_one[1] padframe/mprj_io_analog_en[1] padframe/mprj_io_analog_pol[1]
+ padframe/mprj_io_analog_sel[1] padframe/mprj_io_dm[3] padframe/mprj_io_dm[4] padframe/mprj_io_dm[5]
+ padframe/mprj_io_holdover[1] padframe/mprj_io_ib_mode_sel[1] padframe/mprj_io_in[1]
+ padframe/mprj_io_inp_dis[1] padframe/mprj_io_out[1] padframe/mprj_io_oeb[1] padframe/mprj_io_slow_sel[1]
+ padframe/mprj_io_vtrip_sel[1] gpio_control_bidir_1\[1\]/resetn gpio_control_in_1a\[0\]/resetn
+ gpio_control_bidir_1\[1\]/serial_clock gpio_control_in_1a\[0\]/serial_clock gpio_control_bidir_1\[1\]/serial_data_in
+ gpio_control_in_1a\[0\]/serial_data_in gpio_control_bidir_1\[1\]/serial_load gpio_control_in_1a\[0\]/serial_load
+ mprj/io_in[1] mprj/io_oeb[1] mprj/io_out[1] gpio_defaults_block_1/VPWR vccd1_core
+ gpio_defaults_block_1/VGND vssd1_core housekeeping/mgmt_gpio_in[17] gpio_control_block
Xspare_logic\[2\] spare_logic\[2\]/spare_xfq[0] spare_logic\[2\]/spare_xfq[1] spare_logic\[2\]/spare_xfqn[0]
+ spare_logic\[2\]/spare_xfqn[1] spare_logic\[2\]/spare_xi[0] spare_logic\[2\]/spare_xi[1]
+ spare_logic\[2\]/spare_xi[2] spare_logic\[2\]/spare_xi[3] spare_logic\[2\]/spare_xib
+ spare_logic\[2\]/spare_xmx[0] spare_logic\[2\]/spare_xmx[1] spare_logic\[2\]/spare_xna[0]
+ spare_logic\[2\]/spare_xna[1] spare_logic\[2\]/spare_xno[0] spare_logic\[2\]/spare_xno[1]
+ spare_logic\[2\]/spare_xz[0] spare_logic\[2\]/spare_xz[10] spare_logic\[2\]/spare_xz[11]
+ spare_logic\[2\]/spare_xz[12] spare_logic\[2\]/spare_xz[13] spare_logic\[2\]/spare_xz[14]
+ spare_logic\[2\]/spare_xz[15] spare_logic\[2\]/spare_xz[16] spare_logic\[2\]/spare_xz[17]
+ spare_logic\[2\]/spare_xz[18] spare_logic\[2\]/spare_xz[19] spare_logic\[2\]/spare_xz[1]
+ spare_logic\[2\]/spare_xz[20] spare_logic\[2\]/spare_xz[21] spare_logic\[2\]/spare_xz[22]
+ spare_logic\[2\]/spare_xz[23] spare_logic\[2\]/spare_xz[24] spare_logic\[2\]/spare_xz[25]
+ spare_logic\[2\]/spare_xz[26] spare_logic\[2\]/spare_xz[2] spare_logic\[2\]/spare_xz[3]
+ spare_logic\[2\]/spare_xz[4] spare_logic\[2\]/spare_xz[5] spare_logic\[2\]/spare_xz[6]
+ spare_logic\[2\]/spare_xz[7] spare_logic\[2\]/spare_xz[8] spare_logic\[2\]/spare_xz[9]
+ soc/VPWR soc/VGND spare_logic_block
Xhousekeeping soc/VGND soc/VPWR soc/debug_in soc/debug_mode soc/debug_oeb soc/debug_out
+ soc/irq[3] soc/irq[4] soc/irq[5] user_id_value/mask_rev[0] user_id_value/mask_rev[10]
+ user_id_value/mask_rev[11] user_id_value/mask_rev[12] user_id_value/mask_rev[13]
+ user_id_value/mask_rev[14] user_id_value/mask_rev[15] user_id_value/mask_rev[16]
+ user_id_value/mask_rev[17] user_id_value/mask_rev[18] user_id_value/mask_rev[19]
+ user_id_value/mask_rev[1] user_id_value/mask_rev[20] user_id_value/mask_rev[21]
+ user_id_value/mask_rev[22] user_id_value/mask_rev[23] user_id_value/mask_rev[24]
+ user_id_value/mask_rev[25] user_id_value/mask_rev[26] user_id_value/mask_rev[27]
+ user_id_value/mask_rev[28] user_id_value/mask_rev[29] user_id_value/mask_rev[2]
+ user_id_value/mask_rev[30] user_id_value/mask_rev[31] user_id_value/mask_rev[3]
+ user_id_value/mask_rev[4] user_id_value/mask_rev[5] user_id_value/mask_rev[6] user_id_value/mask_rev[7]
+ user_id_value/mask_rev[8] user_id_value/mask_rev[9] housekeeping/mgmt_gpio_in[0]
+ sigbuf/mgmt_io_in_buf[3] sigbuf/mgmt_io_in_buf[4] sigbuf/mgmt_io_in_buf[5] sigbuf/mgmt_io_in_buf[6]
+ housekeeping/mgmt_gpio_in[15] housekeeping/mgmt_gpio_in[15] housekeeping/mgmt_gpio_in[17]
+ housekeeping/mgmt_gpio_in[17] gpio_control_in_1a\[0\]/zero gpio_control_in_1a\[0\]/zero
+ housekeeping/mgmt_gpio_in[1] gpio_control_in_1a\[1\]/zero gpio_control_in_1a\[1\]/zero
+ gpio_control_in_1a\[2\]/zero gpio_control_in_1a\[2\]/zero gpio_control_in_1a\[3\]/zero
+ sigbuf/mgmt_io_in_buf[7] sigbuf/mgmt_io_in_buf[8] sigbuf/mgmt_io_in_buf[9] sigbuf/mgmt_io_in_buf[10]
+ sigbuf/mgmt_io_in_buf[11] housekeeping/mgmt_gpio_in[2] sigbuf/mgmt_io_in_buf[12]
+ sigbuf/mgmt_io_in_buf[13] sigbuf/mgmt_io_in_buf[14] sigbuf/mgmt_io_in_buf[15] sigbuf/mgmt_io_in_buf[16]
+ sigbuf/mgmt_io_in_buf[17] sigbuf/mgmt_io_in_buf[18] sigbuf/mgmt_io_in_buf[19] housekeeping/mgmt_gpio_in[3]
+ housekeeping/mgmt_gpio_in[4] housekeeping/mgmt_gpio_in[5] housekeeping/mgmt_gpio_in[6]
+ sigbuf/mgmt_io_in_buf[0] sigbuf/mgmt_io_in_buf[1] sigbuf/mgmt_io_in_buf[2] housekeeping/mgmt_gpio_oeb[0]
+ housekeeping/mgmt_gpio_oeb[10] housekeeping/mgmt_gpio_oeb[11] housekeeping/mgmt_gpio_oeb[12]
+ housekeeping/mgmt_gpio_oeb[13] housekeeping/mgmt_gpio_oeb[14] housekeeping/mgmt_gpio_oeb[15]
+ housekeeping/mgmt_gpio_oeb[16] housekeeping/mgmt_gpio_oeb[17] housekeeping/mgmt_gpio_oeb[18]
+ housekeeping/mgmt_gpio_oeb[19] housekeeping/mgmt_gpio_oeb[1] housekeeping/mgmt_gpio_oeb[20]
+ housekeeping/mgmt_gpio_oeb[21] housekeeping/mgmt_gpio_oeb[22] housekeeping/mgmt_gpio_oeb[23]
+ housekeeping/mgmt_gpio_oeb[24] housekeeping/mgmt_gpio_oeb[25] housekeeping/mgmt_gpio_oeb[26]
+ housekeeping/mgmt_gpio_oeb[27] housekeeping/mgmt_gpio_oeb[28] housekeeping/mgmt_gpio_oeb[29]
+ housekeeping/mgmt_gpio_oeb[2] housekeeping/mgmt_gpio_oeb[30] housekeeping/mgmt_gpio_oeb[31]
+ housekeeping/mgmt_gpio_oeb[32] housekeeping/mgmt_gpio_oeb[33] housekeeping/mgmt_gpio_oeb[34]
+ sigbuf/mgmt_io_oeb_unbuf[0] sigbuf/mgmt_io_oeb_unbuf[1] sigbuf/mgmt_io_oeb_unbuf[2]
+ housekeeping/mgmt_gpio_oeb[3] housekeeping/mgmt_gpio_oeb[4] housekeeping/mgmt_gpio_oeb[5]
+ housekeeping/mgmt_gpio_oeb[6] housekeeping/mgmt_gpio_oeb[7] housekeeping/mgmt_gpio_oeb[8]
+ housekeeping/mgmt_gpio_oeb[9] housekeeping/mgmt_gpio_out[0] sigbuf/mgmt_io_out_unbuf[3]
+ sigbuf/mgmt_io_out_unbuf[4] sigbuf/mgmt_io_out_unbuf[5] sigbuf/mgmt_io_out_unbuf[6]
+ housekeeping/mgmt_gpio_out[14] housekeeping/mgmt_gpio_out[15] housekeeping/mgmt_gpio_out[16]
+ housekeeping/mgmt_gpio_out[17] housekeeping/mgmt_gpio_out[18] housekeeping/mgmt_gpio_out[19]
+ housekeeping/mgmt_gpio_out[1] housekeeping/mgmt_gpio_out[20] housekeeping/mgmt_gpio_out[21]
+ housekeeping/mgmt_gpio_out[22] housekeeping/mgmt_gpio_out[23] housekeeping/mgmt_gpio_out[24]
+ sigbuf/mgmt_io_out_unbuf[7] sigbuf/mgmt_io_out_unbuf[8] sigbuf/mgmt_io_out_unbuf[9]
+ sigbuf/mgmt_io_out_unbuf[10] sigbuf/mgmt_io_out_unbuf[11] housekeeping/mgmt_gpio_out[2]
+ sigbuf/mgmt_io_out_unbuf[12] sigbuf/mgmt_io_out_unbuf[13] sigbuf/mgmt_io_out_unbuf[14]
+ sigbuf/mgmt_io_out_unbuf[15] sigbuf/mgmt_io_out_unbuf[16] sigbuf/mgmt_io_out_unbuf[17]
+ sigbuf/mgmt_io_out_unbuf[18] sigbuf/mgmt_io_out_unbuf[19] housekeeping/mgmt_gpio_out[3]
+ housekeeping/mgmt_gpio_out[4] housekeeping/mgmt_gpio_out[5] housekeeping/mgmt_gpio_out[6]
+ sigbuf/mgmt_io_out_unbuf[0] sigbuf/mgmt_io_out_unbuf[1] sigbuf/mgmt_io_out_unbuf[2]
+ housekeeping/pad_flash_clk flash_clkrst_buffers/in_n[7] housekeeping/pad_flash_csb
+ flash_clkrst_buffers/in_n[6] housekeeping/pad_flash_io0_di flash_clkrst_buffers/in_n[1]
+ flash_clkrst_buffers/in_n[3] flash_clkrst_buffers/in_n[5] housekeeping/pad_flash_io1_di
+ flash_clkrst_buffers/in_n[0] flash_clkrst_buffers/in_n[2] flash_clkrst_buffers/in_n[4]
+ clock_ctrl/sel2[0] clock_ctrl/sel2[1] clock_ctrl/sel2[2] clock_ctrl/ext_clk_sel
+ pll/dco pll/div[0] pll/div[1] pll/div[2] pll/div[3] pll/div[4] pll/enable clock_ctrl/sel[0]
+ clock_ctrl/sel[1] clock_ctrl/sel[2] pll/ext_trim[0] pll/ext_trim[10] pll/ext_trim[11]
+ pll/ext_trim[12] pll/ext_trim[13] pll/ext_trim[14] pll/ext_trim[15] pll/ext_trim[16]
+ pll/ext_trim[17] pll/ext_trim[18] pll/ext_trim[19] pll/ext_trim[1] pll/ext_trim[20]
+ pll/ext_trim[21] pll/ext_trim[22] pll/ext_trim[23] pll/ext_trim[24] pll/ext_trim[25]
+ pll/ext_trim[2] pll/ext_trim[3] pll/ext_trim[4] pll/ext_trim[5] pll/ext_trim[6]
+ pll/ext_trim[7] pll/ext_trim[8] pll/ext_trim[9] por/porb_l housekeeping/pwr_ctrl_out[0]
+ housekeeping/pwr_ctrl_out[1] housekeeping/pwr_ctrl_out[2] housekeeping/pwr_ctrl_out[3]
+ soc/qspi_enabled housekeeping/reset soc/ser_rx soc/ser_tx soc/serial_clock_in housekeeping/serial_data_1
+ soc/serial_data_2_in soc/serial_load_in soc/serial_resetn_in soc/spi_csb soc/spi_enabled
+ soc/spi_sck soc/spi_sdi soc/spi_sdo soc/spi_sdoenb soc/flash_clk soc/flash_csb soc/flash_io0_di
+ soc/flash_io0_do soc/flash_io0_oeb soc/flash_io1_di soc/flash_io1_do soc/flash_io1_oeb
+ soc/flash_io2_di soc/flash_io2_do soc/flash_io2_oeb soc/flash_io3_di soc/flash_io3_do
+ soc/flash_io3_oeb soc/trap soc/uart_enabled clock_ctrl/user_clk housekeeping/usr1_vcc_pwrgood
+ housekeeping/usr1_vdd_pwrgood housekeeping/usr2_vcc_pwrgood housekeeping/usr2_vdd_pwrgood
+ soc/hk_ack_i soc/mprj_adr_o[0] soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12]
+ soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17]
+ soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21]
+ soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26]
+ soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30]
+ soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6]
+ soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9] clock_ctrl/core_clk soc/hk_cyc_o
+ soc/mprj_dat_o[0] soc/mprj_dat_o[10] soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13]
+ soc/mprj_dat_o[14] soc/mprj_dat_o[15] soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18]
+ soc/mprj_dat_o[19] soc/mprj_dat_o[1] soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22]
+ soc/mprj_dat_o[23] soc/mprj_dat_o[24] soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27]
+ soc/mprj_dat_o[28] soc/mprj_dat_o[29] soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31]
+ soc/mprj_dat_o[3] soc/mprj_dat_o[4] soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7]
+ soc/mprj_dat_o[8] soc/mprj_dat_o[9] soc/hk_dat_i[0] soc/hk_dat_i[10] soc/hk_dat_i[11]
+ soc/hk_dat_i[12] soc/hk_dat_i[13] soc/hk_dat_i[14] soc/hk_dat_i[15] soc/hk_dat_i[16]
+ soc/hk_dat_i[17] soc/hk_dat_i[18] soc/hk_dat_i[19] soc/hk_dat_i[1] soc/hk_dat_i[20]
+ soc/hk_dat_i[21] soc/hk_dat_i[22] soc/hk_dat_i[23] soc/hk_dat_i[24] soc/hk_dat_i[25]
+ soc/hk_dat_i[26] soc/hk_dat_i[27] soc/hk_dat_i[28] soc/hk_dat_i[29] soc/hk_dat_i[2]
+ soc/hk_dat_i[30] soc/hk_dat_i[31] soc/hk_dat_i[3] soc/hk_dat_i[4] soc/hk_dat_i[5]
+ soc/hk_dat_i[6] soc/hk_dat_i[7] soc/hk_dat_i[8] soc/hk_dat_i[9] housekeeping/wb_rstn_i
+ soc/mprj_sel_o[0] soc/mprj_sel_o[1] soc/mprj_sel_o[2] soc/mprj_sel_o[3] soc/hk_stb_o
+ soc/mprj_we_o housekeeping
Xgpio_control_in_2\[2\] gpio_defaults_block_27/gpio_defaults[0] gpio_defaults_block_27/gpio_defaults[10]
+ gpio_defaults_block_27/gpio_defaults[11] gpio_defaults_block_27/gpio_defaults[12]
+ gpio_defaults_block_27/gpio_defaults[1] gpio_defaults_block_27/gpio_defaults[2]
+ gpio_defaults_block_27/gpio_defaults[3] gpio_defaults_block_27/gpio_defaults[4]
+ gpio_defaults_block_27/gpio_defaults[5] gpio_defaults_block_27/gpio_defaults[6]
+ gpio_defaults_block_27/gpio_defaults[7] gpio_defaults_block_27/gpio_defaults[8]
+ gpio_defaults_block_27/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[9] padframe/mprj_io_one[16]
+ sigbuf/mgmt_io_out_buf[9] padframe/mprj_io_one[16] padframe/mprj_io_analog_en[16]
+ padframe/mprj_io_analog_pol[16] padframe/mprj_io_analog_sel[16] padframe/mprj_io_dm[48]
+ padframe/mprj_io_dm[49] padframe/mprj_io_dm[50] padframe/mprj_io_holdover[16] padframe/mprj_io_ib_mode_sel[16]
+ padframe/mprj_io_in[16] padframe/mprj_io_inp_dis[16] padframe/mprj_io_out[16] padframe/mprj_io_oeb[16]
+ padframe/mprj_io_slow_sel[16] padframe/mprj_io_vtrip_sel[16] gpio_control_in_2\[2\]/resetn
+ gpio_control_in_2\[1\]/resetn gpio_control_in_2\[2\]/serial_clock gpio_control_in_2\[1\]/serial_clock
+ gpio_control_in_2\[2\]/serial_data_in gpio_control_in_2\[1\]/serial_data_in gpio_control_in_2\[2\]/serial_load
+ gpio_control_in_2\[1\]/serial_load mprj/io_in[16] mprj/io_oeb[16] mprj/io_out[16]
+ gpio_defaults_block_27/VPWR vccd1_core gpio_defaults_block_27/VGND vssd1_core gpio_control_in_2\[2\]/zero
+ gpio_control_block
Xgpio_defaults_block_30 VSUBS sigbuf/vccd gpio_defaults_block_30/gpio_defaults[0]
+ gpio_defaults_block_30/gpio_defaults[10] gpio_defaults_block_30/gpio_defaults[11]
+ gpio_defaults_block_30/gpio_defaults[12] gpio_defaults_block_30/gpio_defaults[1]
+ gpio_defaults_block_30/gpio_defaults[2] gpio_defaults_block_30/gpio_defaults[3]
+ gpio_defaults_block_30/gpio_defaults[4] gpio_defaults_block_30/gpio_defaults[5]
+ gpio_defaults_block_30/gpio_defaults[6] gpio_defaults_block_30/gpio_defaults[7]
+ gpio_defaults_block_30/gpio_defaults[8] gpio_defaults_block_30/gpio_defaults[9]
+ gpio_defaults_block
Xspare_logic\[0\] spare_logic\[0\]/spare_xfq[0] spare_logic\[0\]/spare_xfq[1] spare_logic\[0\]/spare_xfqn[0]
+ spare_logic\[0\]/spare_xfqn[1] spare_logic\[0\]/spare_xi[0] spare_logic\[0\]/spare_xi[1]
+ spare_logic\[0\]/spare_xi[2] spare_logic\[0\]/spare_xi[3] spare_logic\[0\]/spare_xib
+ spare_logic\[0\]/spare_xmx[0] spare_logic\[0\]/spare_xmx[1] spare_logic\[0\]/spare_xna[0]
+ spare_logic\[0\]/spare_xna[1] spare_logic\[0\]/spare_xno[0] spare_logic\[0\]/spare_xno[1]
+ spare_logic\[0\]/spare_xz[0] spare_logic\[0\]/spare_xz[10] spare_logic\[0\]/spare_xz[11]
+ spare_logic\[0\]/spare_xz[12] spare_logic\[0\]/spare_xz[13] spare_logic\[0\]/spare_xz[14]
+ spare_logic\[0\]/spare_xz[15] spare_logic\[0\]/spare_xz[16] spare_logic\[0\]/spare_xz[17]
+ spare_logic\[0\]/spare_xz[18] spare_logic\[0\]/spare_xz[19] spare_logic\[0\]/spare_xz[1]
+ spare_logic\[0\]/spare_xz[20] spare_logic\[0\]/spare_xz[21] spare_logic\[0\]/spare_xz[22]
+ spare_logic\[0\]/spare_xz[23] spare_logic\[0\]/spare_xz[24] spare_logic\[0\]/spare_xz[25]
+ spare_logic\[0\]/spare_xz[26] spare_logic\[0\]/spare_xz[2] spare_logic\[0\]/spare_xz[3]
+ spare_logic\[0\]/spare_xz[4] spare_logic\[0\]/spare_xz[5] spare_logic\[0\]/spare_xz[6]
+ spare_logic\[0\]/spare_xz[7] spare_logic\[0\]/spare_xz[8] spare_logic\[0\]/spare_xz[9]
+ soc/VPWR soc/VGND spare_logic_block
Xflash_clkrst_buffers flash_clkrst_buffers/VGND flash_clkrst_buffers/VPWR flash_clkrst_buffers/in_n[0]
+ housekeeping/wb_rstn_i clock_ctrl/core_clk flash_clkrst_buffers/in_n[1] flash_clkrst_buffers/in_n[2]
+ flash_clkrst_buffers/in_n[3] flash_clkrst_buffers/in_n[4] flash_clkrst_buffers/in_n[5]
+ flash_clkrst_buffers/in_n[6] flash_clkrst_buffers/in_n[7] housekeeping/pad_flash_csb
+ housekeeping/pad_flash_clk padframe/flash_io0_di_core padframe/flash_io1_di_core
+ padframe/clock_core housekeeping/pad_flash_io0_di housekeeping/pad_flash_io1_di
+ pll/osc padframe/flash_io1_do_core soc/resetn_in soc/clk_in padframe/flash_io0_do_core
+ padframe/flash_io1_ieb_core padframe/flash_io0_ieb_core padframe/flash_io1_oeb_core
+ padframe/flash_io0_oeb_core padframe/flash_csb_oeb_core padframe/flash_clk_oeb_core
+ padframe/flash_csb_core padframe/flash_clk_core buff_flash_clkrst
Xgpio_defaults_block_10 gpio_defaults_block_10/VGND gpio_defaults_block_10/VPWR gpio_defaults_block_10/gpio_defaults[0]
+ gpio_defaults_block_10/gpio_defaults[10] gpio_defaults_block_10/gpio_defaults[11]
+ gpio_defaults_block_10/gpio_defaults[12] gpio_defaults_block_10/gpio_defaults[1]
+ gpio_defaults_block_10/gpio_defaults[2] gpio_defaults_block_10/gpio_defaults[3]
+ gpio_defaults_block_10/gpio_defaults[4] gpio_defaults_block_10/gpio_defaults[5]
+ gpio_defaults_block_10/gpio_defaults[6] gpio_defaults_block_10/gpio_defaults[7]
+ gpio_defaults_block_10/gpio_defaults[8] gpio_defaults_block_10/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_defaults_block_31 gpio_defaults_block_31/VGND gpio_defaults_block_31/VPWR gpio_defaults_block_31/gpio_defaults[0]
+ gpio_defaults_block_31/gpio_defaults[10] gpio_defaults_block_31/gpio_defaults[11]
+ gpio_defaults_block_31/gpio_defaults[12] gpio_defaults_block_31/gpio_defaults[1]
+ gpio_defaults_block_31/gpio_defaults[2] gpio_defaults_block_31/gpio_defaults[3]
+ gpio_defaults_block_31/gpio_defaults[4] gpio_defaults_block_31/gpio_defaults[5]
+ gpio_defaults_block_31/gpio_defaults[6] gpio_defaults_block_31/gpio_defaults[7]
+ gpio_defaults_block_31/gpio_defaults[8] gpio_defaults_block_31/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_control_in_1a\[5\] gpio_defaults_block_7/gpio_defaults[0] gpio_defaults_block_7/gpio_defaults[10]
+ gpio_defaults_block_7/gpio_defaults[11] gpio_defaults_block_7/gpio_defaults[12]
+ gpio_defaults_block_7/gpio_defaults[1] gpio_defaults_block_7/gpio_defaults[2] gpio_defaults_block_7/gpio_defaults[3]
+ gpio_defaults_block_7/gpio_defaults[4] gpio_defaults_block_7/gpio_defaults[5] gpio_defaults_block_7/gpio_defaults[6]
+ gpio_defaults_block_7/gpio_defaults[7] gpio_defaults_block_7/gpio_defaults[8] gpio_defaults_block_7/gpio_defaults[9]
+ sigbuf/mgmt_io_in_unbuf[0] padframe/mprj_io_one[7] sigbuf/mgmt_io_out_buf[0] padframe/mprj_io_one[7]
+ padframe/mprj_io_analog_en[7] padframe/mprj_io_analog_pol[7] padframe/mprj_io_analog_sel[7]
+ padframe/mprj_io_dm[21] padframe/mprj_io_dm[22] padframe/mprj_io_dm[23] padframe/mprj_io_holdover[7]
+ padframe/mprj_io_ib_mode_sel[7] padframe/mprj_io_in[7] padframe/mprj_io_inp_dis[7]
+ padframe/mprj_io_out[7] padframe/mprj_io_oeb[7] padframe/mprj_io_slow_sel[7] padframe/mprj_io_vtrip_sel[7]
+ gpio_control_in_1a\[5\]/resetn gpio_control_in_1\[0\]/resetn gpio_control_in_1a\[5\]/serial_clock
+ gpio_control_in_1\[0\]/serial_clock gpio_control_in_1a\[5\]/serial_data_in gpio_control_in_1\[0\]/serial_data_in
+ gpio_control_in_1a\[5\]/serial_load gpio_control_in_1\[0\]/serial_load mprj/io_in[7]
+ mprj/io_oeb[7] mprj/io_out[7] gpio_defaults_block_7/VPWR vccd1_core gpio_defaults_block_7/VGND
+ vssd1_core gpio_control_in_1a\[5\]/zero gpio_control_block
Xgpio_defaults_block_32 gpio_defaults_block_32/VGND gpio_defaults_block_32/VPWR gpio_defaults_block_32/gpio_defaults[0]
+ gpio_defaults_block_32/gpio_defaults[10] gpio_defaults_block_32/gpio_defaults[11]
+ gpio_defaults_block_32/gpio_defaults[12] gpio_defaults_block_32/gpio_defaults[1]
+ gpio_defaults_block_32/gpio_defaults[2] gpio_defaults_block_32/gpio_defaults[3]
+ gpio_defaults_block_32/gpio_defaults[4] gpio_defaults_block_32/gpio_defaults[5]
+ gpio_defaults_block_32/gpio_defaults[6] gpio_defaults_block_32/gpio_defaults[7]
+ gpio_defaults_block_32/gpio_defaults[8] gpio_defaults_block_32/gpio_defaults[9]
+ gpio_defaults_block
Xgpio_control_bidir_2\[2\] gpio_defaults_block_37/gpio_defaults[0] gpio_defaults_block_37/gpio_defaults[10]
+ gpio_defaults_block_37/gpio_defaults[11] gpio_defaults_block_37/gpio_defaults[12]
+ gpio_defaults_block_37/gpio_defaults[1] gpio_defaults_block_37/gpio_defaults[2]
+ gpio_defaults_block_37/gpio_defaults[3] gpio_defaults_block_37/gpio_defaults[4]
+ gpio_defaults_block_37/gpio_defaults[5] gpio_defaults_block_37/gpio_defaults[6]
+ gpio_defaults_block_37/gpio_defaults[7] gpio_defaults_block_37/gpio_defaults[8]
+ gpio_defaults_block_37/gpio_defaults[9] sigbuf/mgmt_io_in_unbuf[19] sigbuf/mgmt_io_oeb_buf[2]
+ sigbuf/mgmt_io_out_buf[19] padframe/mprj_io_one[26] padframe/mprj_io_analog_en[26]
+ padframe/mprj_io_analog_pol[26] padframe/mprj_io_analog_sel[26] padframe/mprj_io_dm[78]
+ padframe/mprj_io_dm[79] padframe/mprj_io_dm[80] padframe/mprj_io_holdover[26] padframe/mprj_io_ib_mode_sel[26]
+ padframe/mprj_io_in[26] padframe/mprj_io_inp_dis[26] padframe/mprj_io_out[26] padframe/mprj_io_oeb[26]
+ padframe/mprj_io_slow_sel[26] padframe/mprj_io_vtrip_sel[26] soc/serial_resetn_out
+ gpio_control_bidir_2\[1\]/resetn soc/serial_clock_out gpio_control_bidir_2\[1\]/serial_clock
+ soc/serial_data_2_out gpio_control_bidir_2\[1\]/serial_data_in soc/serial_load_out
+ gpio_control_bidir_2\[1\]/serial_load mprj/io_in[26] mprj/io_oeb[26] mprj/io_out[26]
+ gpio_defaults_block_37/VPWR vccd1_core gpio_defaults_block_37/VGND vssd1_core gpio_control_bidir_2\[2\]/zero
+ gpio_control_block
.ends

