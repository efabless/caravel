magic
tech sky130A
magscale 1 2
timestamp 1637791793
<< error_p >>
rect 585752 994898 585758 994904
rect 590380 994898 590386 994904
rect 585758 994892 585764 994898
rect 590374 994892 590380 994898
rect 575756 994884 575762 994890
rect 580384 994884 580390 994890
rect 575762 994878 575768 994884
rect 580378 994878 580384 994884
rect 675398 903522 676480 903546
rect 675398 902472 675422 903522
rect 676456 902472 676480 903522
rect 675398 902448 676480 902472
rect 671692 901904 672774 901928
rect 671692 900854 671716 901904
rect 672750 900854 672774 901904
rect 671692 900830 672774 900854
rect 686002 900231 686756 900232
rect 686002 899155 686003 900231
rect 686755 899155 686756 900231
rect 686002 899154 686756 899155
rect 679456 898663 680218 898664
rect 679456 897581 679457 898663
rect 680217 897581 680218 898663
rect 679456 897580 680218 897581
rect 30820 820831 31574 820832
rect 30820 819755 30821 820831
rect 31573 819755 31574 820831
rect 30820 819754 31574 819755
rect 37358 819263 38120 819264
rect 37358 818181 37359 819263
rect 38119 818181 38120 819263
rect 37358 818180 38120 818181
rect 30820 777631 31574 777632
rect 30820 776555 30821 777631
rect 31573 776555 31574 777631
rect 30820 776554 31574 776555
rect 37358 776063 38120 776064
rect 37358 774981 37359 776063
rect 38119 774981 38120 776063
rect 37358 774980 38120 774981
rect 30820 734431 31574 734432
rect 30820 733355 30821 734431
rect 31573 733355 31574 734431
rect 30820 733354 31574 733355
rect 37358 732863 38120 732864
rect 37358 731781 37359 732863
rect 38119 731781 38120 732863
rect 37358 731780 38120 731781
rect 675408 722922 676490 722946
rect 675408 721872 675432 722922
rect 676466 721872 676490 722922
rect 675408 721848 676490 721872
rect 671702 721304 672784 721328
rect 671702 720254 671726 721304
rect 672760 720254 672784 721304
rect 671702 720230 672784 720254
rect 686012 719631 686766 719632
rect 686012 718555 686013 719631
rect 686765 718555 686766 719631
rect 686012 718554 686766 718555
rect 679466 718063 680228 718064
rect 679466 716981 679467 718063
rect 680227 716981 680228 718063
rect 679466 716980 680228 716981
rect 30820 691231 31574 691232
rect 30820 690155 30821 691231
rect 31573 690155 31574 691231
rect 30820 690154 31574 690155
rect 37358 689663 38120 689664
rect 37358 688581 37359 689663
rect 38119 688581 38120 689663
rect 37358 688580 38120 688581
rect 675408 677722 676490 677746
rect 675408 676672 675432 677722
rect 676466 676672 676490 677722
rect 675408 676648 676490 676672
rect 671702 676104 672784 676128
rect 671702 675054 671726 676104
rect 672760 675054 672784 676104
rect 671702 675030 672784 675054
rect 686012 674431 686766 674432
rect 686012 673355 686013 674431
rect 686765 673355 686766 674431
rect 686012 673354 686766 673355
rect 679466 672863 680228 672864
rect 679466 671781 679467 672863
rect 680227 671781 680228 672863
rect 679466 671780 680228 671781
rect 30820 648031 31574 648032
rect 30820 646955 30821 648031
rect 31573 646955 31574 648031
rect 30820 646954 31574 646955
rect 37358 646463 38120 646464
rect 37358 645381 37359 646463
rect 38119 645381 38120 646463
rect 37358 645380 38120 645381
rect 675408 632722 676490 632746
rect 675408 631672 675432 632722
rect 676466 631672 676490 632722
rect 675408 631648 676490 631672
rect 671702 631104 672784 631128
rect 671702 630054 671726 631104
rect 672760 630054 672784 631104
rect 671702 630030 672784 630054
rect 686012 629431 686766 629432
rect 686012 628355 686013 629431
rect 686765 628355 686766 629431
rect 686012 628354 686766 628355
rect 679466 627863 680228 627864
rect 679466 626781 679467 627863
rect 680227 626781 680228 627863
rect 679466 626780 680228 626781
rect 30820 604831 31574 604832
rect 30820 603755 30821 604831
rect 31573 603755 31574 604831
rect 30820 603754 31574 603755
rect 37358 603263 38120 603264
rect 37358 602181 37359 603263
rect 38119 602181 38120 603263
rect 37358 602180 38120 602181
rect 675408 587522 676490 587546
rect 675408 586472 675432 587522
rect 676466 586472 676490 587522
rect 675408 586448 676490 586472
rect 671702 585904 672784 585928
rect 671702 584854 671726 585904
rect 672760 584854 672784 585904
rect 671702 584830 672784 584854
rect 686012 584231 686766 584232
rect 686012 583155 686013 584231
rect 686765 583155 686766 584231
rect 686012 583154 686766 583155
rect 679466 582663 680228 582664
rect 679466 581581 679467 582663
rect 680227 581581 680228 582663
rect 679466 581580 680228 581581
rect 30820 561631 31574 561632
rect 30820 560555 30821 561631
rect 31573 560555 31574 561631
rect 30820 560554 31574 560555
rect 37358 560063 38120 560064
rect 37358 558981 37359 560063
rect 38119 558981 38120 560063
rect 37358 558980 38120 558981
rect 675408 542522 676490 542546
rect 675408 541472 675432 542522
rect 676466 541472 676490 542522
rect 675408 541448 676490 541472
rect 671702 540904 672784 540928
rect 671702 539854 671726 540904
rect 672760 539854 672784 540904
rect 671702 539830 672784 539854
rect 686012 539231 686766 539232
rect 686012 538155 686013 539231
rect 686765 538155 686766 539231
rect 686012 538154 686766 538155
rect 679466 537663 680228 537664
rect 679466 536581 679467 537663
rect 680227 536581 680228 537663
rect 679466 536580 680228 536581
rect 675408 498522 676490 498546
rect 675408 497472 675432 498522
rect 676466 497472 676490 498522
rect 675408 497448 676490 497472
rect 671702 496904 672784 496928
rect 671702 495854 671726 496904
rect 672760 495854 672784 496904
rect 671702 495830 672784 495854
rect 686012 495231 686766 495232
rect 686012 494155 686013 495231
rect 686765 494155 686766 495231
rect 686012 494154 686766 494155
rect 679466 493663 680228 493664
rect 679466 492581 679467 493663
rect 680227 492581 680228 493663
rect 679466 492580 680228 492581
rect 30820 434031 31574 434032
rect 30820 432955 30821 434031
rect 31573 432955 31574 434031
rect 30820 432954 31574 432955
rect 37358 432463 38120 432464
rect 37358 431381 37359 432463
rect 38119 431381 38120 432463
rect 37358 431380 38120 431381
rect 675408 410322 676490 410346
rect 675408 409272 675432 410322
rect 676466 409272 676490 410322
rect 675408 409248 676490 409272
rect 671702 408704 672784 408728
rect 671702 407654 671726 408704
rect 672760 407654 672784 408704
rect 671702 407630 672784 407654
rect 686012 407031 686766 407032
rect 686012 405955 686013 407031
rect 686765 405955 686766 407031
rect 686012 405954 686766 405955
rect 679466 405463 680228 405464
rect 679466 404381 679467 405463
rect 680227 404381 680228 405463
rect 679466 404380 680228 404381
rect 30820 390831 31574 390832
rect 30820 389755 30821 390831
rect 31573 389755 31574 390831
rect 30820 389754 31574 389755
rect 37358 389263 38120 389264
rect 37358 388181 37359 389263
rect 38119 388181 38120 389263
rect 37358 388180 38120 388181
rect 675408 365122 676490 365146
rect 675408 364072 675432 365122
rect 676466 364072 676490 365122
rect 675408 364048 676490 364072
rect 671702 363504 672784 363528
rect 671702 362454 671726 363504
rect 672760 362454 672784 363504
rect 671702 362430 672784 362454
rect 686012 361831 686766 361832
rect 686012 360755 686013 361831
rect 686765 360755 686766 361831
rect 686012 360754 686766 360755
rect 679466 360263 680228 360264
rect 679466 359181 679467 360263
rect 680227 359181 680228 360263
rect 679466 359180 680228 359181
rect 30820 347631 31574 347632
rect 30820 346555 30821 347631
rect 31573 346555 31574 347631
rect 30820 346554 31574 346555
rect 37358 346063 38120 346064
rect 37358 344981 37359 346063
rect 38119 344981 38120 346063
rect 37358 344980 38120 344981
rect 675408 320122 676490 320146
rect 675408 319072 675432 320122
rect 676466 319072 676490 320122
rect 675408 319048 676490 319072
rect 671702 318504 672784 318528
rect 671702 317454 671726 318504
rect 672760 317454 672784 318504
rect 671702 317430 672784 317454
rect 686012 316831 686766 316832
rect 686012 315755 686013 316831
rect 686765 315755 686766 316831
rect 686012 315754 686766 315755
rect 679466 315263 680228 315264
rect 679466 314181 679467 315263
rect 680227 314181 680228 315263
rect 679466 314180 680228 314181
rect 30820 304431 31574 304432
rect 30820 303355 30821 304431
rect 31573 303355 31574 304431
rect 30820 303354 31574 303355
rect 37358 302863 38120 302864
rect 37358 301781 37359 302863
rect 38119 301781 38120 302863
rect 37358 301780 38120 301781
rect 675408 275122 676490 275146
rect 675408 274072 675432 275122
rect 676466 274072 676490 275122
rect 675408 274048 676490 274072
rect 671702 273504 672784 273528
rect 671702 272454 671726 273504
rect 672760 272454 672784 273504
rect 671702 272430 672784 272454
rect 686012 271831 686766 271832
rect 686012 270755 686013 271831
rect 686765 270755 686766 271831
rect 686012 270754 686766 270755
rect 679466 270263 680228 270264
rect 679466 269181 679467 270263
rect 680227 269181 680228 270263
rect 679466 269180 680228 269181
rect 30820 261231 31574 261232
rect 30820 260155 30821 261231
rect 31573 260155 31574 261231
rect 30820 260154 31574 260155
rect 37358 259663 38120 259664
rect 37358 258581 37359 259663
rect 38119 258581 38120 259663
rect 37358 258580 38120 258581
rect 674156 249272 676452 249296
rect 674156 246640 674180 249272
rect 676428 246640 676452 249272
rect 674156 246616 676452 246640
rect 41066 245364 43530 245388
rect 41066 238386 41090 245364
rect 43506 238386 43530 245364
rect 41066 238362 43530 238386
rect 44254 241334 46718 241358
rect 44254 234556 44278 241334
rect 46694 234556 46718 241334
rect 44254 234532 46718 234556
rect 675408 229922 676490 229946
rect 675408 228872 675432 229922
rect 676466 228872 676490 229922
rect 675408 228848 676490 228872
rect 671702 228304 672784 228328
rect 671702 227254 671726 228304
rect 672760 227254 672784 228304
rect 671702 227230 672784 227254
rect 686012 226631 686766 226632
rect 686012 225555 686013 226631
rect 686765 225555 686766 226631
rect 686012 225554 686766 225555
rect 679466 225063 680228 225064
rect 679466 223981 679467 225063
rect 680227 223981 680228 225063
rect 679466 223980 680228 223981
rect 30820 218031 31574 218032
rect 30820 216955 30821 218031
rect 31573 216955 31574 218031
rect 30820 216954 31574 216955
rect 37358 216463 38120 216464
rect 37358 215381 37359 216463
rect 38119 215381 38120 216463
rect 37358 215380 38120 215381
rect 675408 184922 676490 184946
rect 675408 183872 675432 184922
rect 676466 183872 676490 184922
rect 675408 183848 676490 183872
rect 671702 183304 672784 183328
rect 671702 182254 671726 183304
rect 672760 182254 672784 183304
rect 671702 182230 672784 182254
rect 686012 181631 686766 181632
rect 686012 180555 686013 181631
rect 686765 180555 686766 181631
rect 686012 180554 686766 180555
rect 679466 180063 680228 180064
rect 679466 178981 679467 180063
rect 680227 178981 680228 180063
rect 679466 178980 680228 178981
rect 675408 139722 676490 139746
rect 675408 138672 675432 139722
rect 676466 138672 676490 139722
rect 675408 138648 676490 138672
rect 671702 138104 672784 138128
rect 671702 137054 671726 138104
rect 672760 137054 672784 138104
rect 671702 137030 672784 137054
rect 686012 136431 686766 136432
rect 686012 135355 686013 136431
rect 686765 135355 686766 136431
rect 686012 135354 686766 135355
rect 679466 134863 680228 134864
rect 679466 133781 679467 134863
rect 680227 133781 680228 134863
rect 679466 133780 680228 133781
rect 234842 38177 237788 38178
rect 234842 37337 234843 38177
rect 237787 37337 237788 38177
rect 234842 37336 237788 37337
rect 149632 35995 150436 35996
rect 149632 35167 149633 35995
rect 150435 35167 150436 35995
rect 149632 35166 150436 35167
rect 148098 34787 148902 34788
rect 148098 33959 148099 34787
rect 148901 33959 148902 34787
rect 642026 34759 643634 34760
rect 642026 33989 642027 34759
rect 643633 33989 643634 34759
rect 642026 33988 643634 33989
rect 148098 33958 148902 33959
rect 204996 31645 207928 31646
rect 204996 30787 204997 31645
rect 207927 30787 207928 31645
rect 204996 30786 207928 30787
<< metal1 >>
rect 648104 47124 649670 47188
rect 648104 46660 648166 47124
rect 649608 46738 649670 47124
rect 649608 46660 650160 46738
rect 648104 46598 650160 46660
rect 648104 46590 649670 46598
<< via1 >>
rect 648166 46660 649608 47124
<< metal2 >>
rect 648104 47124 649670 47188
rect 648104 46660 648166 47124
rect 649608 46660 649670 47124
rect 648104 46590 649670 46660
<< via2 >>
rect 648166 46660 649608 47124
<< metal3 >>
rect 575700 997314 580479 997678
rect 575700 995032 575762 997314
rect 580384 995032 580479 997314
rect 585678 997328 590458 997678
rect 585678 995032 585758 997328
rect 590380 995032 590458 997328
rect 39852 842324 50002 842458
rect 39852 837800 47908 842324
rect 49694 837800 50002 842324
rect 39852 837678 50002 837800
rect 667172 833206 677818 833301
rect 39852 832392 50002 832479
rect 39852 827868 47908 832392
rect 49694 827868 50002 832392
rect 667172 828630 667284 833206
rect 669732 828630 677818 833206
rect 667172 828521 677818 828630
rect 39852 827699 50002 827868
rect 667172 823212 677818 823322
rect 667172 818636 667270 823212
rect 669718 818636 677818 823212
rect 667172 818542 677818 818636
rect 667062 518582 677700 518701
rect 667062 514056 667336 518582
rect 669706 514056 677700 518582
rect 667062 513921 677700 514056
rect 667062 508592 677700 508722
rect 667062 504066 667350 508592
rect 669720 504066 677700 508592
rect 667062 503942 677700 504066
rect 39924 497732 52292 497858
rect 39924 493250 50364 497732
rect 52092 493250 52292 497732
rect 39924 493078 52292 493250
rect 39924 487742 52292 487879
rect 39924 483260 50352 487742
rect 52080 483260 52292 487742
rect 39924 483099 52292 483260
rect 663914 430390 677712 430501
rect 663914 425684 664134 430390
rect 666540 425748 677712 430390
rect 666540 425684 667110 425748
rect 663914 425562 667110 425684
rect 663914 420462 677712 420522
rect 663914 415856 664112 420462
rect 666528 415856 677712 420462
rect 663914 415742 677712 415856
rect 39456 82706 45844 82744
rect 39456 78242 41946 82706
rect 45672 78242 45844 82706
rect 39456 78151 45844 78242
rect 39456 72802 45844 72900
rect 39456 68338 41922 72802
rect 45648 68338 45844 72802
rect 39456 68256 45844 68338
rect 648104 47124 649670 47188
rect 241690 46616 246049 46686
rect 241690 42842 241740 46616
rect 245986 42842 246049 46616
rect 149600 41148 150458 41207
rect 149600 40988 149618 41148
rect 150440 40988 150458 41148
rect 148068 40752 148926 40782
rect 148068 40592 148086 40752
rect 148908 40592 148926 40752
rect 148068 34788 148926 40592
rect 149600 35996 150458 40988
rect 241690 39426 246049 42842
rect 251300 46630 255702 46686
rect 251300 42856 251392 46630
rect 255638 42856 255702 46630
rect 648104 46660 648166 47124
rect 649608 46660 649670 47124
rect 648104 46590 649670 46660
rect 653462 45026 656910 45156
rect 251300 39426 255702 42856
rect 641954 43988 643694 44026
rect 641954 42198 641994 43988
rect 643660 42198 643694 43988
rect 149600 35166 149632 35996
rect 150436 35166 150458 35996
rect 149600 35114 150458 35166
rect 234814 38178 237814 38242
rect 234814 37336 234842 38178
rect 237788 37336 237814 38178
rect 148068 33958 148098 34788
rect 148902 33958 148926 34788
rect 148068 33900 148926 33958
rect 204958 31646 207958 31734
rect 204958 30786 204996 31646
rect 207928 30786 207958 31646
rect 204958 18004 207958 30786
rect 234814 19380 237814 37336
rect 641954 34760 643694 42198
rect 653462 42634 653578 45026
rect 656772 42634 656910 45026
rect 653462 35808 656910 42634
rect 641954 33988 642026 34760
rect 643634 33988 643694 34760
rect 641954 33920 643694 33988
rect 234814 18544 234884 19380
rect 237754 18544 237814 19380
rect 234814 18466 237814 18544
rect 204958 17128 205020 18004
rect 207872 17128 207958 18004
rect 204958 17038 207958 17128
<< via3 >>
rect 575762 994884 580384 997314
rect 585758 994898 590380 997328
rect 47908 837800 49694 842324
rect 47908 827868 49694 832392
rect 667284 828630 669732 833206
rect 667270 818636 669718 823212
rect 667336 514056 669706 518582
rect 667350 504066 669720 508592
rect 50364 493250 52092 497732
rect 50352 483260 52080 487742
rect 664134 425684 666540 430390
rect 664112 415856 666528 420462
rect 41946 78242 45672 82706
rect 41922 68338 45648 72802
rect 241740 42842 245986 46616
rect 149618 40988 150440 41148
rect 148086 40592 148908 40752
rect 251392 42856 255638 46630
rect 648166 46660 649608 47124
rect 641994 42198 643660 43988
rect 149632 35166 150436 35996
rect 234842 37336 237788 38178
rect 148098 33958 148902 34788
rect 204996 30786 207928 31646
rect 653578 42634 656772 45026
rect 642026 33988 643634 34760
rect 234884 18544 237754 19380
rect 205020 17128 207872 18004
<< metal4 >>
rect 575680 997314 580478 997462
rect 575680 994884 575762 997314
rect 580384 994884 580478 997314
rect 575680 994804 580478 994884
rect 585670 997328 590468 997462
rect 585670 994898 585758 997328
rect 590380 994898 590468 997328
rect 585670 994804 590468 994898
rect 47792 842324 49822 842462
rect 47792 837800 47908 842324
rect 49694 837800 49822 842324
rect 47792 837658 49822 837800
rect 667202 833206 669802 833310
rect 47792 832392 49822 832506
rect 47792 827868 47908 832392
rect 49694 827868 49822 832392
rect 667202 828630 667284 833206
rect 669732 828630 669802 833206
rect 667202 828520 669802 828630
rect 47792 827702 49822 827868
rect 667214 823212 669814 823336
rect 667214 818636 667270 823212
rect 669718 818636 669814 823212
rect 667214 818546 669814 818636
rect 667206 518582 669814 518696
rect 667206 514056 667336 518582
rect 669706 514056 669814 518582
rect 667206 513920 669814 514056
rect 667218 508592 669826 508726
rect 667218 504066 667350 508592
rect 669720 504066 669826 508592
rect 667218 503950 669826 504066
rect 50172 497732 52196 497874
rect 50172 493250 50364 497732
rect 52092 493250 52196 497732
rect 50172 493084 52196 493250
rect 50198 487742 52222 487884
rect 50198 483260 50352 487742
rect 52080 483260 52222 487742
rect 50198 483094 52222 483260
rect 664008 430390 666612 430490
rect 664008 425684 664134 430390
rect 666540 425684 666612 430390
rect 664008 425572 666612 425684
rect 664018 420462 666634 420524
rect 664018 415856 664112 420462
rect 666528 415856 666634 420462
rect 664018 415760 666634 415856
rect 393442 269370 394228 269470
rect 393442 266556 393536 269370
rect 394142 266556 394228 269370
rect 393442 266474 394228 266556
rect 394044 262208 394224 266474
rect 409094 265462 409274 265476
rect 408466 265334 409274 265462
rect 408466 262926 408538 265334
rect 409192 262926 409274 265334
rect 408466 262854 409274 262926
rect 409094 262244 409274 262854
rect 47770 261338 59470 261466
rect 47770 258676 48050 261338
rect 49608 261232 59470 261338
rect 49608 258676 56554 261232
rect 47770 258660 56554 258676
rect 59352 258660 59470 261232
rect 47770 258466 59470 258660
rect 394504 261336 395406 261450
rect 394504 258566 394590 261336
rect 395320 258566 395406 261336
rect 394504 258468 395406 258566
rect 50170 257338 60588 257466
rect 50170 254676 50450 257338
rect 52008 257232 60588 257338
rect 52008 254676 56554 257232
rect 50170 254660 56554 254676
rect 60330 254660 60588 257232
rect 50170 254466 60588 254660
rect 409686 257378 410808 257470
rect 409686 254558 409786 257378
rect 410720 254558 410808 257378
rect 409686 254452 410808 254558
rect 52578 253402 63292 253466
rect 52578 250538 52654 253402
rect 53746 253396 63292 253402
rect 53746 250548 56204 253396
rect 63216 250548 63292 253396
rect 53746 250538 63292 250548
rect 52578 250466 63292 250538
rect 211712 253384 212610 253472
rect 211712 250572 211800 253384
rect 212518 250572 212610 253384
rect 211712 250470 212610 250572
rect 241812 253384 242710 253472
rect 241812 250572 241900 253384
rect 242618 250572 242710 253384
rect 241812 250470 242710 250572
rect 272232 253384 272620 253472
rect 272232 250470 272620 250572
rect 302162 253384 302714 253472
rect 302162 250470 302714 250572
rect 332112 253384 333010 253472
rect 332112 250572 332200 253384
rect 332918 250572 333010 253384
rect 332112 250470 333010 250572
rect 362212 253384 363110 253472
rect 362212 250572 362300 253384
rect 363018 250572 363110 253384
rect 362212 250470 363110 250572
rect 392572 253384 393110 253472
rect 393018 250572 393110 253384
rect 392572 250470 393110 250572
rect 196676 249384 197618 249464
rect 196676 246554 196766 249384
rect 197520 246554 197618 249384
rect 196676 246468 197618 246554
rect 226776 249384 227718 249464
rect 226776 246554 226866 249384
rect 227620 246554 227718 249384
rect 226776 246468 227718 246554
rect 256876 249384 257818 249464
rect 256876 246554 256966 249384
rect 257720 246554 257818 249384
rect 287156 249384 287658 249464
rect 347176 249384 348118 249464
rect 256876 246468 257818 246554
rect 317354 246468 317802 246554
rect 347176 246554 347266 249384
rect 348020 246554 348118 249384
rect 347176 246468 348118 246554
rect 377176 249384 378118 249464
rect 377176 246554 377266 249384
rect 378020 246554 378118 249384
rect 377176 246468 378118 246554
rect 407176 249384 408118 249464
rect 407176 246554 407266 249384
rect 408020 246554 408118 249384
rect 407176 246468 408118 246554
rect 666890 249296 676670 249476
rect 666890 249288 674156 249296
rect 666890 246662 667058 249288
rect 669642 246662 674156 249288
rect 666890 246616 674156 246662
rect 676452 246616 676670 249296
rect 666890 246466 676670 246616
rect 40984 245388 63434 245466
rect 40984 238362 41066 245388
rect 43530 245296 63434 245388
rect 43530 242590 56394 245296
rect 63344 242590 63434 245296
rect 43530 242466 63434 242590
rect 212568 245420 213540 245462
rect 212568 242526 212622 245420
rect 213464 242526 213540 245420
rect 43530 238362 43612 242466
rect 212568 242464 213540 242526
rect 242668 245420 243640 245462
rect 242668 242526 242722 245420
rect 243564 242526 243640 245420
rect 242668 242464 243640 242526
rect 272982 245420 273314 245462
rect 272982 242464 273314 242526
rect 303168 245420 303460 245462
rect 303168 242464 303460 242526
rect 332968 245420 333940 245462
rect 332968 242526 333022 245420
rect 333864 242526 333940 245420
rect 332968 242464 333940 242526
rect 363068 245420 364040 245462
rect 363068 242526 363122 245420
rect 363964 242526 364040 245420
rect 363068 242464 364040 242526
rect 393210 245420 393800 245462
rect 393210 242464 393800 242526
rect 40984 238266 43612 238362
rect 44196 241358 63434 241466
rect 44196 234532 44254 241358
rect 46718 241330 63434 241358
rect 46718 238624 56424 241330
rect 63344 238624 63434 241330
rect 46718 238466 63434 238624
rect 197542 241402 198398 241470
rect 197542 238534 197632 241402
rect 198322 238534 198398 241402
rect 197542 238480 198398 238534
rect 227642 241402 228498 241470
rect 227642 238534 227732 241402
rect 228422 238534 228498 241402
rect 227642 238480 228498 238534
rect 257742 241402 258598 241470
rect 257742 238534 257832 241402
rect 258522 238534 258598 241402
rect 257742 238480 258598 238534
rect 288068 241402 288566 241470
rect 288068 238480 288566 238534
rect 318226 241402 318574 241470
rect 318226 238480 318574 238534
rect 348042 241402 348898 241470
rect 348042 238534 348132 241402
rect 348822 238534 348898 241402
rect 348042 238480 348898 238534
rect 378042 241402 378898 241470
rect 378042 238534 378132 241402
rect 378822 238534 378898 241402
rect 378042 238480 378898 238534
rect 408410 241402 408734 241470
rect 408410 238480 408734 238534
rect 46718 234532 46802 238466
rect 44196 234466 46802 234532
rect 47786 237372 63250 237466
rect 47786 237366 56424 237372
rect 47786 234588 47980 237366
rect 50678 234594 56424 237366
rect 63122 234594 63250 237372
rect 50678 234588 63250 234594
rect 47786 234466 63250 234588
rect 210866 237386 211814 237474
rect 210866 234540 210958 237386
rect 211722 234540 211814 237386
rect 210866 234448 211814 234540
rect 240966 237386 241914 237474
rect 240966 234540 241058 237386
rect 241822 234540 241914 237386
rect 240966 234448 241914 234540
rect 271344 237386 272014 237474
rect 271922 234540 272014 237386
rect 331414 237386 332214 237474
rect 271344 234448 272014 234540
rect 302022 234540 302114 237290
rect 301514 234448 302114 234540
rect 332122 234540 332214 237386
rect 331414 234448 332214 234540
rect 361366 237386 362314 237474
rect 361366 234540 361458 237386
rect 362222 234540 362314 237386
rect 361366 234448 362314 234540
rect 391834 237386 392314 237474
rect 392222 234540 392314 237386
rect 391834 234448 392314 234540
rect 44186 233340 63160 233466
rect 44186 230606 56406 233340
rect 63018 230606 63160 233340
rect 89776 232386 90096 233602
rect 93776 232386 94096 233602
rect 89776 232258 94096 232386
rect 89776 231398 89900 232258
rect 93968 231398 94096 232258
rect 89776 231266 94096 231398
rect 169776 232338 170096 233638
rect 173776 232338 174096 233612
rect 169776 232252 174096 232338
rect 169776 231392 169864 232252
rect 173932 231392 174096 232252
rect 169776 231302 174096 231392
rect 195988 233390 196616 233464
rect 44186 230466 63160 230606
rect 195988 230538 196058 233390
rect 196556 230538 196616 233390
rect 195988 230466 196616 230538
rect 226088 233390 226716 233464
rect 226088 230538 226158 233390
rect 226656 230538 226716 233390
rect 226088 230466 226716 230538
rect 256188 233390 256816 233464
rect 256188 230538 256258 233390
rect 256756 230538 256816 233390
rect 256188 230466 256816 230538
rect 286288 233390 286916 233464
rect 286288 230538 286358 233390
rect 286856 230538 286916 233390
rect 286288 230466 286916 230538
rect 316388 233390 317016 233464
rect 316388 230538 316458 233390
rect 316956 230538 317016 233390
rect 316388 230466 317016 230538
rect 346488 233390 347116 233464
rect 346488 230538 346558 233390
rect 347056 230538 347116 233390
rect 346488 230466 347116 230538
rect 376488 233390 377116 233464
rect 376488 230538 376558 233390
rect 377056 230538 377116 233390
rect 376488 230466 377116 230538
rect 406660 233390 407116 233464
rect 407056 230538 407116 233390
rect 429776 232520 430096 233612
rect 433776 232520 434096 233612
rect 429776 232370 434096 232520
rect 429776 231510 429910 232370
rect 433978 231510 434096 232370
rect 429776 231392 434096 231510
rect 406660 230466 407116 230538
rect 44198 197498 46798 230466
rect 598368 212326 610962 212504
rect 598368 209740 598598 212326
rect 601098 209740 607452 212326
rect 609952 209740 610962 212326
rect 598368 209504 610962 209740
rect 641044 212352 642108 212460
rect 641044 209640 641152 212352
rect 642010 209640 642108 212352
rect 641044 209528 642108 209640
rect 596262 208442 605388 208502
rect 596262 207926 596332 208442
rect 597664 208434 605388 208442
rect 597664 207934 602456 208434
rect 605326 207934 605388 208434
rect 597664 207926 605388 207934
rect 596262 207862 605388 207926
rect 610642 207692 610962 209504
rect 641362 207684 641682 209528
rect 598496 197778 601174 197876
rect 44198 197454 52344 197498
rect 44198 196934 51420 197454
rect 52282 196934 52344 197454
rect 598496 197108 598684 197778
rect 601038 197528 601174 197778
rect 601038 197492 606976 197528
rect 601038 197238 606016 197492
rect 606936 197238 606976 197492
rect 601038 197208 606976 197238
rect 601038 197108 601174 197208
rect 598496 196992 601174 197108
rect 44198 196858 52344 196934
rect 44198 176742 46798 196858
rect 596072 184442 605388 184502
rect 596072 183902 596116 184442
rect 596848 184418 605388 184442
rect 596848 183918 602456 184418
rect 605326 183918 605388 184418
rect 596848 183902 605388 183918
rect 596072 183862 605388 183902
rect 41864 176610 46798 176742
rect 41864 173284 42002 176610
rect 45608 173284 46798 176610
rect 41864 173126 46798 173284
rect 42646 171444 52246 171498
rect 42646 170908 42828 171444
rect 45682 171440 52246 171444
rect 45682 170920 51312 171440
rect 52174 170920 52246 171440
rect 45682 170908 52246 170920
rect 42646 170858 52246 170908
rect 598496 167138 601174 167236
rect 598496 166468 598684 167138
rect 601038 166892 601174 167138
rect 601038 166866 606976 166892
rect 601038 166608 605986 166866
rect 606932 166608 606976 166866
rect 601038 166572 606976 166608
rect 601038 166468 601174 166572
rect 598496 166352 601174 166468
rect 594072 158446 605388 158502
rect 594072 157906 594114 158446
rect 596846 158430 605388 158446
rect 596846 157930 602430 158430
rect 605300 157930 605388 158430
rect 596846 157906 605388 157930
rect 594072 157862 605388 157906
rect 42578 145450 52178 145498
rect 42578 144914 42842 145450
rect 45696 145432 52178 145450
rect 45696 144914 51246 145432
rect 42578 144912 51246 144914
rect 52108 144912 52178 145432
rect 42578 144858 52178 144912
rect 598496 136498 601174 136596
rect 598496 135828 598684 136498
rect 601038 136256 601174 136498
rect 601038 136230 606976 136256
rect 601038 135964 605972 136230
rect 606926 135964 606976 136230
rect 601038 135936 606976 135964
rect 601038 135828 601174 135936
rect 598496 135712 601174 135828
rect 594072 132440 605388 132502
rect 594072 131900 594124 132440
rect 596856 132414 605388 132440
rect 596856 131914 602456 132414
rect 605326 131914 605388 132414
rect 596856 131900 605388 131914
rect 594072 131862 605388 131900
rect 42578 119446 52178 119498
rect 42578 118910 42832 119446
rect 45686 119438 52178 119446
rect 45686 118918 51242 119438
rect 52104 118918 52178 119438
rect 45686 118910 52178 118918
rect 42578 118858 52178 118910
rect 594072 106446 605388 106502
rect 594072 105906 594126 106446
rect 596858 106426 605388 106446
rect 596858 105926 602460 106426
rect 605330 105926 605388 106426
rect 596858 105906 605388 105926
rect 594072 105862 605388 105906
rect 598496 105620 601174 105676
rect 598496 105594 606976 105620
rect 598496 105578 605980 105594
rect 598496 104908 598684 105578
rect 601038 105326 605980 105578
rect 606942 105326 606976 105594
rect 601038 105300 606976 105326
rect 601038 104908 601174 105300
rect 598496 104792 601174 104908
rect 626002 98760 626322 102316
rect 656722 98804 657042 102238
rect 625442 98656 626852 98760
rect 625442 96074 625556 98656
rect 626744 96074 626852 98656
rect 636080 98622 636994 98758
rect 636080 96584 636216 98622
rect 636858 96584 636994 98622
rect 636080 96434 636994 96584
rect 656284 98712 657602 98804
rect 625442 95956 626852 96074
rect 636354 94448 636674 96434
rect 656284 96142 656422 98712
rect 657500 96142 657602 98712
rect 656284 96050 657602 96142
rect 42578 93444 52178 93498
rect 42578 92908 42828 93444
rect 45682 93434 52178 93444
rect 45682 92914 51246 93434
rect 52108 92914 52178 93434
rect 45682 92908 52178 92914
rect 42578 92858 52178 92908
rect 41864 82706 45778 82794
rect 41864 78242 41946 82706
rect 45672 78242 45778 82706
rect 632354 80924 632674 82062
rect 640354 81016 640674 82000
rect 632072 80776 633010 80924
rect 594072 80456 605388 80502
rect 594072 79916 594120 80456
rect 596852 80438 605388 80456
rect 596852 79938 602454 80438
rect 605324 79938 605388 80438
rect 596852 79916 605388 79938
rect 594072 79862 605388 79916
rect 41864 78154 45778 78242
rect 632072 78326 632200 80776
rect 632864 78326 633010 80776
rect 632072 78198 633010 78326
rect 640098 80900 640922 81016
rect 640098 78256 640210 80900
rect 640810 78256 640922 80900
rect 640098 78134 640922 78256
rect 41858 72802 45772 72890
rect 41858 68338 41922 72802
rect 45648 68338 45772 72802
rect 41858 68250 45772 68338
rect 41862 67438 52362 67498
rect 41862 66902 41936 67438
rect 45690 67436 52362 67438
rect 45690 66916 51444 67436
rect 52306 66916 52362 67436
rect 45690 66902 52362 66916
rect 41862 66858 52362 66902
rect 41874 51988 58536 52122
rect 41874 48404 42006 51988
rect 45590 51954 58536 51988
rect 45590 48404 54526 51954
rect 41874 48370 54526 48404
rect 58210 48370 58536 51954
rect 143324 50624 144738 50688
rect 143324 50004 143390 50624
rect 144652 50004 144738 50624
rect 143324 49936 144738 50004
rect 143860 49638 144040 49936
rect 41874 48222 58536 48370
rect 641936 47627 650202 48027
rect 142560 45396 142740 47256
rect 141776 45394 142866 45396
rect 141376 45306 142866 45394
rect 141376 44206 141442 45306
rect 142810 44206 142866 45306
rect 141376 44130 142866 44206
rect 143440 40762 143620 47296
rect 144740 41158 144920 47340
rect 241680 46616 246056 46692
rect 241680 42842 241740 46616
rect 245986 42842 246056 46616
rect 241680 42784 246056 42842
rect 251302 46630 255700 46684
rect 251302 42856 251392 46630
rect 255638 42856 255700 46630
rect 251302 42788 255700 42856
rect 641936 43988 643718 47627
rect 661270 47282 669426 47320
rect 648104 47124 649670 47188
rect 648104 46660 648166 47124
rect 649608 46660 649670 47124
rect 648104 46590 649670 46660
rect 641936 42198 641994 43988
rect 643660 42198 643718 43988
rect 653432 45026 656912 47054
rect 661270 47030 666460 47282
rect 669380 47030 669426 47282
rect 661270 46991 669426 47030
rect 653432 42634 653578 45026
rect 656772 42634 656912 45026
rect 653432 42488 656912 42634
rect 641936 42164 643718 42198
rect 144740 41148 150516 41158
rect 144740 40988 149618 41148
rect 150440 40988 150516 41148
rect 144740 40978 150516 40988
rect 143440 40752 148940 40762
rect 143440 40592 148086 40752
rect 148908 40592 148940 40752
rect 143440 40582 148940 40592
rect 208850 19412 209170 19578
rect 208850 18506 208868 19412
rect 209130 18506 209170 19412
rect 204960 18004 207956 18076
rect 204960 17128 205020 18004
rect 207872 17128 207956 18004
rect 204960 17072 207956 17128
rect 208850 16308 209170 18506
rect 210400 18010 210720 19578
rect 210400 17104 210420 18010
rect 210682 17104 210720 18010
rect 210400 16308 210720 17104
rect 211950 19426 212270 19578
rect 211950 18520 211980 19426
rect 212242 18520 212270 19426
rect 211950 16308 212270 18520
rect 213500 18014 213820 19578
rect 213500 17108 213514 18014
rect 213776 17108 213820 18014
rect 213500 16308 213820 17108
rect 215050 19422 215370 19578
rect 215050 18516 215070 19422
rect 215332 18516 215370 19422
rect 215050 16308 215370 18516
rect 216600 18018 216920 19578
rect 216600 17112 216622 18018
rect 216884 17112 216920 18018
rect 216600 16308 216920 17112
rect 218150 19422 218470 19578
rect 218150 18516 218164 19422
rect 218426 18516 218470 19422
rect 218150 16308 218470 18516
rect 219700 18010 220020 19578
rect 219700 17104 219726 18010
rect 219988 17104 220020 18010
rect 219700 16308 220020 17104
rect 221250 19434 221570 19578
rect 221250 18528 221272 19434
rect 221534 18528 221570 19434
rect 221250 16308 221570 18528
rect 222800 18036 223120 19578
rect 234818 19380 237824 19480
rect 234818 18544 234884 19380
rect 237754 18544 237824 19380
rect 234818 18470 237824 18544
rect 222800 17130 222828 18036
rect 223090 17130 223120 18036
rect 222800 16308 223120 17130
<< via4 >>
rect 575762 994884 580384 997314
rect 585758 994898 590380 997328
rect 47908 837800 49694 842324
rect 47908 827868 49694 832392
rect 667284 828630 669732 833206
rect 667270 818636 669718 823212
rect 667336 514056 669706 518582
rect 667350 504066 669720 508592
rect 50364 493250 52092 497732
rect 50352 483260 52080 487742
rect 664134 425684 666540 430390
rect 664112 415856 666528 420462
rect 393536 266556 394142 269370
rect 408538 262926 409192 265334
rect 48050 258676 49608 261338
rect 56554 258660 59352 261232
rect 394590 258566 395320 261336
rect 50450 254676 52008 257338
rect 56554 254660 60330 257232
rect 409786 254558 410720 257378
rect 52654 250538 53746 253402
rect 56204 250548 63216 253396
rect 211800 250572 212518 253384
rect 241900 250572 242618 253384
rect 272232 250572 272620 253384
rect 302162 250572 302714 253384
rect 332200 250572 332918 253384
rect 362300 250572 363018 253384
rect 392572 250572 393018 253384
rect 196766 246554 197520 249384
rect 226866 246554 227620 249384
rect 256966 246554 257720 249384
rect 287156 246790 287658 249384
rect 317354 246554 317802 249324
rect 347266 246554 348020 249384
rect 377266 246554 378020 249384
rect 407266 246554 408020 249384
rect 667058 246662 669642 249288
rect 674156 246616 676452 249296
rect 41066 238362 43530 245388
rect 56394 242590 63344 245296
rect 212622 242526 213464 245420
rect 242722 242526 243564 245420
rect 272982 242526 273314 245420
rect 303168 242526 303460 245420
rect 333022 242526 333864 245420
rect 363122 242526 363964 245420
rect 393210 242526 393800 245420
rect 44254 234532 46718 241358
rect 56424 238624 63344 241330
rect 197632 238534 198322 241402
rect 227732 238534 228422 241402
rect 257832 238534 258522 241402
rect 288068 238534 288566 241402
rect 318226 238534 318574 241402
rect 348132 238534 348822 241402
rect 378132 238534 378822 241402
rect 408410 238534 408734 241402
rect 47980 234588 50678 237366
rect 56424 234594 63122 237372
rect 210958 234540 211722 237386
rect 241058 234540 241822 237386
rect 271344 234540 271922 237386
rect 301514 234540 302022 237290
rect 331414 234540 332122 237386
rect 361458 234540 362222 237386
rect 391834 234540 392222 237386
rect 56406 230606 63018 233340
rect 89900 231398 93968 232258
rect 169864 231392 173932 232252
rect 196058 230538 196556 233390
rect 226158 230538 226656 233390
rect 256258 230538 256756 233390
rect 286358 230538 286856 233390
rect 316458 230538 316956 233390
rect 346558 230538 347056 233390
rect 376558 230538 377056 233390
rect 406660 230538 407056 233390
rect 429910 231510 433978 232370
rect 598598 209740 601098 212326
rect 607452 209740 609952 212326
rect 641152 209640 642010 212352
rect 596332 207926 597664 208442
rect 602456 207934 605326 208434
rect 51420 196934 52282 197454
rect 598684 197108 601038 197778
rect 606016 197238 606936 197492
rect 596116 183902 596848 184442
rect 602456 183918 605326 184418
rect 42002 173284 45608 176610
rect 42828 170908 45682 171444
rect 51312 170920 52174 171440
rect 598684 166468 601038 167138
rect 605986 166608 606932 166866
rect 594114 157906 596846 158446
rect 602430 157930 605300 158430
rect 42842 144914 45696 145450
rect 51246 144912 52108 145432
rect 598684 135828 601038 136498
rect 605972 135964 606926 136230
rect 594124 131900 596856 132440
rect 602456 131914 605326 132414
rect 42832 118910 45686 119446
rect 51242 118918 52104 119438
rect 594126 105906 596858 106446
rect 602460 105926 605330 106426
rect 598684 104908 601038 105578
rect 605980 105326 606942 105594
rect 625556 96074 626744 98656
rect 636216 96584 636858 98622
rect 656422 96142 657500 98712
rect 42828 92908 45682 93444
rect 51246 92914 52108 93434
rect 41946 78242 45672 82706
rect 594120 79916 596852 80456
rect 602454 79938 605324 80438
rect 632200 78326 632864 80776
rect 640210 78256 640810 80900
rect 41922 68338 45648 72802
rect 41936 66902 45690 67438
rect 51444 66916 52306 67436
rect 42006 48404 45590 51988
rect 54526 48370 58210 51954
rect 143390 50004 144652 50624
rect 141442 44206 142810 45306
rect 241740 42842 245986 46616
rect 251392 42856 255638 46630
rect 648166 46660 649608 47124
rect 666460 47030 669380 47282
rect 208868 18506 209130 19412
rect 205020 17128 207872 18004
rect 210420 17104 210682 18010
rect 211980 18520 212242 19426
rect 213514 17108 213776 18014
rect 215070 18516 215332 19422
rect 216622 17112 216884 18018
rect 218164 18516 218426 19422
rect 219726 17104 219988 18010
rect 221272 18528 221534 19434
rect 234884 18544 237754 19380
rect 222828 17130 223090 18036
<< metal5 >>
rect 575640 997328 666620 997396
rect 575640 997314 585758 997328
rect 575640 994884 575762 997314
rect 580384 994898 585758 997314
rect 590380 994898 666620 997328
rect 580384 994884 666620 994898
rect 575640 994796 666620 994884
rect 47798 842324 49798 842560
rect 47798 837800 47908 842324
rect 49694 837800 49798 842324
rect 47798 832392 49798 837800
rect 47798 827868 47908 832392
rect 49694 827868 49798 832392
rect 47798 261338 49798 827868
rect 47798 258676 48050 261338
rect 49608 258676 49798 261338
rect 47798 258484 49798 258676
rect 50198 497732 52198 497992
rect 50198 493250 50364 497732
rect 52092 493250 52198 497732
rect 50198 487742 52198 493250
rect 50198 483260 50352 487742
rect 52080 483260 52198 487742
rect 50198 257338 52198 483260
rect 50198 254676 50450 257338
rect 52008 254676 52198 257338
rect 50198 254498 52198 254676
rect 52598 253402 53798 822658
rect 52598 250538 52654 253402
rect 53746 250538 53798 253402
rect 47836 237366 50836 237612
rect 47836 234588 47980 237366
rect 50678 234588 50836 237366
rect 47836 210498 50836 234588
rect 52598 217742 53798 250538
rect 54198 249466 55398 824290
rect 664020 430390 666620 994796
rect 664020 425684 664134 430390
rect 666540 425684 666620 430390
rect 664020 420462 666620 425684
rect 664020 415856 664112 420462
rect 666528 415856 666620 420462
rect 664020 269466 666620 415856
rect 58222 269370 666620 269466
rect 58222 266556 393536 269370
rect 394142 266556 666620 269370
rect 58222 266466 666620 266556
rect 667220 833206 669820 833474
rect 667220 828630 667284 833206
rect 669732 828630 669820 833206
rect 667220 823212 669820 828630
rect 667220 818636 667270 823212
rect 669718 818636 669820 823212
rect 667220 518582 669820 818636
rect 667220 514056 667336 518582
rect 669706 514056 669820 518582
rect 667220 508592 669820 514056
rect 667220 504066 667350 508592
rect 669720 504066 669820 508592
rect 667220 265466 669820 504066
rect 58222 265334 669820 265466
rect 58222 262926 408538 265334
rect 409192 262926 669820 265334
rect 58222 262466 669820 262926
rect 56370 261336 651174 261466
rect 56370 261232 394590 261336
rect 56370 258660 56554 261232
rect 59352 258660 394590 261232
rect 56370 258566 394590 258660
rect 395320 258566 651174 261336
rect 56370 258466 651174 258566
rect 56370 257378 651174 257466
rect 56370 257232 409786 257378
rect 56370 254660 56554 257232
rect 60330 254660 409786 257232
rect 56370 254558 409786 254660
rect 410720 254558 651174 257378
rect 56370 254466 651174 254558
rect 56126 253396 670986 253466
rect 56126 250548 56204 253396
rect 63216 253384 670986 253396
rect 63216 250572 211800 253384
rect 212518 250572 241900 253384
rect 242618 250572 272232 253384
rect 272620 250572 302162 253384
rect 302714 250572 332200 253384
rect 332918 250572 362300 253384
rect 363018 250572 392572 253384
rect 393018 250572 670986 253384
rect 63216 250548 670986 250572
rect 56126 250466 670986 250548
rect 54198 249384 669890 249466
rect 54198 246554 196766 249384
rect 197520 246554 226866 249384
rect 227620 246554 256966 249384
rect 257720 246790 287156 249384
rect 287658 249324 347266 249384
rect 287658 246790 317354 249324
rect 257720 246554 317354 246790
rect 317802 246554 347266 249324
rect 348020 246554 377266 249384
rect 378020 246554 407266 249384
rect 408020 249288 669890 249384
rect 408020 246662 667058 249288
rect 669642 246662 669890 249288
rect 408020 246554 669890 246662
rect 54198 246466 669890 246554
rect 54198 219342 55398 246466
rect 56278 245420 650946 245466
rect 56278 245296 212622 245420
rect 56278 242590 56394 245296
rect 63344 242590 212622 245296
rect 56278 242526 212622 242590
rect 213464 242526 242722 245420
rect 243564 242526 272982 245420
rect 273314 242526 303168 245420
rect 303460 242526 333022 245420
rect 333864 242526 363122 245420
rect 363964 242526 393210 245420
rect 393800 242526 650946 245420
rect 56278 242466 650946 242526
rect 56278 241402 650946 241466
rect 56278 241330 197632 241402
rect 56278 238624 56424 241330
rect 63344 238624 197632 241330
rect 56278 238534 197632 238624
rect 198322 238534 227732 241402
rect 228422 238534 257832 241402
rect 258522 238534 288068 241402
rect 288566 238534 318226 241402
rect 318574 238534 348132 241402
rect 348822 238534 378132 241402
rect 378822 238534 408410 241402
rect 408734 238534 650946 241402
rect 56278 238466 650946 238534
rect 56288 237386 605390 237466
rect 56288 237372 210958 237386
rect 56288 234594 56424 237372
rect 63122 234594 210958 237372
rect 56288 234540 210958 234594
rect 211722 234540 241058 237386
rect 241822 234540 271344 237386
rect 271922 237290 331414 237386
rect 271922 234540 301514 237290
rect 302022 234540 331414 237290
rect 332122 234540 361458 237386
rect 362222 234540 391834 237386
rect 392222 234540 605390 237386
rect 56288 234466 605390 234540
rect 56296 233390 601374 233466
rect 56296 233340 196058 233390
rect 56296 230606 56406 233340
rect 63018 232258 196058 233340
rect 63018 231398 89900 232258
rect 93968 232252 196058 232258
rect 93968 231398 169864 232252
rect 63018 231392 169864 231398
rect 173932 231392 196058 232252
rect 63018 230606 196058 231392
rect 56296 230538 196058 230606
rect 196556 230538 226158 233390
rect 226656 230538 256258 233390
rect 256756 230538 286358 233390
rect 286856 230538 316458 233390
rect 316956 230538 346558 233390
rect 347056 230538 376558 233390
rect 377056 230538 406660 233390
rect 407056 232370 601374 233390
rect 407056 231510 429910 232370
rect 433978 231510 601374 232370
rect 407056 230538 601374 231510
rect 56296 230466 601374 230538
rect 598374 212326 601374 230466
rect 47836 209858 53232 210498
rect 574646 209858 596910 210498
rect 47836 184498 50836 209858
rect 596270 208502 596910 209858
rect 598374 209740 598598 212326
rect 601098 209740 601374 212326
rect 596270 208442 597742 208502
rect 596270 207926 596332 208442
rect 597664 207926 597742 208442
rect 596270 207862 597742 207926
rect 598374 197778 601374 209740
rect 598374 197498 598684 197778
rect 51344 197454 53216 197498
rect 51344 196934 51420 197454
rect 52282 196934 53216 197454
rect 51344 196858 53216 196934
rect 574646 197108 598684 197498
rect 601038 197108 601374 197778
rect 574646 196858 601374 197108
rect 47836 183858 53212 184498
rect 574646 184442 596910 184498
rect 574646 183902 596116 184442
rect 596848 183902 596910 184442
rect 574646 183858 596910 183902
rect 41768 176610 45768 176874
rect 41768 173284 42002 176610
rect 45608 173284 45768 176610
rect 41768 171444 45768 173284
rect 41768 170908 42828 171444
rect 45682 170908 45768 171444
rect 41768 145450 45768 170908
rect 47836 166788 50836 183858
rect 598374 171498 601374 196858
rect 51246 171440 53240 171498
rect 51246 170920 51312 171440
rect 52174 170920 53240 171440
rect 51246 170858 53240 170920
rect 574646 170858 601374 171498
rect 41768 144914 42842 145450
rect 45696 144914 45768 145450
rect 41768 119446 45768 144914
rect 41768 118910 42832 119446
rect 45686 118910 45768 119446
rect 41768 93444 45768 118910
rect 41768 92908 42828 93444
rect 45682 92908 45768 93444
rect 41768 82706 45768 92908
rect 41768 78242 41946 82706
rect 45672 78242 45768 82706
rect 41768 72802 45768 78242
rect 41768 68338 41922 72802
rect 45648 68338 45768 72802
rect 41768 67438 45768 68338
rect 41768 66902 41936 67438
rect 45690 66902 45768 67438
rect 41768 51988 45768 66902
rect 41768 48404 42006 51988
rect 45590 48404 45768 51988
rect 41768 48074 45768 48404
rect 46836 158498 50836 166788
rect 598374 167138 601374 170858
rect 598374 166468 598684 167138
rect 601038 166468 601374 167138
rect 46836 157858 53220 158498
rect 574646 158446 596910 158498
rect 574646 157906 594114 158446
rect 596846 157906 596910 158446
rect 574646 157858 596910 157906
rect 46836 132498 50836 157858
rect 598374 145498 601374 166468
rect 51178 145432 53266 145498
rect 51178 144912 51246 145432
rect 52108 144912 53266 145432
rect 51178 144858 53266 144912
rect 574646 144858 601374 145498
rect 598374 136498 601374 144858
rect 598374 135828 598684 136498
rect 601038 135828 601374 136498
rect 46836 131858 53206 132498
rect 574646 132440 596910 132498
rect 574646 131900 594124 132440
rect 596856 131900 596910 132440
rect 574646 131858 596910 131900
rect 46836 106498 50836 131858
rect 598374 119498 601374 135828
rect 51178 119438 53266 119498
rect 51178 118918 51242 119438
rect 52104 118918 53266 119438
rect 51178 118858 53266 118918
rect 574646 118858 601374 119498
rect 46836 105858 53222 106498
rect 574646 106446 596910 106498
rect 574646 105906 594126 106446
rect 596858 105906 596910 106446
rect 574646 105858 596910 105906
rect 46836 80498 50836 105858
rect 598374 105578 601374 118858
rect 598374 104908 598684 105578
rect 601038 104908 601374 105578
rect 598374 93498 601374 104908
rect 51178 93434 53266 93498
rect 51178 92914 51246 93434
rect 52108 92914 53266 93434
rect 51178 92858 53266 92914
rect 574646 92858 601374 93498
rect 46836 79858 53168 80498
rect 574646 80456 596910 80498
rect 574646 79916 594120 80456
rect 596852 79916 596910 80456
rect 574646 79858 596910 79916
rect 46836 46788 50836 79858
rect 598374 67498 601374 92858
rect 51362 67436 53172 67498
rect 51362 66916 51444 67436
rect 52306 66916 53172 67436
rect 51362 66858 53172 66916
rect 574754 66858 601374 67498
rect 598374 52222 601374 66858
rect 54374 51954 601374 52222
rect 54374 48370 54526 51954
rect 58210 50624 601374 51954
rect 58210 50004 143390 50624
rect 144652 50004 601374 50624
rect 58210 48370 601374 50004
rect 54374 48222 601374 48370
rect 602390 224536 605390 234466
rect 648666 225872 651190 226192
rect 602390 224192 641044 224536
rect 602390 223872 641990 224192
rect 602390 223336 641044 223872
rect 602390 208434 605390 223336
rect 649990 222192 651190 225872
rect 648662 221872 651190 222192
rect 649990 212504 651190 221872
rect 607252 212352 669426 212504
rect 607252 212326 641152 212352
rect 607252 209740 607452 212326
rect 609952 209740 641152 212326
rect 607252 209640 641152 209740
rect 642010 209640 669426 212352
rect 607252 209504 669426 209640
rect 602390 207934 602456 208434
rect 605326 207934 605390 208434
rect 602390 184418 605390 207934
rect 666426 197528 669426 209504
rect 605976 197492 607594 197528
rect 605976 197238 606016 197492
rect 606936 197238 607594 197492
rect 605976 197208 607594 197238
rect 665238 197208 669426 197528
rect 602390 183918 602456 184418
rect 605326 183918 605390 184418
rect 602390 182210 605390 183918
rect 602390 181890 607594 182210
rect 602390 158430 605390 181890
rect 666426 166892 669426 197208
rect 605952 166866 607594 166892
rect 605952 166608 605986 166866
rect 606932 166608 607594 166866
rect 605952 166572 607594 166608
rect 665206 166572 669426 166892
rect 602390 157930 602430 158430
rect 605300 157930 605390 158430
rect 602390 151574 605390 157930
rect 602390 151254 607594 151574
rect 602390 132414 605390 151254
rect 666426 136256 669426 166572
rect 605940 136230 607594 136256
rect 605940 135964 605972 136230
rect 606926 135964 607594 136230
rect 605940 135936 607594 135964
rect 665164 135936 669426 136256
rect 602390 131914 602456 132414
rect 605326 131914 605390 132414
rect 602390 120938 605390 131914
rect 602390 120618 607610 120938
rect 602390 106426 605390 120618
rect 602390 105926 602460 106426
rect 605330 105926 605390 106426
rect 602390 98956 605390 105926
rect 666426 105620 669426 135936
rect 605940 105594 607594 105620
rect 605940 105326 605980 105594
rect 606942 105326 607594 105594
rect 605940 105300 607594 105326
rect 665176 105300 669426 105620
rect 602390 98712 657728 98956
rect 602390 98656 656422 98712
rect 602390 96074 625556 98656
rect 626744 98622 656422 98656
rect 626744 96584 636216 98622
rect 636858 96584 656422 98622
rect 626744 96142 656422 96584
rect 657500 96142 657728 98712
rect 626744 96074 657728 96142
rect 602390 95956 657728 96074
rect 602390 80438 605390 95956
rect 624824 89474 627824 95956
rect 643544 93474 646544 93588
rect 641906 93154 646544 93474
rect 624824 89154 629362 89474
rect 624824 89012 627824 89154
rect 643544 85474 646544 93154
rect 650994 92590 653994 95956
rect 666426 93406 669426 105300
rect 662522 93086 669426 93406
rect 650994 92270 657754 92590
rect 650994 90958 653994 92270
rect 666426 91774 669426 93086
rect 662484 91454 669426 91774
rect 650994 90638 657784 90958
rect 650994 90522 653994 90638
rect 666426 90142 669426 91454
rect 662504 89822 669426 90142
rect 641968 85154 646544 85474
rect 643544 81082 646544 85154
rect 666426 81082 669426 89822
rect 602390 79938 602454 80438
rect 605324 79938 605390 80438
rect 602390 47188 605390 79938
rect 632002 80900 669426 81082
rect 632002 80776 640210 80900
rect 632002 78326 632200 80776
rect 632864 78326 640210 80776
rect 632002 78256 640210 78326
rect 640810 78256 669426 80900
rect 632002 78082 669426 78256
rect 666426 47282 669426 78082
rect 602390 47124 649668 47188
rect 602390 46788 648166 47124
rect 46836 46660 648166 46788
rect 649608 46660 649668 47124
rect 666426 47030 666460 47282
rect 669380 47030 669426 47282
rect 666426 46978 669426 47030
rect 46836 46630 649668 46660
rect 46836 46616 251392 46630
rect 46836 45306 241740 46616
rect 46836 44206 141442 45306
rect 142810 44206 241740 45306
rect 46836 42842 241740 44206
rect 245986 42856 251392 46616
rect 255638 46588 649668 46630
rect 255638 45788 605390 46588
rect 255638 42856 605396 45788
rect 245986 42842 605396 42856
rect 46836 42788 605396 42842
rect 205820 19434 237824 19472
rect 205820 19426 221272 19434
rect 205820 19412 211980 19426
rect 205820 18506 208868 19412
rect 209130 18520 211980 19412
rect 212242 19422 221272 19426
rect 212242 18520 215070 19422
rect 209130 18516 215070 18520
rect 215332 18516 218164 19422
rect 218426 18528 221272 19422
rect 221534 19380 237824 19434
rect 221534 18544 234884 19380
rect 237754 18544 237824 19380
rect 221534 18528 237824 18544
rect 218426 18516 237824 18528
rect 209130 18506 237824 18516
rect 205820 18472 237824 18506
rect 204580 18036 224806 18072
rect 204580 18018 222828 18036
rect 204580 18014 216622 18018
rect 204580 18010 213514 18014
rect 204580 18004 210420 18010
rect 204580 17128 205020 18004
rect 207872 17128 210420 18004
rect 204580 17104 210420 17128
rect 210682 17108 213514 18010
rect 213776 17112 216622 18014
rect 216884 18010 222828 18018
rect 216884 17112 219726 18010
rect 213776 17108 219726 17112
rect 210682 17104 219726 17108
rect 219988 17130 222828 18010
rect 223090 17130 224806 18036
rect 219988 17104 224806 17130
rect 204580 17072 224806 17104
rect 204580 14000 205380 17072
rect 225246 15690 226046 18472
rect 224498 15370 226046 15690
rect 204580 13680 205930 14000
rect 204580 10620 205380 13680
rect 225246 12310 226046 15370
rect 224464 11990 226046 12310
rect 204580 10300 205808 10620
rect 204580 8096 205380 10300
rect 225246 8930 226046 11990
rect 224586 8610 226046 8930
rect 225246 7838 226046 8610
<< comment >>
rect 0 1037400 717600 1037600
rect 0 200 200 1037400
rect 717400 200 717600 1037400
rect 0 0 717600 200
use gpio_control_power_routing  gpio_control_power_routing_1
timestamp 1637447660
transform 1 0 -10 0 1 43200
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_0
timestamp 1637447660
transform 1 0 -10 0 1 0
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_13
timestamp 1637595202
transform -1 0 717846 0 1 -36400
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_14
timestamp 1637595202
transform -1 0 717846 0 1 -81600
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_11
timestamp 1637595202
transform -1 0 717846 0 1 53800
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_12
timestamp 1637595202
transform -1 0 717846 0 1 8600
box 6032 203748 46226 221470
use gpio_control_power_routing  gpio_control_power_routing_4
timestamp 1637447660
transform 1 0 -10 0 1 172800
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_3
timestamp 1637447660
transform 1 0 -10 0 1 129600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_2
timestamp 1637447660
transform 1 0 -10 0 1 86400
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_8
timestamp 1637595202
transform -1 0 717846 0 1 189000
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_9
timestamp 1637595202
transform -1 0 717846 0 1 143800
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_10
timestamp 1637595202
transform -1 0 717846 0 1 98800
box 6032 203748 46226 221470
use gpio_control_power_routing  gpio_control_power_routing_5
timestamp 1637447660
transform 1 0 -10 0 1 216000
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_6
timestamp 1637447660
transform 1 0 -10 0 1 343600
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_6
timestamp 1637595202
transform -1 0 717846 0 1 321200
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_7
timestamp 1637595202
transform -1 0 717846 0 1 277200
box 6032 203748 46226 221470
use gpio_control_power_routing  gpio_control_power_routing_9
timestamp 1637447660
transform 1 0 -10 0 1 473200
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_8
timestamp 1637447660
transform 1 0 -10 0 1 430000
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_7
timestamp 1637447660
transform 1 0 -10 0 1 386800
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_3
timestamp 1637595202
transform -1 0 717846 0 1 456400
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_4
timestamp 1637595202
transform -1 0 717846 0 1 411400
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_5
timestamp 1637595202
transform -1 0 717846 0 1 366200
box 6032 203748 46226 221470
use gpio_control_power_routing  gpio_control_power_routing_12
timestamp 1637447660
transform 1 0 -10 0 1 602800
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_10
timestamp 1637447660
transform 1 0 -10 0 1 516400
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_11
timestamp 1637447660
transform 1 0 -10 0 1 559600
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_2
timestamp 1637595202
transform -1 0 717846 0 1 501600
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_0
timestamp 1637595202
transform -1 0 717836 0 1 682200
box 6032 203748 46226 221470
<< labels >>
flabel metal5 54316 219436 55324 219998 0 FreeSans 1600 0 0 0 vccd1_core
flabel metal5 52692 217826 53700 218388 0 FreeSans 1600 0 0 0 vssd1_core
flabel metal5 184480 230750 189228 233134 0 FreeSans 16000 0 0 0 vccd_core
flabel metal5 184522 234770 189540 236910 0 FreeSans 16000 0 0 0 vssd_core
flabel metal5 182216 238830 190118 240864 0 FreeSans 16000 0 0 0 vccd2_core
flabel metal5 182126 242838 190088 244986 0 FreeSans 16000 0 0 0 vssd2_core
flabel metal5 181918 254572 189876 257076 0 FreeSans 16000 0 0 0 vdda2_core
flabel metal5 181918 258660 189876 261164 0 FreeSans 16000 0 0 0 vssa2_core
flabel metal5 621960 246802 629984 249230 0 FreeSans 16000 0 0 0 vccd1_core
flabel metal5 621948 250708 629990 253036 0 FreeSans 16000 0 0 0 vssd1_core
flabel metal5 621550 262640 629508 265144 0 FreeSans 16000 0 0 0 vdda1_core
flabel metal5 621514 266692 629472 269196 0 FreeSans 16000 0 0 0 vssa1_core
flabel metal5 590480 230750 595228 233134 0 FreeSans 16000 0 0 0 vccd_core
flabel metal5 590522 234770 595540 236910 0 FreeSans 16000 0 0 0 vssd_core
flabel metal5 42966 171382 45564 172780 0 FreeSans 3200 0 0 0 vccd_core
flabel metal5 664092 267180 666518 267904 0 FreeSans 3200 0 0 0 vssa1_core
flabel metal5 667280 263142 669706 263866 0 FreeSans 3200 0 0 0 vdda1_core
flabel metal5 634330 96284 638114 98514 0 FreeSans 16000 0 0 0 vssd_core
flabel metal5 633452 78554 637236 80784 0 FreeSans 16000 0 0 0 vccd_core
flabel metal5 206106 18628 207168 19326 0 FreeSans 4800 0 0 0 vccd_core
flabel metal5 206018 17180 207080 17878 0 FreeSans 4800 0 0 0 vssd_core
flabel metal5 182024 250550 190042 253308 0 FreeSans 16000 0 0 0 vssd1_core
flabel metal5 182160 246638 190178 249396 0 FreeSans 16000 0 0 0 vccd1_core
flabel metal5 181852 266620 189870 269378 0 FreeSans 16000 0 0 0 vssa1_core
flabel metal5 181950 262574 189968 265332 0 FreeSans 16000 0 0 0 vdda1_core
flabel metal5 47904 265444 49660 265998 0 FreeSans 3200 0 0 0 vssa2_core
flabel metal5 50338 265444 52094 265998 0 FreeSans 3200 0 0 0 vdda2_core
flabel metal5 621512 258708 630212 261250 0 FreeSans 16000 0 0 0 vssa2_core
flabel metal5 621598 254668 630298 257210 0 FreeSans 16000 0 0 0 vdda2_core
flabel metal5 621936 242776 630636 245318 0 FreeSans 16000 0 0 0 vssd2_core
flabel metal5 621794 238736 630494 241278 0 FreeSans 16000 0 0 0 vccd2_core
<< end >>
