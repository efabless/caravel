magic
tech sky130A
magscale 1 2
timestamp 1665916077
<< checkpaint >>
rect 4762 32640 713074 1032956
<< metal1 >>
rect 648104 47110 649670 47188
rect 648104 46674 648189 47110
rect 649585 46738 649670 47110
rect 649585 46674 650160 46738
rect 648104 46598 650160 46674
rect 648104 46590 649670 46598
<< via1 >>
rect 648189 46674 649585 47110
<< metal2 >>
rect 648104 47120 649670 47188
rect 648104 46664 648179 47120
rect 649595 46738 649670 47120
rect 649595 46664 650160 46738
rect 648104 46598 650160 46664
rect 648104 46590 649670 46598
<< via2 >>
rect 648179 47110 649595 47120
rect 648179 46674 648189 47110
rect 648189 46674 649585 47110
rect 649585 46674 649595 47110
rect 648179 46664 649595 46674
<< metal3 >>
rect 575700 997047 580479 997678
rect 575700 995143 575814 997047
rect 580358 995143 580479 997047
rect 575700 995032 580479 995143
rect 585678 997053 590458 997678
rect 585678 995149 585784 997053
rect 590328 995149 590458 997053
rect 585678 995032 590458 995149
rect 44198 953072 61996 953124
rect 44198 953015 61461 953072
rect 44198 951991 44314 953015
rect 46698 951991 61461 953015
rect 44198 951968 61461 951991
rect 61925 951968 61996 953072
rect 44198 951924 61996 951968
rect 40984 951480 61032 951524
rect 40984 951433 60497 951480
rect 40984 950409 41104 951433
rect 43488 950409 60497 951433
rect 40984 950376 60497 950409
rect 60961 950376 61032 951480
rect 40984 950324 61032 950376
rect 55372 949682 58218 949982
rect 55372 949629 63922 949682
rect 55372 948782 63379 949629
rect 57038 948525 63379 948782
rect 63843 948525 63922 949629
rect 57038 948482 63922 948525
rect 53768 948182 56610 948382
rect 53768 948121 62944 948182
rect 53768 947182 62411 948121
rect 55432 947017 62411 947182
rect 62875 947017 62944 948121
rect 55432 946982 62944 947017
rect 650616 946337 675364 946382
rect 650616 945233 650656 946337
rect 651200 945233 675364 946337
rect 650616 945182 675364 945233
rect 651580 944733 671668 944782
rect 651580 943629 651614 944733
rect 652158 943629 671668 944733
rect 651580 943582 671668 943629
rect 650616 901137 675830 901182
rect 650616 900033 650656 901137
rect 651200 901105 675830 901137
rect 651200 900081 674765 901105
rect 675709 900081 675830 901105
rect 651200 900033 675830 900081
rect 650616 899982 675830 900033
rect 651580 899533 672676 899582
rect 651580 898429 651614 899533
rect 652158 899497 672676 899533
rect 652158 898473 671569 899497
rect 672593 898473 672676 899497
rect 652158 898429 672676 898473
rect 651580 898382 672676 898429
rect 650616 856137 675264 856182
rect 650616 855033 650656 856137
rect 651200 856096 675264 856137
rect 651200 855072 674136 856096
rect 675160 855072 675264 856096
rect 651200 855033 675264 855072
rect 650616 854982 675264 855033
rect 651580 854533 672708 854582
rect 651580 853429 651614 854533
rect 652158 854494 672708 854533
rect 652158 853470 671592 854494
rect 672616 853470 672708 854494
rect 652158 853429 672708 853470
rect 651580 853382 672708 853429
rect 39852 842294 50002 842458
rect 39852 837830 47929 842294
rect 49673 837830 50002 842294
rect 39852 837678 50002 837830
rect 667172 833190 677818 833301
rect 39852 832362 50002 832479
rect 39852 827898 47929 832362
rect 49673 827898 50002 832362
rect 667172 828646 667316 833190
rect 669700 828646 677818 833190
rect 667172 828521 677818 828646
rect 39852 827699 50002 827898
rect 44198 827272 61996 827324
rect 44198 827215 61461 827272
rect 44198 826191 44314 827215
rect 46698 826191 61461 827215
rect 44198 826168 61461 826191
rect 61925 826168 61996 827272
rect 44198 826124 61996 826168
rect 40984 825680 61032 825724
rect 40984 825633 60497 825680
rect 40984 824609 41104 825633
rect 43488 824609 60497 825633
rect 40984 824576 60497 824609
rect 60961 824576 61032 825680
rect 40984 824524 61032 824576
rect 55372 824129 63922 824182
rect 55372 823025 63379 824129
rect 63843 823025 63922 824129
rect 55372 822982 63922 823025
rect 667172 823196 677818 823322
rect 53768 822521 62944 822582
rect 53768 821417 62411 822521
rect 62875 821417 62944 822521
rect 53768 821382 62944 821417
rect 667172 818652 667302 823196
rect 669686 818652 677818 823196
rect 667172 818542 677818 818652
rect 44198 785672 61996 785724
rect 44198 785615 61461 785672
rect 44198 784591 44314 785615
rect 46698 784591 61461 785615
rect 44198 784568 61461 784591
rect 61925 784568 61996 785672
rect 44198 784524 61996 784568
rect 40984 784080 61032 784124
rect 40984 784033 60497 784080
rect 40984 783009 41104 784033
rect 43488 783009 60497 784033
rect 40984 782976 60497 783009
rect 60961 782976 61032 784080
rect 40984 782924 61032 782976
rect 56078 782129 63922 782182
rect 56078 781025 63379 782129
rect 63843 781025 63922 782129
rect 56078 780982 63922 781025
rect 55372 779782 57370 780982
rect 53768 779321 62944 779382
rect 53768 778217 62411 779321
rect 62875 778217 62944 779321
rect 53768 778182 62944 778217
rect 650616 767937 675364 767982
rect 650616 766833 650656 767937
rect 651200 766833 675364 767937
rect 650616 766782 675364 766833
rect 651580 766333 671668 766382
rect 651580 765229 651614 766333
rect 652158 765229 671668 766333
rect 651580 765182 671668 765229
rect 44198 740872 61996 740924
rect 44198 740815 61461 740872
rect 44198 739791 44314 740815
rect 46698 739791 61461 740815
rect 44198 739768 61461 739791
rect 61925 739768 61996 740872
rect 44198 739724 61996 739768
rect 40984 739280 61032 739324
rect 40984 739233 60497 739280
rect 40984 738209 41104 739233
rect 43488 738209 60497 739233
rect 40984 738176 60497 738209
rect 60961 738176 61032 739280
rect 40984 738124 61032 738176
rect 55372 737729 63922 737782
rect 55372 736625 63379 737729
rect 63843 736625 63922 737729
rect 55372 736582 63922 736625
rect 53768 736121 62944 736182
rect 53768 735017 62411 736121
rect 62875 735017 62944 736121
rect 53768 734982 62944 735017
rect 650616 722937 675364 722982
rect 650616 721833 650656 722937
rect 651200 721833 675364 722937
rect 650616 721782 675364 721833
rect 651580 721333 671668 721382
rect 651580 720229 651614 721333
rect 652158 720229 671668 721333
rect 651580 720182 671668 720229
rect 44198 697672 61996 697724
rect 44198 697615 61461 697672
rect 44198 696591 44314 697615
rect 46698 696591 61461 697615
rect 44198 696568 61461 696591
rect 61925 696568 61996 697672
rect 44198 696524 61996 696568
rect 40984 696080 61032 696124
rect 40984 696033 60497 696080
rect 40984 695009 41104 696033
rect 43488 695009 60497 696033
rect 40984 694976 60497 695009
rect 60961 694976 61032 696080
rect 40984 694924 61032 694976
rect 55372 694529 63922 694582
rect 55372 693425 63379 694529
rect 63843 693425 63922 694529
rect 55372 693382 63922 693425
rect 53768 692921 62944 692982
rect 53768 691817 62411 692921
rect 62875 691817 62944 692921
rect 53768 691782 62944 691817
rect 650616 677737 675364 677782
rect 650616 676633 650656 677737
rect 651200 676633 675364 677737
rect 650616 676582 675364 676633
rect 651580 676133 671668 676182
rect 651580 675029 651614 676133
rect 652158 675029 671668 676133
rect 651580 674982 671668 675029
rect 44198 654472 61996 654524
rect 44198 654415 61461 654472
rect 44198 653391 44314 654415
rect 46698 653391 61461 654415
rect 44198 653368 61461 653391
rect 61925 653368 61996 654472
rect 44198 653324 61996 653368
rect 40984 652880 61032 652924
rect 40984 652833 60497 652880
rect 40984 651809 41104 652833
rect 43488 651809 60497 652833
rect 40984 651776 60497 651809
rect 60961 651776 61032 652880
rect 40984 651724 61032 651776
rect 55372 651329 63922 651382
rect 55372 650225 63379 651329
rect 63843 650225 63922 651329
rect 55372 650182 63922 650225
rect 53768 649721 62944 649782
rect 53768 648617 62411 649721
rect 62875 648617 62944 649721
rect 53768 648582 62944 648617
rect 650616 632737 675364 632782
rect 650616 631633 650656 632737
rect 651200 631633 675364 632737
rect 650616 631582 675364 631633
rect 659310 629982 671668 631182
rect 651580 629933 660600 629982
rect 651580 628829 651614 629933
rect 652158 628829 660600 629933
rect 651580 628782 660600 628829
rect 44198 612332 61996 612384
rect 44198 612275 61461 612332
rect 44198 611251 44314 612275
rect 46698 611251 61461 612275
rect 44198 611228 61461 611251
rect 61925 611228 61996 612332
rect 44198 611184 61996 611228
rect 40984 610740 61032 610784
rect 40984 610693 60497 610740
rect 40984 609669 41104 610693
rect 43488 609669 60497 610693
rect 40984 609636 60497 609669
rect 60961 609636 61032 610740
rect 40984 609584 61032 609636
rect 55372 608129 63922 608182
rect 55372 607025 63379 608129
rect 63843 607025 63922 608129
rect 55372 606982 63922 607025
rect 53768 606521 62944 606582
rect 53768 605417 62411 606521
rect 62875 605417 62944 606521
rect 53768 605382 62944 605417
rect 650616 587537 675364 587582
rect 650616 586433 650656 587537
rect 651200 586433 675364 587537
rect 650616 586382 675364 586433
rect 651580 585933 671668 585982
rect 651580 584829 651614 585933
rect 652158 584829 671668 585933
rect 651580 584782 671668 584829
rect 44198 568072 61996 568124
rect 44198 568015 61461 568072
rect 44198 566991 44314 568015
rect 46698 566991 61461 568015
rect 44198 566968 61461 566991
rect 61925 566968 61996 568072
rect 44198 566924 61996 566968
rect 40984 566480 61032 566524
rect 40984 566433 60497 566480
rect 40984 565409 41104 566433
rect 43488 565409 60497 566433
rect 40984 565376 60497 565409
rect 60961 565376 61032 566480
rect 40984 565324 61032 565376
rect 55372 564929 63922 564982
rect 55372 563825 63379 564929
rect 63843 563825 63922 564929
rect 55372 563782 63922 563825
rect 53768 563321 62944 563382
rect 53768 562217 62411 563321
rect 62875 562217 62944 563321
rect 53768 562182 62944 562217
rect 650616 542537 675364 542582
rect 650616 541433 650656 542537
rect 651200 541433 675364 542537
rect 650616 541382 675364 541433
rect 651580 540933 671668 540982
rect 651580 539829 651614 540933
rect 652158 539829 671668 540933
rect 651580 539782 671668 539829
rect 667062 518551 677700 518701
rect 667062 514087 667369 518551
rect 669673 514087 677700 518551
rect 667062 513921 677700 514087
rect 667062 508561 677700 508722
rect 667062 504097 667383 508561
rect 669687 504097 677700 508561
rect 667062 503942 677700 504097
rect 650616 499137 659758 499182
rect 650616 498033 650656 499137
rect 651200 498582 659758 499137
rect 651200 498033 675364 498582
rect 650616 497982 675364 498033
rect 39924 497723 52292 497858
rect 39924 493259 50396 497723
rect 52060 493259 52292 497723
rect 658568 497382 675364 497982
rect 651580 496933 671668 496982
rect 651580 495829 651614 496933
rect 652158 495829 671668 496933
rect 651580 495782 671668 495829
rect 39924 493078 52292 493259
rect 39924 487733 52292 487879
rect 39924 483269 50384 487733
rect 52048 483269 52292 487733
rect 39924 483099 52292 483269
rect 44198 440472 61996 440524
rect 44198 440415 61461 440472
rect 44198 439391 44314 440415
rect 46698 439391 61461 440415
rect 44198 439368 61461 439391
rect 61925 439368 61996 440472
rect 44198 439324 61996 439368
rect 40984 438880 61032 438924
rect 40984 438833 60497 438880
rect 40984 437809 41104 438833
rect 43488 437809 60497 438833
rect 40984 437776 60497 437809
rect 60961 437776 61032 438880
rect 40984 437724 61032 437776
rect 55372 437329 63922 437382
rect 55372 436225 63379 437329
rect 63843 436225 63922 437329
rect 55372 436182 63922 436225
rect 53768 435721 62944 435782
rect 53768 434617 62411 435721
rect 62875 434617 62944 435721
rect 53768 434582 62944 434617
rect 663914 430389 677712 430501
rect 663914 425685 664145 430389
rect 666529 425748 677712 430389
rect 666529 425685 667110 425748
rect 663914 425562 667110 425685
rect 663914 420431 677712 420522
rect 663914 415887 664128 420431
rect 666512 415887 677712 420431
rect 663914 415742 677712 415887
rect 650616 410337 675364 410382
rect 650616 409233 650656 410337
rect 651200 409233 675364 410337
rect 650616 409182 675364 409233
rect 651580 408733 671668 408782
rect 651580 407629 651614 408733
rect 652158 407629 671668 408733
rect 651580 407582 671668 407629
rect 44198 397272 61996 397324
rect 44198 397215 61461 397272
rect 44198 396191 44314 397215
rect 46698 396191 61461 397215
rect 44198 396168 61461 396191
rect 61925 396168 61996 397272
rect 44198 396124 61996 396168
rect 40984 395680 61032 395724
rect 40984 395633 60497 395680
rect 40984 394609 41104 395633
rect 43488 394609 60497 395633
rect 40984 394576 60497 394609
rect 60961 394576 61032 395680
rect 40984 394524 61032 394576
rect 55372 394129 63922 394182
rect 55372 393025 63379 394129
rect 63843 393025 63922 394129
rect 55372 392982 63922 393025
rect 53768 392521 62944 392582
rect 53768 391417 62411 392521
rect 62875 391417 62944 392521
rect 53768 391382 62944 391417
rect 650616 366537 665664 366582
rect 650616 365433 650656 366537
rect 651200 365433 665664 366537
rect 650616 365382 665664 365433
rect 664464 365182 665664 365382
rect 664464 363982 675364 365182
rect 651580 363533 671668 363582
rect 651580 362429 651614 363533
rect 652158 362429 671668 363533
rect 651580 362382 671668 362429
rect 44198 355072 61996 355124
rect 44198 355015 61461 355072
rect 44198 353991 44314 355015
rect 46698 353991 61461 355015
rect 44198 353968 61461 353991
rect 61925 353968 61996 355072
rect 44198 353924 61996 353968
rect 40984 353480 61032 353524
rect 40984 353433 60497 353480
rect 40984 352409 41104 353433
rect 43488 352409 60497 353433
rect 40984 352376 60497 352409
rect 60961 352376 61032 353480
rect 40984 352324 61032 352376
rect 55968 351729 63922 351782
rect 55968 350982 63379 351729
rect 55372 350625 63379 350982
rect 63843 350625 63922 351729
rect 55372 350582 63922 350625
rect 55372 349782 57264 350582
rect 53768 349321 62944 349382
rect 53768 348217 62411 349321
rect 62875 348217 62944 349321
rect 53768 348182 62944 348217
rect 650616 320137 676922 320182
rect 650616 319033 650656 320137
rect 651200 319033 676922 320137
rect 650616 318982 676922 319033
rect 651580 318533 673726 318582
rect 651580 317429 651614 318533
rect 652158 317429 673726 318533
rect 651580 317382 673726 317429
rect 44198 310872 61996 310924
rect 44198 310815 61461 310872
rect 44198 309791 44314 310815
rect 46698 309791 61461 310815
rect 44198 309768 61461 309791
rect 61925 309768 61996 310872
rect 44198 309724 61996 309768
rect 40984 309280 61032 309324
rect 40984 309233 60497 309280
rect 40984 308209 41104 309233
rect 43488 308209 60497 309233
rect 40984 308176 60497 308209
rect 60961 308176 61032 309280
rect 40984 308124 61032 308176
rect 55432 307729 63922 307782
rect 55432 306625 63379 307729
rect 63843 306625 63922 307729
rect 55432 306582 63922 306625
rect 53790 306121 62944 306182
rect 53790 305017 62411 306121
rect 62875 305017 62944 306121
rect 53790 304982 62944 305017
rect 39456 82706 45844 82744
rect 39456 78242 41977 82706
rect 45641 78242 45844 82706
rect 39456 78151 45844 78242
rect 39456 72802 45844 72900
rect 39456 68338 41953 72802
rect 45617 68338 45844 72802
rect 39456 68256 45844 68338
rect 648104 47124 649670 47188
rect 241690 46601 246049 46686
rect 241690 42857 241751 46601
rect 245975 42857 246049 46601
rect 149600 41140 150458 41207
rect 149600 40996 149637 41140
rect 150421 40996 150458 41140
rect 148068 40744 148926 40782
rect 148068 40600 148105 40744
rect 148889 40600 148926 40744
rect 148068 34765 148926 40600
rect 149600 35973 150458 40996
rect 241690 39426 246049 42857
rect 251300 46615 255702 46686
rect 251300 42871 251403 46615
rect 255627 42871 255702 46615
rect 648104 46660 648175 47124
rect 649599 46844 649670 47124
rect 649599 46660 650158 46844
rect 648104 46598 650158 46660
rect 648104 46590 649670 46598
rect 653462 45022 656910 45156
rect 251300 39426 255702 42871
rect 641954 43965 643694 44026
rect 641954 42221 641995 43965
rect 643659 42221 643694 43965
rect 149600 35189 149642 35973
rect 150426 35189 150458 35973
rect 149600 35114 150458 35189
rect 148068 33981 148108 34765
rect 148892 33981 148926 34765
rect 148068 33900 148926 33981
rect 641954 34726 643694 42221
rect 653462 42638 653583 45022
rect 656767 42638 656910 45022
rect 653462 35808 656910 42638
rect 641954 34022 642038 34726
rect 643622 34022 643694 34726
rect 641954 33920 643694 34022
<< via3 >>
rect 575814 995143 580358 997047
rect 585784 995149 590328 997053
rect 44314 951991 46698 953015
rect 61461 951968 61925 953072
rect 41104 950409 43488 951433
rect 60497 950376 60961 951480
rect 63379 948525 63843 949629
rect 62411 947017 62875 948121
rect 650656 945233 651200 946337
rect 651614 943629 652158 944733
rect 650656 900033 651200 901137
rect 674765 900081 675709 901105
rect 651614 898429 652158 899533
rect 671569 898473 672593 899497
rect 650656 855033 651200 856137
rect 674136 855072 675160 856096
rect 651614 853429 652158 854533
rect 671592 853470 672616 854494
rect 47929 837830 49673 842294
rect 47929 827898 49673 832362
rect 667316 828646 669700 833190
rect 44314 826191 46698 827215
rect 61461 826168 61925 827272
rect 41104 824609 43488 825633
rect 60497 824576 60961 825680
rect 63379 823025 63843 824129
rect 62411 821417 62875 822521
rect 667302 818652 669686 823196
rect 44314 784591 46698 785615
rect 61461 784568 61925 785672
rect 41104 783009 43488 784033
rect 60497 782976 60961 784080
rect 63379 781025 63843 782129
rect 62411 778217 62875 779321
rect 650656 766833 651200 767937
rect 651614 765229 652158 766333
rect 44314 739791 46698 740815
rect 61461 739768 61925 740872
rect 41104 738209 43488 739233
rect 60497 738176 60961 739280
rect 63379 736625 63843 737729
rect 62411 735017 62875 736121
rect 650656 721833 651200 722937
rect 651614 720229 652158 721333
rect 44314 696591 46698 697615
rect 61461 696568 61925 697672
rect 41104 695009 43488 696033
rect 60497 694976 60961 696080
rect 63379 693425 63843 694529
rect 62411 691817 62875 692921
rect 650656 676633 651200 677737
rect 651614 675029 652158 676133
rect 44314 653391 46698 654415
rect 61461 653368 61925 654472
rect 41104 651809 43488 652833
rect 60497 651776 60961 652880
rect 63379 650225 63843 651329
rect 62411 648617 62875 649721
rect 650656 631633 651200 632737
rect 651614 628829 652158 629933
rect 44314 611251 46698 612275
rect 61461 611228 61925 612332
rect 41104 609669 43488 610693
rect 60497 609636 60961 610740
rect 63379 607025 63843 608129
rect 62411 605417 62875 606521
rect 650656 586433 651200 587537
rect 651614 584829 652158 585933
rect 44314 566991 46698 568015
rect 61461 566968 61925 568072
rect 41104 565409 43488 566433
rect 60497 565376 60961 566480
rect 63379 563825 63843 564929
rect 62411 562217 62875 563321
rect 650656 541433 651200 542537
rect 651614 539829 652158 540933
rect 667369 514087 669673 518551
rect 667383 504097 669687 508561
rect 650656 498033 651200 499137
rect 50396 493259 52060 497723
rect 651614 495829 652158 496933
rect 50384 483269 52048 487733
rect 44314 439391 46698 440415
rect 61461 439368 61925 440472
rect 41104 437809 43488 438833
rect 60497 437776 60961 438880
rect 63379 436225 63843 437329
rect 62411 434617 62875 435721
rect 664145 425685 666529 430389
rect 664128 415887 666512 420431
rect 650656 409233 651200 410337
rect 651614 407629 652158 408733
rect 44314 396191 46698 397215
rect 61461 396168 61925 397272
rect 41104 394609 43488 395633
rect 60497 394576 60961 395680
rect 63379 393025 63843 394129
rect 62411 391417 62875 392521
rect 650656 365433 651200 366537
rect 651614 362429 652158 363533
rect 44314 353991 46698 355015
rect 61461 353968 61925 355072
rect 41104 352409 43488 353433
rect 60497 352376 60961 353480
rect 63379 350625 63843 351729
rect 62411 348217 62875 349321
rect 650656 319033 651200 320137
rect 651614 317429 652158 318533
rect 44314 309791 46698 310815
rect 61461 309768 61925 310872
rect 41104 308209 43488 309233
rect 60497 308176 60961 309280
rect 63379 306625 63843 307729
rect 62411 305017 62875 306121
rect 41977 78242 45641 82706
rect 41953 68338 45617 72802
rect 241751 42857 245975 46601
rect 149637 40996 150421 41140
rect 148105 40600 148889 40744
rect 251403 42871 255627 46615
rect 648175 47120 649599 47124
rect 648175 46664 648179 47120
rect 648179 46664 649595 47120
rect 649595 46664 649599 47120
rect 648175 46660 649599 46664
rect 641995 42221 643659 43965
rect 149642 35189 150426 35973
rect 148108 33981 148892 34765
rect 653583 42638 656767 45022
rect 642038 34022 643622 34726
<< metal4 >>
rect 575680 997047 580478 997130
rect 575680 995143 575814 997047
rect 580358 995143 580478 997047
rect 575680 993177 580478 995143
rect 575680 991021 575875 993177
rect 580271 991021 580478 993177
rect 575680 990788 580478 991021
rect 585670 997053 590468 997144
rect 585670 995149 585784 997053
rect 590328 995149 590468 997053
rect 670816 996692 673426 996696
rect 670808 996544 676654 996692
rect 670808 995668 671036 996544
rect 676392 995668 676654 996544
rect 670808 995492 676654 995668
rect 585670 993191 590468 995149
rect 585670 991035 585871 993191
rect 590267 991035 590468 993191
rect 585670 990802 590468 991035
rect 670816 992520 673426 995492
rect 670816 990364 671042 992520
rect 673198 990364 673426 992520
rect 47796 990126 56582 990310
rect 670816 990200 673426 990364
rect 47796 990125 55829 990126
rect 47796 989889 47874 990125
rect 48110 989889 48194 990125
rect 48430 989889 48514 990125
rect 48750 989889 48834 990125
rect 49070 989889 49154 990125
rect 49390 989889 49474 990125
rect 49710 989890 55829 990125
rect 56065 989890 56149 990126
rect 56385 989890 56582 990126
rect 49710 989889 56582 989890
rect 47796 989692 56582 989889
rect 50194 989166 56434 989348
rect 50194 989161 55833 989166
rect 50194 988925 50280 989161
rect 50516 988925 50600 989161
rect 50836 988925 50920 989161
rect 51156 988925 51240 989161
rect 51476 988925 51560 989161
rect 51796 988925 51880 989161
rect 52116 988930 55833 989161
rect 56069 988930 56153 989166
rect 56389 988930 56434 989166
rect 52116 988925 56434 988930
rect 50194 988736 56434 988925
rect 658380 987247 669826 987436
rect 658380 987242 667281 987247
rect 658380 987006 658577 987242
rect 658813 987006 658897 987242
rect 659133 987006 659217 987242
rect 659453 987006 659537 987242
rect 659773 987006 659857 987242
rect 660093 987006 660177 987242
rect 660413 987006 660497 987242
rect 660733 987006 660817 987242
rect 661053 987006 661137 987242
rect 661373 987006 661457 987242
rect 661693 987006 661777 987242
rect 662013 987006 662097 987242
rect 662333 987006 662417 987242
rect 662653 987006 662737 987242
rect 662973 987011 667281 987242
rect 667517 987011 667601 987247
rect 667837 987011 667921 987247
rect 668157 987011 668241 987247
rect 668477 987011 668561 987247
rect 668797 987011 668881 987247
rect 669117 987011 669201 987247
rect 669437 987011 669521 987247
rect 669757 987011 669826 987247
rect 662973 987006 669826 987011
rect 658380 986812 669826 987006
rect 40993 986441 56414 986468
rect 40993 985885 41066 986441
rect 43542 986279 56414 986441
rect 43542 986043 55813 986279
rect 56049 986043 56133 986279
rect 56369 986043 56414 986279
rect 43542 985885 56414 986043
rect 40993 985854 56414 985885
rect 44200 985486 56440 985526
rect 44200 984930 44269 985486
rect 46745 985475 56440 985486
rect 46745 984930 55828 985475
rect 44200 984919 55828 984930
rect 56384 984919 56440 985475
rect 44200 984874 56440 984919
rect 52596 984517 56404 984548
rect 52596 984357 55811 984517
rect 52596 984121 52759 984357
rect 52995 984121 53079 984357
rect 53315 984121 53399 984357
rect 53635 984121 55811 984357
rect 52596 983961 55811 984121
rect 56367 983961 56404 984517
rect 52596 983928 56404 983961
rect 658316 984521 673430 984570
rect 658316 984356 670883 984521
rect 658316 984120 658391 984356
rect 658627 984120 658711 984356
rect 658947 984120 659031 984356
rect 659267 984120 659351 984356
rect 659587 984120 659671 984356
rect 659907 984120 659991 984356
rect 660227 984120 660311 984356
rect 660547 984120 660631 984356
rect 660867 984120 660951 984356
rect 661187 984120 661271 984356
rect 661507 984120 661591 984356
rect 661827 984120 661911 984356
rect 662147 984120 662231 984356
rect 662467 984120 662551 984356
rect 662787 984120 662871 984356
rect 663107 984120 670883 984356
rect 658316 983965 670883 984120
rect 673359 983965 673430 984521
rect 658316 983928 673430 983965
rect 658288 983559 676624 983602
rect 658288 983400 674081 983559
rect 658288 983164 658373 983400
rect 658609 983164 658693 983400
rect 658929 983164 659013 983400
rect 659249 983164 659333 983400
rect 659569 983164 659653 983400
rect 659889 983164 659973 983400
rect 660209 983164 660293 983400
rect 660529 983164 660613 983400
rect 660849 983164 660933 983400
rect 661169 983164 661253 983400
rect 661489 983164 661573 983400
rect 661809 983164 661893 983400
rect 662129 983164 662213 983400
rect 662449 983164 662533 983400
rect 662769 983164 662853 983400
rect 663089 983164 674081 983400
rect 658288 983003 674081 983164
rect 676557 983003 676624 983559
rect 658288 982960 676624 983003
rect 44200 953015 46792 953126
rect 44200 951991 44314 953015
rect 46698 951991 46792 953015
rect 44200 951922 46792 951991
rect 61424 953072 61962 953080
rect 61424 951968 61461 953072
rect 61925 951968 61962 953072
rect 61424 951960 61962 951968
rect 40994 951433 43588 951522
rect 40994 950409 41104 951433
rect 43488 950409 43588 951433
rect 40994 950326 43588 950409
rect 60460 951480 60998 951488
rect 60460 950376 60497 951480
rect 60961 950376 60998 951480
rect 60460 950368 60998 950376
rect 63350 949629 63872 949632
rect 63350 948525 63379 949629
rect 63843 948525 63872 949629
rect 63350 948522 63872 948525
rect 62382 948121 62904 948124
rect 62382 947017 62411 948121
rect 62875 947017 62904 948121
rect 62382 947014 62904 947017
rect 650654 946337 651202 946346
rect 650654 945233 650656 946337
rect 651200 945233 651202 946337
rect 650654 945224 651202 945233
rect 651602 944733 652170 944750
rect 651602 943629 651614 944733
rect 652158 943629 652170 944733
rect 651602 943612 652170 943629
rect 650654 901137 651202 901146
rect 650654 900033 650656 901137
rect 651200 900033 651202 901137
rect 650654 900024 651202 900033
rect 674630 901105 675830 901182
rect 674630 900081 674765 901105
rect 675709 900081 675830 901105
rect 674630 899982 675830 900081
rect 651602 899533 652170 899550
rect 651602 898429 651614 899533
rect 652158 898429 652170 899533
rect 651602 898412 652170 898429
rect 671476 899497 672676 899582
rect 671476 898473 671569 899497
rect 672593 898473 672676 899497
rect 671476 898382 672676 898473
rect 650654 856137 651202 856146
rect 650654 855033 650656 856137
rect 651200 855033 651202 856137
rect 650654 855024 651202 855033
rect 674054 856096 675254 856182
rect 674054 855072 674136 856096
rect 675160 855072 675254 856096
rect 674054 854982 675254 855072
rect 651602 854533 652170 854550
rect 651602 853429 651614 854533
rect 652158 853429 652170 854533
rect 651602 853412 652170 853429
rect 671508 854494 672708 854582
rect 671508 853470 671592 854494
rect 672616 853470 672708 854494
rect 671508 853382 672708 853470
rect 47792 842294 49822 842462
rect 47792 837830 47929 842294
rect 49673 837830 49822 842294
rect 47792 837658 49822 837830
rect 667202 833190 669802 833310
rect 47792 832362 49822 832506
rect 47792 827898 47929 832362
rect 49673 827898 49822 832362
rect 667202 828646 667316 833190
rect 669700 828646 669802 833190
rect 667202 828520 669802 828646
rect 47792 827702 49822 827898
rect 44200 827215 46792 827326
rect 44200 826191 44314 827215
rect 46698 826191 46792 827215
rect 44200 826122 46792 826191
rect 61424 827272 61962 827280
rect 61424 826168 61461 827272
rect 61925 826168 61962 827272
rect 61424 826160 61962 826168
rect 40994 825633 43588 825722
rect 40994 824609 41104 825633
rect 43488 824609 43588 825633
rect 40994 824526 43588 824609
rect 60460 825680 60998 825688
rect 60460 824576 60497 825680
rect 60961 824576 60998 825680
rect 60460 824568 60998 824576
rect 63350 824129 63872 824132
rect 63350 823025 63379 824129
rect 63843 823025 63872 824129
rect 63350 823022 63872 823025
rect 667214 823196 669814 823336
rect 62382 822521 62904 822524
rect 62382 821417 62411 822521
rect 62875 821417 62904 822521
rect 62382 821414 62904 821417
rect 667214 818652 667302 823196
rect 669686 818652 669814 823196
rect 667214 818546 669814 818652
rect 44200 785615 46792 785726
rect 44200 784591 44314 785615
rect 46698 784591 46792 785615
rect 44200 784522 46792 784591
rect 61424 785672 61962 785680
rect 61424 784568 61461 785672
rect 61925 784568 61962 785672
rect 61424 784560 61962 784568
rect 40994 784033 43588 784122
rect 40994 783009 41104 784033
rect 43488 783009 43588 784033
rect 40994 782926 43588 783009
rect 60460 784080 60998 784088
rect 60460 782976 60497 784080
rect 60961 782976 60998 784080
rect 60460 782968 60998 782976
rect 63350 782129 63872 782132
rect 63350 781025 63379 782129
rect 63843 781025 63872 782129
rect 63350 781022 63872 781025
rect 62382 779321 62904 779324
rect 62382 778217 62411 779321
rect 62875 778217 62904 779321
rect 62382 778214 62904 778217
rect 650654 767937 651202 767946
rect 650654 766833 650656 767937
rect 651200 766833 651202 767937
rect 650654 766824 651202 766833
rect 651602 766333 652170 766350
rect 651602 765229 651614 766333
rect 652158 765229 652170 766333
rect 651602 765212 652170 765229
rect 44200 740815 46792 740926
rect 44200 739791 44314 740815
rect 46698 739791 46792 740815
rect 44200 739722 46792 739791
rect 61424 740872 61962 740880
rect 61424 739768 61461 740872
rect 61925 739768 61962 740872
rect 61424 739760 61962 739768
rect 40994 739233 43588 739322
rect 40994 738209 41104 739233
rect 43488 738209 43588 739233
rect 40994 738126 43588 738209
rect 60460 739280 60998 739288
rect 60460 738176 60497 739280
rect 60961 738176 60998 739280
rect 60460 738168 60998 738176
rect 63350 737729 63872 737732
rect 63350 736625 63379 737729
rect 63843 736625 63872 737729
rect 63350 736622 63872 736625
rect 62382 736121 62904 736124
rect 62382 735017 62411 736121
rect 62875 735017 62904 736121
rect 62382 735014 62904 735017
rect 650654 722937 651202 722946
rect 650654 721833 650656 722937
rect 651200 721833 651202 722937
rect 650654 721824 651202 721833
rect 651602 721333 652170 721350
rect 651602 720229 651614 721333
rect 652158 720229 652170 721333
rect 651602 720212 652170 720229
rect 44200 697615 46792 697726
rect 44200 696591 44314 697615
rect 46698 696591 46792 697615
rect 44200 696522 46792 696591
rect 61424 697672 61962 697680
rect 61424 696568 61461 697672
rect 61925 696568 61962 697672
rect 61424 696560 61962 696568
rect 40994 696033 43588 696122
rect 40994 695009 41104 696033
rect 43488 695009 43588 696033
rect 40994 694926 43588 695009
rect 60460 696080 60998 696088
rect 60460 694976 60497 696080
rect 60961 694976 60998 696080
rect 60460 694968 60998 694976
rect 63350 694529 63872 694532
rect 63350 693425 63379 694529
rect 63843 693425 63872 694529
rect 63350 693422 63872 693425
rect 62382 692921 62904 692924
rect 62382 691817 62411 692921
rect 62875 691817 62904 692921
rect 62382 691814 62904 691817
rect 650654 677737 651202 677746
rect 650654 676633 650656 677737
rect 651200 676633 651202 677737
rect 650654 676624 651202 676633
rect 651602 676133 652170 676150
rect 651602 675029 651614 676133
rect 652158 675029 652170 676133
rect 651602 675012 652170 675029
rect 44200 654415 46792 654526
rect 44200 653391 44314 654415
rect 46698 653391 46792 654415
rect 44200 653322 46792 653391
rect 61424 654472 61962 654480
rect 61424 653368 61461 654472
rect 61925 653368 61962 654472
rect 61424 653360 61962 653368
rect 40994 652833 43588 652922
rect 40994 651809 41104 652833
rect 43488 651809 43588 652833
rect 40994 651726 43588 651809
rect 60460 652880 60998 652888
rect 60460 651776 60497 652880
rect 60961 651776 60998 652880
rect 60460 651768 60998 651776
rect 63350 651329 63872 651332
rect 63350 650225 63379 651329
rect 63843 650225 63872 651329
rect 63350 650222 63872 650225
rect 62382 649721 62904 649724
rect 62382 648617 62411 649721
rect 62875 648617 62904 649721
rect 62382 648614 62904 648617
rect 650654 632737 651202 632746
rect 650654 631633 650656 632737
rect 651200 631633 651202 632737
rect 650654 631624 651202 631633
rect 651602 629933 652170 629950
rect 651602 628829 651614 629933
rect 652158 628829 652170 629933
rect 651602 628812 652170 628829
rect 44200 612275 46792 612386
rect 44200 611251 44314 612275
rect 46698 611251 46792 612275
rect 44200 611182 46792 611251
rect 61424 612332 61962 612340
rect 61424 611228 61461 612332
rect 61925 611228 61962 612332
rect 61424 611220 61962 611228
rect 40994 610693 43588 610782
rect 40994 609669 41104 610693
rect 43488 609669 43588 610693
rect 40994 609586 43588 609669
rect 60460 610740 60998 610748
rect 60460 609636 60497 610740
rect 60961 609636 60998 610740
rect 60460 609628 60998 609636
rect 63350 608129 63872 608132
rect 63350 607025 63379 608129
rect 63843 607025 63872 608129
rect 63350 607022 63872 607025
rect 62382 606521 62904 606524
rect 62382 605417 62411 606521
rect 62875 605417 62904 606521
rect 62382 605414 62904 605417
rect 650654 587537 651202 587546
rect 650654 586433 650656 587537
rect 651200 586433 651202 587537
rect 650654 586424 651202 586433
rect 651602 585933 652170 585950
rect 651602 584829 651614 585933
rect 652158 584829 652170 585933
rect 651602 584812 652170 584829
rect 44200 568015 46792 568126
rect 44200 566991 44314 568015
rect 46698 566991 46792 568015
rect 44200 566922 46792 566991
rect 61424 568072 61962 568080
rect 61424 566968 61461 568072
rect 61925 566968 61962 568072
rect 61424 566960 61962 566968
rect 40994 566433 43588 566522
rect 40994 565409 41104 566433
rect 43488 565409 43588 566433
rect 40994 565326 43588 565409
rect 60460 566480 60998 566488
rect 60460 565376 60497 566480
rect 60961 565376 60998 566480
rect 60460 565368 60998 565376
rect 63350 564929 63872 564932
rect 63350 563825 63379 564929
rect 63843 563825 63872 564929
rect 63350 563822 63872 563825
rect 62382 563321 62904 563324
rect 62382 562217 62411 563321
rect 62875 562217 62904 563321
rect 62382 562214 62904 562217
rect 650654 542537 651202 542546
rect 650654 541433 650656 542537
rect 651200 541433 651202 542537
rect 650654 541424 651202 541433
rect 651602 540933 652170 540950
rect 651602 539829 651614 540933
rect 652158 539829 652170 540933
rect 651602 539812 652170 539829
rect 667206 518551 669814 518696
rect 667206 514087 667369 518551
rect 669673 514087 669814 518551
rect 667206 513920 669814 514087
rect 667218 508561 669826 508726
rect 667218 504097 667383 508561
rect 669687 504097 669826 508561
rect 667218 503950 669826 504097
rect 650654 499137 651202 499146
rect 650654 498033 650656 499137
rect 651200 498033 651202 499137
rect 650654 498024 651202 498033
rect 50172 497723 52196 497874
rect 50172 493259 50396 497723
rect 52060 493259 52196 497723
rect 651602 496933 652170 496950
rect 651602 495829 651614 496933
rect 652158 495829 652170 496933
rect 651602 495812 652170 495829
rect 50172 493084 52196 493259
rect 50198 487733 52222 487884
rect 50198 483269 50384 487733
rect 52048 483269 52222 487733
rect 50198 483094 52222 483269
rect 44200 440415 46792 440526
rect 44200 439391 44314 440415
rect 46698 439391 46792 440415
rect 44200 439322 46792 439391
rect 61424 440472 61962 440480
rect 61424 439368 61461 440472
rect 61925 439368 61962 440472
rect 61424 439360 61962 439368
rect 40994 438833 43588 438922
rect 40994 437809 41104 438833
rect 43488 437809 43588 438833
rect 40994 437726 43588 437809
rect 60460 438880 60998 438888
rect 60460 437776 60497 438880
rect 60961 437776 60998 438880
rect 60460 437768 60998 437776
rect 63350 437329 63872 437332
rect 63350 436225 63379 437329
rect 63843 436225 63872 437329
rect 63350 436222 63872 436225
rect 62382 435721 62904 435724
rect 62382 434617 62411 435721
rect 62875 434617 62904 435721
rect 62382 434614 62904 434617
rect 664008 430389 666612 430490
rect 664008 425685 664145 430389
rect 666529 425685 666612 430389
rect 664008 425572 666612 425685
rect 664018 420431 666634 420524
rect 664018 415887 664128 420431
rect 666512 415887 666634 420431
rect 664018 415760 666634 415887
rect 650654 410337 651202 410346
rect 650654 409233 650656 410337
rect 651200 409233 651202 410337
rect 650654 409224 651202 409233
rect 651602 408733 652170 408750
rect 651602 407629 651614 408733
rect 652158 407629 652170 408733
rect 651602 407612 652170 407629
rect 44200 397215 46792 397326
rect 44200 396191 44314 397215
rect 46698 396191 46792 397215
rect 44200 396122 46792 396191
rect 61424 397272 61962 397280
rect 61424 396168 61461 397272
rect 61925 396168 61962 397272
rect 61424 396160 61962 396168
rect 40994 395633 43588 395722
rect 40994 394609 41104 395633
rect 43488 394609 43588 395633
rect 40994 394526 43588 394609
rect 60460 395680 60998 395688
rect 60460 394576 60497 395680
rect 60961 394576 60998 395680
rect 60460 394568 60998 394576
rect 63350 394129 63872 394132
rect 63350 393025 63379 394129
rect 63843 393025 63872 394129
rect 63350 393022 63872 393025
rect 62382 392521 62904 392524
rect 62382 391417 62411 392521
rect 62875 391417 62904 392521
rect 62382 391414 62904 391417
rect 650654 366537 651202 366546
rect 650654 365433 650656 366537
rect 651200 365433 651202 366537
rect 650654 365424 651202 365433
rect 651602 363533 652170 363550
rect 651602 362429 651614 363533
rect 652158 362429 652170 363533
rect 651602 362412 652170 362429
rect 44200 355015 46792 355126
rect 44200 353991 44314 355015
rect 46698 353991 46792 355015
rect 44200 353922 46792 353991
rect 61424 355072 61962 355080
rect 61424 353968 61461 355072
rect 61925 353968 61962 355072
rect 61424 353960 61962 353968
rect 40994 353433 43588 353522
rect 40994 352409 41104 353433
rect 43488 352409 43588 353433
rect 40994 352326 43588 352409
rect 60460 353480 60998 353488
rect 60460 352376 60497 353480
rect 60961 352376 60998 353480
rect 60460 352368 60998 352376
rect 63350 351729 63872 351732
rect 63350 350625 63379 351729
rect 63843 350625 63872 351729
rect 63350 350622 63872 350625
rect 62382 349321 62904 349324
rect 62382 348217 62411 349321
rect 62875 348217 62904 349321
rect 62382 348214 62904 348217
rect 650654 320137 651202 320146
rect 650654 319033 650656 320137
rect 651200 319033 651202 320137
rect 650654 319024 651202 319033
rect 651602 318533 652170 318550
rect 651602 317429 651614 318533
rect 652158 317429 652170 318533
rect 651602 317412 652170 317429
rect 44200 310815 46792 310926
rect 44200 309791 44314 310815
rect 46698 309791 46792 310815
rect 44200 309722 46792 309791
rect 61424 310872 61962 310880
rect 61424 309768 61461 310872
rect 61925 309768 61962 310872
rect 61424 309760 61962 309768
rect 40994 309233 43588 309322
rect 40994 308209 41104 309233
rect 43488 308209 43588 309233
rect 40994 308126 43588 308209
rect 60460 309280 60998 309288
rect 60460 308176 60497 309280
rect 60961 308176 60998 309280
rect 60460 308168 60998 308176
rect 63350 307729 63872 307732
rect 63350 306625 63379 307729
rect 63843 306625 63872 307729
rect 63350 306622 63872 306625
rect 62382 306121 62904 306124
rect 62382 305017 62411 306121
rect 62875 305017 62904 306121
rect 62382 305014 62904 305017
rect 658882 278346 676628 278406
rect 658882 278211 674086 278346
rect 52582 277886 53800 278046
rect 44195 277173 46802 277284
rect 44195 275977 44257 277173
rect 46733 276484 46802 277173
rect 52582 277010 52753 277886
rect 53629 277446 53800 277886
rect 658882 277975 658984 278211
rect 659220 277975 659304 278211
rect 659540 277975 659624 278211
rect 659860 277975 659944 278211
rect 660180 277975 660264 278211
rect 660500 277975 660584 278211
rect 660820 277975 660904 278211
rect 661140 277975 661224 278211
rect 661460 277975 661544 278211
rect 661780 277975 661864 278211
rect 662100 277975 662184 278211
rect 662420 277975 662504 278211
rect 662740 277975 662824 278211
rect 663060 277975 674086 278211
rect 53629 277415 56416 277446
rect 53629 277010 55806 277415
rect 52582 276859 55806 277010
rect 56362 276859 56416 277415
rect 52582 276822 56416 276859
rect 46733 276288 56432 276484
rect 46733 276052 55816 276288
rect 56052 276052 56136 276288
rect 56372 276052 56432 276288
rect 46733 275977 56432 276052
rect 44195 275858 56432 275977
rect 42746 275416 56448 275532
rect 42746 269420 42901 275416
rect 43457 275334 56448 275416
rect 43457 275098 55824 275334
rect 56060 275098 56144 275334
rect 56380 275098 56448 275334
rect 43457 274906 56448 275098
rect 43457 269420 43610 274906
rect 50186 273332 52198 273438
rect 50186 272136 50273 273332
rect 52109 272638 52198 273332
rect 52109 272613 56406 272638
rect 52109 272136 55802 272613
rect 50186 272057 55802 272136
rect 56358 272057 56406 272613
rect 50186 272026 56406 272057
rect 47792 271650 56616 271688
rect 47792 271579 55856 271650
rect 47792 270383 47879 271579
rect 49715 271094 55856 271579
rect 56412 271094 56616 271650
rect 49715 271082 56616 271094
rect 49715 271058 57202 271082
rect 49715 270383 49802 271058
rect 47792 270258 49802 270383
rect 42746 269278 43610 269420
rect 56572 261466 57202 271058
rect 57542 264698 58162 272042
rect 58502 269364 59122 272992
rect 58502 269128 58689 269364
rect 58925 269128 59122 269364
rect 58502 269044 59122 269128
rect 58502 268808 58689 269044
rect 58925 268808 59122 269044
rect 58502 268724 59122 268808
rect 58502 268488 58689 268724
rect 58925 268488 59122 268724
rect 58502 268404 59122 268488
rect 58502 268168 58689 268404
rect 58925 268168 59122 268404
rect 58502 268084 59122 268168
rect 58502 267848 58689 268084
rect 58925 267848 59122 268084
rect 58502 267764 59122 267848
rect 58502 267528 58689 267764
rect 58925 267528 59122 267764
rect 58502 267444 59122 267528
rect 58502 267208 58689 267444
rect 58925 267208 59122 267444
rect 58502 267124 59122 267208
rect 58502 266888 58689 267124
rect 58925 266888 59122 267124
rect 58502 266804 59122 266888
rect 58502 266568 58689 266804
rect 58925 266568 59122 266804
rect 58502 266408 59122 266568
rect 59462 266618 60082 273952
rect 60422 267578 61042 274922
rect 61382 268538 62002 275876
rect 62342 269498 62962 276834
rect 63302 270458 63922 277792
rect 63302 269838 67172 270458
rect 62342 268878 66212 269498
rect 61382 267918 65252 268538
rect 60422 266958 64292 267578
rect 59462 265998 63332 266618
rect 62712 265360 63332 265998
rect 62712 265124 62897 265360
rect 63133 265124 63332 265360
rect 62712 265040 63332 265124
rect 62712 264804 62897 265040
rect 63133 264804 63332 265040
rect 62712 264720 63332 264804
rect 57542 264078 61412 264698
rect 47770 261245 59470 261466
rect 47770 258769 48071 261245
rect 49587 261184 59470 261245
rect 49587 258769 56555 261184
rect 47770 258708 56555 258769
rect 59351 258708 59470 261184
rect 47770 258466 59470 258708
rect 60792 257466 61412 264078
rect 62712 264484 62897 264720
rect 63133 264484 63332 264720
rect 62712 264400 63332 264484
rect 62712 264164 62897 264400
rect 63133 264164 63332 264400
rect 62712 264080 63332 264164
rect 62712 263844 62897 264080
rect 63133 263844 63332 264080
rect 62712 263760 63332 263844
rect 62712 263524 62897 263760
rect 63133 263524 63332 263760
rect 62712 263440 63332 263524
rect 62712 263204 62897 263440
rect 63133 263204 63332 263440
rect 62712 263120 63332 263204
rect 62712 262884 62897 263120
rect 63133 262884 63332 263120
rect 62712 262800 63332 262884
rect 62712 262564 62897 262800
rect 63133 262564 63332 262800
rect 62712 262402 63332 262564
rect 50170 257362 61412 257466
rect 50170 257245 60980 257362
rect 50170 254769 50471 257245
rect 51987 257184 60980 257245
rect 51987 254769 56564 257184
rect 50170 254708 56564 254769
rect 60320 257126 60980 257184
rect 61216 257126 61412 257362
rect 60320 257042 61412 257126
rect 60320 256806 60980 257042
rect 61216 256806 61412 257042
rect 60320 256722 61412 256806
rect 60320 256486 60980 256722
rect 61216 256486 61412 256722
rect 60320 256402 61412 256486
rect 60320 256166 60980 256402
rect 61216 256166 61412 256402
rect 60320 256082 61412 256166
rect 60320 255846 60980 256082
rect 61216 255846 61412 256082
rect 60320 255762 61412 255846
rect 60320 255526 60980 255762
rect 61216 255526 61412 255762
rect 60320 255442 61412 255526
rect 60320 255206 60980 255442
rect 61216 255206 61412 255442
rect 60320 255122 61412 255206
rect 60320 254886 60980 255122
rect 61216 254886 61412 255122
rect 60320 254802 61412 254886
rect 60320 254708 60980 254802
rect 50170 254566 60980 254708
rect 61216 254566 61412 254802
rect 50170 254466 61412 254566
rect 60792 254422 61412 254466
rect 52578 253370 63292 253466
rect 52578 253368 56232 253370
rect 52578 250572 52762 253368
rect 53638 250574 56232 253368
rect 63188 250574 63292 253370
rect 53638 250572 63292 250574
rect 52578 250466 63292 250572
rect 63672 245466 64292 266958
rect 40984 245370 64292 245466
rect 40984 245353 63863 245370
rect 40984 238397 41220 245353
rect 43376 245181 63863 245353
rect 43376 242705 56551 245181
rect 63187 245134 63863 245181
rect 64099 245134 64292 245370
rect 63187 245050 64292 245134
rect 63187 244814 63863 245050
rect 64099 244814 64292 245050
rect 63187 244730 64292 244814
rect 63187 244494 63863 244730
rect 64099 244494 64292 244730
rect 63187 244410 64292 244494
rect 63187 244174 63863 244410
rect 64099 244174 64292 244410
rect 63187 244090 64292 244174
rect 63187 243854 63863 244090
rect 64099 243854 64292 244090
rect 63187 243770 64292 243854
rect 63187 243534 63863 243770
rect 64099 243534 64292 243770
rect 63187 243450 64292 243534
rect 63187 243214 63863 243450
rect 64099 243214 64292 243450
rect 63187 243130 64292 243214
rect 63187 242894 63863 243130
rect 64099 242894 64292 243130
rect 63187 242810 64292 242894
rect 63187 242705 63863 242810
rect 43376 242574 63863 242705
rect 64099 242574 64292 242810
rect 43376 242466 64292 242574
rect 43376 238397 43612 242466
rect 63672 242358 64292 242466
rect 64632 241466 65252 267918
rect 65592 253358 66212 268878
rect 65592 253122 65775 253358
rect 66011 253122 66212 253358
rect 65592 253038 66212 253122
rect 65592 252802 65775 253038
rect 66011 252802 66212 253038
rect 65592 252718 66212 252802
rect 65592 252482 65775 252718
rect 66011 252482 66212 252718
rect 65592 252398 66212 252482
rect 65592 252162 65775 252398
rect 66011 252162 66212 252398
rect 65592 252078 66212 252162
rect 65592 251842 65775 252078
rect 66011 251842 66212 252078
rect 65592 251758 66212 251842
rect 65592 251522 65775 251758
rect 66011 251522 66212 251758
rect 65592 251438 66212 251522
rect 65592 251202 65775 251438
rect 66011 251202 66212 251438
rect 65592 251118 66212 251202
rect 65592 250882 65775 251118
rect 66011 250882 66212 251118
rect 65592 250798 66212 250882
rect 65592 250562 65775 250798
rect 66011 250562 66212 250798
rect 65592 250386 66212 250562
rect 66552 249370 67172 269838
rect 390772 269361 391558 269470
rect 390772 266565 390891 269361
rect 391447 266565 391558 269361
rect 390772 266474 391558 266565
rect 405822 269361 406608 269470
rect 405822 266565 405941 269361
rect 406497 266565 406608 269361
rect 405822 266474 406608 266565
rect 383994 265462 384174 265476
rect 383366 265208 384174 265462
rect 383366 263052 383487 265208
rect 384043 263052 384174 265208
rect 383366 262854 384174 263052
rect 383994 262244 384174 262854
rect 391374 262208 391554 266474
rect 399044 265462 399224 265476
rect 398416 265208 399224 265462
rect 398416 263052 398537 265208
rect 399093 263052 399224 265208
rect 398416 262854 399224 263052
rect 399044 262244 399224 262854
rect 406424 262208 406604 266474
rect 391944 261189 392846 261450
rect 391944 258713 392117 261189
rect 392673 258713 392846 261189
rect 391944 258468 392846 258713
rect 407064 261189 407966 261450
rect 407064 258713 407237 261189
rect 407793 258713 407966 261189
rect 407064 258468 407966 258713
rect 384586 257366 385708 257470
rect 384586 254570 384715 257366
rect 385591 254570 385708 257366
rect 384586 254452 385708 254570
rect 399686 257366 400808 257470
rect 399686 254570 399815 257366
rect 400691 254570 400808 257366
rect 399686 254452 400808 254570
rect 276722 253376 277260 253472
rect 276722 253140 276827 253376
rect 277063 253140 277260 253376
rect 276722 253056 277260 253140
rect 276722 252820 276827 253056
rect 277063 252820 277260 253056
rect 276722 252736 277260 252820
rect 276722 252500 276827 252736
rect 277063 252500 277260 252736
rect 276722 252416 277260 252500
rect 276722 252180 276827 252416
rect 277063 252180 277260 252416
rect 276722 252096 277260 252180
rect 276722 251860 276827 252096
rect 277063 251860 277260 252096
rect 276722 251776 277260 251860
rect 276722 251540 276827 251776
rect 277063 251540 277260 251776
rect 276722 251456 277260 251540
rect 276722 251220 276827 251456
rect 277063 251220 277260 251456
rect 276722 251136 277260 251220
rect 276722 250900 276827 251136
rect 277063 250900 277260 251136
rect 276722 250816 277260 250900
rect 276722 250580 276827 250816
rect 277063 250580 277260 250816
rect 276722 250470 277260 250580
rect 291722 253376 292260 253472
rect 291722 253140 291827 253376
rect 292063 253140 292260 253376
rect 291722 253056 292260 253140
rect 291722 252820 291827 253056
rect 292063 252820 292260 253056
rect 291722 252736 292260 252820
rect 291722 252500 291827 252736
rect 292063 252500 292260 252736
rect 291722 252416 292260 252500
rect 291722 252180 291827 252416
rect 292063 252180 292260 252416
rect 291722 252096 292260 252180
rect 291722 251860 291827 252096
rect 292063 251860 292260 252096
rect 291722 251776 292260 251860
rect 291722 251540 291827 251776
rect 292063 251540 292260 251776
rect 291722 251456 292260 251540
rect 291722 251220 291827 251456
rect 292063 251220 292260 251456
rect 291722 251136 292260 251220
rect 291722 250900 291827 251136
rect 292063 250900 292260 251136
rect 291722 250816 292260 250900
rect 291722 250580 291827 250816
rect 292063 250580 292260 250816
rect 291722 250470 292260 250580
rect 306762 253376 307300 253472
rect 306762 253140 306867 253376
rect 307103 253140 307300 253376
rect 306762 253056 307300 253140
rect 306762 252820 306867 253056
rect 307103 252820 307300 253056
rect 306762 252736 307300 252820
rect 306762 252500 306867 252736
rect 307103 252500 307300 252736
rect 306762 252416 307300 252500
rect 306762 252180 306867 252416
rect 307103 252180 307300 252416
rect 306762 252096 307300 252180
rect 306762 251860 306867 252096
rect 307103 251860 307300 252096
rect 306762 251776 307300 251860
rect 306762 251540 306867 251776
rect 307103 251540 307300 251776
rect 306762 251456 307300 251540
rect 306762 251220 306867 251456
rect 307103 251220 307300 251456
rect 306762 251136 307300 251220
rect 306762 250900 306867 251136
rect 307103 250900 307300 251136
rect 306762 250816 307300 250900
rect 306762 250580 306867 250816
rect 307103 250580 307300 250816
rect 306762 250470 307300 250580
rect 321882 253376 322420 253472
rect 321882 253140 321987 253376
rect 322223 253140 322420 253376
rect 321882 253056 322420 253140
rect 321882 252820 321987 253056
rect 322223 252820 322420 253056
rect 321882 252736 322420 252820
rect 321882 252500 321987 252736
rect 322223 252500 322420 252736
rect 321882 252416 322420 252500
rect 321882 252180 321987 252416
rect 322223 252180 322420 252416
rect 321882 252096 322420 252180
rect 321882 251860 321987 252096
rect 322223 251860 322420 252096
rect 321882 251776 322420 251860
rect 321882 251540 321987 251776
rect 322223 251540 322420 251776
rect 321882 251456 322420 251540
rect 321882 251220 321987 251456
rect 322223 251220 322420 251456
rect 321882 251136 322420 251220
rect 321882 250900 321987 251136
rect 322223 250900 322420 251136
rect 321882 250816 322420 250900
rect 321882 250580 321987 250816
rect 322223 250580 322420 250816
rect 321882 250470 322420 250580
rect 66552 249134 66739 249370
rect 66975 249134 67172 249370
rect 650618 249375 651238 277798
rect 658882 277774 674086 277975
rect 658856 277340 673450 277456
rect 658856 277266 670886 277340
rect 658856 277030 658965 277266
rect 659201 277030 659285 277266
rect 659521 277030 659605 277266
rect 659841 277030 659925 277266
rect 660161 277030 660245 277266
rect 660481 277030 660565 277266
rect 660801 277030 660885 277266
rect 661121 277030 661205 277266
rect 661441 277030 661525 277266
rect 661761 277030 661845 277266
rect 662081 277030 662165 277266
rect 662401 277030 662485 277266
rect 662721 277030 662805 277266
rect 663041 277030 670886 277266
rect 651578 253357 652198 276844
rect 658856 276816 670886 277030
rect 670818 276144 670886 276816
rect 673362 276144 673450 277340
rect 674016 276830 674086 277774
rect 676562 276830 676628 278346
rect 674016 276774 676628 276830
rect 670818 276016 673450 276144
rect 651578 250561 651614 253357
rect 652170 250561 652198 253357
rect 651578 250392 652198 250561
rect 66552 249050 67172 249134
rect 66552 248814 66739 249050
rect 66975 248814 67172 249050
rect 66552 248730 67172 248814
rect 66552 248494 66739 248730
rect 66975 248494 67172 248730
rect 66552 248410 67172 248494
rect 66552 248174 66739 248410
rect 66975 248174 67172 248410
rect 66552 248090 67172 248174
rect 66552 247854 66739 248090
rect 66975 247854 67172 248090
rect 66552 247770 67172 247854
rect 66552 247534 66739 247770
rect 66975 247534 67172 247770
rect 66552 247450 67172 247534
rect 66552 247214 66739 247450
rect 66975 247214 67172 247450
rect 66552 247130 67172 247214
rect 66552 246894 66739 247130
rect 66975 246894 67172 247130
rect 66552 246810 67172 246894
rect 66552 246574 66739 246810
rect 66975 246574 67172 246810
rect 66552 246348 67172 246574
rect 269364 249177 269812 249324
rect 269364 248941 269470 249177
rect 269706 248941 269812 249177
rect 269364 248857 269812 248941
rect 269364 248621 269470 248857
rect 269706 248621 269812 248857
rect 269364 248537 269812 248621
rect 269364 248301 269470 248537
rect 269706 248301 269812 248537
rect 269364 248217 269812 248301
rect 269364 247981 269470 248217
rect 269706 247981 269812 248217
rect 269364 247897 269812 247981
rect 269364 247661 269470 247897
rect 269706 247661 269812 247897
rect 269364 247577 269812 247661
rect 269364 247341 269470 247577
rect 269706 247341 269812 247577
rect 269364 247257 269812 247341
rect 269364 247021 269470 247257
rect 269706 247021 269812 247257
rect 269364 246937 269812 247021
rect 269364 246701 269470 246937
rect 269706 246701 269812 246937
rect 269364 246468 269812 246701
rect 284354 249177 284802 249324
rect 284354 248941 284460 249177
rect 284696 248941 284802 249177
rect 284354 248857 284802 248941
rect 284354 248621 284460 248857
rect 284696 248621 284802 248857
rect 284354 248537 284802 248621
rect 284354 248301 284460 248537
rect 284696 248301 284802 248537
rect 284354 248217 284802 248301
rect 284354 247981 284460 248217
rect 284696 247981 284802 248217
rect 284354 247897 284802 247981
rect 284354 247661 284460 247897
rect 284696 247661 284802 247897
rect 284354 247577 284802 247661
rect 284354 247341 284460 247577
rect 284696 247341 284802 247577
rect 284354 247257 284802 247341
rect 284354 247021 284460 247257
rect 284696 247021 284802 247257
rect 284354 246937 284802 247021
rect 284354 246701 284460 246937
rect 284696 246701 284802 246937
rect 284354 246468 284802 246701
rect 299354 249177 299802 249324
rect 299354 248941 299460 249177
rect 299696 248941 299802 249177
rect 299354 248857 299802 248941
rect 299354 248621 299460 248857
rect 299696 248621 299802 248857
rect 299354 248537 299802 248621
rect 299354 248301 299460 248537
rect 299696 248301 299802 248537
rect 299354 248217 299802 248301
rect 299354 247981 299460 248217
rect 299696 247981 299802 248217
rect 299354 247897 299802 247981
rect 299354 247661 299460 247897
rect 299696 247661 299802 247897
rect 299354 247577 299802 247661
rect 299354 247341 299460 247577
rect 299696 247341 299802 247577
rect 299354 247257 299802 247341
rect 299354 247021 299460 247257
rect 299696 247021 299802 247257
rect 299354 246937 299802 247021
rect 299354 246701 299460 246937
rect 299696 246701 299802 246937
rect 299354 246468 299802 246701
rect 314614 249177 315062 249324
rect 314614 248941 314720 249177
rect 314956 248941 315062 249177
rect 314614 248857 315062 248941
rect 314614 248621 314720 248857
rect 314956 248621 315062 248857
rect 314614 248537 315062 248621
rect 314614 248301 314720 248537
rect 314956 248301 315062 248537
rect 314614 248217 315062 248301
rect 314614 247981 314720 248217
rect 314956 247981 315062 248217
rect 314614 247897 315062 247981
rect 314614 247661 314720 247897
rect 314956 247661 315062 247897
rect 314614 247577 315062 247661
rect 314614 247341 314720 247577
rect 314956 247341 315062 247577
rect 314614 247257 315062 247341
rect 314614 247021 314720 247257
rect 314956 247021 315062 247257
rect 314614 246937 315062 247021
rect 314614 246701 314720 246937
rect 314956 246701 315062 246937
rect 314614 246468 315062 246701
rect 650618 246579 650648 249375
rect 651204 246579 651238 249375
rect 650618 246296 651238 246579
rect 199062 245373 199394 245464
rect 199062 245137 199110 245373
rect 199346 245137 199394 245373
rect 199062 245053 199394 245137
rect 199062 244817 199110 245053
rect 199346 244817 199394 245053
rect 199062 244733 199394 244817
rect 199062 244497 199110 244733
rect 199346 244497 199394 244733
rect 199062 244413 199394 244497
rect 199062 244177 199110 244413
rect 199346 244177 199394 244413
rect 199062 244093 199394 244177
rect 199062 243857 199110 244093
rect 199346 243857 199394 244093
rect 199062 243773 199394 243857
rect 199062 243537 199110 243773
rect 199346 243537 199394 243773
rect 199062 243453 199394 243537
rect 199062 243217 199110 243453
rect 199346 243217 199394 243453
rect 199062 243133 199394 243217
rect 199062 242897 199110 243133
rect 199346 242897 199394 243133
rect 199062 242813 199394 242897
rect 199062 242577 199110 242813
rect 199346 242577 199394 242813
rect 199062 242466 199394 242577
rect 209122 245375 209454 245466
rect 209122 245139 209170 245375
rect 209406 245139 209454 245375
rect 209122 245055 209454 245139
rect 209122 244819 209170 245055
rect 209406 244819 209454 245055
rect 209122 244735 209454 244819
rect 209122 244499 209170 244735
rect 209406 244499 209454 244735
rect 209122 244415 209454 244499
rect 209122 244179 209170 244415
rect 209406 244179 209454 244415
rect 209122 244095 209454 244179
rect 209122 243859 209170 244095
rect 209406 243859 209454 244095
rect 209122 243775 209454 243859
rect 209122 243539 209170 243775
rect 209406 243539 209454 243775
rect 209122 243455 209454 243539
rect 209122 243219 209170 243455
rect 209406 243219 209454 243455
rect 209122 243135 209454 243219
rect 209122 242899 209170 243135
rect 209406 242899 209454 243135
rect 209122 242815 209454 242899
rect 209122 242579 209170 242815
rect 209406 242579 209454 242815
rect 209122 242468 209454 242579
rect 40984 238266 43612 238397
rect 44196 241366 65252 241466
rect 44196 241263 64813 241366
rect 44196 234627 44408 241263
rect 46564 241215 64813 241263
rect 46564 238739 56566 241215
rect 63202 241130 64813 241215
rect 65049 241130 65252 241366
rect 63202 241046 65252 241130
rect 63202 240810 64813 241046
rect 65049 240810 65252 241046
rect 63202 240726 65252 240810
rect 63202 240490 64813 240726
rect 65049 240490 65252 240726
rect 63202 240406 65252 240490
rect 63202 240170 64813 240406
rect 65049 240170 65252 240406
rect 63202 240086 65252 240170
rect 63202 239850 64813 240086
rect 65049 239850 65252 240086
rect 63202 239766 65252 239850
rect 63202 239530 64813 239766
rect 65049 239530 65252 239766
rect 63202 239446 65252 239530
rect 63202 239210 64813 239446
rect 65049 239210 65252 239446
rect 63202 239126 65252 239210
rect 63202 238890 64813 239126
rect 65049 238890 65252 239126
rect 63202 238806 65252 238890
rect 63202 238739 64813 238806
rect 46564 238570 64813 238739
rect 65049 238570 65252 238806
rect 46564 238466 65252 238570
rect 194882 241373 195214 241464
rect 194882 241137 194930 241373
rect 195166 241137 195214 241373
rect 194882 241053 195214 241137
rect 194882 240817 194930 241053
rect 195166 240817 195214 241053
rect 194882 240733 195214 240817
rect 194882 240497 194930 240733
rect 195166 240497 195214 240733
rect 194882 240413 195214 240497
rect 194882 240177 194930 240413
rect 195166 240177 195214 240413
rect 194882 240093 195214 240177
rect 194882 239857 194930 240093
rect 195166 239857 195214 240093
rect 194882 239773 195214 239857
rect 194882 239537 194930 239773
rect 195166 239537 195214 239773
rect 194882 239453 195214 239537
rect 194882 239217 194930 239453
rect 195166 239217 195214 239453
rect 194882 239133 195214 239217
rect 194882 238897 194930 239133
rect 195166 238897 195214 239133
rect 194882 238813 195214 238897
rect 194882 238577 194930 238813
rect 195166 238577 195214 238813
rect 194882 238466 195214 238577
rect 205002 241373 205334 241464
rect 205002 241137 205050 241373
rect 205286 241137 205334 241373
rect 205002 241053 205334 241137
rect 205002 240817 205050 241053
rect 205286 240817 205334 241053
rect 205002 240733 205334 240817
rect 205002 240497 205050 240733
rect 205286 240497 205334 240733
rect 205002 240413 205334 240497
rect 205002 240177 205050 240413
rect 205286 240177 205334 240413
rect 205002 240093 205334 240177
rect 205002 239857 205050 240093
rect 205286 239857 205334 240093
rect 205002 239773 205334 239857
rect 205002 239537 205050 239773
rect 205286 239537 205334 239773
rect 205002 239453 205334 239537
rect 205002 239217 205050 239453
rect 205286 239217 205334 239453
rect 205002 239133 205334 239217
rect 205002 238897 205050 239133
rect 205286 238897 205334 239133
rect 205002 238813 205334 238897
rect 205002 238577 205050 238813
rect 205286 238577 205334 238813
rect 205002 238466 205334 238577
rect 652538 241371 653158 275876
rect 653498 245373 654118 274916
rect 658950 274452 669812 274574
rect 658950 274365 667448 274452
rect 658950 274129 659185 274365
rect 659421 274129 659505 274365
rect 659741 274129 659825 274365
rect 660061 274129 660145 274365
rect 660381 274129 660465 274365
rect 660701 274129 660785 274365
rect 661021 274129 661105 274365
rect 661341 274129 661425 274365
rect 661661 274129 661745 274365
rect 661981 274129 662065 274365
rect 662301 274129 662385 274365
rect 662621 274129 662705 274365
rect 662941 274129 667448 274365
rect 654458 265359 655078 273956
rect 658950 273938 667448 274129
rect 667216 273256 667448 273938
rect 669604 273256 669812 274452
rect 667216 273138 669812 273256
rect 655418 269361 656038 273004
rect 655418 269125 655607 269361
rect 655843 269125 656038 269361
rect 655418 269041 656038 269125
rect 655418 268805 655607 269041
rect 655843 268805 656038 269041
rect 655418 268721 656038 268805
rect 655418 268485 655607 268721
rect 655843 268485 656038 268721
rect 655418 268401 656038 268485
rect 655418 268165 655607 268401
rect 655843 268165 656038 268401
rect 655418 268081 656038 268165
rect 655418 267845 655607 268081
rect 655843 267845 656038 268081
rect 655418 267761 656038 267845
rect 655418 267525 655607 267761
rect 655843 267525 656038 267761
rect 655418 267441 656038 267525
rect 655418 267205 655607 267441
rect 655843 267205 656038 267441
rect 655418 267121 656038 267205
rect 655418 266885 655607 267121
rect 655843 266885 656038 267121
rect 655418 266801 656038 266885
rect 655418 266565 655607 266801
rect 655843 266565 656038 266801
rect 655418 266386 656038 266565
rect 654458 265123 654649 265359
rect 654885 265123 655078 265359
rect 654458 265039 655078 265123
rect 654458 264803 654649 265039
rect 654885 264803 655078 265039
rect 654458 264719 655078 264803
rect 654458 264483 654649 264719
rect 654885 264483 655078 264719
rect 654458 264399 655078 264483
rect 654458 264163 654649 264399
rect 654885 264163 655078 264399
rect 654458 264079 655078 264163
rect 654458 263843 654649 264079
rect 654885 263843 655078 264079
rect 654458 263759 655078 263843
rect 654458 263523 654649 263759
rect 654885 263523 655078 263759
rect 654458 263439 655078 263523
rect 654458 263203 654649 263439
rect 654885 263203 655078 263439
rect 654458 263119 655078 263203
rect 654458 262883 654649 263119
rect 654885 262883 655078 263119
rect 654458 262799 655078 262883
rect 654458 262563 654649 262799
rect 654885 262563 655078 262799
rect 654458 262362 655078 262563
rect 656378 257355 656998 272036
rect 657338 261373 657958 271082
rect 657338 261137 657523 261373
rect 657759 261137 657958 261373
rect 657338 261053 657958 261137
rect 657338 260817 657523 261053
rect 657759 260817 657958 261053
rect 657338 260733 657958 260817
rect 657338 260497 657523 260733
rect 657759 260497 657958 260733
rect 657338 260413 657958 260497
rect 657338 260177 657523 260413
rect 657759 260177 657958 260413
rect 657338 260093 657958 260177
rect 657338 259857 657523 260093
rect 657759 259857 657958 260093
rect 657338 259773 657958 259857
rect 657338 259537 657523 259773
rect 657759 259537 657958 259773
rect 657338 259453 657958 259537
rect 657338 259217 657523 259453
rect 657759 259217 657958 259453
rect 657338 259133 657958 259217
rect 657338 258897 657523 259133
rect 657759 258897 657958 259133
rect 657338 258813 657958 258897
rect 657338 258577 657523 258813
rect 657759 258577 657958 258813
rect 657338 258390 657958 258577
rect 656378 257119 656561 257355
rect 656797 257119 656998 257355
rect 656378 257035 656998 257119
rect 656378 256799 656561 257035
rect 656797 256799 656998 257035
rect 656378 256715 656998 256799
rect 656378 256479 656561 256715
rect 656797 256479 656998 256715
rect 656378 256395 656998 256479
rect 656378 256159 656561 256395
rect 656797 256159 656998 256395
rect 656378 256075 656998 256159
rect 656378 255839 656561 256075
rect 656797 255839 656998 256075
rect 656378 255755 656998 255839
rect 656378 255519 656561 255755
rect 656797 255519 656998 255755
rect 656378 255435 656998 255519
rect 656378 255199 656561 255435
rect 656797 255199 656998 255435
rect 656378 255115 656998 255199
rect 656378 254879 656561 255115
rect 656797 254879 656998 255115
rect 656378 254795 656998 254879
rect 656378 254559 656561 254795
rect 656797 254559 656998 254795
rect 656378 254386 656998 254559
rect 666890 249213 676670 249476
rect 666890 246737 667112 249213
rect 669588 249194 676670 249213
rect 669588 246737 674226 249194
rect 666890 246718 674226 246737
rect 676382 246718 676670 249194
rect 666890 246466 676670 246718
rect 653498 245137 653679 245373
rect 653915 245137 654118 245373
rect 653498 245053 654118 245137
rect 653498 244817 653679 245053
rect 653915 244817 654118 245053
rect 653498 244733 654118 244817
rect 653498 244497 653679 244733
rect 653915 244497 654118 244733
rect 653498 244413 654118 244497
rect 653498 244177 653679 244413
rect 653915 244177 654118 244413
rect 653498 244093 654118 244177
rect 653498 243857 653679 244093
rect 653915 243857 654118 244093
rect 653498 243773 654118 243857
rect 653498 243537 653679 243773
rect 653915 243537 654118 243773
rect 653498 243453 654118 243537
rect 653498 243217 653679 243453
rect 653915 243217 654118 243453
rect 653498 243133 654118 243217
rect 653498 242897 653679 243133
rect 653915 242897 654118 243133
rect 653498 242813 654118 242897
rect 653498 242577 653679 242813
rect 653915 242577 654118 242813
rect 653498 242362 654118 242577
rect 652538 241135 652721 241371
rect 652957 241135 653158 241371
rect 652538 241051 653158 241135
rect 652538 240815 652721 241051
rect 652957 240815 653158 241051
rect 652538 240731 653158 240815
rect 652538 240495 652721 240731
rect 652957 240495 653158 240731
rect 652538 240411 653158 240495
rect 652538 240175 652721 240411
rect 652957 240175 653158 240411
rect 652538 240091 653158 240175
rect 652538 239855 652721 240091
rect 652957 239855 653158 240091
rect 652538 239771 653158 239855
rect 652538 239535 652721 239771
rect 652957 239535 653158 239771
rect 652538 239451 653158 239535
rect 652538 239215 652721 239451
rect 652957 239215 653158 239451
rect 652538 239131 653158 239215
rect 652538 238895 652721 239131
rect 652957 238895 653158 239131
rect 652538 238811 653158 238895
rect 652538 238575 652721 238811
rect 652957 238575 653158 238811
rect 46564 234627 46802 238466
rect 64632 238400 65252 238466
rect 652538 238266 653158 238575
rect 44196 234466 46802 234627
rect 47786 237221 63250 237466
rect 47786 237215 56455 237221
rect 47786 234739 48091 237215
rect 50567 234745 56455 237215
rect 63091 234745 63250 237221
rect 50567 234739 63250 234745
rect 47786 234466 63250 234739
rect 140444 237361 140924 237474
rect 140444 237125 140520 237361
rect 140756 237125 140924 237361
rect 140444 237041 140924 237125
rect 140444 236805 140520 237041
rect 140756 236805 140924 237041
rect 140444 236721 140924 236805
rect 140444 236485 140520 236721
rect 140756 236485 140924 236721
rect 140444 236401 140924 236485
rect 140444 236165 140520 236401
rect 140756 236165 140924 236401
rect 140444 236081 140924 236165
rect 140444 235845 140520 236081
rect 140756 235845 140924 236081
rect 140444 235761 140924 235845
rect 140444 235525 140520 235761
rect 140756 235525 140924 235761
rect 140444 235441 140924 235525
rect 140444 235205 140520 235441
rect 140756 235205 140924 235441
rect 140444 235121 140924 235205
rect 140444 234885 140520 235121
rect 140756 234885 140924 235121
rect 140444 234801 140924 234885
rect 140444 234565 140520 234801
rect 140756 234565 140924 234801
rect 140444 234448 140924 234565
rect 155524 237361 156004 237474
rect 155524 237125 155600 237361
rect 155836 237125 156004 237361
rect 155524 237041 156004 237125
rect 155524 236805 155600 237041
rect 155836 236805 156004 237041
rect 155524 236721 156004 236805
rect 155524 236485 155600 236721
rect 155836 236485 156004 236721
rect 155524 236401 156004 236485
rect 155524 236165 155600 236401
rect 155836 236165 156004 236401
rect 155524 236081 156004 236165
rect 155524 235845 155600 236081
rect 155836 235845 156004 236081
rect 155524 235761 156004 235845
rect 155524 235525 155600 235761
rect 155836 235525 156004 235761
rect 155524 235441 156004 235525
rect 155524 235205 155600 235441
rect 155836 235205 156004 235441
rect 155524 235121 156004 235205
rect 155524 234885 155600 235121
rect 155836 234885 156004 235121
rect 155524 234801 156004 234885
rect 155524 234565 155600 234801
rect 155836 234565 156004 234801
rect 155524 234448 156004 234565
rect 170574 237361 171054 237474
rect 170574 237125 170650 237361
rect 170886 237125 171054 237361
rect 170574 237041 171054 237125
rect 170574 236805 170650 237041
rect 170886 236805 171054 237041
rect 170574 236721 171054 236805
rect 170574 236485 170650 236721
rect 170886 236485 171054 236721
rect 170574 236401 171054 236485
rect 170574 236165 170650 236401
rect 170886 236165 171054 236401
rect 170574 236081 171054 236165
rect 170574 235845 170650 236081
rect 170886 235845 171054 236081
rect 170574 235761 171054 235845
rect 170574 235525 170650 235761
rect 170886 235525 171054 235761
rect 170574 235441 171054 235525
rect 170574 235205 170650 235441
rect 170886 235205 171054 235441
rect 170574 235121 171054 235205
rect 170574 234885 170650 235121
rect 170886 234885 171054 235121
rect 170574 234801 171054 234885
rect 170574 234565 170650 234801
rect 170886 234565 171054 234801
rect 170574 234448 171054 234565
rect 185584 237361 186064 237474
rect 185584 237125 185660 237361
rect 185896 237125 186064 237361
rect 185584 237041 186064 237125
rect 185584 236805 185660 237041
rect 185896 236805 186064 237041
rect 185584 236721 186064 236805
rect 185584 236485 185660 236721
rect 185896 236485 186064 236721
rect 185584 236401 186064 236485
rect 185584 236165 185660 236401
rect 185896 236165 186064 236401
rect 185584 236081 186064 236165
rect 185584 235845 185660 236081
rect 185896 235845 186064 236081
rect 185584 235761 186064 235845
rect 185584 235525 185660 235761
rect 185896 235525 186064 235761
rect 185584 235441 186064 235525
rect 185584 235205 185660 235441
rect 185896 235205 186064 235441
rect 185584 235121 186064 235205
rect 185584 234885 185660 235121
rect 185896 234885 186064 235121
rect 185584 234801 186064 234885
rect 185584 234565 185660 234801
rect 185896 234565 186064 234801
rect 185584 234448 186064 234565
rect 215724 237361 216204 237474
rect 215724 237125 215800 237361
rect 216036 237125 216204 237361
rect 215724 237041 216204 237125
rect 215724 236805 215800 237041
rect 216036 236805 216204 237041
rect 215724 236721 216204 236805
rect 215724 236485 215800 236721
rect 216036 236485 216204 236721
rect 215724 236401 216204 236485
rect 215724 236165 215800 236401
rect 216036 236165 216204 236401
rect 215724 236081 216204 236165
rect 215724 235845 215800 236081
rect 216036 235845 216204 236081
rect 215724 235761 216204 235845
rect 215724 235525 215800 235761
rect 216036 235525 216204 235761
rect 215724 235441 216204 235525
rect 215724 235205 215800 235441
rect 216036 235205 216204 235441
rect 215724 235121 216204 235205
rect 215724 234885 215800 235121
rect 216036 234885 216204 235121
rect 215724 234801 216204 234885
rect 215724 234565 215800 234801
rect 216036 234565 216204 234801
rect 215724 234448 216204 234565
rect 230774 237361 231254 237474
rect 230774 237125 230850 237361
rect 231086 237125 231254 237361
rect 230774 237041 231254 237125
rect 230774 236805 230850 237041
rect 231086 236805 231254 237041
rect 230774 236721 231254 236805
rect 230774 236485 230850 236721
rect 231086 236485 231254 236721
rect 230774 236401 231254 236485
rect 230774 236165 230850 236401
rect 231086 236165 231254 236401
rect 230774 236081 231254 236165
rect 230774 235845 230850 236081
rect 231086 235845 231254 236081
rect 230774 235761 231254 235845
rect 230774 235525 230850 235761
rect 231086 235525 231254 235761
rect 230774 235441 231254 235525
rect 230774 235205 230850 235441
rect 231086 235205 231254 235441
rect 230774 235121 231254 235205
rect 230774 234885 230850 235121
rect 231086 234885 231254 235121
rect 230774 234801 231254 234885
rect 230774 234565 230850 234801
rect 231086 234565 231254 234801
rect 230774 234448 231254 234565
rect 245824 237361 246304 237474
rect 245824 237125 245900 237361
rect 246136 237125 246304 237361
rect 245824 237041 246304 237125
rect 245824 236805 245900 237041
rect 246136 236805 246304 237041
rect 245824 236721 246304 236805
rect 245824 236485 245900 236721
rect 246136 236485 246304 236721
rect 245824 236401 246304 236485
rect 245824 236165 245900 236401
rect 246136 236165 246304 236401
rect 245824 236081 246304 236165
rect 245824 235845 245900 236081
rect 246136 235845 246304 236081
rect 245824 235761 246304 235845
rect 245824 235525 245900 235761
rect 246136 235525 246304 235761
rect 245824 235441 246304 235525
rect 245824 235205 245900 235441
rect 246136 235205 246304 235441
rect 245824 235121 246304 235205
rect 245824 234885 245900 235121
rect 246136 234885 246304 235121
rect 245824 234801 246304 234885
rect 245824 234565 245900 234801
rect 246136 234565 246304 234801
rect 245824 234448 246304 234565
rect 260874 237361 261354 237474
rect 260874 237125 260950 237361
rect 261186 237125 261354 237361
rect 260874 237041 261354 237125
rect 260874 236805 260950 237041
rect 261186 236805 261354 237041
rect 260874 236721 261354 236805
rect 260874 236485 260950 236721
rect 261186 236485 261354 236721
rect 260874 236401 261354 236485
rect 260874 236165 260950 236401
rect 261186 236165 261354 236401
rect 260874 236081 261354 236165
rect 260874 235845 260950 236081
rect 261186 235845 261354 236081
rect 260874 235761 261354 235845
rect 260874 235525 260950 235761
rect 261186 235525 261354 235761
rect 260874 235441 261354 235525
rect 260874 235205 260950 235441
rect 261186 235205 261354 235441
rect 260874 235121 261354 235205
rect 260874 234885 260950 235121
rect 261186 234885 261354 235121
rect 260874 234801 261354 234885
rect 260874 234565 260950 234801
rect 261186 234565 261354 234801
rect 260874 234448 261354 234565
rect 275924 237361 276404 237474
rect 275924 237125 276000 237361
rect 276236 237125 276404 237361
rect 275924 237041 276404 237125
rect 275924 236805 276000 237041
rect 276236 236805 276404 237041
rect 275924 236721 276404 236805
rect 275924 236485 276000 236721
rect 276236 236485 276404 236721
rect 275924 236401 276404 236485
rect 275924 236165 276000 236401
rect 276236 236165 276404 236401
rect 275924 236081 276404 236165
rect 275924 235845 276000 236081
rect 276236 235845 276404 236081
rect 275924 235761 276404 235845
rect 275924 235525 276000 235761
rect 276236 235525 276404 235761
rect 275924 235441 276404 235525
rect 275924 235205 276000 235441
rect 276236 235205 276404 235441
rect 275924 235121 276404 235205
rect 275924 234885 276000 235121
rect 276236 234885 276404 235121
rect 275924 234801 276404 234885
rect 275924 234565 276000 234801
rect 276236 234565 276404 234801
rect 275924 234448 276404 234565
rect 290974 237361 291454 237474
rect 290974 237125 291050 237361
rect 291286 237125 291454 237361
rect 290974 237041 291454 237125
rect 290974 236805 291050 237041
rect 291286 236805 291454 237041
rect 290974 236721 291454 236805
rect 290974 236485 291050 236721
rect 291286 236485 291454 236721
rect 290974 236401 291454 236485
rect 290974 236165 291050 236401
rect 291286 236165 291454 236401
rect 290974 236081 291454 236165
rect 290974 235845 291050 236081
rect 291286 235845 291454 236081
rect 290974 235761 291454 235845
rect 290974 235525 291050 235761
rect 291286 235525 291454 235761
rect 290974 235441 291454 235525
rect 290974 235205 291050 235441
rect 291286 235205 291454 235441
rect 290974 235121 291454 235205
rect 290974 234885 291050 235121
rect 291286 234885 291454 235121
rect 290974 234801 291454 234885
rect 290974 234565 291050 234801
rect 291286 234565 291454 234801
rect 290974 234448 291454 234565
rect 305984 237361 306464 237474
rect 305984 237125 306060 237361
rect 306296 237125 306464 237361
rect 305984 237041 306464 237125
rect 305984 236805 306060 237041
rect 306296 236805 306464 237041
rect 305984 236721 306464 236805
rect 305984 236485 306060 236721
rect 306296 236485 306464 236721
rect 305984 236401 306464 236485
rect 305984 236165 306060 236401
rect 306296 236165 306464 236401
rect 305984 236081 306464 236165
rect 305984 235845 306060 236081
rect 306296 235845 306464 236081
rect 305984 235761 306464 235845
rect 305984 235525 306060 235761
rect 306296 235525 306464 235761
rect 305984 235441 306464 235525
rect 305984 235205 306060 235441
rect 306296 235205 306464 235441
rect 305984 235121 306464 235205
rect 305984 234885 306060 235121
rect 306296 234885 306464 235121
rect 305984 234801 306464 234885
rect 305984 234565 306060 234801
rect 306296 234565 306464 234801
rect 305984 234448 306464 234565
rect 321174 237361 321654 237474
rect 321174 237125 321250 237361
rect 321486 237125 321654 237361
rect 321174 237041 321654 237125
rect 321174 236805 321250 237041
rect 321486 236805 321654 237041
rect 321174 236721 321654 236805
rect 321174 236485 321250 236721
rect 321486 236485 321654 236721
rect 321174 236401 321654 236485
rect 321174 236165 321250 236401
rect 321486 236165 321654 236401
rect 321174 236081 321654 236165
rect 321174 235845 321250 236081
rect 321486 235845 321654 236081
rect 321174 235761 321654 235845
rect 321174 235525 321250 235761
rect 321486 235525 321654 235761
rect 321174 235441 321654 235525
rect 321174 235205 321250 235441
rect 321486 235205 321654 235441
rect 321174 235121 321654 235205
rect 321174 234885 321250 235121
rect 321486 234885 321654 235121
rect 321174 234801 321654 234885
rect 321174 234565 321250 234801
rect 321486 234565 321654 234801
rect 321174 234448 321654 234565
rect 336124 237361 336604 237474
rect 336124 237125 336200 237361
rect 336436 237125 336604 237361
rect 336124 237041 336604 237125
rect 336124 236805 336200 237041
rect 336436 236805 336604 237041
rect 336124 236721 336604 236805
rect 336124 236485 336200 236721
rect 336436 236485 336604 236721
rect 336124 236401 336604 236485
rect 336124 236165 336200 236401
rect 336436 236165 336604 236401
rect 336124 236081 336604 236165
rect 336124 235845 336200 236081
rect 336436 235845 336604 236081
rect 336124 235761 336604 235845
rect 336124 235525 336200 235761
rect 336436 235525 336604 235761
rect 336124 235441 336604 235525
rect 336124 235205 336200 235441
rect 336436 235205 336604 235441
rect 336124 235121 336604 235205
rect 336124 234885 336200 235121
rect 336436 234885 336604 235121
rect 336124 234801 336604 234885
rect 336124 234565 336200 234801
rect 336436 234565 336604 234801
rect 336124 234448 336604 234565
rect 351274 237361 351754 237474
rect 351274 237125 351350 237361
rect 351586 237125 351754 237361
rect 351274 237041 351754 237125
rect 351274 236805 351350 237041
rect 351586 236805 351754 237041
rect 351274 236721 351754 236805
rect 351274 236485 351350 236721
rect 351586 236485 351754 236721
rect 351274 236401 351754 236485
rect 351274 236165 351350 236401
rect 351586 236165 351754 236401
rect 351274 236081 351754 236165
rect 351274 235845 351350 236081
rect 351586 235845 351754 236081
rect 351274 235761 351754 235845
rect 351274 235525 351350 235761
rect 351586 235525 351754 235761
rect 351274 235441 351754 235525
rect 351274 235205 351350 235441
rect 351586 235205 351754 235441
rect 351274 235121 351754 235205
rect 351274 234885 351350 235121
rect 351586 234885 351754 235121
rect 351274 234801 351754 234885
rect 351274 234565 351350 234801
rect 351586 234565 351754 234801
rect 351274 234448 351754 234565
rect 366224 237361 366704 237474
rect 366224 237125 366300 237361
rect 366536 237125 366704 237361
rect 366224 237041 366704 237125
rect 366224 236805 366300 237041
rect 366536 236805 366704 237041
rect 366224 236721 366704 236805
rect 366224 236485 366300 236721
rect 366536 236485 366704 236721
rect 366224 236401 366704 236485
rect 366224 236165 366300 236401
rect 366536 236165 366704 236401
rect 366224 236081 366704 236165
rect 366224 235845 366300 236081
rect 366536 235845 366704 236081
rect 366224 235761 366704 235845
rect 366224 235525 366300 235761
rect 366536 235525 366704 235761
rect 366224 235441 366704 235525
rect 366224 235205 366300 235441
rect 366536 235205 366704 235441
rect 366224 235121 366704 235205
rect 366224 234885 366300 235121
rect 366536 234885 366704 235121
rect 366224 234801 366704 234885
rect 366224 234565 366300 234801
rect 366536 234565 366704 234801
rect 366224 234448 366704 234565
rect 381074 237361 381554 237474
rect 381074 237125 381150 237361
rect 381386 237125 381554 237361
rect 381074 237041 381554 237125
rect 381074 236805 381150 237041
rect 381386 236805 381554 237041
rect 381074 236721 381554 236805
rect 381074 236485 381150 236721
rect 381386 236485 381554 236721
rect 381074 236401 381554 236485
rect 381074 236165 381150 236401
rect 381386 236165 381554 236401
rect 381074 236081 381554 236165
rect 381074 235845 381150 236081
rect 381386 235845 381554 236081
rect 381074 235761 381554 235845
rect 381074 235525 381150 235761
rect 381386 235525 381554 235761
rect 381074 235441 381554 235525
rect 381074 235205 381150 235441
rect 381386 235205 381554 235441
rect 381074 235121 381554 235205
rect 381074 234885 381150 235121
rect 381386 234885 381554 235121
rect 381074 234801 381554 234885
rect 381074 234565 381150 234801
rect 381386 234565 381554 234801
rect 381074 234448 381554 234565
rect 396244 237361 396724 237474
rect 396244 237125 396320 237361
rect 396556 237125 396724 237361
rect 396244 237041 396724 237125
rect 396244 236805 396320 237041
rect 396556 236805 396724 237041
rect 396244 236721 396724 236805
rect 396244 236485 396320 236721
rect 396556 236485 396724 236721
rect 396244 236401 396724 236485
rect 396244 236165 396320 236401
rect 396556 236165 396724 236401
rect 396244 236081 396724 236165
rect 396244 235845 396320 236081
rect 396556 235845 396724 236081
rect 396244 235761 396724 235845
rect 396244 235525 396320 235761
rect 396556 235525 396724 235761
rect 396244 235441 396724 235525
rect 396244 235205 396320 235441
rect 396556 235205 396724 235441
rect 396244 235121 396724 235205
rect 396244 234885 396320 235121
rect 396556 234885 396724 235121
rect 396244 234801 396724 234885
rect 396244 234565 396320 234801
rect 396556 234565 396724 234801
rect 396244 234448 396724 234565
rect 411374 237361 411854 237474
rect 411374 237125 411450 237361
rect 411686 237125 411854 237361
rect 411374 237041 411854 237125
rect 411374 236805 411450 237041
rect 411686 236805 411854 237041
rect 411374 236721 411854 236805
rect 411374 236485 411450 236721
rect 411686 236485 411854 236721
rect 411374 236401 411854 236485
rect 411374 236165 411450 236401
rect 411686 236165 411854 236401
rect 411374 236081 411854 236165
rect 411374 235845 411450 236081
rect 411686 235845 411854 236081
rect 411374 235761 411854 235845
rect 411374 235525 411450 235761
rect 411686 235525 411854 235761
rect 411374 235441 411854 235525
rect 411374 235205 411450 235441
rect 411686 235205 411854 235441
rect 411374 235121 411854 235205
rect 411374 234885 411450 235121
rect 411686 234885 411854 235121
rect 411374 234801 411854 234885
rect 411374 234565 411450 234801
rect 411686 234565 411854 234801
rect 411374 234448 411854 234565
rect 426424 237361 426904 237474
rect 426424 237125 426500 237361
rect 426736 237125 426904 237361
rect 426424 237041 426904 237125
rect 426424 236805 426500 237041
rect 426736 236805 426904 237041
rect 426424 236721 426904 236805
rect 426424 236485 426500 236721
rect 426736 236485 426904 236721
rect 426424 236401 426904 236485
rect 426424 236165 426500 236401
rect 426736 236165 426904 236401
rect 426424 236081 426904 236165
rect 426424 235845 426500 236081
rect 426736 235845 426904 236081
rect 426424 235761 426904 235845
rect 426424 235525 426500 235761
rect 426736 235525 426904 235761
rect 426424 235441 426904 235525
rect 426424 235205 426500 235441
rect 426736 235205 426904 235441
rect 426424 235121 426904 235205
rect 426424 234885 426500 235121
rect 426736 234885 426904 235121
rect 426424 234801 426904 234885
rect 426424 234565 426500 234801
rect 426736 234565 426904 234801
rect 426424 234448 426904 234565
rect 441474 237361 441954 237474
rect 441474 237125 441550 237361
rect 441786 237125 441954 237361
rect 441474 237041 441954 237125
rect 441474 236805 441550 237041
rect 441786 236805 441954 237041
rect 441474 236721 441954 236805
rect 441474 236485 441550 236721
rect 441786 236485 441954 236721
rect 441474 236401 441954 236485
rect 441474 236165 441550 236401
rect 441786 236165 441954 236401
rect 441474 236081 441954 236165
rect 441474 235845 441550 236081
rect 441786 235845 441954 236081
rect 441474 235761 441954 235845
rect 441474 235525 441550 235761
rect 441786 235525 441954 235761
rect 441474 235441 441954 235525
rect 441474 235205 441550 235441
rect 441786 235205 441954 235441
rect 441474 235121 441954 235205
rect 441474 234885 441550 235121
rect 441786 234885 441954 235121
rect 441474 234801 441954 234885
rect 441474 234565 441550 234801
rect 441786 234565 441954 234801
rect 441474 234448 441954 234565
rect 456524 237361 457004 237474
rect 456524 237125 456600 237361
rect 456836 237125 457004 237361
rect 456524 237041 457004 237125
rect 456524 236805 456600 237041
rect 456836 236805 457004 237041
rect 456524 236721 457004 236805
rect 456524 236485 456600 236721
rect 456836 236485 457004 236721
rect 456524 236401 457004 236485
rect 456524 236165 456600 236401
rect 456836 236165 457004 236401
rect 456524 236081 457004 236165
rect 456524 235845 456600 236081
rect 456836 235845 457004 236081
rect 456524 235761 457004 235845
rect 456524 235525 456600 235761
rect 456836 235525 457004 235761
rect 456524 235441 457004 235525
rect 456524 235205 456600 235441
rect 456836 235205 457004 235441
rect 456524 235121 457004 235205
rect 456524 234885 456600 235121
rect 456836 234885 457004 235121
rect 456524 234801 457004 234885
rect 456524 234565 456600 234801
rect 456836 234565 457004 234801
rect 456524 234448 457004 234565
rect 471574 237361 472054 237474
rect 471574 237125 471650 237361
rect 471886 237125 472054 237361
rect 471574 237041 472054 237125
rect 471574 236805 471650 237041
rect 471886 236805 472054 237041
rect 471574 236721 472054 236805
rect 471574 236485 471650 236721
rect 471886 236485 472054 236721
rect 471574 236401 472054 236485
rect 471574 236165 471650 236401
rect 471886 236165 472054 236401
rect 471574 236081 472054 236165
rect 471574 235845 471650 236081
rect 471886 235845 472054 236081
rect 471574 235761 472054 235845
rect 471574 235525 471650 235761
rect 471886 235525 472054 235761
rect 471574 235441 472054 235525
rect 471574 235205 471650 235441
rect 471886 235205 472054 235441
rect 471574 235121 472054 235205
rect 471574 234885 471650 235121
rect 471886 234885 472054 235121
rect 471574 234801 472054 234885
rect 471574 234565 471650 234801
rect 471886 234565 472054 234801
rect 471574 234448 472054 234565
rect 486624 237361 487104 237474
rect 486624 237125 486700 237361
rect 486936 237125 487104 237361
rect 486624 237041 487104 237125
rect 486624 236805 486700 237041
rect 486936 236805 487104 237041
rect 486624 236721 487104 236805
rect 486624 236485 486700 236721
rect 486936 236485 487104 236721
rect 486624 236401 487104 236485
rect 486624 236165 486700 236401
rect 486936 236165 487104 236401
rect 486624 236081 487104 236165
rect 486624 235845 486700 236081
rect 486936 235845 487104 236081
rect 486624 235761 487104 235845
rect 486624 235525 486700 235761
rect 486936 235525 487104 235761
rect 486624 235441 487104 235525
rect 486624 235205 486700 235441
rect 486936 235205 487104 235441
rect 486624 235121 487104 235205
rect 486624 234885 486700 235121
rect 486936 234885 487104 235121
rect 486624 234801 487104 234885
rect 486624 234565 486700 234801
rect 486936 234565 487104 234801
rect 486624 234448 487104 234565
rect 501674 237361 502154 237474
rect 501674 237125 501750 237361
rect 501986 237125 502154 237361
rect 501674 237041 502154 237125
rect 501674 236805 501750 237041
rect 501986 236805 502154 237041
rect 501674 236721 502154 236805
rect 501674 236485 501750 236721
rect 501986 236485 502154 236721
rect 501674 236401 502154 236485
rect 501674 236165 501750 236401
rect 501986 236165 502154 236401
rect 501674 236081 502154 236165
rect 501674 235845 501750 236081
rect 501986 235845 502154 236081
rect 501674 235761 502154 235845
rect 501674 235525 501750 235761
rect 501986 235525 502154 235761
rect 501674 235441 502154 235525
rect 501674 235205 501750 235441
rect 501986 235205 502154 235441
rect 501674 235121 502154 235205
rect 501674 234885 501750 235121
rect 501986 234885 502154 235121
rect 501674 234801 502154 234885
rect 501674 234565 501750 234801
rect 501986 234565 502154 234801
rect 501674 234448 502154 234565
rect 44186 233211 63160 233466
rect 44186 230735 56554 233211
rect 62870 230735 63160 233211
rect 44186 230466 63160 230735
rect 133060 233362 133516 233464
rect 133060 233126 133140 233362
rect 133376 233126 133516 233362
rect 133060 233042 133516 233126
rect 133060 232806 133140 233042
rect 133376 232806 133516 233042
rect 133060 232722 133516 232806
rect 133060 232486 133140 232722
rect 133376 232486 133516 232722
rect 133060 232402 133516 232486
rect 133060 232166 133140 232402
rect 133376 232166 133516 232402
rect 133060 232082 133516 232166
rect 133060 231846 133140 232082
rect 133376 231846 133516 232082
rect 133060 231762 133516 231846
rect 133060 231526 133140 231762
rect 133376 231526 133516 231762
rect 133060 231442 133516 231526
rect 133060 231206 133140 231442
rect 133376 231206 133516 231442
rect 133060 231122 133516 231206
rect 133060 230886 133140 231122
rect 133376 230886 133516 231122
rect 133060 230802 133516 230886
rect 133060 230566 133140 230802
rect 133376 230566 133516 230802
rect 133060 230466 133516 230566
rect 148110 233362 148566 233464
rect 148110 233126 148190 233362
rect 148426 233126 148566 233362
rect 148110 233042 148566 233126
rect 148110 232806 148190 233042
rect 148426 232806 148566 233042
rect 148110 232722 148566 232806
rect 148110 232486 148190 232722
rect 148426 232486 148566 232722
rect 148110 232402 148566 232486
rect 148110 232166 148190 232402
rect 148426 232166 148566 232402
rect 148110 232082 148566 232166
rect 148110 231846 148190 232082
rect 148426 231846 148566 232082
rect 148110 231762 148566 231846
rect 148110 231526 148190 231762
rect 148426 231526 148566 231762
rect 148110 231442 148566 231526
rect 148110 231206 148190 231442
rect 148426 231206 148566 231442
rect 148110 231122 148566 231206
rect 148110 230886 148190 231122
rect 148426 230886 148566 231122
rect 148110 230802 148566 230886
rect 148110 230566 148190 230802
rect 148426 230566 148566 230802
rect 148110 230466 148566 230566
rect 163160 233362 163616 233464
rect 163160 233126 163240 233362
rect 163476 233126 163616 233362
rect 163160 233042 163616 233126
rect 163160 232806 163240 233042
rect 163476 232806 163616 233042
rect 163160 232722 163616 232806
rect 163160 232486 163240 232722
rect 163476 232486 163616 232722
rect 163160 232402 163616 232486
rect 163160 232166 163240 232402
rect 163476 232166 163616 232402
rect 163160 232082 163616 232166
rect 163160 231846 163240 232082
rect 163476 231846 163616 232082
rect 163160 231762 163616 231846
rect 163160 231526 163240 231762
rect 163476 231526 163616 231762
rect 163160 231442 163616 231526
rect 163160 231206 163240 231442
rect 163476 231206 163616 231442
rect 163160 231122 163616 231206
rect 163160 230886 163240 231122
rect 163476 230886 163616 231122
rect 163160 230802 163616 230886
rect 163160 230566 163240 230802
rect 163476 230566 163616 230802
rect 163160 230466 163616 230566
rect 178210 233362 178666 233464
rect 178210 233126 178290 233362
rect 178526 233126 178666 233362
rect 178210 233042 178666 233126
rect 178210 232806 178290 233042
rect 178526 232806 178666 233042
rect 178210 232722 178666 232806
rect 178210 232486 178290 232722
rect 178526 232486 178666 232722
rect 178210 232402 178666 232486
rect 178210 232166 178290 232402
rect 178526 232166 178666 232402
rect 178210 232082 178666 232166
rect 178210 231846 178290 232082
rect 178526 231846 178666 232082
rect 178210 231762 178666 231846
rect 178210 231526 178290 231762
rect 178526 231526 178666 231762
rect 178210 231442 178666 231526
rect 178210 231206 178290 231442
rect 178526 231206 178666 231442
rect 178210 231122 178666 231206
rect 178210 230886 178290 231122
rect 178526 230886 178666 231122
rect 178210 230802 178666 230886
rect 178210 230566 178290 230802
rect 178526 230566 178666 230802
rect 178210 230466 178666 230566
rect 193260 233362 193716 233464
rect 193260 233126 193340 233362
rect 193576 233126 193716 233362
rect 193260 233042 193716 233126
rect 193260 232806 193340 233042
rect 193576 232806 193716 233042
rect 193260 232722 193716 232806
rect 193260 232486 193340 232722
rect 193576 232486 193716 232722
rect 193260 232402 193716 232486
rect 193260 232166 193340 232402
rect 193576 232166 193716 232402
rect 193260 232082 193716 232166
rect 193260 231846 193340 232082
rect 193576 231846 193716 232082
rect 193260 231762 193716 231846
rect 193260 231526 193340 231762
rect 193576 231526 193716 231762
rect 193260 231442 193716 231526
rect 193260 231206 193340 231442
rect 193576 231206 193716 231442
rect 193260 231122 193716 231206
rect 193260 230886 193340 231122
rect 193576 230886 193716 231122
rect 193260 230802 193716 230886
rect 193260 230566 193340 230802
rect 193576 230566 193716 230802
rect 193260 230466 193716 230566
rect 208310 233362 208766 233464
rect 208310 233126 208390 233362
rect 208626 233126 208766 233362
rect 208310 233042 208766 233126
rect 208310 232806 208390 233042
rect 208626 232806 208766 233042
rect 208310 232722 208766 232806
rect 208310 232486 208390 232722
rect 208626 232486 208766 232722
rect 208310 232402 208766 232486
rect 208310 232166 208390 232402
rect 208626 232166 208766 232402
rect 208310 232082 208766 232166
rect 208310 231846 208390 232082
rect 208626 231846 208766 232082
rect 208310 231762 208766 231846
rect 208310 231526 208390 231762
rect 208626 231526 208766 231762
rect 208310 231442 208766 231526
rect 208310 231206 208390 231442
rect 208626 231206 208766 231442
rect 208310 231122 208766 231206
rect 208310 230886 208390 231122
rect 208626 230886 208766 231122
rect 208310 230802 208766 230886
rect 208310 230566 208390 230802
rect 208626 230566 208766 230802
rect 208310 230466 208766 230566
rect 223360 233362 223816 233464
rect 223360 233126 223440 233362
rect 223676 233126 223816 233362
rect 223360 233042 223816 233126
rect 223360 232806 223440 233042
rect 223676 232806 223816 233042
rect 223360 232722 223816 232806
rect 223360 232486 223440 232722
rect 223676 232486 223816 232722
rect 223360 232402 223816 232486
rect 223360 232166 223440 232402
rect 223676 232166 223816 232402
rect 223360 232082 223816 232166
rect 223360 231846 223440 232082
rect 223676 231846 223816 232082
rect 223360 231762 223816 231846
rect 223360 231526 223440 231762
rect 223676 231526 223816 231762
rect 223360 231442 223816 231526
rect 223360 231206 223440 231442
rect 223676 231206 223816 231442
rect 223360 231122 223816 231206
rect 223360 230886 223440 231122
rect 223676 230886 223816 231122
rect 223360 230802 223816 230886
rect 223360 230566 223440 230802
rect 223676 230566 223816 230802
rect 223360 230466 223816 230566
rect 238410 233362 238866 233464
rect 238410 233126 238490 233362
rect 238726 233126 238866 233362
rect 238410 233042 238866 233126
rect 238410 232806 238490 233042
rect 238726 232806 238866 233042
rect 238410 232722 238866 232806
rect 238410 232486 238490 232722
rect 238726 232486 238866 232722
rect 238410 232402 238866 232486
rect 238410 232166 238490 232402
rect 238726 232166 238866 232402
rect 238410 232082 238866 232166
rect 238410 231846 238490 232082
rect 238726 231846 238866 232082
rect 238410 231762 238866 231846
rect 238410 231526 238490 231762
rect 238726 231526 238866 231762
rect 238410 231442 238866 231526
rect 238410 231206 238490 231442
rect 238726 231206 238866 231442
rect 238410 231122 238866 231206
rect 238410 230886 238490 231122
rect 238726 230886 238866 231122
rect 238410 230802 238866 230886
rect 238410 230566 238490 230802
rect 238726 230566 238866 230802
rect 238410 230466 238866 230566
rect 253460 233362 253916 233464
rect 253460 233126 253540 233362
rect 253776 233126 253916 233362
rect 253460 233042 253916 233126
rect 253460 232806 253540 233042
rect 253776 232806 253916 233042
rect 253460 232722 253916 232806
rect 253460 232486 253540 232722
rect 253776 232486 253916 232722
rect 253460 232402 253916 232486
rect 253460 232166 253540 232402
rect 253776 232166 253916 232402
rect 253460 232082 253916 232166
rect 253460 231846 253540 232082
rect 253776 231846 253916 232082
rect 253460 231762 253916 231846
rect 253460 231526 253540 231762
rect 253776 231526 253916 231762
rect 253460 231442 253916 231526
rect 253460 231206 253540 231442
rect 253776 231206 253916 231442
rect 253460 231122 253916 231206
rect 253460 230886 253540 231122
rect 253776 230886 253916 231122
rect 253460 230802 253916 230886
rect 253460 230566 253540 230802
rect 253776 230566 253916 230802
rect 253460 230466 253916 230566
rect 268510 233362 268966 233464
rect 268510 233126 268590 233362
rect 268826 233126 268966 233362
rect 268510 233042 268966 233126
rect 268510 232806 268590 233042
rect 268826 232806 268966 233042
rect 268510 232722 268966 232806
rect 268510 232486 268590 232722
rect 268826 232486 268966 232722
rect 268510 232402 268966 232486
rect 268510 232166 268590 232402
rect 268826 232166 268966 232402
rect 268510 232082 268966 232166
rect 268510 231846 268590 232082
rect 268826 231846 268966 232082
rect 268510 231762 268966 231846
rect 268510 231526 268590 231762
rect 268826 231526 268966 231762
rect 268510 231442 268966 231526
rect 268510 231206 268590 231442
rect 268826 231206 268966 231442
rect 268510 231122 268966 231206
rect 268510 230886 268590 231122
rect 268826 230886 268966 231122
rect 268510 230802 268966 230886
rect 268510 230566 268590 230802
rect 268826 230566 268966 230802
rect 268510 230466 268966 230566
rect 283560 233362 284016 233464
rect 283560 233126 283640 233362
rect 283876 233126 284016 233362
rect 283560 233042 284016 233126
rect 283560 232806 283640 233042
rect 283876 232806 284016 233042
rect 283560 232722 284016 232806
rect 283560 232486 283640 232722
rect 283876 232486 284016 232722
rect 283560 232402 284016 232486
rect 283560 232166 283640 232402
rect 283876 232166 284016 232402
rect 283560 232082 284016 232166
rect 283560 231846 283640 232082
rect 283876 231846 284016 232082
rect 283560 231762 284016 231846
rect 283560 231526 283640 231762
rect 283876 231526 284016 231762
rect 283560 231442 284016 231526
rect 283560 231206 283640 231442
rect 283876 231206 284016 231442
rect 283560 231122 284016 231206
rect 283560 230886 283640 231122
rect 283876 230886 284016 231122
rect 283560 230802 284016 230886
rect 283560 230566 283640 230802
rect 283876 230566 284016 230802
rect 283560 230466 284016 230566
rect 298610 233362 299066 233464
rect 298610 233126 298690 233362
rect 298926 233126 299066 233362
rect 298610 233042 299066 233126
rect 298610 232806 298690 233042
rect 298926 232806 299066 233042
rect 298610 232722 299066 232806
rect 298610 232486 298690 232722
rect 298926 232486 299066 232722
rect 298610 232402 299066 232486
rect 298610 232166 298690 232402
rect 298926 232166 299066 232402
rect 298610 232082 299066 232166
rect 298610 231846 298690 232082
rect 298926 231846 299066 232082
rect 298610 231762 299066 231846
rect 298610 231526 298690 231762
rect 298926 231526 299066 231762
rect 298610 231442 299066 231526
rect 298610 231206 298690 231442
rect 298926 231206 299066 231442
rect 298610 231122 299066 231206
rect 298610 230886 298690 231122
rect 298926 230886 299066 231122
rect 298610 230802 299066 230886
rect 298610 230566 298690 230802
rect 298926 230566 299066 230802
rect 298610 230466 299066 230566
rect 313660 233362 314116 233464
rect 313660 233126 313740 233362
rect 313976 233126 314116 233362
rect 313660 233042 314116 233126
rect 313660 232806 313740 233042
rect 313976 232806 314116 233042
rect 313660 232722 314116 232806
rect 313660 232486 313740 232722
rect 313976 232486 314116 232722
rect 313660 232402 314116 232486
rect 313660 232166 313740 232402
rect 313976 232166 314116 232402
rect 313660 232082 314116 232166
rect 313660 231846 313740 232082
rect 313976 231846 314116 232082
rect 313660 231762 314116 231846
rect 313660 231526 313740 231762
rect 313976 231526 314116 231762
rect 313660 231442 314116 231526
rect 313660 231206 313740 231442
rect 313976 231206 314116 231442
rect 313660 231122 314116 231206
rect 313660 230886 313740 231122
rect 313976 230886 314116 231122
rect 313660 230802 314116 230886
rect 313660 230566 313740 230802
rect 313976 230566 314116 230802
rect 313660 230466 314116 230566
rect 328710 233362 329166 233464
rect 328710 233126 328790 233362
rect 329026 233126 329166 233362
rect 328710 233042 329166 233126
rect 328710 232806 328790 233042
rect 329026 232806 329166 233042
rect 328710 232722 329166 232806
rect 328710 232486 328790 232722
rect 329026 232486 329166 232722
rect 328710 232402 329166 232486
rect 328710 232166 328790 232402
rect 329026 232166 329166 232402
rect 328710 232082 329166 232166
rect 328710 231846 328790 232082
rect 329026 231846 329166 232082
rect 328710 231762 329166 231846
rect 328710 231526 328790 231762
rect 329026 231526 329166 231762
rect 328710 231442 329166 231526
rect 328710 231206 328790 231442
rect 329026 231206 329166 231442
rect 328710 231122 329166 231206
rect 328710 230886 328790 231122
rect 329026 230886 329166 231122
rect 328710 230802 329166 230886
rect 328710 230566 328790 230802
rect 329026 230566 329166 230802
rect 328710 230466 329166 230566
rect 343760 233362 344216 233464
rect 343760 233126 343840 233362
rect 344076 233126 344216 233362
rect 343760 233042 344216 233126
rect 343760 232806 343840 233042
rect 344076 232806 344216 233042
rect 343760 232722 344216 232806
rect 343760 232486 343840 232722
rect 344076 232486 344216 232722
rect 343760 232402 344216 232486
rect 343760 232166 343840 232402
rect 344076 232166 344216 232402
rect 343760 232082 344216 232166
rect 343760 231846 343840 232082
rect 344076 231846 344216 232082
rect 343760 231762 344216 231846
rect 343760 231526 343840 231762
rect 344076 231526 344216 231762
rect 343760 231442 344216 231526
rect 343760 231206 343840 231442
rect 344076 231206 344216 231442
rect 343760 231122 344216 231206
rect 343760 230886 343840 231122
rect 344076 230886 344216 231122
rect 343760 230802 344216 230886
rect 343760 230566 343840 230802
rect 344076 230566 344216 230802
rect 343760 230466 344216 230566
rect 358810 233362 359266 233464
rect 358810 233126 358890 233362
rect 359126 233126 359266 233362
rect 358810 233042 359266 233126
rect 358810 232806 358890 233042
rect 359126 232806 359266 233042
rect 358810 232722 359266 232806
rect 358810 232486 358890 232722
rect 359126 232486 359266 232722
rect 358810 232402 359266 232486
rect 358810 232166 358890 232402
rect 359126 232166 359266 232402
rect 358810 232082 359266 232166
rect 358810 231846 358890 232082
rect 359126 231846 359266 232082
rect 358810 231762 359266 231846
rect 358810 231526 358890 231762
rect 359126 231526 359266 231762
rect 358810 231442 359266 231526
rect 358810 231206 358890 231442
rect 359126 231206 359266 231442
rect 358810 231122 359266 231206
rect 358810 230886 358890 231122
rect 359126 230886 359266 231122
rect 358810 230802 359266 230886
rect 358810 230566 358890 230802
rect 359126 230566 359266 230802
rect 358810 230466 359266 230566
rect 373860 233362 374316 233464
rect 373860 233126 373940 233362
rect 374176 233126 374316 233362
rect 373860 233042 374316 233126
rect 373860 232806 373940 233042
rect 374176 232806 374316 233042
rect 373860 232722 374316 232806
rect 373860 232486 373940 232722
rect 374176 232486 374316 232722
rect 373860 232402 374316 232486
rect 373860 232166 373940 232402
rect 374176 232166 374316 232402
rect 373860 232082 374316 232166
rect 373860 231846 373940 232082
rect 374176 231846 374316 232082
rect 373860 231762 374316 231846
rect 373860 231526 373940 231762
rect 374176 231526 374316 231762
rect 373860 231442 374316 231526
rect 373860 231206 373940 231442
rect 374176 231206 374316 231442
rect 373860 231122 374316 231206
rect 373860 230886 373940 231122
rect 374176 230886 374316 231122
rect 373860 230802 374316 230886
rect 373860 230566 373940 230802
rect 374176 230566 374316 230802
rect 373860 230466 374316 230566
rect 388910 233362 389366 233464
rect 388910 233126 388990 233362
rect 389226 233126 389366 233362
rect 388910 233042 389366 233126
rect 388910 232806 388990 233042
rect 389226 232806 389366 233042
rect 388910 232722 389366 232806
rect 388910 232486 388990 232722
rect 389226 232486 389366 232722
rect 388910 232402 389366 232486
rect 388910 232166 388990 232402
rect 389226 232166 389366 232402
rect 388910 232082 389366 232166
rect 388910 231846 388990 232082
rect 389226 231846 389366 232082
rect 388910 231762 389366 231846
rect 388910 231526 388990 231762
rect 389226 231526 389366 231762
rect 388910 231442 389366 231526
rect 388910 231206 388990 231442
rect 389226 231206 389366 231442
rect 388910 231122 389366 231206
rect 388910 230886 388990 231122
rect 389226 230886 389366 231122
rect 388910 230802 389366 230886
rect 388910 230566 388990 230802
rect 389226 230566 389366 230802
rect 388910 230466 389366 230566
rect 403960 233362 404416 233464
rect 403960 233126 404040 233362
rect 404276 233126 404416 233362
rect 403960 233042 404416 233126
rect 403960 232806 404040 233042
rect 404276 232806 404416 233042
rect 403960 232722 404416 232806
rect 403960 232486 404040 232722
rect 404276 232486 404416 232722
rect 403960 232402 404416 232486
rect 403960 232166 404040 232402
rect 404276 232166 404416 232402
rect 403960 232082 404416 232166
rect 403960 231846 404040 232082
rect 404276 231846 404416 232082
rect 403960 231762 404416 231846
rect 403960 231526 404040 231762
rect 404276 231526 404416 231762
rect 403960 231442 404416 231526
rect 403960 231206 404040 231442
rect 404276 231206 404416 231442
rect 403960 231122 404416 231206
rect 403960 230886 404040 231122
rect 404276 230886 404416 231122
rect 403960 230802 404416 230886
rect 403960 230566 404040 230802
rect 404276 230566 404416 230802
rect 403960 230466 404416 230566
rect 419010 233362 419466 233464
rect 419010 233126 419090 233362
rect 419326 233126 419466 233362
rect 419010 233042 419466 233126
rect 419010 232806 419090 233042
rect 419326 232806 419466 233042
rect 419010 232722 419466 232806
rect 419010 232486 419090 232722
rect 419326 232486 419466 232722
rect 419010 232402 419466 232486
rect 419010 232166 419090 232402
rect 419326 232166 419466 232402
rect 419010 232082 419466 232166
rect 419010 231846 419090 232082
rect 419326 231846 419466 232082
rect 419010 231762 419466 231846
rect 419010 231526 419090 231762
rect 419326 231526 419466 231762
rect 419010 231442 419466 231526
rect 419010 231206 419090 231442
rect 419326 231206 419466 231442
rect 419010 231122 419466 231206
rect 419010 230886 419090 231122
rect 419326 230886 419466 231122
rect 419010 230802 419466 230886
rect 419010 230566 419090 230802
rect 419326 230566 419466 230802
rect 419010 230466 419466 230566
rect 434060 233362 434516 233464
rect 434060 233126 434140 233362
rect 434376 233126 434516 233362
rect 434060 233042 434516 233126
rect 434060 232806 434140 233042
rect 434376 232806 434516 233042
rect 434060 232722 434516 232806
rect 434060 232486 434140 232722
rect 434376 232486 434516 232722
rect 434060 232402 434516 232486
rect 434060 232166 434140 232402
rect 434376 232166 434516 232402
rect 434060 232082 434516 232166
rect 434060 231846 434140 232082
rect 434376 231846 434516 232082
rect 434060 231762 434516 231846
rect 434060 231526 434140 231762
rect 434376 231526 434516 231762
rect 434060 231442 434516 231526
rect 434060 231206 434140 231442
rect 434376 231206 434516 231442
rect 434060 231122 434516 231206
rect 434060 230886 434140 231122
rect 434376 230886 434516 231122
rect 434060 230802 434516 230886
rect 434060 230566 434140 230802
rect 434376 230566 434516 230802
rect 434060 230466 434516 230566
rect 449110 233362 449566 233464
rect 449110 233126 449190 233362
rect 449426 233126 449566 233362
rect 449110 233042 449566 233126
rect 449110 232806 449190 233042
rect 449426 232806 449566 233042
rect 449110 232722 449566 232806
rect 449110 232486 449190 232722
rect 449426 232486 449566 232722
rect 449110 232402 449566 232486
rect 449110 232166 449190 232402
rect 449426 232166 449566 232402
rect 449110 232082 449566 232166
rect 449110 231846 449190 232082
rect 449426 231846 449566 232082
rect 449110 231762 449566 231846
rect 449110 231526 449190 231762
rect 449426 231526 449566 231762
rect 449110 231442 449566 231526
rect 449110 231206 449190 231442
rect 449426 231206 449566 231442
rect 449110 231122 449566 231206
rect 449110 230886 449190 231122
rect 449426 230886 449566 231122
rect 449110 230802 449566 230886
rect 449110 230566 449190 230802
rect 449426 230566 449566 230802
rect 449110 230466 449566 230566
rect 464160 233362 464616 233464
rect 464160 233126 464240 233362
rect 464476 233126 464616 233362
rect 464160 233042 464616 233126
rect 464160 232806 464240 233042
rect 464476 232806 464616 233042
rect 464160 232722 464616 232806
rect 464160 232486 464240 232722
rect 464476 232486 464616 232722
rect 464160 232402 464616 232486
rect 464160 232166 464240 232402
rect 464476 232166 464616 232402
rect 464160 232082 464616 232166
rect 464160 231846 464240 232082
rect 464476 231846 464616 232082
rect 464160 231762 464616 231846
rect 464160 231526 464240 231762
rect 464476 231526 464616 231762
rect 464160 231442 464616 231526
rect 464160 231206 464240 231442
rect 464476 231206 464616 231442
rect 464160 231122 464616 231206
rect 464160 230886 464240 231122
rect 464476 230886 464616 231122
rect 464160 230802 464616 230886
rect 464160 230566 464240 230802
rect 464476 230566 464616 230802
rect 464160 230466 464616 230566
rect 479210 233362 479666 233464
rect 479210 233126 479290 233362
rect 479526 233126 479666 233362
rect 479210 233042 479666 233126
rect 479210 232806 479290 233042
rect 479526 232806 479666 233042
rect 479210 232722 479666 232806
rect 479210 232486 479290 232722
rect 479526 232486 479666 232722
rect 479210 232402 479666 232486
rect 479210 232166 479290 232402
rect 479526 232166 479666 232402
rect 479210 232082 479666 232166
rect 479210 231846 479290 232082
rect 479526 231846 479666 232082
rect 479210 231762 479666 231846
rect 479210 231526 479290 231762
rect 479526 231526 479666 231762
rect 479210 231442 479666 231526
rect 479210 231206 479290 231442
rect 479526 231206 479666 231442
rect 479210 231122 479666 231206
rect 479210 230886 479290 231122
rect 479526 230886 479666 231122
rect 479210 230802 479666 230886
rect 479210 230566 479290 230802
rect 479526 230566 479666 230802
rect 479210 230466 479666 230566
rect 494260 233362 494716 233464
rect 494260 233126 494340 233362
rect 494576 233126 494716 233362
rect 494260 233042 494716 233126
rect 494260 232806 494340 233042
rect 494576 232806 494716 233042
rect 494260 232722 494716 232806
rect 494260 232486 494340 232722
rect 494576 232486 494716 232722
rect 494260 232402 494716 232486
rect 494260 232166 494340 232402
rect 494576 232166 494716 232402
rect 494260 232082 494716 232166
rect 494260 231846 494340 232082
rect 494576 231846 494716 232082
rect 494260 231762 494716 231846
rect 494260 231526 494340 231762
rect 494576 231526 494716 231762
rect 494260 231442 494716 231526
rect 494260 231206 494340 231442
rect 494576 231206 494716 231442
rect 494260 231122 494716 231206
rect 494260 230886 494340 231122
rect 494576 230886 494716 231122
rect 494260 230802 494716 230886
rect 494260 230566 494340 230802
rect 494576 230566 494716 230802
rect 494260 230466 494716 230566
rect 44198 197498 46798 230466
rect 584368 212271 596962 212504
rect 584368 209795 584610 212271
rect 587086 209795 593464 212271
rect 595940 209795 596962 212271
rect 584368 209504 596962 209795
rect 627044 212234 628108 212460
rect 627044 209758 627303 212234
rect 627859 209758 628108 212234
rect 627044 209528 628108 209758
rect 582262 208302 591388 208502
rect 582262 208066 582400 208302
rect 582636 208066 582720 208302
rect 582956 208066 583040 208302
rect 583276 208066 583360 208302
rect 583596 208066 588493 208302
rect 588729 208066 588813 208302
rect 589049 208066 589133 208302
rect 589369 208066 589453 208302
rect 589689 208066 589773 208302
rect 590009 208066 590093 208302
rect 590329 208066 590413 208302
rect 590649 208066 590733 208302
rect 590969 208066 591053 208302
rect 591289 208066 591388 208302
rect 582262 207862 591388 208066
rect 596642 207692 596962 209504
rect 627362 207684 627682 209528
rect 584496 197721 587174 197876
rect 44198 197312 52344 197498
rect 44198 197076 51573 197312
rect 51809 197076 51893 197312
rect 52129 197076 52344 197312
rect 44198 196858 52344 197076
rect 584496 197165 584783 197721
rect 586939 197528 587174 197721
rect 586939 197483 592976 197528
rect 586939 197247 592038 197483
rect 592274 197247 592358 197483
rect 592594 197247 592678 197483
rect 592914 197247 592976 197483
rect 586939 197208 592976 197247
rect 586939 197165 587174 197208
rect 584496 196992 587174 197165
rect 44198 176742 46798 196858
rect 582072 184290 591388 184502
rect 582072 184054 582204 184290
rect 582440 184054 582524 184290
rect 582760 184286 591388 184290
rect 582760 184054 588493 184286
rect 582072 184050 588493 184054
rect 588729 184050 588813 184286
rect 589049 184050 589133 184286
rect 589369 184050 589453 184286
rect 589689 184050 589773 184286
rect 590009 184050 590093 184286
rect 590329 184050 590413 184286
rect 590649 184050 590733 184286
rect 590969 184050 591053 184286
rect 591289 184050 591388 184286
rect 582072 183862 591388 184050
rect 41864 176505 46798 176742
rect 41864 173389 42087 176505
rect 45523 173389 46798 176505
rect 41864 173126 46798 173389
rect 42646 171298 52246 171498
rect 42646 171294 51465 171298
rect 42646 171058 42857 171294
rect 43093 171058 43177 171294
rect 43413 171058 43497 171294
rect 43733 171058 43817 171294
rect 44053 171058 44137 171294
rect 44373 171058 44457 171294
rect 44693 171058 44777 171294
rect 45013 171058 45097 171294
rect 45333 171058 45417 171294
rect 45653 171062 51465 171294
rect 51701 171062 51785 171298
rect 52021 171062 52246 171298
rect 45653 171058 52246 171062
rect 42646 170858 52246 171058
rect 584496 167081 587174 167236
rect 584496 166525 584783 167081
rect 586939 166892 587174 167081
rect 586939 166855 592976 166892
rect 586939 166619 592021 166855
rect 592257 166619 592341 166855
rect 592577 166619 592661 166855
rect 592897 166619 592976 166855
rect 586939 166572 592976 166619
rect 586939 166525 587174 166572
rect 584496 166352 587174 166525
rect 580072 158298 591388 158502
rect 580072 158294 588467 158298
rect 580072 158058 580242 158294
rect 580478 158058 580562 158294
rect 580798 158058 580882 158294
rect 581118 158058 581202 158294
rect 581438 158058 581522 158294
rect 581758 158058 581842 158294
rect 582078 158058 582162 158294
rect 582398 158058 582482 158294
rect 582718 158062 588467 158294
rect 588703 158062 588787 158298
rect 589023 158062 589107 158298
rect 589343 158062 589427 158298
rect 589663 158062 589747 158298
rect 589983 158062 590067 158298
rect 590303 158062 590387 158298
rect 590623 158062 590707 158298
rect 590943 158062 591027 158298
rect 591263 158062 591388 158298
rect 582718 158058 591388 158062
rect 580072 157862 591388 158058
rect 42578 145300 52178 145498
rect 42578 145064 42871 145300
rect 43107 145064 43191 145300
rect 43427 145064 43511 145300
rect 43747 145064 43831 145300
rect 44067 145064 44151 145300
rect 44387 145064 44471 145300
rect 44707 145064 44791 145300
rect 45027 145064 45111 145300
rect 45347 145064 45431 145300
rect 45667 145290 52178 145300
rect 45667 145064 51399 145290
rect 42578 145054 51399 145064
rect 51635 145054 51719 145290
rect 51955 145054 52178 145290
rect 42578 144858 52178 145054
rect 584496 136441 587174 136596
rect 584496 135885 584783 136441
rect 586939 136256 587174 136441
rect 586939 136215 592976 136256
rect 586939 135979 592011 136215
rect 592247 135979 592331 136215
rect 592567 135979 592651 136215
rect 592887 135979 592976 136215
rect 586939 135936 592976 135979
rect 586939 135885 587174 135936
rect 584496 135712 587174 135885
rect 580072 132288 591388 132502
rect 580072 132052 580252 132288
rect 580488 132052 580572 132288
rect 580808 132052 580892 132288
rect 581128 132052 581212 132288
rect 581448 132052 581532 132288
rect 581768 132052 581852 132288
rect 582088 132052 582172 132288
rect 582408 132052 582492 132288
rect 582728 132282 591388 132288
rect 582728 132052 588493 132282
rect 580072 132046 588493 132052
rect 588729 132046 588813 132282
rect 589049 132046 589133 132282
rect 589369 132046 589453 132282
rect 589689 132046 589773 132282
rect 590009 132046 590093 132282
rect 590329 132046 590413 132282
rect 590649 132046 590733 132282
rect 590969 132046 591053 132282
rect 591289 132046 591388 132282
rect 580072 131862 591388 132046
rect 42578 119296 52178 119498
rect 42578 119060 42861 119296
rect 43097 119060 43181 119296
rect 43417 119060 43501 119296
rect 43737 119060 43821 119296
rect 44057 119060 44141 119296
rect 44377 119060 44461 119296
rect 44697 119060 44781 119296
rect 45017 119060 45101 119296
rect 45337 119060 45421 119296
rect 45657 119060 51395 119296
rect 51631 119060 51715 119296
rect 51951 119060 52178 119296
rect 42578 118858 52178 119060
rect 580072 106294 591388 106502
rect 580072 106058 580254 106294
rect 580490 106058 580574 106294
rect 580810 106058 580894 106294
rect 581130 106058 581214 106294
rect 581450 106058 581534 106294
rect 581770 106058 581854 106294
rect 582090 106058 582174 106294
rect 582410 106058 582494 106294
rect 582730 106058 588497 106294
rect 588733 106058 588817 106294
rect 589053 106058 589137 106294
rect 589373 106058 589457 106294
rect 589693 106058 589777 106294
rect 590013 106058 590097 106294
rect 590333 106058 590417 106294
rect 590653 106058 590737 106294
rect 590973 106058 591057 106294
rect 591293 106058 591388 106294
rect 580072 105862 591388 106058
rect 584496 105620 587174 105676
rect 584496 105578 592976 105620
rect 584496 105521 592023 105578
rect 584496 104965 584783 105521
rect 586939 105342 592023 105521
rect 592259 105342 592343 105578
rect 592579 105342 592663 105578
rect 592899 105342 592976 105578
rect 586939 105300 592976 105342
rect 586939 104965 587174 105300
rect 584496 104792 587174 104965
rect 597302 98760 597622 102316
rect 628022 98804 628342 102238
rect 596742 98603 598152 98760
rect 596742 96127 597012 98603
rect 597888 96127 598152 98603
rect 596742 95956 598152 96127
rect 627584 98665 628902 98804
rect 627584 96189 627823 98665
rect 628699 96189 628902 98665
rect 636080 98521 636994 98758
rect 636080 96685 636259 98521
rect 636815 96685 636994 98521
rect 636080 96434 636994 96685
rect 627584 96050 628902 96189
rect 636354 94448 636674 96434
rect 42578 93294 52178 93498
rect 42578 93058 42857 93294
rect 43093 93058 43177 93294
rect 43413 93058 43497 93294
rect 43733 93058 43817 93294
rect 44053 93058 44137 93294
rect 44373 93058 44457 93294
rect 44693 93058 44777 93294
rect 45013 93058 45097 93294
rect 45333 93058 45417 93294
rect 45653 93292 52178 93294
rect 45653 93058 51399 93292
rect 42578 93056 51399 93058
rect 51635 93056 51719 93292
rect 51955 93056 52178 93292
rect 42578 92858 52178 93056
rect 41864 82706 45778 82794
rect 41864 78242 41977 82706
rect 45641 78242 45778 82706
rect 632354 80924 632674 82062
rect 640354 81016 640674 82000
rect 632072 80629 633010 80924
rect 580072 80306 591388 80502
rect 580072 80304 588491 80306
rect 580072 80068 580248 80304
rect 580484 80068 580568 80304
rect 580804 80068 580888 80304
rect 581124 80068 581208 80304
rect 581444 80068 581528 80304
rect 581764 80068 581848 80304
rect 582084 80068 582168 80304
rect 582404 80068 582488 80304
rect 582724 80070 588491 80304
rect 588727 80070 588811 80306
rect 589047 80070 589131 80306
rect 589367 80070 589451 80306
rect 589687 80070 589771 80306
rect 590007 80070 590091 80306
rect 590327 80070 590411 80306
rect 590647 80070 590731 80306
rect 590967 80070 591051 80306
rect 591287 80070 591388 80306
rect 582724 80068 591388 80070
rect 580072 79862 591388 80068
rect 41864 78154 45778 78242
rect 632072 78473 632254 80629
rect 632810 78473 633010 80629
rect 632072 78198 633010 78473
rect 640098 80816 640922 81016
rect 640098 78340 640232 80816
rect 640788 78340 640922 80816
rect 640098 78134 640922 78340
rect 629888 77193 630208 77374
rect 629888 76957 629919 77193
rect 630155 76957 630208 77193
rect 629888 76873 630208 76957
rect 629888 76637 629919 76873
rect 630155 76637 630208 76873
rect 629888 76553 630208 76637
rect 629888 76317 629919 76553
rect 630155 76317 630208 76553
rect 629888 74104 630208 76317
rect 631438 75791 631758 77374
rect 631438 75555 631471 75791
rect 631707 75555 631758 75791
rect 631438 75471 631758 75555
rect 631438 75235 631471 75471
rect 631707 75235 631758 75471
rect 631438 75151 631758 75235
rect 631438 74915 631471 75151
rect 631707 74915 631758 75151
rect 631438 74104 631758 74915
rect 632988 77207 633308 77374
rect 632988 76971 633031 77207
rect 633267 76971 633308 77207
rect 632988 76887 633308 76971
rect 632988 76651 633031 76887
rect 633267 76651 633308 76887
rect 632988 76567 633308 76651
rect 632988 76331 633031 76567
rect 633267 76331 633308 76567
rect 632988 74104 633308 76331
rect 634538 75795 634858 77374
rect 634538 75559 634565 75795
rect 634801 75559 634858 75795
rect 634538 75475 634858 75559
rect 634538 75239 634565 75475
rect 634801 75239 634858 75475
rect 634538 75155 634858 75239
rect 634538 74919 634565 75155
rect 634801 74919 634858 75155
rect 634538 74104 634858 74919
rect 636088 77203 636408 77374
rect 636088 76967 636121 77203
rect 636357 76967 636408 77203
rect 636088 76883 636408 76967
rect 636088 76647 636121 76883
rect 636357 76647 636408 76883
rect 636088 76563 636408 76647
rect 636088 76327 636121 76563
rect 636357 76327 636408 76563
rect 636088 74104 636408 76327
rect 637638 75799 637958 77374
rect 637638 75563 637673 75799
rect 637909 75563 637958 75799
rect 637638 75479 637958 75563
rect 637638 75243 637673 75479
rect 637909 75243 637958 75479
rect 637638 75159 637958 75243
rect 637638 74923 637673 75159
rect 637909 74923 637958 75159
rect 637638 74104 637958 74923
rect 639188 77203 639508 77374
rect 639188 76967 639215 77203
rect 639451 76967 639508 77203
rect 639188 76883 639508 76967
rect 639188 76647 639215 76883
rect 639451 76647 639508 76883
rect 639188 76563 639508 76647
rect 639188 76327 639215 76563
rect 639451 76327 639508 76563
rect 639188 74104 639508 76327
rect 640738 75791 641058 77374
rect 640738 75555 640777 75791
rect 641013 75555 641058 75791
rect 640738 75471 641058 75555
rect 640738 75235 640777 75471
rect 641013 75235 641058 75471
rect 640738 75151 641058 75235
rect 640738 74915 640777 75151
rect 641013 74915 641058 75151
rect 640738 74104 641058 74915
rect 642288 77215 642608 77374
rect 642288 76979 642323 77215
rect 642559 76979 642608 77215
rect 642288 76895 642608 76979
rect 642288 76659 642323 76895
rect 642559 76659 642608 76895
rect 642288 76575 642608 76659
rect 642288 76339 642323 76575
rect 642559 76339 642608 76575
rect 642288 74104 642608 76339
rect 643838 75817 644158 77374
rect 643838 75581 643879 75817
rect 644115 75581 644158 75817
rect 643838 75497 644158 75581
rect 643838 75261 643879 75497
rect 644115 75261 644158 75497
rect 643838 75177 644158 75261
rect 643838 74941 643879 75177
rect 644115 74941 644158 75177
rect 643838 74104 644158 74941
rect 41858 72802 45772 72890
rect 41858 68338 41953 72802
rect 45617 68338 45772 72802
rect 41858 68250 45772 68338
rect 41862 67294 52362 67498
rect 41862 67288 51597 67294
rect 41862 67052 42095 67288
rect 42331 67052 42415 67288
rect 42651 67052 42735 67288
rect 42971 67052 43055 67288
rect 43291 67052 43375 67288
rect 43611 67052 43695 67288
rect 43931 67052 44015 67288
rect 44251 67052 44335 67288
rect 44571 67052 44655 67288
rect 44891 67052 44975 67288
rect 45211 67052 45295 67288
rect 45531 67058 51597 67288
rect 51833 67058 51917 67294
rect 52153 67058 52362 67294
rect 45531 67052 52362 67058
rect 41862 66858 52362 67052
rect 41874 51914 58536 52122
rect 41874 48478 42080 51914
rect 45516 51880 58536 51914
rect 45516 48478 54650 51880
rect 41874 48444 54650 48478
rect 58086 48444 58536 51880
rect 143324 50592 144738 50688
rect 143324 50036 143423 50592
rect 144619 50036 144738 50592
rect 143324 49936 144738 50036
rect 143860 49638 144040 49936
rect 41874 48222 58536 48444
rect 641936 47627 650202 48027
rect 142560 45396 142740 47256
rect 141776 45394 142866 45396
rect 141376 45194 142866 45394
rect 141376 44318 141528 45194
rect 142724 44318 142866 45194
rect 141376 44130 142866 44318
rect 143440 40762 143620 47296
rect 144740 41158 144920 47340
rect 241680 46607 246056 46692
rect 241680 46601 241825 46607
rect 245901 46601 246056 46607
rect 241680 42857 241751 46601
rect 245975 42857 246056 46601
rect 241680 42851 241825 42857
rect 245901 42851 246056 42857
rect 241680 42784 246056 42851
rect 251302 46621 255700 46684
rect 251302 46615 251477 46621
rect 255553 46615 255700 46621
rect 251302 42871 251403 46615
rect 255627 42871 255700 46615
rect 251302 42865 251477 42871
rect 255553 42865 255700 42871
rect 251302 42788 255700 42865
rect 641936 43965 643718 47627
rect 661270 47274 669426 47320
rect 648104 47124 649670 47188
rect 648104 46660 648175 47124
rect 649599 46660 649670 47124
rect 648104 46590 649670 46660
rect 641936 42221 641995 43965
rect 643659 42221 643718 43965
rect 653432 45022 656912 47054
rect 661270 47038 666522 47274
rect 666758 47038 666842 47274
rect 667078 47038 667162 47274
rect 667398 47038 667482 47274
rect 667718 47038 667802 47274
rect 668038 47038 668122 47274
rect 668358 47038 668442 47274
rect 668678 47038 668762 47274
rect 668998 47038 669082 47274
rect 669318 47038 669426 47274
rect 661270 46991 669426 47038
rect 653432 42638 653583 45022
rect 656767 42638 656912 45022
rect 653432 42488 656912 42638
rect 641936 42164 643718 42221
rect 144740 41140 150516 41158
rect 144740 40996 149637 41140
rect 150421 40996 150516 41140
rect 144740 40978 150516 40996
rect 143440 40744 148940 40762
rect 143440 40600 148105 40744
rect 148889 40600 148940 40744
rect 143440 40582 148940 40600
rect 149632 35973 150436 35996
rect 149632 35189 149642 35973
rect 150426 35189 150436 35973
rect 149632 35166 150436 35189
rect 148098 34765 148902 34788
rect 148098 33981 148108 34765
rect 148892 33981 148902 34765
rect 642026 34726 643634 34760
rect 642026 34022 642038 34726
rect 643622 34022 643634 34726
rect 642026 33988 643634 34022
rect 148098 33958 148902 33981
<< via4 >>
rect 575875 991021 580271 993177
rect 671036 995668 676392 996544
rect 585871 991035 590267 993191
rect 671042 990364 673198 992520
rect 47874 989889 48110 990125
rect 48194 989889 48430 990125
rect 48514 989889 48750 990125
rect 48834 989889 49070 990125
rect 49154 989889 49390 990125
rect 49474 989889 49710 990125
rect 55829 989890 56065 990126
rect 56149 989890 56385 990126
rect 50280 988925 50516 989161
rect 50600 988925 50836 989161
rect 50920 988925 51156 989161
rect 51240 988925 51476 989161
rect 51560 988925 51796 989161
rect 51880 988925 52116 989161
rect 55833 988930 56069 989166
rect 56153 988930 56389 989166
rect 658577 987006 658813 987242
rect 658897 987006 659133 987242
rect 659217 987006 659453 987242
rect 659537 987006 659773 987242
rect 659857 987006 660093 987242
rect 660177 987006 660413 987242
rect 660497 987006 660733 987242
rect 660817 987006 661053 987242
rect 661137 987006 661373 987242
rect 661457 987006 661693 987242
rect 661777 987006 662013 987242
rect 662097 987006 662333 987242
rect 662417 987006 662653 987242
rect 662737 987006 662973 987242
rect 667281 987011 667517 987247
rect 667601 987011 667837 987247
rect 667921 987011 668157 987247
rect 668241 987011 668477 987247
rect 668561 987011 668797 987247
rect 668881 987011 669117 987247
rect 669201 987011 669437 987247
rect 669521 987011 669757 987247
rect 41066 985885 43542 986441
rect 55813 986043 56049 986279
rect 56133 986043 56369 986279
rect 44269 984930 46745 985486
rect 55828 984919 56384 985475
rect 52759 984121 52995 984357
rect 53079 984121 53315 984357
rect 53399 984121 53635 984357
rect 55811 983961 56367 984517
rect 658391 984120 658627 984356
rect 658711 984120 658947 984356
rect 659031 984120 659267 984356
rect 659351 984120 659587 984356
rect 659671 984120 659907 984356
rect 659991 984120 660227 984356
rect 660311 984120 660547 984356
rect 660631 984120 660867 984356
rect 660951 984120 661187 984356
rect 661271 984120 661507 984356
rect 661591 984120 661827 984356
rect 661911 984120 662147 984356
rect 662231 984120 662467 984356
rect 662551 984120 662787 984356
rect 662871 984120 663107 984356
rect 670883 983965 673359 984521
rect 658373 983164 658609 983400
rect 658693 983164 658929 983400
rect 659013 983164 659249 983400
rect 659333 983164 659569 983400
rect 659653 983164 659889 983400
rect 659973 983164 660209 983400
rect 660293 983164 660529 983400
rect 660613 983164 660849 983400
rect 660933 983164 661169 983400
rect 661253 983164 661489 983400
rect 661573 983164 661809 983400
rect 661893 983164 662129 983400
rect 662213 983164 662449 983400
rect 662533 983164 662769 983400
rect 662853 983164 663089 983400
rect 674081 983003 676557 983559
rect 44428 952065 46584 952941
rect 41218 950483 43374 951359
rect 674799 900155 675675 901031
rect 671643 898547 672519 899423
rect 674210 855146 675086 856022
rect 671666 853544 672542 854420
rect 48043 837864 49559 842260
rect 48043 827932 49559 832328
rect 667430 828720 669586 833116
rect 44428 826265 46584 827141
rect 41218 824683 43374 825559
rect 667416 818726 669572 823122
rect 44428 784665 46584 785541
rect 41218 783083 43374 783959
rect 44428 739865 46584 740741
rect 41218 738283 43374 739159
rect 44428 696665 46584 697541
rect 41218 695083 43374 695959
rect 44428 653465 46584 654341
rect 41218 651883 43374 652759
rect 44428 611325 46584 612201
rect 41218 609743 43374 610619
rect 44428 567065 46584 567941
rect 41218 565483 43374 566359
rect 667443 514121 669599 518517
rect 667457 504131 669613 508527
rect 50470 493293 51986 497689
rect 50458 483303 51974 487699
rect 44428 439465 46584 440341
rect 41218 437883 43374 438759
rect 664259 425839 666415 430235
rect 664242 415961 666398 420357
rect 44428 396265 46584 397141
rect 41218 394683 43374 395559
rect 44428 354065 46584 354941
rect 41218 352483 43374 353359
rect 44428 309865 46584 310741
rect 41218 308283 43374 309159
rect 44257 275977 46733 277173
rect 52753 277010 53629 277886
rect 658984 277975 659220 278211
rect 659304 277975 659540 278211
rect 659624 277975 659860 278211
rect 659944 277975 660180 278211
rect 660264 277975 660500 278211
rect 660584 277975 660820 278211
rect 660904 277975 661140 278211
rect 661224 277975 661460 278211
rect 661544 277975 661780 278211
rect 661864 277975 662100 278211
rect 662184 277975 662420 278211
rect 662504 277975 662740 278211
rect 662824 277975 663060 278211
rect 55806 276859 56362 277415
rect 55816 276052 56052 276288
rect 56136 276052 56372 276288
rect 42901 269420 43457 275416
rect 55824 275098 56060 275334
rect 56144 275098 56380 275334
rect 50273 272136 52109 273332
rect 55802 272057 56358 272613
rect 47879 270383 49715 271579
rect 55856 271094 56412 271650
rect 58689 269128 58925 269364
rect 58689 268808 58925 269044
rect 58689 268488 58925 268724
rect 58689 268168 58925 268404
rect 58689 267848 58925 268084
rect 58689 267528 58925 267764
rect 58689 267208 58925 267444
rect 58689 266888 58925 267124
rect 58689 266568 58925 266804
rect 62897 265124 63133 265360
rect 62897 264804 63133 265040
rect 48071 258769 49587 261245
rect 56555 258708 59351 261184
rect 62897 264484 63133 264720
rect 62897 264164 63133 264400
rect 62897 263844 63133 264080
rect 62897 263524 63133 263760
rect 62897 263204 63133 263440
rect 62897 262884 63133 263120
rect 62897 262564 63133 262800
rect 50471 254769 51987 257245
rect 56564 254708 60320 257184
rect 60980 257126 61216 257362
rect 60980 256806 61216 257042
rect 60980 256486 61216 256722
rect 60980 256166 61216 256402
rect 60980 255846 61216 256082
rect 60980 255526 61216 255762
rect 60980 255206 61216 255442
rect 60980 254886 61216 255122
rect 60980 254566 61216 254802
rect 52762 250572 53638 253368
rect 56232 250574 63188 253370
rect 41220 238397 43376 245353
rect 56551 242705 63187 245181
rect 63863 245134 64099 245370
rect 63863 244814 64099 245050
rect 63863 244494 64099 244730
rect 63863 244174 64099 244410
rect 63863 243854 64099 244090
rect 63863 243534 64099 243770
rect 63863 243214 64099 243450
rect 63863 242894 64099 243130
rect 63863 242574 64099 242810
rect 65775 253122 66011 253358
rect 65775 252802 66011 253038
rect 65775 252482 66011 252718
rect 65775 252162 66011 252398
rect 65775 251842 66011 252078
rect 65775 251522 66011 251758
rect 65775 251202 66011 251438
rect 65775 250882 66011 251118
rect 65775 250562 66011 250798
rect 390891 266565 391447 269361
rect 405941 266565 406497 269361
rect 383487 263052 384043 265208
rect 398537 263052 399093 265208
rect 392117 258713 392673 261189
rect 407237 258713 407793 261189
rect 384715 254570 385591 257366
rect 399815 254570 400691 257366
rect 276827 253140 277063 253376
rect 276827 252820 277063 253056
rect 276827 252500 277063 252736
rect 276827 252180 277063 252416
rect 276827 251860 277063 252096
rect 276827 251540 277063 251776
rect 276827 251220 277063 251456
rect 276827 250900 277063 251136
rect 276827 250580 277063 250816
rect 291827 253140 292063 253376
rect 291827 252820 292063 253056
rect 291827 252500 292063 252736
rect 291827 252180 292063 252416
rect 291827 251860 292063 252096
rect 291827 251540 292063 251776
rect 291827 251220 292063 251456
rect 291827 250900 292063 251136
rect 291827 250580 292063 250816
rect 306867 253140 307103 253376
rect 306867 252820 307103 253056
rect 306867 252500 307103 252736
rect 306867 252180 307103 252416
rect 306867 251860 307103 252096
rect 306867 251540 307103 251776
rect 306867 251220 307103 251456
rect 306867 250900 307103 251136
rect 306867 250580 307103 250816
rect 321987 253140 322223 253376
rect 321987 252820 322223 253056
rect 321987 252500 322223 252736
rect 321987 252180 322223 252416
rect 321987 251860 322223 252096
rect 321987 251540 322223 251776
rect 321987 251220 322223 251456
rect 321987 250900 322223 251136
rect 321987 250580 322223 250816
rect 66739 249134 66975 249370
rect 658965 277030 659201 277266
rect 659285 277030 659521 277266
rect 659605 277030 659841 277266
rect 659925 277030 660161 277266
rect 660245 277030 660481 277266
rect 660565 277030 660801 277266
rect 660885 277030 661121 277266
rect 661205 277030 661441 277266
rect 661525 277030 661761 277266
rect 661845 277030 662081 277266
rect 662165 277030 662401 277266
rect 662485 277030 662721 277266
rect 662805 277030 663041 277266
rect 670886 276144 673362 277340
rect 674086 276830 676562 278346
rect 651614 250561 652170 253357
rect 66739 248814 66975 249050
rect 66739 248494 66975 248730
rect 66739 248174 66975 248410
rect 66739 247854 66975 248090
rect 66739 247534 66975 247770
rect 66739 247214 66975 247450
rect 66739 246894 66975 247130
rect 66739 246574 66975 246810
rect 269470 248941 269706 249177
rect 269470 248621 269706 248857
rect 269470 248301 269706 248537
rect 269470 247981 269706 248217
rect 269470 247661 269706 247897
rect 269470 247341 269706 247577
rect 269470 247021 269706 247257
rect 269470 246701 269706 246937
rect 284460 248941 284696 249177
rect 284460 248621 284696 248857
rect 284460 248301 284696 248537
rect 284460 247981 284696 248217
rect 284460 247661 284696 247897
rect 284460 247341 284696 247577
rect 284460 247021 284696 247257
rect 284460 246701 284696 246937
rect 299460 248941 299696 249177
rect 299460 248621 299696 248857
rect 299460 248301 299696 248537
rect 299460 247981 299696 248217
rect 299460 247661 299696 247897
rect 299460 247341 299696 247577
rect 299460 247021 299696 247257
rect 299460 246701 299696 246937
rect 314720 248941 314956 249177
rect 314720 248621 314956 248857
rect 314720 248301 314956 248537
rect 314720 247981 314956 248217
rect 314720 247661 314956 247897
rect 314720 247341 314956 247577
rect 314720 247021 314956 247257
rect 314720 246701 314956 246937
rect 650648 246579 651204 249375
rect 199110 245137 199346 245373
rect 199110 244817 199346 245053
rect 199110 244497 199346 244733
rect 199110 244177 199346 244413
rect 199110 243857 199346 244093
rect 199110 243537 199346 243773
rect 199110 243217 199346 243453
rect 199110 242897 199346 243133
rect 199110 242577 199346 242813
rect 209170 245139 209406 245375
rect 209170 244819 209406 245055
rect 209170 244499 209406 244735
rect 209170 244179 209406 244415
rect 209170 243859 209406 244095
rect 209170 243539 209406 243775
rect 209170 243219 209406 243455
rect 209170 242899 209406 243135
rect 209170 242579 209406 242815
rect 44408 234627 46564 241263
rect 56566 238739 63202 241215
rect 64813 241130 65049 241366
rect 64813 240810 65049 241046
rect 64813 240490 65049 240726
rect 64813 240170 65049 240406
rect 64813 239850 65049 240086
rect 64813 239530 65049 239766
rect 64813 239210 65049 239446
rect 64813 238890 65049 239126
rect 64813 238570 65049 238806
rect 194930 241137 195166 241373
rect 194930 240817 195166 241053
rect 194930 240497 195166 240733
rect 194930 240177 195166 240413
rect 194930 239857 195166 240093
rect 194930 239537 195166 239773
rect 194930 239217 195166 239453
rect 194930 238897 195166 239133
rect 194930 238577 195166 238813
rect 205050 241137 205286 241373
rect 205050 240817 205286 241053
rect 205050 240497 205286 240733
rect 205050 240177 205286 240413
rect 205050 239857 205286 240093
rect 205050 239537 205286 239773
rect 205050 239217 205286 239453
rect 205050 238897 205286 239133
rect 205050 238577 205286 238813
rect 659185 274129 659421 274365
rect 659505 274129 659741 274365
rect 659825 274129 660061 274365
rect 660145 274129 660381 274365
rect 660465 274129 660701 274365
rect 660785 274129 661021 274365
rect 661105 274129 661341 274365
rect 661425 274129 661661 274365
rect 661745 274129 661981 274365
rect 662065 274129 662301 274365
rect 662385 274129 662621 274365
rect 662705 274129 662941 274365
rect 667448 273256 669604 274452
rect 655607 269125 655843 269361
rect 655607 268805 655843 269041
rect 655607 268485 655843 268721
rect 655607 268165 655843 268401
rect 655607 267845 655843 268081
rect 655607 267525 655843 267761
rect 655607 267205 655843 267441
rect 655607 266885 655843 267121
rect 655607 266565 655843 266801
rect 654649 265123 654885 265359
rect 654649 264803 654885 265039
rect 654649 264483 654885 264719
rect 654649 264163 654885 264399
rect 654649 263843 654885 264079
rect 654649 263523 654885 263759
rect 654649 263203 654885 263439
rect 654649 262883 654885 263119
rect 654649 262563 654885 262799
rect 657523 261137 657759 261373
rect 657523 260817 657759 261053
rect 657523 260497 657759 260733
rect 657523 260177 657759 260413
rect 657523 259857 657759 260093
rect 657523 259537 657759 259773
rect 657523 259217 657759 259453
rect 657523 258897 657759 259133
rect 657523 258577 657759 258813
rect 656561 257119 656797 257355
rect 656561 256799 656797 257035
rect 656561 256479 656797 256715
rect 656561 256159 656797 256395
rect 656561 255839 656797 256075
rect 656561 255519 656797 255755
rect 656561 255199 656797 255435
rect 656561 254879 656797 255115
rect 656561 254559 656797 254795
rect 667112 246737 669588 249213
rect 674226 246718 676382 249194
rect 653679 245137 653915 245373
rect 653679 244817 653915 245053
rect 653679 244497 653915 244733
rect 653679 244177 653915 244413
rect 653679 243857 653915 244093
rect 653679 243537 653915 243773
rect 653679 243217 653915 243453
rect 653679 242897 653915 243133
rect 653679 242577 653915 242813
rect 652721 241135 652957 241371
rect 652721 240815 652957 241051
rect 652721 240495 652957 240731
rect 652721 240175 652957 240411
rect 652721 239855 652957 240091
rect 652721 239535 652957 239771
rect 652721 239215 652957 239451
rect 652721 238895 652957 239131
rect 652721 238575 652957 238811
rect 48091 234739 50567 237215
rect 56455 234745 63091 237221
rect 140520 237125 140756 237361
rect 140520 236805 140756 237041
rect 140520 236485 140756 236721
rect 140520 236165 140756 236401
rect 140520 235845 140756 236081
rect 140520 235525 140756 235761
rect 140520 235205 140756 235441
rect 140520 234885 140756 235121
rect 140520 234565 140756 234801
rect 155600 237125 155836 237361
rect 155600 236805 155836 237041
rect 155600 236485 155836 236721
rect 155600 236165 155836 236401
rect 155600 235845 155836 236081
rect 155600 235525 155836 235761
rect 155600 235205 155836 235441
rect 155600 234885 155836 235121
rect 155600 234565 155836 234801
rect 170650 237125 170886 237361
rect 170650 236805 170886 237041
rect 170650 236485 170886 236721
rect 170650 236165 170886 236401
rect 170650 235845 170886 236081
rect 170650 235525 170886 235761
rect 170650 235205 170886 235441
rect 170650 234885 170886 235121
rect 170650 234565 170886 234801
rect 185660 237125 185896 237361
rect 185660 236805 185896 237041
rect 185660 236485 185896 236721
rect 185660 236165 185896 236401
rect 185660 235845 185896 236081
rect 185660 235525 185896 235761
rect 185660 235205 185896 235441
rect 185660 234885 185896 235121
rect 185660 234565 185896 234801
rect 215800 237125 216036 237361
rect 215800 236805 216036 237041
rect 215800 236485 216036 236721
rect 215800 236165 216036 236401
rect 215800 235845 216036 236081
rect 215800 235525 216036 235761
rect 215800 235205 216036 235441
rect 215800 234885 216036 235121
rect 215800 234565 216036 234801
rect 230850 237125 231086 237361
rect 230850 236805 231086 237041
rect 230850 236485 231086 236721
rect 230850 236165 231086 236401
rect 230850 235845 231086 236081
rect 230850 235525 231086 235761
rect 230850 235205 231086 235441
rect 230850 234885 231086 235121
rect 230850 234565 231086 234801
rect 245900 237125 246136 237361
rect 245900 236805 246136 237041
rect 245900 236485 246136 236721
rect 245900 236165 246136 236401
rect 245900 235845 246136 236081
rect 245900 235525 246136 235761
rect 245900 235205 246136 235441
rect 245900 234885 246136 235121
rect 245900 234565 246136 234801
rect 260950 237125 261186 237361
rect 260950 236805 261186 237041
rect 260950 236485 261186 236721
rect 260950 236165 261186 236401
rect 260950 235845 261186 236081
rect 260950 235525 261186 235761
rect 260950 235205 261186 235441
rect 260950 234885 261186 235121
rect 260950 234565 261186 234801
rect 276000 237125 276236 237361
rect 276000 236805 276236 237041
rect 276000 236485 276236 236721
rect 276000 236165 276236 236401
rect 276000 235845 276236 236081
rect 276000 235525 276236 235761
rect 276000 235205 276236 235441
rect 276000 234885 276236 235121
rect 276000 234565 276236 234801
rect 291050 237125 291286 237361
rect 291050 236805 291286 237041
rect 291050 236485 291286 236721
rect 291050 236165 291286 236401
rect 291050 235845 291286 236081
rect 291050 235525 291286 235761
rect 291050 235205 291286 235441
rect 291050 234885 291286 235121
rect 291050 234565 291286 234801
rect 306060 237125 306296 237361
rect 306060 236805 306296 237041
rect 306060 236485 306296 236721
rect 306060 236165 306296 236401
rect 306060 235845 306296 236081
rect 306060 235525 306296 235761
rect 306060 235205 306296 235441
rect 306060 234885 306296 235121
rect 306060 234565 306296 234801
rect 321250 237125 321486 237361
rect 321250 236805 321486 237041
rect 321250 236485 321486 236721
rect 321250 236165 321486 236401
rect 321250 235845 321486 236081
rect 321250 235525 321486 235761
rect 321250 235205 321486 235441
rect 321250 234885 321486 235121
rect 321250 234565 321486 234801
rect 336200 237125 336436 237361
rect 336200 236805 336436 237041
rect 336200 236485 336436 236721
rect 336200 236165 336436 236401
rect 336200 235845 336436 236081
rect 336200 235525 336436 235761
rect 336200 235205 336436 235441
rect 336200 234885 336436 235121
rect 336200 234565 336436 234801
rect 351350 237125 351586 237361
rect 351350 236805 351586 237041
rect 351350 236485 351586 236721
rect 351350 236165 351586 236401
rect 351350 235845 351586 236081
rect 351350 235525 351586 235761
rect 351350 235205 351586 235441
rect 351350 234885 351586 235121
rect 351350 234565 351586 234801
rect 366300 237125 366536 237361
rect 366300 236805 366536 237041
rect 366300 236485 366536 236721
rect 366300 236165 366536 236401
rect 366300 235845 366536 236081
rect 366300 235525 366536 235761
rect 366300 235205 366536 235441
rect 366300 234885 366536 235121
rect 366300 234565 366536 234801
rect 381150 237125 381386 237361
rect 381150 236805 381386 237041
rect 381150 236485 381386 236721
rect 381150 236165 381386 236401
rect 381150 235845 381386 236081
rect 381150 235525 381386 235761
rect 381150 235205 381386 235441
rect 381150 234885 381386 235121
rect 381150 234565 381386 234801
rect 396320 237125 396556 237361
rect 396320 236805 396556 237041
rect 396320 236485 396556 236721
rect 396320 236165 396556 236401
rect 396320 235845 396556 236081
rect 396320 235525 396556 235761
rect 396320 235205 396556 235441
rect 396320 234885 396556 235121
rect 396320 234565 396556 234801
rect 411450 237125 411686 237361
rect 411450 236805 411686 237041
rect 411450 236485 411686 236721
rect 411450 236165 411686 236401
rect 411450 235845 411686 236081
rect 411450 235525 411686 235761
rect 411450 235205 411686 235441
rect 411450 234885 411686 235121
rect 411450 234565 411686 234801
rect 426500 237125 426736 237361
rect 426500 236805 426736 237041
rect 426500 236485 426736 236721
rect 426500 236165 426736 236401
rect 426500 235845 426736 236081
rect 426500 235525 426736 235761
rect 426500 235205 426736 235441
rect 426500 234885 426736 235121
rect 426500 234565 426736 234801
rect 441550 237125 441786 237361
rect 441550 236805 441786 237041
rect 441550 236485 441786 236721
rect 441550 236165 441786 236401
rect 441550 235845 441786 236081
rect 441550 235525 441786 235761
rect 441550 235205 441786 235441
rect 441550 234885 441786 235121
rect 441550 234565 441786 234801
rect 456600 237125 456836 237361
rect 456600 236805 456836 237041
rect 456600 236485 456836 236721
rect 456600 236165 456836 236401
rect 456600 235845 456836 236081
rect 456600 235525 456836 235761
rect 456600 235205 456836 235441
rect 456600 234885 456836 235121
rect 456600 234565 456836 234801
rect 471650 237125 471886 237361
rect 471650 236805 471886 237041
rect 471650 236485 471886 236721
rect 471650 236165 471886 236401
rect 471650 235845 471886 236081
rect 471650 235525 471886 235761
rect 471650 235205 471886 235441
rect 471650 234885 471886 235121
rect 471650 234565 471886 234801
rect 486700 237125 486936 237361
rect 486700 236805 486936 237041
rect 486700 236485 486936 236721
rect 486700 236165 486936 236401
rect 486700 235845 486936 236081
rect 486700 235525 486936 235761
rect 486700 235205 486936 235441
rect 486700 234885 486936 235121
rect 486700 234565 486936 234801
rect 501750 237125 501986 237361
rect 501750 236805 501986 237041
rect 501750 236485 501986 236721
rect 501750 236165 501986 236401
rect 501750 235845 501986 236081
rect 501750 235525 501986 235761
rect 501750 235205 501986 235441
rect 501750 234885 501986 235121
rect 501750 234565 501986 234801
rect 56554 230735 62870 233211
rect 133140 233126 133376 233362
rect 133140 232806 133376 233042
rect 133140 232486 133376 232722
rect 133140 232166 133376 232402
rect 133140 231846 133376 232082
rect 133140 231526 133376 231762
rect 133140 231206 133376 231442
rect 133140 230886 133376 231122
rect 133140 230566 133376 230802
rect 148190 233126 148426 233362
rect 148190 232806 148426 233042
rect 148190 232486 148426 232722
rect 148190 232166 148426 232402
rect 148190 231846 148426 232082
rect 148190 231526 148426 231762
rect 148190 231206 148426 231442
rect 148190 230886 148426 231122
rect 148190 230566 148426 230802
rect 163240 233126 163476 233362
rect 163240 232806 163476 233042
rect 163240 232486 163476 232722
rect 163240 232166 163476 232402
rect 163240 231846 163476 232082
rect 163240 231526 163476 231762
rect 163240 231206 163476 231442
rect 163240 230886 163476 231122
rect 163240 230566 163476 230802
rect 178290 233126 178526 233362
rect 178290 232806 178526 233042
rect 178290 232486 178526 232722
rect 178290 232166 178526 232402
rect 178290 231846 178526 232082
rect 178290 231526 178526 231762
rect 178290 231206 178526 231442
rect 178290 230886 178526 231122
rect 178290 230566 178526 230802
rect 193340 233126 193576 233362
rect 193340 232806 193576 233042
rect 193340 232486 193576 232722
rect 193340 232166 193576 232402
rect 193340 231846 193576 232082
rect 193340 231526 193576 231762
rect 193340 231206 193576 231442
rect 193340 230886 193576 231122
rect 193340 230566 193576 230802
rect 208390 233126 208626 233362
rect 208390 232806 208626 233042
rect 208390 232486 208626 232722
rect 208390 232166 208626 232402
rect 208390 231846 208626 232082
rect 208390 231526 208626 231762
rect 208390 231206 208626 231442
rect 208390 230886 208626 231122
rect 208390 230566 208626 230802
rect 223440 233126 223676 233362
rect 223440 232806 223676 233042
rect 223440 232486 223676 232722
rect 223440 232166 223676 232402
rect 223440 231846 223676 232082
rect 223440 231526 223676 231762
rect 223440 231206 223676 231442
rect 223440 230886 223676 231122
rect 223440 230566 223676 230802
rect 238490 233126 238726 233362
rect 238490 232806 238726 233042
rect 238490 232486 238726 232722
rect 238490 232166 238726 232402
rect 238490 231846 238726 232082
rect 238490 231526 238726 231762
rect 238490 231206 238726 231442
rect 238490 230886 238726 231122
rect 238490 230566 238726 230802
rect 253540 233126 253776 233362
rect 253540 232806 253776 233042
rect 253540 232486 253776 232722
rect 253540 232166 253776 232402
rect 253540 231846 253776 232082
rect 253540 231526 253776 231762
rect 253540 231206 253776 231442
rect 253540 230886 253776 231122
rect 253540 230566 253776 230802
rect 268590 233126 268826 233362
rect 268590 232806 268826 233042
rect 268590 232486 268826 232722
rect 268590 232166 268826 232402
rect 268590 231846 268826 232082
rect 268590 231526 268826 231762
rect 268590 231206 268826 231442
rect 268590 230886 268826 231122
rect 268590 230566 268826 230802
rect 283640 233126 283876 233362
rect 283640 232806 283876 233042
rect 283640 232486 283876 232722
rect 283640 232166 283876 232402
rect 283640 231846 283876 232082
rect 283640 231526 283876 231762
rect 283640 231206 283876 231442
rect 283640 230886 283876 231122
rect 283640 230566 283876 230802
rect 298690 233126 298926 233362
rect 298690 232806 298926 233042
rect 298690 232486 298926 232722
rect 298690 232166 298926 232402
rect 298690 231846 298926 232082
rect 298690 231526 298926 231762
rect 298690 231206 298926 231442
rect 298690 230886 298926 231122
rect 298690 230566 298926 230802
rect 313740 233126 313976 233362
rect 313740 232806 313976 233042
rect 313740 232486 313976 232722
rect 313740 232166 313976 232402
rect 313740 231846 313976 232082
rect 313740 231526 313976 231762
rect 313740 231206 313976 231442
rect 313740 230886 313976 231122
rect 313740 230566 313976 230802
rect 328790 233126 329026 233362
rect 328790 232806 329026 233042
rect 328790 232486 329026 232722
rect 328790 232166 329026 232402
rect 328790 231846 329026 232082
rect 328790 231526 329026 231762
rect 328790 231206 329026 231442
rect 328790 230886 329026 231122
rect 328790 230566 329026 230802
rect 343840 233126 344076 233362
rect 343840 232806 344076 233042
rect 343840 232486 344076 232722
rect 343840 232166 344076 232402
rect 343840 231846 344076 232082
rect 343840 231526 344076 231762
rect 343840 231206 344076 231442
rect 343840 230886 344076 231122
rect 343840 230566 344076 230802
rect 358890 233126 359126 233362
rect 358890 232806 359126 233042
rect 358890 232486 359126 232722
rect 358890 232166 359126 232402
rect 358890 231846 359126 232082
rect 358890 231526 359126 231762
rect 358890 231206 359126 231442
rect 358890 230886 359126 231122
rect 358890 230566 359126 230802
rect 373940 233126 374176 233362
rect 373940 232806 374176 233042
rect 373940 232486 374176 232722
rect 373940 232166 374176 232402
rect 373940 231846 374176 232082
rect 373940 231526 374176 231762
rect 373940 231206 374176 231442
rect 373940 230886 374176 231122
rect 373940 230566 374176 230802
rect 388990 233126 389226 233362
rect 388990 232806 389226 233042
rect 388990 232486 389226 232722
rect 388990 232166 389226 232402
rect 388990 231846 389226 232082
rect 388990 231526 389226 231762
rect 388990 231206 389226 231442
rect 388990 230886 389226 231122
rect 388990 230566 389226 230802
rect 404040 233126 404276 233362
rect 404040 232806 404276 233042
rect 404040 232486 404276 232722
rect 404040 232166 404276 232402
rect 404040 231846 404276 232082
rect 404040 231526 404276 231762
rect 404040 231206 404276 231442
rect 404040 230886 404276 231122
rect 404040 230566 404276 230802
rect 419090 233126 419326 233362
rect 419090 232806 419326 233042
rect 419090 232486 419326 232722
rect 419090 232166 419326 232402
rect 419090 231846 419326 232082
rect 419090 231526 419326 231762
rect 419090 231206 419326 231442
rect 419090 230886 419326 231122
rect 419090 230566 419326 230802
rect 434140 233126 434376 233362
rect 434140 232806 434376 233042
rect 434140 232486 434376 232722
rect 434140 232166 434376 232402
rect 434140 231846 434376 232082
rect 434140 231526 434376 231762
rect 434140 231206 434376 231442
rect 434140 230886 434376 231122
rect 434140 230566 434376 230802
rect 449190 233126 449426 233362
rect 449190 232806 449426 233042
rect 449190 232486 449426 232722
rect 449190 232166 449426 232402
rect 449190 231846 449426 232082
rect 449190 231526 449426 231762
rect 449190 231206 449426 231442
rect 449190 230886 449426 231122
rect 449190 230566 449426 230802
rect 464240 233126 464476 233362
rect 464240 232806 464476 233042
rect 464240 232486 464476 232722
rect 464240 232166 464476 232402
rect 464240 231846 464476 232082
rect 464240 231526 464476 231762
rect 464240 231206 464476 231442
rect 464240 230886 464476 231122
rect 464240 230566 464476 230802
rect 479290 233126 479526 233362
rect 479290 232806 479526 233042
rect 479290 232486 479526 232722
rect 479290 232166 479526 232402
rect 479290 231846 479526 232082
rect 479290 231526 479526 231762
rect 479290 231206 479526 231442
rect 479290 230886 479526 231122
rect 479290 230566 479526 230802
rect 494340 233126 494576 233362
rect 494340 232806 494576 233042
rect 494340 232486 494576 232722
rect 494340 232166 494576 232402
rect 494340 231846 494576 232082
rect 494340 231526 494576 231762
rect 494340 231206 494576 231442
rect 494340 230886 494576 231122
rect 494340 230566 494576 230802
rect 584610 209795 587086 212271
rect 593464 209795 595940 212271
rect 627303 209758 627859 212234
rect 582400 208066 582636 208302
rect 582720 208066 582956 208302
rect 583040 208066 583276 208302
rect 583360 208066 583596 208302
rect 588493 208066 588729 208302
rect 588813 208066 589049 208302
rect 589133 208066 589369 208302
rect 589453 208066 589689 208302
rect 589773 208066 590009 208302
rect 590093 208066 590329 208302
rect 590413 208066 590649 208302
rect 590733 208066 590969 208302
rect 591053 208066 591289 208302
rect 51573 197076 51809 197312
rect 51893 197076 52129 197312
rect 584783 197165 586939 197721
rect 592038 197247 592274 197483
rect 592358 197247 592594 197483
rect 592678 197247 592914 197483
rect 582204 184054 582440 184290
rect 582524 184054 582760 184290
rect 588493 184050 588729 184286
rect 588813 184050 589049 184286
rect 589133 184050 589369 184286
rect 589453 184050 589689 184286
rect 589773 184050 590009 184286
rect 590093 184050 590329 184286
rect 590413 184050 590649 184286
rect 590733 184050 590969 184286
rect 591053 184050 591289 184286
rect 42087 173389 45523 176505
rect 42857 171058 43093 171294
rect 43177 171058 43413 171294
rect 43497 171058 43733 171294
rect 43817 171058 44053 171294
rect 44137 171058 44373 171294
rect 44457 171058 44693 171294
rect 44777 171058 45013 171294
rect 45097 171058 45333 171294
rect 45417 171058 45653 171294
rect 51465 171062 51701 171298
rect 51785 171062 52021 171298
rect 584783 166525 586939 167081
rect 592021 166619 592257 166855
rect 592341 166619 592577 166855
rect 592661 166619 592897 166855
rect 580242 158058 580478 158294
rect 580562 158058 580798 158294
rect 580882 158058 581118 158294
rect 581202 158058 581438 158294
rect 581522 158058 581758 158294
rect 581842 158058 582078 158294
rect 582162 158058 582398 158294
rect 582482 158058 582718 158294
rect 588467 158062 588703 158298
rect 588787 158062 589023 158298
rect 589107 158062 589343 158298
rect 589427 158062 589663 158298
rect 589747 158062 589983 158298
rect 590067 158062 590303 158298
rect 590387 158062 590623 158298
rect 590707 158062 590943 158298
rect 591027 158062 591263 158298
rect 42871 145064 43107 145300
rect 43191 145064 43427 145300
rect 43511 145064 43747 145300
rect 43831 145064 44067 145300
rect 44151 145064 44387 145300
rect 44471 145064 44707 145300
rect 44791 145064 45027 145300
rect 45111 145064 45347 145300
rect 45431 145064 45667 145300
rect 51399 145054 51635 145290
rect 51719 145054 51955 145290
rect 584783 135885 586939 136441
rect 592011 135979 592247 136215
rect 592331 135979 592567 136215
rect 592651 135979 592887 136215
rect 580252 132052 580488 132288
rect 580572 132052 580808 132288
rect 580892 132052 581128 132288
rect 581212 132052 581448 132288
rect 581532 132052 581768 132288
rect 581852 132052 582088 132288
rect 582172 132052 582408 132288
rect 582492 132052 582728 132288
rect 588493 132046 588729 132282
rect 588813 132046 589049 132282
rect 589133 132046 589369 132282
rect 589453 132046 589689 132282
rect 589773 132046 590009 132282
rect 590093 132046 590329 132282
rect 590413 132046 590649 132282
rect 590733 132046 590969 132282
rect 591053 132046 591289 132282
rect 42861 119060 43097 119296
rect 43181 119060 43417 119296
rect 43501 119060 43737 119296
rect 43821 119060 44057 119296
rect 44141 119060 44377 119296
rect 44461 119060 44697 119296
rect 44781 119060 45017 119296
rect 45101 119060 45337 119296
rect 45421 119060 45657 119296
rect 51395 119060 51631 119296
rect 51715 119060 51951 119296
rect 580254 106058 580490 106294
rect 580574 106058 580810 106294
rect 580894 106058 581130 106294
rect 581214 106058 581450 106294
rect 581534 106058 581770 106294
rect 581854 106058 582090 106294
rect 582174 106058 582410 106294
rect 582494 106058 582730 106294
rect 588497 106058 588733 106294
rect 588817 106058 589053 106294
rect 589137 106058 589373 106294
rect 589457 106058 589693 106294
rect 589777 106058 590013 106294
rect 590097 106058 590333 106294
rect 590417 106058 590653 106294
rect 590737 106058 590973 106294
rect 591057 106058 591293 106294
rect 584783 104965 586939 105521
rect 592023 105342 592259 105578
rect 592343 105342 592579 105578
rect 592663 105342 592899 105578
rect 597012 96127 597888 98603
rect 627823 96189 628699 98665
rect 636259 96685 636815 98521
rect 42857 93058 43093 93294
rect 43177 93058 43413 93294
rect 43497 93058 43733 93294
rect 43817 93058 44053 93294
rect 44137 93058 44373 93294
rect 44457 93058 44693 93294
rect 44777 93058 45013 93294
rect 45097 93058 45333 93294
rect 45417 93058 45653 93294
rect 51399 93056 51635 93292
rect 51719 93056 51955 93292
rect 42091 78276 45527 82672
rect 580248 80068 580484 80304
rect 580568 80068 580804 80304
rect 580888 80068 581124 80304
rect 581208 80068 581444 80304
rect 581528 80068 581764 80304
rect 581848 80068 582084 80304
rect 582168 80068 582404 80304
rect 582488 80068 582724 80304
rect 588491 80070 588727 80306
rect 588811 80070 589047 80306
rect 589131 80070 589367 80306
rect 589451 80070 589687 80306
rect 589771 80070 590007 80306
rect 590091 80070 590327 80306
rect 590411 80070 590647 80306
rect 590731 80070 590967 80306
rect 591051 80070 591287 80306
rect 632254 78473 632810 80629
rect 640232 78340 640788 80816
rect 629919 76957 630155 77193
rect 629919 76637 630155 76873
rect 629919 76317 630155 76553
rect 631471 75555 631707 75791
rect 631471 75235 631707 75471
rect 631471 74915 631707 75151
rect 633031 76971 633267 77207
rect 633031 76651 633267 76887
rect 633031 76331 633267 76567
rect 634565 75559 634801 75795
rect 634565 75239 634801 75475
rect 634565 74919 634801 75155
rect 636121 76967 636357 77203
rect 636121 76647 636357 76883
rect 636121 76327 636357 76563
rect 637673 75563 637909 75799
rect 637673 75243 637909 75479
rect 637673 74923 637909 75159
rect 639215 76967 639451 77203
rect 639215 76647 639451 76883
rect 639215 76327 639451 76563
rect 640777 75555 641013 75791
rect 640777 75235 641013 75471
rect 640777 74915 641013 75151
rect 642323 76979 642559 77215
rect 642323 76659 642559 76895
rect 642323 76339 642559 76575
rect 643879 75581 644115 75817
rect 643879 75261 644115 75497
rect 643879 74941 644115 75177
rect 42067 68372 45503 72768
rect 42095 67052 42331 67288
rect 42415 67052 42651 67288
rect 42735 67052 42971 67288
rect 43055 67052 43291 67288
rect 43375 67052 43611 67288
rect 43695 67052 43931 67288
rect 44015 67052 44251 67288
rect 44335 67052 44571 67288
rect 44655 67052 44891 67288
rect 44975 67052 45211 67288
rect 45295 67052 45531 67288
rect 51597 67058 51833 67294
rect 51917 67058 52153 67294
rect 42080 48478 45516 51914
rect 54650 48444 58086 51880
rect 143423 50036 144619 50592
rect 141528 44318 142724 45194
rect 241825 46601 245901 46607
rect 241825 42857 245901 46601
rect 241825 42851 245901 42857
rect 251477 46615 255553 46621
rect 251477 42871 255553 46615
rect 251477 42865 255553 42871
rect 648289 46774 648525 47010
rect 648609 46774 648845 47010
rect 648929 46774 649165 47010
rect 649249 46774 649485 47010
rect 666522 47038 666758 47274
rect 666842 47038 667078 47274
rect 667162 47038 667398 47274
rect 667482 47038 667718 47274
rect 667802 47038 668038 47274
rect 668122 47038 668358 47274
rect 668442 47038 668678 47274
rect 668762 47038 668998 47274
rect 669082 47038 669318 47274
<< metal5 >>
rect 52598 996544 676660 996702
rect 52598 995668 671036 996544
rect 676392 995668 676660 996544
rect 52598 995502 676660 995668
rect 47798 990125 49798 990466
rect 47798 989889 47874 990125
rect 48110 989889 48194 990125
rect 48430 989889 48514 990125
rect 48750 989889 48834 990125
rect 49070 989889 49154 990125
rect 49390 989889 49474 990125
rect 49710 989889 49798 990125
rect 41034 986441 43574 986448
rect 41034 985885 41066 986441
rect 43542 985885 43574 986441
rect 41034 985878 43574 985885
rect 44242 985486 46772 985498
rect 44242 984930 44269 985486
rect 46745 984930 46772 985486
rect 44242 984918 46772 984930
rect 44278 952941 46734 953030
rect 44278 952065 44428 952941
rect 46584 952065 46734 952941
rect 44278 951976 46734 952065
rect 41068 951359 43524 951448
rect 41068 950483 41218 951359
rect 43374 950483 43524 951359
rect 41068 950394 43524 950483
rect 47798 842260 49798 989889
rect 47798 837864 48043 842260
rect 49559 837864 49798 842260
rect 47798 832328 49798 837864
rect 47798 827932 48043 832328
rect 49559 827932 49798 832328
rect 44278 827141 46734 827230
rect 44278 826265 44428 827141
rect 46584 826265 46734 827141
rect 44278 826176 46734 826265
rect 41068 825559 43524 825648
rect 41068 824683 41218 825559
rect 43374 824683 43524 825559
rect 41068 824594 43524 824683
rect 44278 785541 46734 785630
rect 44278 784665 44428 785541
rect 46584 784665 46734 785541
rect 44278 784576 46734 784665
rect 41068 783959 43524 784048
rect 41068 783083 41218 783959
rect 43374 783083 43524 783959
rect 41068 782994 43524 783083
rect 44278 740741 46734 740830
rect 44278 739865 44428 740741
rect 46584 739865 46734 740741
rect 44278 739776 46734 739865
rect 41068 739159 43524 739248
rect 41068 738283 41218 739159
rect 43374 738283 43524 739159
rect 41068 738194 43524 738283
rect 44278 697541 46734 697630
rect 44278 696665 44428 697541
rect 46584 696665 46734 697541
rect 44278 696576 46734 696665
rect 41068 695959 43524 696048
rect 41068 695083 41218 695959
rect 43374 695083 43524 695959
rect 41068 694994 43524 695083
rect 44278 654341 46734 654430
rect 44278 653465 44428 654341
rect 46584 653465 46734 654341
rect 44278 653376 46734 653465
rect 41068 652759 43524 652848
rect 41068 651883 41218 652759
rect 43374 651883 43524 652759
rect 41068 651794 43524 651883
rect 44278 612201 46734 612290
rect 44278 611325 44428 612201
rect 46584 611325 46734 612201
rect 44278 611236 46734 611325
rect 41068 610619 43524 610708
rect 41068 609743 41218 610619
rect 43374 609743 43524 610619
rect 41068 609654 43524 609743
rect 44278 567941 46734 568030
rect 44278 567065 44428 567941
rect 46584 567065 46734 567941
rect 44278 566976 46734 567065
rect 41068 566359 43524 566448
rect 41068 565483 41218 566359
rect 43374 565483 43524 566359
rect 41068 565394 43524 565483
rect 44278 440341 46734 440430
rect 44278 439465 44428 440341
rect 46584 439465 46734 440341
rect 44278 439376 46734 439465
rect 41068 438759 43524 438848
rect 41068 437883 41218 438759
rect 43374 437883 43524 438759
rect 41068 437794 43524 437883
rect 44278 397141 46734 397230
rect 44278 396265 44428 397141
rect 46584 396265 46734 397141
rect 44278 396176 46734 396265
rect 41068 395559 43524 395648
rect 41068 394683 41218 395559
rect 43374 394683 43524 395559
rect 41068 394594 43524 394683
rect 44278 354941 46734 355030
rect 44278 354065 44428 354941
rect 46584 354065 46734 354941
rect 44278 353976 46734 354065
rect 41068 353359 43524 353448
rect 41068 352483 41218 353359
rect 43374 352483 43524 353359
rect 41068 352394 43524 352483
rect 44278 310741 46734 310830
rect 44278 309865 44428 310741
rect 46584 309865 46734 310741
rect 44278 309776 46734 309865
rect 41068 309159 43524 309248
rect 41068 308283 41218 309159
rect 43374 308283 43524 309159
rect 41068 308194 43524 308283
rect 44228 277173 46762 277262
rect 44228 275977 44257 277173
rect 46733 275977 46762 277173
rect 44228 275888 46762 275977
rect 42830 275416 43528 275458
rect 42830 269420 42901 275416
rect 43457 269420 43528 275416
rect 42830 269378 43528 269420
rect 47798 271579 49798 827932
rect 47798 270383 47879 271579
rect 49715 270383 49798 271579
rect 47798 261245 49798 270383
rect 47798 258769 48071 261245
rect 49587 258769 49798 261245
rect 47798 258484 49798 258769
rect 50198 989161 52198 990466
rect 50198 988925 50280 989161
rect 50516 988925 50600 989161
rect 50836 988925 50920 989161
rect 51156 988925 51240 989161
rect 51476 988925 51560 989161
rect 51796 988925 51880 989161
rect 52116 988925 52198 989161
rect 50198 497689 52198 988925
rect 50198 493293 50470 497689
rect 51986 493293 52198 497689
rect 50198 487699 52198 493293
rect 50198 483303 50458 487699
rect 51974 483303 52198 487699
rect 50198 273332 52198 483303
rect 50198 272136 50273 273332
rect 52109 272136 52198 273332
rect 50198 257245 52198 272136
rect 50198 254769 50471 257245
rect 51987 254769 52198 257245
rect 50198 254498 52198 254769
rect 52598 984357 53798 995502
rect 52598 984121 52759 984357
rect 52995 984121 53079 984357
rect 53315 984121 53399 984357
rect 53635 984121 53798 984357
rect 52598 277886 53798 984121
rect 52598 277010 52753 277886
rect 53629 277010 53798 277886
rect 52598 253368 53798 277010
rect 52598 250572 52762 253368
rect 53638 250572 53798 253368
rect 41066 245353 43530 245388
rect 41066 238397 41220 245353
rect 43376 238397 43530 245353
rect 41066 238362 43530 238397
rect 44254 241263 46718 241358
rect 44254 234627 44408 241263
rect 46564 234627 46718 241263
rect 44254 234532 46718 234627
rect 47836 237215 50836 237612
rect 47836 234739 48091 237215
rect 50567 234739 50836 237215
rect 47836 210498 50836 234739
rect 52598 217742 53798 250572
rect 54198 993902 676620 995102
rect 54198 983588 55398 993902
rect 575640 993191 666620 993396
rect 575640 993177 585871 993191
rect 575640 991021 575875 993177
rect 580271 991035 585871 993177
rect 590267 991035 666620 993191
rect 674020 992696 676620 993902
rect 580271 991021 666620 991035
rect 575640 990796 666620 991021
rect 55776 990126 56596 990308
rect 55776 989890 55829 990126
rect 56065 989890 56149 990126
rect 56385 989890 56596 990126
rect 55776 989688 56596 989890
rect 55776 989166 57552 989348
rect 55776 988930 55833 989166
rect 56069 988930 56153 989166
rect 56389 988930 57552 989166
rect 55776 988728 57552 988930
rect 664020 988388 666620 990796
rect 670976 992520 673264 992530
rect 670976 990364 671042 992520
rect 673198 990364 673264 992520
rect 670976 990354 673264 990364
rect 656038 987768 666620 988388
rect 655078 987242 663178 987428
rect 655078 987006 658577 987242
rect 658813 987006 658897 987242
rect 659133 987006 659217 987242
rect 659453 987006 659537 987242
rect 659773 987006 659857 987242
rect 660093 987006 660177 987242
rect 660413 987006 660497 987242
rect 660733 987006 660817 987242
rect 661053 987006 661137 987242
rect 661373 987006 661457 987242
rect 661693 987006 661777 987242
rect 662013 987006 662097 987242
rect 662333 987006 662417 987242
rect 662653 987006 662737 987242
rect 662973 987006 663178 987242
rect 655078 986808 663178 987006
rect 55776 986279 60436 986468
rect 55776 986043 55813 986279
rect 56049 986043 56133 986279
rect 56369 986043 60436 986279
rect 55776 985848 60436 986043
rect 55776 985475 61398 985508
rect 55776 984919 55828 985475
rect 56384 984919 61398 985475
rect 55776 984888 61398 984919
rect 55776 984517 62358 984548
rect 55776 983961 55811 984517
rect 56367 983961 62358 984517
rect 55776 983928 62358 983961
rect 652180 984356 663178 984548
rect 652180 984120 658391 984356
rect 658627 984120 658711 984356
rect 658947 984120 659031 984356
rect 659267 984120 659351 984356
rect 659587 984120 659671 984356
rect 659907 984120 659991 984356
rect 660227 984120 660311 984356
rect 660547 984120 660631 984356
rect 660867 984120 660951 984356
rect 661187 984120 661271 984356
rect 661507 984120 661591 984356
rect 661827 984120 661911 984356
rect 662147 984120 662231 984356
rect 662467 984120 662551 984356
rect 662787 984120 662871 984356
rect 663107 984120 663178 984356
rect 652180 983928 663178 984120
rect 54198 982968 63316 983588
rect 651228 983400 663178 983588
rect 651228 983164 658373 983400
rect 658609 983164 658693 983400
rect 658929 983164 659013 983400
rect 659249 983164 659333 983400
rect 659569 983164 659653 983400
rect 659889 983164 659973 983400
rect 660209 983164 660293 983400
rect 660529 983164 660613 983400
rect 660849 983164 660933 983400
rect 661169 983164 661253 983400
rect 661489 983164 661573 983400
rect 661809 983164 661893 983400
rect 662129 983164 662213 983400
rect 662449 983164 662533 983400
rect 662769 983164 662853 983400
rect 663089 983164 663178 983400
rect 651228 982968 663178 983164
rect 54198 278404 55398 982968
rect 664020 430235 666620 987768
rect 664020 425839 664259 430235
rect 666415 425839 666620 430235
rect 664020 420357 666620 425839
rect 664020 415961 664242 420357
rect 666398 415961 666620 420357
rect 54198 277784 63312 278404
rect 651226 278211 663158 278404
rect 651226 277975 658984 278211
rect 659220 277975 659304 278211
rect 659540 277975 659624 278211
rect 659860 277975 659944 278211
rect 660180 277975 660264 278211
rect 660500 277975 660584 278211
rect 660820 277975 660904 278211
rect 661140 277975 661224 278211
rect 661460 277975 661544 278211
rect 661780 277975 661864 278211
rect 662100 277975 662184 278211
rect 662420 277975 662504 278211
rect 662740 277975 662824 278211
rect 663060 277975 663158 278211
rect 651226 277784 663158 277975
rect 54198 249466 55398 277784
rect 55754 277415 62352 277444
rect 55754 276859 55806 277415
rect 56362 276859 62352 277415
rect 55754 276824 62352 276859
rect 652188 277266 663158 277444
rect 652188 277030 658965 277266
rect 659201 277030 659285 277266
rect 659521 277030 659605 277266
rect 659841 277030 659925 277266
rect 660161 277030 660245 277266
rect 660481 277030 660565 277266
rect 660801 277030 660885 277266
rect 661121 277030 661205 277266
rect 661441 277030 661525 277266
rect 661761 277030 661845 277266
rect 662081 277030 662165 277266
rect 662401 277030 662485 277266
rect 662721 277030 662805 277266
rect 663041 277030 663158 277266
rect 652188 276824 663158 277030
rect 55754 276288 61388 276484
rect 55754 276052 55816 276288
rect 56052 276052 56136 276288
rect 56372 276052 61388 276288
rect 55754 275864 61388 276052
rect 55754 275334 60428 275524
rect 55754 275098 55824 275334
rect 56060 275098 56144 275334
rect 56380 275098 60428 275334
rect 55754 274904 60428 275098
rect 655060 274365 663158 274564
rect 655060 274129 659185 274365
rect 659421 274129 659505 274365
rect 659741 274129 659825 274365
rect 660061 274129 660145 274365
rect 660381 274129 660465 274365
rect 660701 274129 660785 274365
rect 661021 274129 661105 274365
rect 661341 274129 661425 274365
rect 661661 274129 661745 274365
rect 661981 274129 662065 274365
rect 662301 274129 662385 274365
rect 662621 274129 662705 274365
rect 662941 274129 663158 274365
rect 655060 273944 663158 274129
rect 664020 273604 666620 415961
rect 656026 272984 666620 273604
rect 55754 272613 57546 272644
rect 55754 272057 55802 272613
rect 56358 272057 57546 272613
rect 55754 272024 57546 272057
rect 55754 271650 56590 271684
rect 55754 271094 55856 271650
rect 56412 271094 56590 271650
rect 55754 271064 56590 271094
rect 664020 269466 666620 272984
rect 58388 269364 666620 269466
rect 58388 269128 58689 269364
rect 58925 269361 666620 269364
rect 58925 269128 390891 269361
rect 58388 269044 390891 269128
rect 58388 268808 58689 269044
rect 58925 268808 390891 269044
rect 58388 268724 390891 268808
rect 58388 268488 58689 268724
rect 58925 268488 390891 268724
rect 58388 268404 390891 268488
rect 58388 268168 58689 268404
rect 58925 268168 390891 268404
rect 58388 268084 390891 268168
rect 58388 267848 58689 268084
rect 58925 267848 390891 268084
rect 58388 267764 390891 267848
rect 58388 267528 58689 267764
rect 58925 267528 390891 267764
rect 58388 267444 390891 267528
rect 58388 267208 58689 267444
rect 58925 267208 390891 267444
rect 58388 267124 390891 267208
rect 58388 266888 58689 267124
rect 58925 266888 390891 267124
rect 58388 266804 390891 266888
rect 58388 266568 58689 266804
rect 58925 266568 390891 266804
rect 58388 266565 390891 266568
rect 391447 266565 405941 269361
rect 406497 269125 655607 269361
rect 655843 269125 666620 269361
rect 406497 269041 666620 269125
rect 406497 268805 655607 269041
rect 655843 268805 666620 269041
rect 406497 268721 666620 268805
rect 406497 268485 655607 268721
rect 655843 268485 666620 268721
rect 406497 268401 666620 268485
rect 406497 268165 655607 268401
rect 655843 268165 666620 268401
rect 406497 268081 666620 268165
rect 406497 267845 655607 268081
rect 655843 267845 666620 268081
rect 406497 267761 666620 267845
rect 406497 267525 655607 267761
rect 655843 267525 666620 267761
rect 406497 267441 666620 267525
rect 406497 267205 655607 267441
rect 655843 267205 666620 267441
rect 406497 267121 666620 267205
rect 406497 266885 655607 267121
rect 655843 266885 666620 267121
rect 406497 266801 666620 266885
rect 406497 266565 655607 266801
rect 655843 266565 666620 266801
rect 58388 266466 666620 266565
rect 667220 987247 669820 987566
rect 667220 987011 667281 987247
rect 667517 987011 667601 987247
rect 667837 987011 667921 987247
rect 668157 987011 668241 987247
rect 668477 987011 668561 987247
rect 668797 987011 668881 987247
rect 669117 987011 669201 987247
rect 669437 987011 669521 987247
rect 669757 987011 669820 987247
rect 667220 833116 669820 987011
rect 670858 984521 673384 984536
rect 670858 983965 670883 984521
rect 673359 983965 673384 984521
rect 670858 983950 673384 983965
rect 674056 983559 676582 983574
rect 674056 983003 674081 983559
rect 676557 983003 676582 983559
rect 674056 982988 676582 983003
rect 674734 901031 675740 901112
rect 674734 900155 674799 901031
rect 675675 900155 675740 901031
rect 674734 900074 675740 900155
rect 671566 899423 672596 899504
rect 671566 898547 671643 899423
rect 672519 898547 672596 899423
rect 671566 898466 672596 898547
rect 674116 856022 675180 856116
rect 674116 855146 674210 856022
rect 675086 855146 675180 856022
rect 674116 855052 675180 855146
rect 671570 854420 672638 854522
rect 671570 853544 671666 854420
rect 672542 853544 672638 854420
rect 671570 853442 672638 853544
rect 667220 828720 667430 833116
rect 669586 828720 669820 833116
rect 667220 823122 669820 828720
rect 667220 818726 667416 823122
rect 669572 818726 669820 823122
rect 667220 518517 669820 818726
rect 667220 514121 667443 518517
rect 669599 514121 669820 518517
rect 667220 508527 669820 514121
rect 667220 504131 667457 508527
rect 669613 504131 669820 508527
rect 667220 274452 669820 504131
rect 674084 278346 676564 278356
rect 670884 277340 673364 277410
rect 670884 276144 670886 277340
rect 673362 276144 673364 277340
rect 674084 276830 674086 278346
rect 676562 276830 676564 278346
rect 674084 276820 676564 276830
rect 670884 276074 673364 276144
rect 667220 273256 667448 274452
rect 669604 273256 669820 274452
rect 667220 265466 669820 273256
rect 62534 265360 669820 265466
rect 62534 265124 62897 265360
rect 63133 265359 669820 265360
rect 63133 265208 654649 265359
rect 63133 265124 383487 265208
rect 62534 265040 383487 265124
rect 62534 264804 62897 265040
rect 63133 264804 383487 265040
rect 62534 264720 383487 264804
rect 62534 264484 62897 264720
rect 63133 264484 383487 264720
rect 62534 264400 383487 264484
rect 62534 264164 62897 264400
rect 63133 264164 383487 264400
rect 62534 264080 383487 264164
rect 62534 263844 62897 264080
rect 63133 263844 383487 264080
rect 62534 263760 383487 263844
rect 62534 263524 62897 263760
rect 63133 263524 383487 263760
rect 62534 263440 383487 263524
rect 62534 263204 62897 263440
rect 63133 263204 383487 263440
rect 62534 263120 383487 263204
rect 62534 262884 62897 263120
rect 63133 263052 383487 263120
rect 384043 263052 398537 265208
rect 399093 265123 654649 265208
rect 654885 265123 669820 265359
rect 399093 265039 669820 265123
rect 399093 264803 654649 265039
rect 654885 264803 669820 265039
rect 399093 264719 669820 264803
rect 399093 264483 654649 264719
rect 654885 264483 669820 264719
rect 399093 264399 669820 264483
rect 399093 264163 654649 264399
rect 654885 264163 669820 264399
rect 399093 264079 669820 264163
rect 399093 263843 654649 264079
rect 654885 263843 669820 264079
rect 399093 263759 669820 263843
rect 399093 263523 654649 263759
rect 654885 263523 669820 263759
rect 399093 263439 669820 263523
rect 399093 263203 654649 263439
rect 654885 263203 669820 263439
rect 399093 263119 669820 263203
rect 399093 263052 654649 263119
rect 63133 262884 654649 263052
rect 62534 262883 654649 262884
rect 654885 262883 669820 263119
rect 62534 262800 669820 262883
rect 62534 262564 62897 262800
rect 63133 262799 669820 262800
rect 63133 262564 654649 262799
rect 62534 262563 654649 262564
rect 654885 262563 669820 262799
rect 62534 262466 669820 262563
rect 56370 261373 658090 261466
rect 56370 261189 657523 261373
rect 56370 261184 392117 261189
rect 56370 258708 56555 261184
rect 59351 258713 392117 261184
rect 392673 258713 407237 261189
rect 407793 261137 657523 261189
rect 657759 261137 658090 261373
rect 407793 261053 658090 261137
rect 407793 260817 657523 261053
rect 657759 260817 658090 261053
rect 407793 260733 658090 260817
rect 407793 260497 657523 260733
rect 657759 260497 658090 260733
rect 407793 260413 658090 260497
rect 407793 260177 657523 260413
rect 657759 260177 658090 260413
rect 407793 260093 658090 260177
rect 407793 259857 657523 260093
rect 657759 259857 658090 260093
rect 407793 259773 658090 259857
rect 407793 259537 657523 259773
rect 657759 259537 658090 259773
rect 407793 259453 658090 259537
rect 407793 259217 657523 259453
rect 657759 259217 658090 259453
rect 407793 259133 658090 259217
rect 407793 258897 657523 259133
rect 657759 258897 658090 259133
rect 407793 258813 658090 258897
rect 407793 258713 657523 258813
rect 59351 258708 657523 258713
rect 56370 258577 657523 258708
rect 657759 258577 658090 258813
rect 56370 258466 658090 258577
rect 56370 257366 657076 257466
rect 56370 257362 384715 257366
rect 56370 257184 60980 257362
rect 56370 254708 56564 257184
rect 60320 257126 60980 257184
rect 61216 257126 384715 257362
rect 60320 257042 384715 257126
rect 60320 256806 60980 257042
rect 61216 256806 384715 257042
rect 60320 256722 384715 256806
rect 60320 256486 60980 256722
rect 61216 256486 384715 256722
rect 60320 256402 384715 256486
rect 60320 256166 60980 256402
rect 61216 256166 384715 256402
rect 60320 256082 384715 256166
rect 60320 255846 60980 256082
rect 61216 255846 384715 256082
rect 60320 255762 384715 255846
rect 60320 255526 60980 255762
rect 61216 255526 384715 255762
rect 60320 255442 384715 255526
rect 60320 255206 60980 255442
rect 61216 255206 384715 255442
rect 60320 255122 384715 255206
rect 60320 254886 60980 255122
rect 61216 254886 384715 255122
rect 60320 254802 384715 254886
rect 60320 254708 60980 254802
rect 56370 254566 60980 254708
rect 61216 254570 384715 254802
rect 385591 254570 399815 257366
rect 400691 257355 657076 257366
rect 400691 257119 656561 257355
rect 656797 257119 657076 257355
rect 400691 257035 657076 257119
rect 400691 256799 656561 257035
rect 656797 256799 657076 257035
rect 400691 256715 657076 256799
rect 400691 256479 656561 256715
rect 656797 256479 657076 256715
rect 400691 256395 657076 256479
rect 400691 256159 656561 256395
rect 656797 256159 657076 256395
rect 400691 256075 657076 256159
rect 400691 255839 656561 256075
rect 656797 255839 657076 256075
rect 400691 255755 657076 255839
rect 400691 255519 656561 255755
rect 656797 255519 657076 255755
rect 400691 255435 657076 255519
rect 400691 255199 656561 255435
rect 656797 255199 657076 255435
rect 400691 255115 657076 255199
rect 400691 254879 656561 255115
rect 656797 254879 657076 255115
rect 400691 254795 657076 254879
rect 400691 254570 656561 254795
rect 61216 254566 656561 254570
rect 56370 254559 656561 254566
rect 656797 254559 657076 254795
rect 56370 254466 657076 254559
rect 56126 253376 670986 253466
rect 56126 253370 276827 253376
rect 56126 250574 56232 253370
rect 63188 253358 276827 253370
rect 63188 253122 65775 253358
rect 66011 253140 276827 253358
rect 277063 253140 291827 253376
rect 292063 253140 306867 253376
rect 307103 253140 321987 253376
rect 322223 253357 670986 253376
rect 322223 253140 651614 253357
rect 66011 253122 651614 253140
rect 63188 253056 651614 253122
rect 63188 253038 276827 253056
rect 63188 252802 65775 253038
rect 66011 252820 276827 253038
rect 277063 252820 291827 253056
rect 292063 252820 306867 253056
rect 307103 252820 321987 253056
rect 322223 252820 651614 253056
rect 66011 252802 651614 252820
rect 63188 252736 651614 252802
rect 63188 252718 276827 252736
rect 63188 252482 65775 252718
rect 66011 252500 276827 252718
rect 277063 252500 291827 252736
rect 292063 252500 306867 252736
rect 307103 252500 321987 252736
rect 322223 252500 651614 252736
rect 66011 252482 651614 252500
rect 63188 252416 651614 252482
rect 63188 252398 276827 252416
rect 63188 252162 65775 252398
rect 66011 252180 276827 252398
rect 277063 252180 291827 252416
rect 292063 252180 306867 252416
rect 307103 252180 321987 252416
rect 322223 252180 651614 252416
rect 66011 252162 651614 252180
rect 63188 252096 651614 252162
rect 63188 252078 276827 252096
rect 63188 251842 65775 252078
rect 66011 251860 276827 252078
rect 277063 251860 291827 252096
rect 292063 251860 306867 252096
rect 307103 251860 321987 252096
rect 322223 251860 651614 252096
rect 66011 251842 651614 251860
rect 63188 251776 651614 251842
rect 63188 251758 276827 251776
rect 63188 251522 65775 251758
rect 66011 251540 276827 251758
rect 277063 251540 291827 251776
rect 292063 251540 306867 251776
rect 307103 251540 321987 251776
rect 322223 251540 651614 251776
rect 66011 251522 651614 251540
rect 63188 251456 651614 251522
rect 63188 251438 276827 251456
rect 63188 251202 65775 251438
rect 66011 251220 276827 251438
rect 277063 251220 291827 251456
rect 292063 251220 306867 251456
rect 307103 251220 321987 251456
rect 322223 251220 651614 251456
rect 66011 251202 651614 251220
rect 63188 251136 651614 251202
rect 63188 251118 276827 251136
rect 63188 250882 65775 251118
rect 66011 250900 276827 251118
rect 277063 250900 291827 251136
rect 292063 250900 306867 251136
rect 307103 250900 321987 251136
rect 322223 250900 651614 251136
rect 66011 250882 651614 250900
rect 63188 250816 651614 250882
rect 63188 250798 276827 250816
rect 63188 250574 65775 250798
rect 56126 250562 65775 250574
rect 66011 250580 276827 250798
rect 277063 250580 291827 250816
rect 292063 250580 306867 250816
rect 307103 250580 321987 250816
rect 322223 250580 651614 250816
rect 66011 250562 651614 250580
rect 56126 250561 651614 250562
rect 652170 250561 670986 253357
rect 56126 250466 670986 250561
rect 54198 249375 669890 249466
rect 54198 249370 650648 249375
rect 54198 249134 66739 249370
rect 66975 249177 650648 249370
rect 66975 249134 269470 249177
rect 54198 249050 269470 249134
rect 54198 248814 66739 249050
rect 66975 248941 269470 249050
rect 269706 248941 284460 249177
rect 284696 248941 299460 249177
rect 299696 248941 314720 249177
rect 314956 248941 650648 249177
rect 66975 248857 650648 248941
rect 66975 248814 269470 248857
rect 54198 248730 269470 248814
rect 54198 248494 66739 248730
rect 66975 248621 269470 248730
rect 269706 248621 284460 248857
rect 284696 248621 299460 248857
rect 299696 248621 314720 248857
rect 314956 248621 650648 248857
rect 66975 248537 650648 248621
rect 66975 248494 269470 248537
rect 54198 248410 269470 248494
rect 54198 248174 66739 248410
rect 66975 248301 269470 248410
rect 269706 248301 284460 248537
rect 284696 248301 299460 248537
rect 299696 248301 314720 248537
rect 314956 248301 650648 248537
rect 66975 248217 650648 248301
rect 66975 248174 269470 248217
rect 54198 248090 269470 248174
rect 54198 247854 66739 248090
rect 66975 247981 269470 248090
rect 269706 247981 284460 248217
rect 284696 247981 299460 248217
rect 299696 247981 314720 248217
rect 314956 247981 650648 248217
rect 66975 247897 650648 247981
rect 66975 247854 269470 247897
rect 54198 247770 269470 247854
rect 54198 247534 66739 247770
rect 66975 247661 269470 247770
rect 269706 247661 284460 247897
rect 284696 247661 299460 247897
rect 299696 247661 314720 247897
rect 314956 247661 650648 247897
rect 66975 247577 650648 247661
rect 66975 247534 269470 247577
rect 54198 247450 269470 247534
rect 54198 247214 66739 247450
rect 66975 247341 269470 247450
rect 269706 247341 284460 247577
rect 284696 247341 299460 247577
rect 299696 247341 314720 247577
rect 314956 247341 650648 247577
rect 66975 247257 650648 247341
rect 66975 247214 269470 247257
rect 54198 247130 269470 247214
rect 54198 246894 66739 247130
rect 66975 247021 269470 247130
rect 269706 247021 284460 247257
rect 284696 247021 299460 247257
rect 299696 247021 314720 247257
rect 314956 247021 650648 247257
rect 66975 246937 650648 247021
rect 66975 246894 269470 246937
rect 54198 246810 269470 246894
rect 54198 246574 66739 246810
rect 66975 246701 269470 246810
rect 269706 246701 284460 246937
rect 284696 246701 299460 246937
rect 299696 246701 314720 246937
rect 314956 246701 650648 246937
rect 66975 246579 650648 246701
rect 651204 249213 669890 249375
rect 651204 246737 667112 249213
rect 669588 246737 669890 249213
rect 651204 246579 669890 246737
rect 674156 249194 676452 249296
rect 674156 246718 674226 249194
rect 676382 246718 676452 249194
rect 674156 246616 676452 246718
rect 66975 246574 669890 246579
rect 54198 246466 669890 246574
rect 54198 219342 55398 246466
rect 56278 245375 654222 245466
rect 56278 245373 209170 245375
rect 56278 245370 199110 245373
rect 56278 245181 63863 245370
rect 56278 242705 56551 245181
rect 63187 245134 63863 245181
rect 64099 245137 199110 245370
rect 199346 245139 209170 245373
rect 209406 245373 654222 245375
rect 209406 245139 653679 245373
rect 199346 245137 653679 245139
rect 653915 245137 654222 245373
rect 64099 245134 654222 245137
rect 63187 245055 654222 245134
rect 63187 245053 209170 245055
rect 63187 245050 199110 245053
rect 63187 244814 63863 245050
rect 64099 244817 199110 245050
rect 199346 244819 209170 245053
rect 209406 245053 654222 245055
rect 209406 244819 653679 245053
rect 199346 244817 653679 244819
rect 653915 244817 654222 245053
rect 64099 244814 654222 244817
rect 63187 244735 654222 244814
rect 63187 244733 209170 244735
rect 63187 244730 199110 244733
rect 63187 244494 63863 244730
rect 64099 244497 199110 244730
rect 199346 244499 209170 244733
rect 209406 244733 654222 244735
rect 209406 244499 653679 244733
rect 199346 244497 653679 244499
rect 653915 244497 654222 244733
rect 64099 244494 654222 244497
rect 63187 244415 654222 244494
rect 63187 244413 209170 244415
rect 63187 244410 199110 244413
rect 63187 244174 63863 244410
rect 64099 244177 199110 244410
rect 199346 244179 209170 244413
rect 209406 244413 654222 244415
rect 209406 244179 653679 244413
rect 199346 244177 653679 244179
rect 653915 244177 654222 244413
rect 64099 244174 654222 244177
rect 63187 244095 654222 244174
rect 63187 244093 209170 244095
rect 63187 244090 199110 244093
rect 63187 243854 63863 244090
rect 64099 243857 199110 244090
rect 199346 243859 209170 244093
rect 209406 244093 654222 244095
rect 209406 243859 653679 244093
rect 199346 243857 653679 243859
rect 653915 243857 654222 244093
rect 64099 243854 654222 243857
rect 63187 243775 654222 243854
rect 63187 243773 209170 243775
rect 63187 243770 199110 243773
rect 63187 243534 63863 243770
rect 64099 243537 199110 243770
rect 199346 243539 209170 243773
rect 209406 243773 654222 243775
rect 209406 243539 653679 243773
rect 199346 243537 653679 243539
rect 653915 243537 654222 243773
rect 64099 243534 654222 243537
rect 63187 243455 654222 243534
rect 63187 243453 209170 243455
rect 63187 243450 199110 243453
rect 63187 243214 63863 243450
rect 64099 243217 199110 243450
rect 199346 243219 209170 243453
rect 209406 243453 654222 243455
rect 209406 243219 653679 243453
rect 199346 243217 653679 243219
rect 653915 243217 654222 243453
rect 64099 243214 654222 243217
rect 63187 243135 654222 243214
rect 63187 243133 209170 243135
rect 63187 243130 199110 243133
rect 63187 242894 63863 243130
rect 64099 242897 199110 243130
rect 199346 242899 209170 243133
rect 209406 243133 654222 243135
rect 209406 242899 653679 243133
rect 199346 242897 653679 242899
rect 653915 242897 654222 243133
rect 64099 242894 654222 242897
rect 63187 242815 654222 242894
rect 63187 242813 209170 242815
rect 63187 242810 199110 242813
rect 63187 242705 63863 242810
rect 56278 242574 63863 242705
rect 64099 242577 199110 242810
rect 199346 242579 209170 242813
rect 209406 242813 654222 242815
rect 209406 242579 653679 242813
rect 199346 242577 653679 242579
rect 653915 242577 654222 242813
rect 64099 242574 654222 242577
rect 56278 242466 654222 242574
rect 56278 241373 653306 241466
rect 56278 241366 194930 241373
rect 56278 241215 64813 241366
rect 56278 238739 56566 241215
rect 63202 241130 64813 241215
rect 65049 241137 194930 241366
rect 195166 241137 205050 241373
rect 205286 241371 653306 241373
rect 205286 241137 652721 241371
rect 65049 241135 652721 241137
rect 652957 241135 653306 241371
rect 65049 241130 653306 241135
rect 63202 241053 653306 241130
rect 63202 241046 194930 241053
rect 63202 240810 64813 241046
rect 65049 240817 194930 241046
rect 195166 240817 205050 241053
rect 205286 241051 653306 241053
rect 205286 240817 652721 241051
rect 65049 240815 652721 240817
rect 652957 240815 653306 241051
rect 65049 240810 653306 240815
rect 63202 240733 653306 240810
rect 63202 240726 194930 240733
rect 63202 240490 64813 240726
rect 65049 240497 194930 240726
rect 195166 240497 205050 240733
rect 205286 240731 653306 240733
rect 205286 240497 652721 240731
rect 65049 240495 652721 240497
rect 652957 240495 653306 240731
rect 65049 240490 653306 240495
rect 63202 240413 653306 240490
rect 63202 240406 194930 240413
rect 63202 240170 64813 240406
rect 65049 240177 194930 240406
rect 195166 240177 205050 240413
rect 205286 240411 653306 240413
rect 205286 240177 652721 240411
rect 65049 240175 652721 240177
rect 652957 240175 653306 240411
rect 65049 240170 653306 240175
rect 63202 240093 653306 240170
rect 63202 240086 194930 240093
rect 63202 239850 64813 240086
rect 65049 239857 194930 240086
rect 195166 239857 205050 240093
rect 205286 240091 653306 240093
rect 205286 239857 652721 240091
rect 65049 239855 652721 239857
rect 652957 239855 653306 240091
rect 65049 239850 653306 239855
rect 63202 239773 653306 239850
rect 63202 239766 194930 239773
rect 63202 239530 64813 239766
rect 65049 239537 194930 239766
rect 195166 239537 205050 239773
rect 205286 239771 653306 239773
rect 205286 239537 652721 239771
rect 65049 239535 652721 239537
rect 652957 239535 653306 239771
rect 65049 239530 653306 239535
rect 63202 239453 653306 239530
rect 63202 239446 194930 239453
rect 63202 239210 64813 239446
rect 65049 239217 194930 239446
rect 195166 239217 205050 239453
rect 205286 239451 653306 239453
rect 205286 239217 652721 239451
rect 65049 239215 652721 239217
rect 652957 239215 653306 239451
rect 65049 239210 653306 239215
rect 63202 239133 653306 239210
rect 63202 239126 194930 239133
rect 63202 238890 64813 239126
rect 65049 238897 194930 239126
rect 195166 238897 205050 239133
rect 205286 239131 653306 239133
rect 205286 238897 652721 239131
rect 65049 238895 652721 238897
rect 652957 238895 653306 239131
rect 65049 238890 653306 238895
rect 63202 238813 653306 238890
rect 63202 238806 194930 238813
rect 63202 238739 64813 238806
rect 56278 238570 64813 238739
rect 65049 238577 194930 238806
rect 195166 238577 205050 238813
rect 205286 238811 653306 238813
rect 205286 238577 652721 238811
rect 65049 238575 652721 238577
rect 652957 238575 653306 238811
rect 65049 238570 653306 238575
rect 56278 238466 653306 238570
rect 56288 237361 591390 237466
rect 56288 237221 140520 237361
rect 56288 234745 56455 237221
rect 63091 237125 140520 237221
rect 140756 237125 155600 237361
rect 155836 237125 170650 237361
rect 170886 237125 185660 237361
rect 185896 237125 215800 237361
rect 216036 237125 230850 237361
rect 231086 237125 245900 237361
rect 246136 237125 260950 237361
rect 261186 237125 276000 237361
rect 276236 237125 291050 237361
rect 291286 237125 306060 237361
rect 306296 237125 321250 237361
rect 321486 237125 336200 237361
rect 336436 237125 351350 237361
rect 351586 237125 366300 237361
rect 366536 237125 381150 237361
rect 381386 237125 396320 237361
rect 396556 237125 411450 237361
rect 411686 237125 426500 237361
rect 426736 237125 441550 237361
rect 441786 237125 456600 237361
rect 456836 237125 471650 237361
rect 471886 237125 486700 237361
rect 486936 237125 501750 237361
rect 501986 237125 591390 237361
rect 63091 237041 591390 237125
rect 63091 236805 140520 237041
rect 140756 236805 155600 237041
rect 155836 236805 170650 237041
rect 170886 236805 185660 237041
rect 185896 236805 215800 237041
rect 216036 236805 230850 237041
rect 231086 236805 245900 237041
rect 246136 236805 260950 237041
rect 261186 236805 276000 237041
rect 276236 236805 291050 237041
rect 291286 236805 306060 237041
rect 306296 236805 321250 237041
rect 321486 236805 336200 237041
rect 336436 236805 351350 237041
rect 351586 236805 366300 237041
rect 366536 236805 381150 237041
rect 381386 236805 396320 237041
rect 396556 236805 411450 237041
rect 411686 236805 426500 237041
rect 426736 236805 441550 237041
rect 441786 236805 456600 237041
rect 456836 236805 471650 237041
rect 471886 236805 486700 237041
rect 486936 236805 501750 237041
rect 501986 236805 591390 237041
rect 63091 236721 591390 236805
rect 63091 236485 140520 236721
rect 140756 236485 155600 236721
rect 155836 236485 170650 236721
rect 170886 236485 185660 236721
rect 185896 236485 215800 236721
rect 216036 236485 230850 236721
rect 231086 236485 245900 236721
rect 246136 236485 260950 236721
rect 261186 236485 276000 236721
rect 276236 236485 291050 236721
rect 291286 236485 306060 236721
rect 306296 236485 321250 236721
rect 321486 236485 336200 236721
rect 336436 236485 351350 236721
rect 351586 236485 366300 236721
rect 366536 236485 381150 236721
rect 381386 236485 396320 236721
rect 396556 236485 411450 236721
rect 411686 236485 426500 236721
rect 426736 236485 441550 236721
rect 441786 236485 456600 236721
rect 456836 236485 471650 236721
rect 471886 236485 486700 236721
rect 486936 236485 501750 236721
rect 501986 236485 591390 236721
rect 63091 236401 591390 236485
rect 63091 236165 140520 236401
rect 140756 236165 155600 236401
rect 155836 236165 170650 236401
rect 170886 236165 185660 236401
rect 185896 236165 215800 236401
rect 216036 236165 230850 236401
rect 231086 236165 245900 236401
rect 246136 236165 260950 236401
rect 261186 236165 276000 236401
rect 276236 236165 291050 236401
rect 291286 236165 306060 236401
rect 306296 236165 321250 236401
rect 321486 236165 336200 236401
rect 336436 236165 351350 236401
rect 351586 236165 366300 236401
rect 366536 236165 381150 236401
rect 381386 236165 396320 236401
rect 396556 236165 411450 236401
rect 411686 236165 426500 236401
rect 426736 236165 441550 236401
rect 441786 236165 456600 236401
rect 456836 236165 471650 236401
rect 471886 236165 486700 236401
rect 486936 236165 501750 236401
rect 501986 236165 591390 236401
rect 63091 236081 591390 236165
rect 63091 235845 140520 236081
rect 140756 235845 155600 236081
rect 155836 235845 170650 236081
rect 170886 235845 185660 236081
rect 185896 235845 215800 236081
rect 216036 235845 230850 236081
rect 231086 235845 245900 236081
rect 246136 235845 260950 236081
rect 261186 235845 276000 236081
rect 276236 235845 291050 236081
rect 291286 235845 306060 236081
rect 306296 235845 321250 236081
rect 321486 235845 336200 236081
rect 336436 235845 351350 236081
rect 351586 235845 366300 236081
rect 366536 235845 381150 236081
rect 381386 235845 396320 236081
rect 396556 235845 411450 236081
rect 411686 235845 426500 236081
rect 426736 235845 441550 236081
rect 441786 235845 456600 236081
rect 456836 235845 471650 236081
rect 471886 235845 486700 236081
rect 486936 235845 501750 236081
rect 501986 235845 591390 236081
rect 63091 235761 591390 235845
rect 63091 235525 140520 235761
rect 140756 235525 155600 235761
rect 155836 235525 170650 235761
rect 170886 235525 185660 235761
rect 185896 235525 215800 235761
rect 216036 235525 230850 235761
rect 231086 235525 245900 235761
rect 246136 235525 260950 235761
rect 261186 235525 276000 235761
rect 276236 235525 291050 235761
rect 291286 235525 306060 235761
rect 306296 235525 321250 235761
rect 321486 235525 336200 235761
rect 336436 235525 351350 235761
rect 351586 235525 366300 235761
rect 366536 235525 381150 235761
rect 381386 235525 396320 235761
rect 396556 235525 411450 235761
rect 411686 235525 426500 235761
rect 426736 235525 441550 235761
rect 441786 235525 456600 235761
rect 456836 235525 471650 235761
rect 471886 235525 486700 235761
rect 486936 235525 501750 235761
rect 501986 235525 591390 235761
rect 63091 235441 591390 235525
rect 63091 235205 140520 235441
rect 140756 235205 155600 235441
rect 155836 235205 170650 235441
rect 170886 235205 185660 235441
rect 185896 235205 215800 235441
rect 216036 235205 230850 235441
rect 231086 235205 245900 235441
rect 246136 235205 260950 235441
rect 261186 235205 276000 235441
rect 276236 235205 291050 235441
rect 291286 235205 306060 235441
rect 306296 235205 321250 235441
rect 321486 235205 336200 235441
rect 336436 235205 351350 235441
rect 351586 235205 366300 235441
rect 366536 235205 381150 235441
rect 381386 235205 396320 235441
rect 396556 235205 411450 235441
rect 411686 235205 426500 235441
rect 426736 235205 441550 235441
rect 441786 235205 456600 235441
rect 456836 235205 471650 235441
rect 471886 235205 486700 235441
rect 486936 235205 501750 235441
rect 501986 235205 591390 235441
rect 63091 235121 591390 235205
rect 63091 234885 140520 235121
rect 140756 234885 155600 235121
rect 155836 234885 170650 235121
rect 170886 234885 185660 235121
rect 185896 234885 215800 235121
rect 216036 234885 230850 235121
rect 231086 234885 245900 235121
rect 246136 234885 260950 235121
rect 261186 234885 276000 235121
rect 276236 234885 291050 235121
rect 291286 234885 306060 235121
rect 306296 234885 321250 235121
rect 321486 234885 336200 235121
rect 336436 234885 351350 235121
rect 351586 234885 366300 235121
rect 366536 234885 381150 235121
rect 381386 234885 396320 235121
rect 396556 234885 411450 235121
rect 411686 234885 426500 235121
rect 426736 234885 441550 235121
rect 441786 234885 456600 235121
rect 456836 234885 471650 235121
rect 471886 234885 486700 235121
rect 486936 234885 501750 235121
rect 501986 234885 591390 235121
rect 63091 234801 591390 234885
rect 63091 234745 140520 234801
rect 56288 234565 140520 234745
rect 140756 234565 155600 234801
rect 155836 234565 170650 234801
rect 170886 234565 185660 234801
rect 185896 234565 215800 234801
rect 216036 234565 230850 234801
rect 231086 234565 245900 234801
rect 246136 234565 260950 234801
rect 261186 234565 276000 234801
rect 276236 234565 291050 234801
rect 291286 234565 306060 234801
rect 306296 234565 321250 234801
rect 321486 234565 336200 234801
rect 336436 234565 351350 234801
rect 351586 234565 366300 234801
rect 366536 234565 381150 234801
rect 381386 234565 396320 234801
rect 396556 234565 411450 234801
rect 411686 234565 426500 234801
rect 426736 234565 441550 234801
rect 441786 234565 456600 234801
rect 456836 234565 471650 234801
rect 471886 234565 486700 234801
rect 486936 234565 501750 234801
rect 501986 234565 591390 234801
rect 56288 234466 591390 234565
rect 56296 233362 587374 233466
rect 56296 233211 133140 233362
rect 56296 230735 56554 233211
rect 62870 233126 133140 233211
rect 133376 233126 148190 233362
rect 148426 233126 163240 233362
rect 163476 233126 178290 233362
rect 178526 233126 193340 233362
rect 193576 233126 208390 233362
rect 208626 233126 223440 233362
rect 223676 233126 238490 233362
rect 238726 233126 253540 233362
rect 253776 233126 268590 233362
rect 268826 233126 283640 233362
rect 283876 233126 298690 233362
rect 298926 233126 313740 233362
rect 313976 233126 328790 233362
rect 329026 233126 343840 233362
rect 344076 233126 358890 233362
rect 359126 233126 373940 233362
rect 374176 233126 388990 233362
rect 389226 233126 404040 233362
rect 404276 233126 419090 233362
rect 419326 233126 434140 233362
rect 434376 233126 449190 233362
rect 449426 233126 464240 233362
rect 464476 233126 479290 233362
rect 479526 233126 494340 233362
rect 494576 233126 587374 233362
rect 62870 233042 587374 233126
rect 62870 232806 133140 233042
rect 133376 232806 148190 233042
rect 148426 232806 163240 233042
rect 163476 232806 178290 233042
rect 178526 232806 193340 233042
rect 193576 232806 208390 233042
rect 208626 232806 223440 233042
rect 223676 232806 238490 233042
rect 238726 232806 253540 233042
rect 253776 232806 268590 233042
rect 268826 232806 283640 233042
rect 283876 232806 298690 233042
rect 298926 232806 313740 233042
rect 313976 232806 328790 233042
rect 329026 232806 343840 233042
rect 344076 232806 358890 233042
rect 359126 232806 373940 233042
rect 374176 232806 388990 233042
rect 389226 232806 404040 233042
rect 404276 232806 419090 233042
rect 419326 232806 434140 233042
rect 434376 232806 449190 233042
rect 449426 232806 464240 233042
rect 464476 232806 479290 233042
rect 479526 232806 494340 233042
rect 494576 232806 587374 233042
rect 62870 232722 587374 232806
rect 62870 232486 133140 232722
rect 133376 232486 148190 232722
rect 148426 232486 163240 232722
rect 163476 232486 178290 232722
rect 178526 232486 193340 232722
rect 193576 232486 208390 232722
rect 208626 232486 223440 232722
rect 223676 232486 238490 232722
rect 238726 232486 253540 232722
rect 253776 232486 268590 232722
rect 268826 232486 283640 232722
rect 283876 232486 298690 232722
rect 298926 232486 313740 232722
rect 313976 232486 328790 232722
rect 329026 232486 343840 232722
rect 344076 232486 358890 232722
rect 359126 232486 373940 232722
rect 374176 232486 388990 232722
rect 389226 232486 404040 232722
rect 404276 232486 419090 232722
rect 419326 232486 434140 232722
rect 434376 232486 449190 232722
rect 449426 232486 464240 232722
rect 464476 232486 479290 232722
rect 479526 232486 494340 232722
rect 494576 232486 587374 232722
rect 62870 232402 587374 232486
rect 62870 232166 133140 232402
rect 133376 232166 148190 232402
rect 148426 232166 163240 232402
rect 163476 232166 178290 232402
rect 178526 232166 193340 232402
rect 193576 232166 208390 232402
rect 208626 232166 223440 232402
rect 223676 232166 238490 232402
rect 238726 232166 253540 232402
rect 253776 232166 268590 232402
rect 268826 232166 283640 232402
rect 283876 232166 298690 232402
rect 298926 232166 313740 232402
rect 313976 232166 328790 232402
rect 329026 232166 343840 232402
rect 344076 232166 358890 232402
rect 359126 232166 373940 232402
rect 374176 232166 388990 232402
rect 389226 232166 404040 232402
rect 404276 232166 419090 232402
rect 419326 232166 434140 232402
rect 434376 232166 449190 232402
rect 449426 232166 464240 232402
rect 464476 232166 479290 232402
rect 479526 232166 494340 232402
rect 494576 232166 587374 232402
rect 62870 232082 587374 232166
rect 62870 231846 133140 232082
rect 133376 231846 148190 232082
rect 148426 231846 163240 232082
rect 163476 231846 178290 232082
rect 178526 231846 193340 232082
rect 193576 231846 208390 232082
rect 208626 231846 223440 232082
rect 223676 231846 238490 232082
rect 238726 231846 253540 232082
rect 253776 231846 268590 232082
rect 268826 231846 283640 232082
rect 283876 231846 298690 232082
rect 298926 231846 313740 232082
rect 313976 231846 328790 232082
rect 329026 231846 343840 232082
rect 344076 231846 358890 232082
rect 359126 231846 373940 232082
rect 374176 231846 388990 232082
rect 389226 231846 404040 232082
rect 404276 231846 419090 232082
rect 419326 231846 434140 232082
rect 434376 231846 449190 232082
rect 449426 231846 464240 232082
rect 464476 231846 479290 232082
rect 479526 231846 494340 232082
rect 494576 231846 587374 232082
rect 62870 231762 587374 231846
rect 62870 231526 133140 231762
rect 133376 231526 148190 231762
rect 148426 231526 163240 231762
rect 163476 231526 178290 231762
rect 178526 231526 193340 231762
rect 193576 231526 208390 231762
rect 208626 231526 223440 231762
rect 223676 231526 238490 231762
rect 238726 231526 253540 231762
rect 253776 231526 268590 231762
rect 268826 231526 283640 231762
rect 283876 231526 298690 231762
rect 298926 231526 313740 231762
rect 313976 231526 328790 231762
rect 329026 231526 343840 231762
rect 344076 231526 358890 231762
rect 359126 231526 373940 231762
rect 374176 231526 388990 231762
rect 389226 231526 404040 231762
rect 404276 231526 419090 231762
rect 419326 231526 434140 231762
rect 434376 231526 449190 231762
rect 449426 231526 464240 231762
rect 464476 231526 479290 231762
rect 479526 231526 494340 231762
rect 494576 231526 587374 231762
rect 62870 231442 587374 231526
rect 62870 231206 133140 231442
rect 133376 231206 148190 231442
rect 148426 231206 163240 231442
rect 163476 231206 178290 231442
rect 178526 231206 193340 231442
rect 193576 231206 208390 231442
rect 208626 231206 223440 231442
rect 223676 231206 238490 231442
rect 238726 231206 253540 231442
rect 253776 231206 268590 231442
rect 268826 231206 283640 231442
rect 283876 231206 298690 231442
rect 298926 231206 313740 231442
rect 313976 231206 328790 231442
rect 329026 231206 343840 231442
rect 344076 231206 358890 231442
rect 359126 231206 373940 231442
rect 374176 231206 388990 231442
rect 389226 231206 404040 231442
rect 404276 231206 419090 231442
rect 419326 231206 434140 231442
rect 434376 231206 449190 231442
rect 449426 231206 464240 231442
rect 464476 231206 479290 231442
rect 479526 231206 494340 231442
rect 494576 231206 587374 231442
rect 62870 231122 587374 231206
rect 62870 230886 133140 231122
rect 133376 230886 148190 231122
rect 148426 230886 163240 231122
rect 163476 230886 178290 231122
rect 178526 230886 193340 231122
rect 193576 230886 208390 231122
rect 208626 230886 223440 231122
rect 223676 230886 238490 231122
rect 238726 230886 253540 231122
rect 253776 230886 268590 231122
rect 268826 230886 283640 231122
rect 283876 230886 298690 231122
rect 298926 230886 313740 231122
rect 313976 230886 328790 231122
rect 329026 230886 343840 231122
rect 344076 230886 358890 231122
rect 359126 230886 373940 231122
rect 374176 230886 388990 231122
rect 389226 230886 404040 231122
rect 404276 230886 419090 231122
rect 419326 230886 434140 231122
rect 434376 230886 449190 231122
rect 449426 230886 464240 231122
rect 464476 230886 479290 231122
rect 479526 230886 494340 231122
rect 494576 230886 587374 231122
rect 62870 230802 587374 230886
rect 62870 230735 133140 230802
rect 56296 230566 133140 230735
rect 133376 230566 148190 230802
rect 148426 230566 163240 230802
rect 163476 230566 178290 230802
rect 178526 230566 193340 230802
rect 193576 230566 208390 230802
rect 208626 230566 223440 230802
rect 223676 230566 238490 230802
rect 238726 230566 253540 230802
rect 253776 230566 268590 230802
rect 268826 230566 283640 230802
rect 283876 230566 298690 230802
rect 298926 230566 313740 230802
rect 313976 230566 328790 230802
rect 329026 230566 343840 230802
rect 344076 230566 358890 230802
rect 359126 230566 373940 230802
rect 374176 230566 388990 230802
rect 389226 230566 404040 230802
rect 404276 230566 419090 230802
rect 419326 230566 434140 230802
rect 434376 230566 449190 230802
rect 449426 230566 464240 230802
rect 464476 230566 479290 230802
rect 479526 230566 494340 230802
rect 494576 230566 587374 230802
rect 56296 230466 587374 230566
rect 584374 212271 587374 230466
rect 47836 209858 53232 210498
rect 574646 209858 582910 210498
rect 47836 184498 50836 209858
rect 582270 208502 582910 209858
rect 584374 209795 584610 212271
rect 587086 209795 587374 212271
rect 582270 208302 583742 208502
rect 582270 208066 582400 208302
rect 582636 208066 582720 208302
rect 582956 208066 583040 208302
rect 583276 208066 583360 208302
rect 583596 208066 583742 208302
rect 582270 207862 583742 208066
rect 584374 197721 587374 209795
rect 584374 197498 584783 197721
rect 51344 197312 53216 197498
rect 51344 197076 51573 197312
rect 51809 197076 51893 197312
rect 52129 197076 53216 197312
rect 51344 196858 53216 197076
rect 574646 197165 584783 197498
rect 586939 197165 587374 197721
rect 574646 196858 587374 197165
rect 47836 183858 53212 184498
rect 574646 184290 582910 184498
rect 574646 184054 582204 184290
rect 582440 184054 582524 184290
rect 582760 184054 582910 184290
rect 574646 183858 582910 184054
rect 41768 176505 45768 176874
rect 41768 173389 42087 176505
rect 45523 173389 45768 176505
rect 41768 171294 45768 173389
rect 41768 171058 42857 171294
rect 43093 171058 43177 171294
rect 43413 171058 43497 171294
rect 43733 171058 43817 171294
rect 44053 171058 44137 171294
rect 44373 171058 44457 171294
rect 44693 171058 44777 171294
rect 45013 171058 45097 171294
rect 45333 171058 45417 171294
rect 45653 171058 45768 171294
rect 41768 145300 45768 171058
rect 47836 166788 50836 183858
rect 584374 171498 587374 196858
rect 51246 171298 53240 171498
rect 51246 171062 51465 171298
rect 51701 171062 51785 171298
rect 52021 171062 53240 171298
rect 51246 170858 53240 171062
rect 574646 170858 587374 171498
rect 41768 145064 42871 145300
rect 43107 145064 43191 145300
rect 43427 145064 43511 145300
rect 43747 145064 43831 145300
rect 44067 145064 44151 145300
rect 44387 145064 44471 145300
rect 44707 145064 44791 145300
rect 45027 145064 45111 145300
rect 45347 145064 45431 145300
rect 45667 145064 45768 145300
rect 41768 119296 45768 145064
rect 41768 119060 42861 119296
rect 43097 119060 43181 119296
rect 43417 119060 43501 119296
rect 43737 119060 43821 119296
rect 44057 119060 44141 119296
rect 44377 119060 44461 119296
rect 44697 119060 44781 119296
rect 45017 119060 45101 119296
rect 45337 119060 45421 119296
rect 45657 119060 45768 119296
rect 41768 93294 45768 119060
rect 41768 93058 42857 93294
rect 43093 93058 43177 93294
rect 43413 93058 43497 93294
rect 43733 93058 43817 93294
rect 44053 93058 44137 93294
rect 44373 93058 44457 93294
rect 44693 93058 44777 93294
rect 45013 93058 45097 93294
rect 45333 93058 45417 93294
rect 45653 93058 45768 93294
rect 41768 82672 45768 93058
rect 41768 78276 42091 82672
rect 45527 78276 45768 82672
rect 41768 72768 45768 78276
rect 41768 68372 42067 72768
rect 45503 68372 45768 72768
rect 41768 67288 45768 68372
rect 41768 67052 42095 67288
rect 42331 67052 42415 67288
rect 42651 67052 42735 67288
rect 42971 67052 43055 67288
rect 43291 67052 43375 67288
rect 43611 67052 43695 67288
rect 43931 67052 44015 67288
rect 44251 67052 44335 67288
rect 44571 67052 44655 67288
rect 44891 67052 44975 67288
rect 45211 67052 45295 67288
rect 45531 67052 45768 67288
rect 41768 51914 45768 67052
rect 41768 48478 42080 51914
rect 45516 48478 45768 51914
rect 41768 48074 45768 48478
rect 46836 158498 50836 166788
rect 584374 167081 587374 170858
rect 584374 166525 584783 167081
rect 586939 166525 587374 167081
rect 46836 157858 53220 158498
rect 574646 158294 582910 158498
rect 574646 158058 580242 158294
rect 580478 158058 580562 158294
rect 580798 158058 580882 158294
rect 581118 158058 581202 158294
rect 581438 158058 581522 158294
rect 581758 158058 581842 158294
rect 582078 158058 582162 158294
rect 582398 158058 582482 158294
rect 582718 158058 582910 158294
rect 574646 157858 582910 158058
rect 46836 132498 50836 157858
rect 584374 145498 587374 166525
rect 51178 145290 53266 145498
rect 51178 145054 51399 145290
rect 51635 145054 51719 145290
rect 51955 145054 53266 145290
rect 51178 144858 53266 145054
rect 574646 144858 587374 145498
rect 584374 136441 587374 144858
rect 584374 135885 584783 136441
rect 586939 135885 587374 136441
rect 46836 131858 53206 132498
rect 574646 132288 582910 132498
rect 574646 132052 580252 132288
rect 580488 132052 580572 132288
rect 580808 132052 580892 132288
rect 581128 132052 581212 132288
rect 581448 132052 581532 132288
rect 581768 132052 581852 132288
rect 582088 132052 582172 132288
rect 582408 132052 582492 132288
rect 582728 132052 582910 132288
rect 574646 131858 582910 132052
rect 46836 106498 50836 131858
rect 584374 119498 587374 135885
rect 51178 119296 53266 119498
rect 51178 119060 51395 119296
rect 51631 119060 51715 119296
rect 51951 119060 53266 119296
rect 51178 118858 53266 119060
rect 574646 118858 587374 119498
rect 46836 105858 53222 106498
rect 574646 106294 582910 106498
rect 574646 106058 580254 106294
rect 580490 106058 580574 106294
rect 580810 106058 580894 106294
rect 581130 106058 581214 106294
rect 581450 106058 581534 106294
rect 581770 106058 581854 106294
rect 582090 106058 582174 106294
rect 582410 106058 582494 106294
rect 582730 106058 582910 106294
rect 574646 105858 582910 106058
rect 46836 80498 50836 105858
rect 584374 105521 587374 118858
rect 584374 104965 584783 105521
rect 586939 104965 587374 105521
rect 584374 93498 587374 104965
rect 51178 93292 53266 93498
rect 51178 93056 51399 93292
rect 51635 93056 51719 93292
rect 51955 93056 53266 93292
rect 51178 92858 53266 93056
rect 574646 92858 587374 93498
rect 46836 79858 53168 80498
rect 574646 80304 582910 80498
rect 574646 80068 580248 80304
rect 580484 80068 580568 80304
rect 580804 80068 580888 80304
rect 581124 80068 581208 80304
rect 581444 80068 581528 80304
rect 581764 80068 581848 80304
rect 582084 80068 582168 80304
rect 582404 80068 582488 80304
rect 582724 80068 582910 80304
rect 574646 79858 582910 80068
rect 46836 46788 50836 79858
rect 584374 67498 587374 92858
rect 51362 67294 53172 67498
rect 51362 67058 51597 67294
rect 51833 67058 51917 67294
rect 52153 67058 53172 67294
rect 51362 66858 53172 67058
rect 574754 66858 587374 67498
rect 584374 52222 587374 66858
rect 54374 51880 587374 52222
rect 54374 48444 54650 51880
rect 58086 50592 587374 51880
rect 58086 50036 143423 50592
rect 144619 50036 587374 50592
rect 58086 48444 587374 50036
rect 54374 48222 587374 48444
rect 588390 226084 591390 234466
rect 588390 224192 640366 226084
rect 648608 225872 651358 226192
rect 588390 224082 641998 224192
rect 588390 208302 591390 224082
rect 639466 223872 641998 224082
rect 650224 222192 651358 225872
rect 648640 221872 651358 222192
rect 650224 212504 651358 221872
rect 593252 212271 669426 212504
rect 593252 209795 593464 212271
rect 595940 212234 669426 212271
rect 595940 209795 627303 212234
rect 593252 209758 627303 209795
rect 627859 209758 669426 212234
rect 593252 209504 669426 209758
rect 588390 208066 588493 208302
rect 588729 208066 588813 208302
rect 589049 208066 589133 208302
rect 589369 208066 589453 208302
rect 589689 208066 589773 208302
rect 590009 208066 590093 208302
rect 590329 208066 590413 208302
rect 590649 208066 590733 208302
rect 590969 208066 591053 208302
rect 591289 208066 591390 208302
rect 588390 184286 591390 208066
rect 666426 197528 669426 209504
rect 591976 197483 593594 197528
rect 591976 197247 592038 197483
rect 592274 197247 592358 197483
rect 592594 197247 592678 197483
rect 592914 197247 593594 197483
rect 591976 197208 593594 197247
rect 665238 197208 669426 197528
rect 588390 184050 588493 184286
rect 588729 184050 588813 184286
rect 589049 184050 589133 184286
rect 589369 184050 589453 184286
rect 589689 184050 589773 184286
rect 590009 184050 590093 184286
rect 590329 184050 590413 184286
rect 590649 184050 590733 184286
rect 590969 184050 591053 184286
rect 591289 184050 591390 184286
rect 588390 182210 591390 184050
rect 588390 181890 593594 182210
rect 588390 158298 591390 181890
rect 666426 166892 669426 197208
rect 591952 166855 593594 166892
rect 591952 166619 592021 166855
rect 592257 166619 592341 166855
rect 592577 166619 592661 166855
rect 592897 166619 593594 166855
rect 591952 166572 593594 166619
rect 665206 166572 669426 166892
rect 588390 158062 588467 158298
rect 588703 158062 588787 158298
rect 589023 158062 589107 158298
rect 589343 158062 589427 158298
rect 589663 158062 589747 158298
rect 589983 158062 590067 158298
rect 590303 158062 590387 158298
rect 590623 158062 590707 158298
rect 590943 158062 591027 158298
rect 591263 158062 591390 158298
rect 588390 151574 591390 158062
rect 588390 151254 593594 151574
rect 588390 132282 591390 151254
rect 666426 136256 669426 166572
rect 591940 136215 593594 136256
rect 591940 135979 592011 136215
rect 592247 135979 592331 136215
rect 592567 135979 592651 136215
rect 592887 135979 593594 136215
rect 591940 135936 593594 135979
rect 665164 135936 669426 136256
rect 588390 132046 588493 132282
rect 588729 132046 588813 132282
rect 589049 132046 589133 132282
rect 589369 132046 589453 132282
rect 589689 132046 589773 132282
rect 590009 132046 590093 132282
rect 590329 132046 590413 132282
rect 590649 132046 590733 132282
rect 590969 132046 591053 132282
rect 591289 132046 591390 132282
rect 588390 120938 591390 132046
rect 588390 120618 593610 120938
rect 588390 106294 591390 120618
rect 588390 106058 588497 106294
rect 588733 106058 588817 106294
rect 589053 106058 589137 106294
rect 589373 106058 589457 106294
rect 589693 106058 589777 106294
rect 590013 106058 590097 106294
rect 590333 106058 590417 106294
rect 590653 106058 590737 106294
rect 590973 106058 591057 106294
rect 591293 106058 591390 106294
rect 588390 98956 591390 106058
rect 666426 105620 669426 135936
rect 591940 105578 593594 105620
rect 591940 105342 592023 105578
rect 592259 105342 592343 105578
rect 592579 105342 592663 105578
rect 592899 105342 593594 105578
rect 591940 105300 593594 105342
rect 665176 105300 669426 105620
rect 588390 98665 657728 98956
rect 588390 98603 627823 98665
rect 588390 96127 597012 98603
rect 597888 96189 627823 98603
rect 628699 98521 657728 98665
rect 628699 96685 636259 98521
rect 636815 96685 657728 98521
rect 628699 96189 657728 96685
rect 597888 96127 657728 96189
rect 588390 95956 657728 96127
rect 588390 80306 591390 95956
rect 624824 89474 627824 95956
rect 643544 93474 646544 93588
rect 641906 93154 646544 93474
rect 624824 89154 629362 89474
rect 624824 89012 627824 89154
rect 588390 80070 588491 80306
rect 588727 80070 588811 80306
rect 589047 80070 589131 80306
rect 589367 80070 589451 80306
rect 589687 80070 589771 80306
rect 590007 80070 590091 80306
rect 590327 80070 590411 80306
rect 590647 80070 590731 80306
rect 590967 80070 591051 80306
rect 591287 80070 591390 80306
rect 588390 47188 591390 80070
rect 625618 75868 627034 89012
rect 643544 85474 646544 93154
rect 650994 92590 653994 95956
rect 666426 93406 669426 105300
rect 662522 93086 669426 93406
rect 650994 92270 657754 92590
rect 650994 90958 653994 92270
rect 666426 91774 669426 93086
rect 662484 91454 669426 91774
rect 650994 90638 657784 90958
rect 650994 90522 653994 90638
rect 666426 90142 669426 91454
rect 662504 89822 669426 90142
rect 641968 85154 646544 85474
rect 643544 81082 646544 85154
rect 666426 81082 669426 89822
rect 632002 80816 669426 81082
rect 632002 80629 640232 80816
rect 632002 78473 632254 80629
rect 632810 78473 640232 80629
rect 632002 78340 640232 78473
rect 640788 78340 669426 80816
rect 632002 78082 669426 78340
rect 645256 77268 647084 78082
rect 629786 77215 647084 77268
rect 629786 77207 642323 77215
rect 629786 77193 633031 77207
rect 629786 76957 629919 77193
rect 630155 76971 633031 77193
rect 633267 77203 642323 77207
rect 633267 76971 636121 77203
rect 630155 76967 636121 76971
rect 636357 76967 639215 77203
rect 639451 76979 642323 77203
rect 642559 76979 647084 77215
rect 639451 76967 647084 76979
rect 630155 76957 647084 76967
rect 629786 76895 647084 76957
rect 629786 76887 642323 76895
rect 629786 76873 633031 76887
rect 629786 76637 629919 76873
rect 630155 76651 633031 76873
rect 633267 76883 642323 76887
rect 633267 76651 636121 76883
rect 630155 76647 636121 76651
rect 636357 76647 639215 76883
rect 639451 76659 642323 76883
rect 642559 76659 647084 76895
rect 639451 76647 647084 76659
rect 630155 76637 647084 76647
rect 629786 76575 647084 76637
rect 629786 76567 642323 76575
rect 629786 76553 633031 76567
rect 629786 76317 629919 76553
rect 630155 76331 633031 76553
rect 633267 76563 642323 76567
rect 633267 76331 636121 76563
rect 630155 76327 636121 76331
rect 636357 76327 639215 76563
rect 639451 76339 642323 76563
rect 642559 76339 647084 76575
rect 639451 76327 647084 76339
rect 630155 76317 647084 76327
rect 629786 76268 647084 76317
rect 625618 75817 644188 75868
rect 625618 75799 643879 75817
rect 625618 75795 637673 75799
rect 625618 75791 634565 75795
rect 625618 75555 631471 75791
rect 631707 75559 634565 75791
rect 634801 75563 637673 75795
rect 637909 75791 643879 75799
rect 637909 75563 640777 75791
rect 634801 75559 640777 75563
rect 631707 75555 640777 75559
rect 641013 75581 643879 75791
rect 644115 75581 644188 75817
rect 641013 75555 644188 75581
rect 625618 75497 644188 75555
rect 625618 75479 643879 75497
rect 625618 75475 637673 75479
rect 625618 75471 634565 75475
rect 625618 75235 631471 75471
rect 631707 75239 634565 75471
rect 634801 75243 637673 75475
rect 637909 75471 643879 75479
rect 637909 75243 640777 75471
rect 634801 75239 640777 75243
rect 631707 75235 640777 75239
rect 641013 75261 643879 75471
rect 644115 75261 644188 75497
rect 641013 75235 644188 75261
rect 625618 75177 644188 75235
rect 625618 75159 643879 75177
rect 625618 75155 637673 75159
rect 625618 75151 634565 75155
rect 625618 74915 631471 75151
rect 631707 74919 634565 75151
rect 634801 74923 637673 75155
rect 637909 75151 643879 75159
rect 637909 74923 640777 75151
rect 634801 74919 640777 74923
rect 631707 74915 640777 74919
rect 641013 74941 643879 75151
rect 644115 74941 644188 75177
rect 641013 74915 644188 74941
rect 625618 74868 644188 74915
rect 625618 71796 626418 74868
rect 646284 73486 647084 76268
rect 645536 73166 647084 73486
rect 625618 71476 626968 71796
rect 625618 68416 626418 71476
rect 646284 70106 647084 73166
rect 645502 69786 647084 70106
rect 625618 68096 626846 68416
rect 646284 66726 647084 69786
rect 645624 66406 647084 66726
rect 666426 47274 669426 78082
rect 588390 47010 649668 47188
rect 588390 46788 648289 47010
rect 46836 46774 648289 46788
rect 648525 46774 648609 47010
rect 648845 46774 648929 47010
rect 649165 46774 649249 47010
rect 649485 46774 649668 47010
rect 666426 47038 666522 47274
rect 666758 47038 666842 47274
rect 667078 47038 667162 47274
rect 667398 47038 667482 47274
rect 667718 47038 667802 47274
rect 668038 47038 668122 47274
rect 668358 47038 668442 47274
rect 668678 47038 668762 47274
rect 668998 47038 669082 47274
rect 669318 47038 669426 47274
rect 666426 46978 669426 47038
rect 46836 46621 649668 46774
rect 46836 46607 251477 46621
rect 46836 45194 241825 46607
rect 46836 44318 141528 45194
rect 142724 44318 241825 45194
rect 46836 42851 241825 44318
rect 245901 42865 251477 46607
rect 255553 46588 649668 46621
rect 255553 42865 591396 46588
rect 245901 42851 591396 42865
rect 46836 42788 591396 42851
use gpio_control_power_routing  gpio_control_power_routing_0
timestamp 1493648132
transform 1 0 -10 0 1 728600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_1
timestamp 1493648132
transform 1 0 -10 0 1 602800
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_2
timestamp 1493648132
transform 1 0 -10 0 1 559600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_3
timestamp 1493648132
transform 1 0 -10 0 1 516400
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_4
timestamp 1493648132
transform 1 0 -10 0 1 473200
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_5
timestamp 1493648132
transform 1 0 -10 0 1 430000
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_6
timestamp 1493648132
transform 1 0 -10 0 1 386800
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_7
timestamp 1493648132
transform 1 0 -10 0 1 343600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_8
timestamp 1493648132
transform 1 0 -10 0 1 216000
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_9
timestamp 1493648132
transform 1 0 -10 0 1 172800
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_10
timestamp 1493648132
transform 1 0 -10 0 1 129600
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_11
timestamp 1493648132
transform 1 0 -10 0 1 86400
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_12
timestamp 1493648132
transform 1 0 -10 0 1 43200
box 6032 203748 55470 221470
use gpio_control_power_routing  gpio_control_power_routing_13
timestamp 1493648132
transform 1 0 -10 0 1 0
box 6032 203748 55470 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_0
timestamp 1493648132
transform -1 0 717836 0 1 725000
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_1
timestamp 1493648132
transform -1 0 717846 0 1 456400
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_2
timestamp 1493648132
transform -1 0 717846 0 1 501600
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_3
timestamp 1493648132
transform -1 0 717846 0 1 546600
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_4
timestamp 1493648132
transform -1 0 717846 0 1 321200
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_5
timestamp 1493648132
transform -1 0 717846 0 1 366200
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_6
timestamp 1493648132
transform -1 0 717846 0 1 411400
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_7
timestamp 1493648132
transform -1 0 717846 0 1 189000
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_8
timestamp 1493648132
transform -1 0 717846 0 1 277200
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_9
timestamp 1493648132
transform -1 0 717846 0 1 53800
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_10
timestamp 1493648132
transform -1 0 717846 0 1 98800
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_11
timestamp 1493648132
transform -1 0 717846 0 1 143800
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_12
timestamp 1493648132
transform -1 0 717846 0 1 -81600
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_13
timestamp 1493648132
transform -1 0 717846 0 1 -36400
box 6032 203748 46226 221470
use gpio_control_power_routing_right  gpio_control_power_routing_right_14
timestamp 1493648132
transform -1 0 717846 0 1 8600
box 6032 203748 46226 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_0
timestamp 1493648132
transform 0 1 346600 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_1
timestamp 1493648132
transform 0 1 295200 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_2
timestamp 1493648132
transform 0 1 218200 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_3
timestamp 1493648132
transform 0 1 150800 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_4
timestamp 1493648132
transform 0 1 100400 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_5
timestamp 1493648132
transform 0 1 48800 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_6
timestamp 1493648132
transform 0 1 -2600 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_7
timestamp 1493648132
transform 0 1 -54000 -1 0 1037728
box 6032 203748 43870 221470
use gpio_control_power_routing_top  gpio_control_power_routing_top_8
timestamp 1493648132
transform 0 1 -105400 -1 0 1037728
box 6032 203748 43870 221470
<< labels >>
flabel metal5 s 576480 230750 581228 233134 0 FreeSans 20000 0 0 0 vccd_core
port 1 nsew
flabel metal5 s 576522 234770 581540 236910 0 FreeSans 20000 0 0 0 vssd_core
port 2 nsew
flabel metal5 s 118216 238830 126118 240864 0 FreeSans 20000 0 0 0 vccd2_core
port 3 nsew
flabel metal5 s 118126 242838 126088 244986 0 FreeSans 20000 0 0 0 vssd2_core
port 4 nsew
flabel metal5 s 117918 254572 125876 257076 0 FreeSans 20000 0 0 0 vdda2_core
port 5 nsew
flabel metal5 s 117918 258660 125876 261164 0 FreeSans 20000 0 0 0 vssa2_core
port 6 nsew
flabel metal5 s 118024 250550 126042 253308 0 FreeSans 20000 0 0 0 vssd1_core
port 7 nsew
flabel metal5 s 118160 246638 126178 249396 0 FreeSans 20000 0 0 0 vccd1_core
port 8 nsew
flabel metal5 s 117852 266620 125870 269378 0 FreeSans 20000 0 0 0 vssa1_core
port 9 nsew
flabel metal5 s 117950 262574 125968 265332 0 FreeSans 20000 0 0 0 vdda1_core
port 10 nsew
flabel metal5 s 120522 234770 125540 236910 0 FreeSans 20000 0 0 0 vssd_core
port 2 nsew
flabel metal5 s 120480 230750 125228 233134 0 FreeSans 20000 0 0 0 vccd_core
port 1 nsew
flabel metal5 s 54316 219436 55324 219998 0 FreeSans 2000 0 0 0 vccd1_core
port 8 nsew
flabel metal5 s 52692 217826 53700 218388 0 FreeSans 2000 0 0 0 vssd1_core
port 7 nsew
flabel metal5 s 621960 246802 629984 249230 0 FreeSans 20000 0 0 0 vccd1_core
port 8 nsew
flabel metal5 s 621948 250708 629990 253036 0 FreeSans 20000 0 0 0 vssd1_core
port 7 nsew
flabel metal5 s 621550 262640 629508 265144 0 FreeSans 20000 0 0 0 vdda1_core
port 10 nsew
flabel metal5 s 621514 266692 629472 269196 0 FreeSans 20000 0 0 0 vssa1_core
port 9 nsew
flabel metal5 s 42966 171382 45564 172780 0 FreeSans 4000 0 0 0 vccd_core
port 1 nsew
flabel metal5 s 664092 267180 666518 267904 0 FreeSans 4000 0 0 0 vssa1_core
port 9 nsew
flabel metal5 s 667280 263142 669706 263866 0 FreeSans 4000 0 0 0 vdda1_core
port 10 nsew
flabel metal5 s 634330 96284 638114 98514 0 FreeSans 20000 0 0 0 vssd_core
port 2 nsew
flabel metal5 s 633452 78554 637236 80784 0 FreeSans 20000 0 0 0 vccd_core
port 1 nsew
flabel metal5 s 47904 265444 49660 265998 0 FreeSans 4000 0 0 0 vssa2_core
port 6 nsew
flabel metal5 s 50338 265444 52094 265998 0 FreeSans 4000 0 0 0 vdda2_core
port 5 nsew
flabel metal5 s 621512 258708 630212 261250 0 FreeSans 20000 0 0 0 vssa2_core
port 6 nsew
flabel metal5 s 621598 254668 630298 257210 0 FreeSans 20000 0 0 0 vdda2_core
port 5 nsew
flabel metal5 s 621936 242776 630636 245318 0 FreeSans 20000 0 0 0 vssd2_core
port 4 nsew
flabel metal5 s 621794 238736 630494 241278 0 FreeSans 20000 0 0 0 vccd2_core
port 3 nsew
flabel metal5 s 627056 74976 628118 75674 0 FreeSans 6000 0 0 0 vssd_core
port 2 nsew
flabel metal5 s 644752 76466 645814 77164 0 FreeSans 6000 0 0 0 vccd_core
port 1 nsew
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
